magic
tech scmos
magscale 1 2
timestamp 1727514457
<< error_s >>
rect 10 5984 6070 5996
rect 10 5724 6070 5736
rect 10 5464 6070 5476
rect 10 5204 6070 5216
rect 10 4944 6070 4956
rect 10 4684 6070 4696
rect 10 4424 6070 4436
rect 10 4164 6070 4176
rect 10 3904 6070 3916
rect 10 3644 6070 3656
rect 10 3384 6070 3396
rect 10 3124 6070 3136
rect 10 2864 6070 2876
rect 10 2604 6070 2616
rect 10 2344 6070 2356
rect 10 2084 6070 2096
rect 10 1824 6070 1836
rect 10 1564 6070 1576
rect 10 1304 6070 1316
rect 10 1044 6070 1056
rect 10 784 6070 796
rect 10 524 6070 536
rect 10 264 6070 276
rect 10 4 6070 16
<< nwell >>
rect 4937 5172 4943 5174
<< metal1 >>
rect -57 5738 3 5998
rect 6050 5982 6137 5998
rect 326 5903 340 5907
rect 326 5893 343 5903
rect 337 5767 343 5893
rect 517 5807 523 5953
rect 540 5903 553 5907
rect 537 5893 553 5903
rect 537 5767 543 5893
rect 677 5807 683 5873
rect 697 5767 703 5893
rect 857 5807 863 5873
rect 2557 5847 2563 5893
rect 2677 5767 2683 5913
rect 2717 5767 2723 5893
rect 3437 5847 3443 5933
rect 3597 5847 3603 5933
rect 3597 5767 3603 5833
rect 3877 5767 3883 5833
rect 4737 5787 4743 5933
rect 4917 5787 4923 5933
rect 5117 5927 5123 5953
rect 5257 5767 5263 5893
rect 5277 5787 5283 5953
rect 5417 5787 5423 5813
rect 5437 5767 5443 5953
rect 3586 5757 3603 5767
rect 3586 5753 3600 5757
rect -57 5722 30 5738
rect -57 5218 3 5722
rect 3706 5693 3707 5700
rect 657 5507 663 5613
rect 837 5527 843 5613
rect 1377 5607 1383 5673
rect 1677 5647 1683 5693
rect 2657 5667 2663 5693
rect 2657 5627 2663 5653
rect 2957 5627 2963 5693
rect 2837 5507 2843 5553
rect 3137 5527 3143 5653
rect 3257 5507 3263 5693
rect 3693 5687 3707 5693
rect 3693 5680 3713 5687
rect 3697 5677 3713 5680
rect 3700 5673 3713 5677
rect 3577 5527 3583 5613
rect 4337 5547 4343 5693
rect 4737 5547 4743 5693
rect 3566 5517 3583 5527
rect 3566 5513 3580 5517
rect 4897 5507 4903 5533
rect 4917 5528 4923 5633
rect 5057 5567 5063 5693
rect 5237 5507 5243 5673
rect 5377 5507 5383 5653
rect 5677 5507 5683 5693
rect 5817 5587 5823 5613
rect 6057 5507 6063 5533
rect 5667 5497 5683 5507
rect 5667 5493 5680 5497
rect 6077 5478 6137 5982
rect 6050 5462 6137 5478
rect 197 5267 203 5433
rect 677 5247 683 5413
rect 837 5327 843 5433
rect 1097 5327 1103 5433
rect 1097 5287 1103 5313
rect 1117 5247 1123 5373
rect 1417 5267 1423 5393
rect 1717 5287 1723 5433
rect 1857 5247 1863 5373
rect 2317 5247 2323 5273
rect 2757 5267 2763 5373
rect 2777 5247 2783 5293
rect 2797 5267 2803 5433
rect 2917 5267 2923 5313
rect 2937 5247 2943 5413
rect 3117 5327 3123 5433
rect 3437 5287 3443 5393
rect 3457 5267 3463 5293
rect 3617 5247 3623 5413
rect 4077 5387 4083 5433
rect 4097 5267 4103 5413
rect 4237 5267 4243 5393
rect 4257 5307 4263 5333
rect 4397 5327 4403 5413
rect 4677 5267 4683 5393
rect 4697 5247 4703 5433
rect 4837 5247 4843 5413
rect 4957 5287 4963 5433
rect 5297 5247 5303 5313
rect 5737 5247 5743 5433
rect 5997 5247 6003 5373
rect 6017 5287 6023 5433
rect 1846 5237 1863 5247
rect 1846 5233 1860 5237
rect 5287 5237 5303 5247
rect 5287 5233 5300 5237
rect -57 5202 30 5218
rect -57 4698 3 5202
rect 1400 5163 1413 5167
rect 1397 5153 1413 5163
rect 657 4987 663 5133
rect 797 4987 803 5053
rect 977 4987 983 5053
rect 1117 5027 1123 5153
rect 1257 5107 1263 5133
rect 1137 4987 1143 5053
rect 1397 4987 1403 5153
rect 1577 5047 1583 5153
rect 2477 5007 2483 5033
rect 2517 5007 2523 5153
rect 2640 5063 2653 5067
rect 2637 5053 2653 5063
rect 2637 5027 2643 5053
rect 3097 5027 3103 5053
rect 3117 4987 3123 5133
rect 3137 5027 3143 5173
rect 3277 5007 3283 5153
rect 3297 5027 3303 5173
rect 3317 5047 3323 5153
rect 3597 5007 3603 5173
rect 3737 5027 3743 5093
rect 4357 4987 4363 5133
rect 4497 5007 4503 5113
rect 4937 5007 4943 5174
rect 5397 4987 5403 5133
rect 5517 5047 5523 5173
rect 5677 5087 5683 5153
rect 5977 5067 5983 5133
rect 6057 5107 6063 5153
rect 5967 5057 5983 5067
rect 5967 5053 5980 5057
rect 797 4977 813 4987
rect 800 4973 813 4977
rect 6077 4958 6137 5462
rect 6050 4942 6137 4958
rect 457 4727 463 4873
rect 597 4747 603 4853
rect 1217 4747 1223 4813
rect 1657 4787 1663 4913
rect 2097 4867 2103 4893
rect 1647 4777 1663 4787
rect 1647 4773 1660 4777
rect 1957 4727 1963 4853
rect 2517 4847 2523 4913
rect 2217 4727 2223 4833
rect 2537 4767 2543 4893
rect 2677 4767 2683 4853
rect 2837 4747 2843 4853
rect 3277 4727 3283 4753
rect 3537 4727 3543 4853
rect 3557 4747 3563 4893
rect 3897 4727 3903 4853
rect 4037 4747 4043 4893
rect 4197 4767 4203 4913
rect 4237 4867 4243 4893
rect 4337 4747 4343 4893
rect 4637 4767 4643 4913
rect 4777 4827 4783 4913
rect 4337 4737 4353 4747
rect 4340 4733 4353 4737
rect 5077 4727 5083 4793
rect 5097 4727 5103 4853
rect 5217 4767 5223 4913
rect 5237 4767 5243 4833
rect 5357 4727 5363 4913
rect 5897 4747 5903 4873
rect 5917 4847 5923 4913
rect 6037 4827 6043 4913
rect 6037 4727 6043 4773
rect 6057 4747 6063 4893
rect -57 4682 30 4698
rect -57 4178 3 4682
rect 2697 4660 2743 4663
rect 2693 4657 2743 4660
rect 600 4643 612 4647
rect 597 4633 612 4643
rect 597 4487 603 4633
rect 1077 4527 1083 4573
rect 1237 4467 1243 4633
rect 1557 4587 1563 4613
rect 1557 4487 1563 4573
rect 1677 4467 1683 4613
rect 2117 4523 2123 4633
rect 2257 4607 2263 4633
rect 2257 4597 2273 4607
rect 2260 4593 2273 4597
rect 2297 4527 2303 4653
rect 2097 4517 2123 4523
rect 1997 4467 2003 4513
rect 2097 4467 2103 4517
rect 2297 4467 2303 4513
rect 2417 4467 2423 4613
rect 2557 4487 2563 4653
rect 2693 4647 2707 4657
rect 2706 4640 2707 4647
rect 2717 4467 2723 4633
rect 2737 4627 2743 4657
rect 4827 4663 4840 4667
rect 4827 4653 4843 4663
rect 2867 4603 2880 4607
rect 2867 4600 2883 4603
rect 2867 4593 2887 4600
rect 2873 4587 2887 4593
rect 2757 4467 2763 4513
rect 2857 4507 2863 4553
rect 2857 4497 2873 4507
rect 2860 4493 2873 4497
rect 2997 4467 3003 4613
rect 3497 4487 3503 4533
rect 3517 4507 3523 4653
rect 3677 4487 3683 4653
rect 3837 4527 3843 4653
rect 3997 4467 4003 4613
rect 4097 4501 4103 4593
rect 4257 4467 4263 4653
rect 4377 4583 4383 4653
rect 4377 4577 4403 4583
rect 4397 4507 4403 4577
rect 4387 4497 4403 4507
rect 4387 4493 4400 4497
rect 4417 4487 4423 4653
rect 4837 4467 4843 4653
rect 4877 4567 4883 4633
rect 4867 4557 4883 4567
rect 4867 4553 4880 4557
rect 5017 4547 5023 4653
rect 4897 4467 4903 4513
rect 5157 4467 5163 4653
rect 5317 4467 5323 4653
rect 5617 4527 5623 4653
rect 5777 4487 5783 4633
rect 5917 4487 5923 4633
rect 5937 4547 5943 4573
rect 6037 4467 6043 4653
rect 2297 4457 2313 4467
rect 2300 4453 2313 4457
rect 5148 4457 5163 4467
rect 5148 4453 5160 4457
rect 6037 4457 6053 4467
rect 6040 4453 6053 4457
rect 6077 4438 6137 4942
rect 6050 4422 6137 4438
rect 2187 4403 2200 4407
rect 2187 4400 2203 4403
rect 2187 4393 2207 4400
rect 197 4207 203 4293
rect 337 4247 343 4373
rect 1577 4307 1583 4393
rect 1197 4247 1203 4273
rect 1737 4207 1743 4393
rect 1931 4373 1937 4393
rect 2193 4387 2207 4393
rect 2193 4380 2194 4387
rect 1877 4307 1883 4373
rect 1917 4367 1937 4373
rect 1917 4347 1923 4367
rect 2957 4347 2963 4393
rect 2180 4303 2193 4307
rect 2177 4293 2193 4303
rect 2177 4207 2183 4293
rect 2737 4207 2743 4333
rect 3217 4247 3223 4373
rect 3877 4247 3883 4393
rect 3917 4247 3923 4333
rect 2777 4207 2783 4233
rect 4797 4207 4803 4353
rect 4937 4267 4943 4393
rect 4967 4303 4980 4307
rect 4967 4293 4983 4303
rect 4977 4247 4983 4293
rect 5137 4207 5143 4353
rect 5277 4267 5283 4333
rect 5717 4207 5723 4393
rect 5737 4247 5743 4333
rect 2768 4197 2783 4207
rect 2768 4193 2780 4197
rect -57 4162 30 4178
rect -57 3658 3 4162
rect 497 4023 503 4113
rect 497 4020 523 4023
rect 497 4017 527 4020
rect 477 3967 483 4013
rect 513 4007 527 4017
rect 857 4007 863 4073
rect 513 4000 514 4007
rect 1557 3947 1563 4133
rect 2177 3947 2183 4093
rect 2317 4087 2323 4133
rect 2497 3967 2503 4133
rect 3057 3967 3063 4133
rect 3797 3947 3803 4093
rect 4237 3947 4243 4093
rect 5277 4087 5283 4133
rect 5277 3947 5283 3993
rect 5297 3967 5303 4133
rect 5457 3967 5463 4093
rect 5597 3947 5603 4113
rect 5777 4007 5783 4093
rect 5917 3947 5923 4133
rect 6077 3918 6137 4422
rect 6050 3902 6137 3918
rect 17 3847 23 3873
rect 317 3727 323 3813
rect 617 3687 623 3873
rect 800 3823 814 3827
rect 797 3813 814 3823
rect 777 3707 783 3753
rect 797 3687 803 3813
rect 1097 3687 1103 3753
rect 1337 3707 1343 3813
rect 2377 3687 2383 3813
rect 2537 3727 2543 3853
rect 2677 3707 2683 3813
rect 3117 3687 3123 3753
rect 3417 3687 3423 3813
rect 3757 3727 3763 3853
rect 4177 3847 4183 3873
rect 3857 3687 3863 3753
rect 3877 3747 3883 3813
rect 4817 3727 4823 3873
rect 4837 3847 4843 3873
rect 5217 3687 5223 3853
rect -57 3642 30 3658
rect -57 3138 3 3642
rect 297 3427 303 3593
rect 577 3487 583 3573
rect 1277 3547 1283 3613
rect 577 3447 583 3473
rect 2417 3427 2423 3473
rect 3057 3427 3063 3613
rect 3357 3447 3363 3613
rect 4277 3467 4283 3613
rect 4437 3467 4443 3613
rect 5357 3427 5363 3613
rect 5957 3447 5963 3553
rect 6077 3398 6137 3902
rect 6050 3382 6137 3398
rect 357 3167 363 3353
rect 637 3207 643 3353
rect 877 3307 883 3353
rect 2637 3307 2643 3353
rect 3057 3187 3063 3233
rect 3077 3207 3083 3353
rect 3237 3207 3243 3353
rect 3257 3187 3263 3293
rect 3817 3247 3823 3353
rect 4117 3207 4123 3293
rect 4697 3207 4703 3293
rect 5477 3167 5483 3353
rect 5617 3187 5623 3353
rect 5897 3307 5903 3353
rect 5757 3207 5763 3293
rect 347 3157 363 3167
rect 347 3153 360 3157
rect -57 3122 30 3138
rect -57 2618 3 3122
rect 217 2967 223 3033
rect 2577 2927 2583 3073
rect 2877 2927 2883 3073
rect 3177 2967 3183 3053
rect 5337 2927 5343 3013
rect 5357 2907 5363 3093
rect 5957 2907 5963 2953
rect 6077 2878 6137 3382
rect 6050 2862 6137 2878
rect 297 2687 303 2813
rect 1657 2647 1663 2673
rect 1777 2667 1783 2793
rect 2077 2647 2083 2793
rect 3377 2667 3383 2773
rect 4737 2707 4743 2773
rect 4877 2647 4883 2773
rect 5437 2647 5443 2773
rect -57 2602 30 2618
rect -57 2098 3 2602
rect 1217 2447 1223 2493
rect 1237 2467 1243 2573
rect 1357 2387 1363 2533
rect 1537 2387 1543 2573
rect 1957 2387 1963 2493
rect 2117 2447 2123 2533
rect 3477 2487 3483 2573
rect 4277 2407 4283 2513
rect 4617 2407 4623 2513
rect 5517 2387 5523 2573
rect 1537 2377 1553 2387
rect 1540 2373 1553 2377
rect 6077 2358 6137 2862
rect 6050 2342 6137 2358
rect 557 2167 563 2273
rect 4097 2267 4103 2313
rect 3377 2187 3383 2253
rect 5197 2247 5203 2293
rect 5937 2127 5943 2253
rect -57 2082 30 2098
rect -57 1578 3 2082
rect 1417 1867 1423 2033
rect 6077 1838 6137 2342
rect 6050 1822 6137 1838
rect 197 1647 203 1793
rect 1317 1647 1323 1673
rect 1617 1647 1623 1733
rect 2997 1607 3003 1693
rect 3037 1627 3043 1753
rect 3417 1667 3423 1713
rect 3437 1627 3443 1793
rect 4537 1607 4543 1693
rect 4777 1647 4783 1793
rect 5357 1647 5363 1773
rect 5657 1647 5663 1753
rect 4767 1617 4793 1623
rect -57 1562 30 1578
rect -57 1058 3 1562
rect 477 1447 483 1493
rect 2637 1347 2643 1473
rect 2817 1387 2823 1513
rect 2957 1367 2963 1533
rect 4597 1347 4603 1433
rect 5897 1347 5903 1533
rect 6077 1318 6137 1822
rect 6050 1302 6137 1318
rect 597 1087 603 1213
rect 2137 1088 2143 1273
rect 2437 1107 2443 1173
rect 2457 1087 2463 1273
rect 2857 1227 2863 1273
rect 3377 1107 3383 1213
rect 4157 1107 4163 1173
rect 5217 1127 5223 1253
rect -57 1042 30 1058
rect -57 538 3 1042
rect 317 887 323 1013
rect 337 847 343 973
rect 497 887 503 973
rect 637 827 643 993
rect 837 927 843 1013
rect 2917 847 2923 953
rect 2937 927 2943 973
rect 3117 887 3123 993
rect 3257 827 3263 973
rect 5237 887 5243 953
rect 6077 798 6137 1302
rect 6050 782 6137 798
rect 3100 763 3113 767
rect 3097 753 3113 763
rect 657 567 663 753
rect 797 607 803 693
rect 1297 567 1303 653
rect 1597 647 1603 753
rect 2537 587 2543 753
rect 2937 647 2943 733
rect 2557 567 2563 593
rect 3097 587 3103 753
rect 3277 567 3283 713
rect 3637 567 3643 733
rect 4037 587 4043 753
rect 4317 607 4323 753
rect 4337 587 4343 733
rect 4357 567 4363 633
rect 4817 607 4823 733
rect 5917 567 5923 633
rect -57 522 30 538
rect -57 18 3 522
rect 617 327 623 493
rect 777 307 783 413
rect 1037 367 1043 473
rect 1717 327 1723 413
rect 2577 327 2583 433
rect 2737 327 2743 413
rect 3497 407 3503 453
rect 5637 327 5643 433
rect 6077 278 6137 782
rect 6050 262 6137 278
rect 157 47 163 233
rect 1797 47 1803 173
rect 2117 87 2123 193
rect 2957 127 2963 233
rect 5117 47 5123 233
rect -57 2 30 18
rect 6077 2 6137 262
<< m2contact >>
rect 513 5953 527 5967
rect 5113 5953 5127 5967
rect 5274 5953 5288 5967
rect 5433 5953 5447 5967
rect 312 5893 326 5907
rect 3433 5933 3447 5947
rect 3593 5933 3607 5947
rect 4733 5933 4747 5947
rect 4913 5933 4927 5947
rect 2673 5913 2687 5927
rect 553 5893 567 5907
rect 693 5893 707 5907
rect 2553 5893 2567 5907
rect 513 5793 527 5807
rect 673 5873 687 5887
rect 673 5793 687 5807
rect 853 5873 867 5887
rect 2553 5833 2567 5847
rect 853 5793 867 5807
rect 2713 5893 2727 5907
rect 3433 5833 3447 5847
rect 3593 5833 3607 5847
rect 3873 5833 3887 5847
rect 5113 5913 5127 5927
rect 5253 5893 5267 5907
rect 4732 5773 4746 5787
rect 4913 5773 4927 5787
rect 5412 5813 5426 5827
rect 5273 5773 5287 5787
rect 5413 5773 5427 5787
rect 333 5753 347 5767
rect 532 5753 546 5767
rect 693 5753 707 5767
rect 2673 5753 2687 5767
rect 2713 5753 2727 5767
rect 3572 5753 3586 5767
rect 3873 5753 3887 5767
rect 5252 5753 5266 5767
rect 5433 5753 5447 5767
rect 1673 5693 1687 5707
rect 2653 5693 2667 5707
rect 2953 5693 2967 5707
rect 3253 5693 3267 5707
rect 3692 5693 3706 5707
rect 4333 5693 4347 5707
rect 4733 5693 4747 5707
rect 5053 5693 5067 5707
rect 5673 5693 5687 5707
rect 1373 5673 1387 5687
rect 653 5613 667 5627
rect 833 5613 847 5627
rect 2653 5653 2667 5667
rect 1673 5633 1687 5647
rect 3133 5653 3147 5667
rect 2653 5613 2667 5627
rect 2953 5613 2967 5627
rect 1373 5593 1387 5607
rect 2833 5553 2847 5567
rect 833 5513 847 5527
rect 3133 5513 3147 5527
rect 3713 5673 3727 5687
rect 3573 5613 3587 5627
rect 4913 5633 4927 5647
rect 4333 5533 4347 5547
rect 4733 5533 4747 5547
rect 4893 5533 4907 5547
rect 3552 5513 3566 5527
rect 5233 5673 5247 5687
rect 5053 5553 5067 5567
rect 4913 5514 4927 5528
rect 5373 5653 5387 5667
rect 5813 5613 5827 5627
rect 5813 5573 5827 5587
rect 6053 5533 6067 5547
rect 653 5493 667 5507
rect 2833 5493 2847 5507
rect 3253 5493 3267 5507
rect 4892 5493 4906 5507
rect 5233 5493 5247 5507
rect 5373 5493 5387 5507
rect 5653 5493 5667 5507
rect 6053 5493 6067 5507
rect 193 5433 207 5447
rect 833 5433 847 5447
rect 1093 5433 1107 5447
rect 1713 5433 1727 5447
rect 2793 5433 2807 5447
rect 3114 5433 3128 5447
rect 4073 5433 4087 5447
rect 4693 5433 4707 5447
rect 4953 5433 4967 5447
rect 5734 5433 5748 5447
rect 6013 5433 6027 5447
rect 673 5413 687 5427
rect 193 5253 207 5267
rect 1413 5393 1427 5407
rect 1113 5373 1127 5387
rect 833 5313 847 5327
rect 1093 5313 1107 5327
rect 1093 5273 1107 5287
rect 1853 5373 1867 5387
rect 2753 5373 2767 5387
rect 1713 5273 1727 5287
rect 1414 5253 1428 5267
rect 2313 5273 2327 5287
rect 2773 5293 2787 5307
rect 2752 5253 2766 5267
rect 2933 5413 2947 5427
rect 2913 5313 2927 5327
rect 2793 5253 2807 5267
rect 2912 5253 2926 5267
rect 3613 5413 3627 5427
rect 3433 5393 3447 5407
rect 3113 5313 3127 5327
rect 3453 5293 3467 5307
rect 3433 5273 3447 5287
rect 3453 5253 3467 5267
rect 4094 5413 4108 5427
rect 4393 5413 4407 5427
rect 4073 5373 4087 5387
rect 4233 5393 4247 5407
rect 4253 5333 4267 5347
rect 4673 5393 4687 5407
rect 4393 5313 4407 5327
rect 4253 5293 4267 5307
rect 4093 5253 4107 5267
rect 4233 5253 4247 5267
rect 4673 5253 4687 5267
rect 4833 5413 4847 5427
rect 5292 5313 5306 5327
rect 4953 5273 4967 5287
rect 5993 5373 6007 5387
rect 6013 5273 6027 5287
rect 673 5233 687 5247
rect 1113 5233 1127 5247
rect 1832 5233 1846 5247
rect 2313 5233 2327 5247
rect 2773 5233 2787 5247
rect 2933 5233 2947 5247
rect 3613 5233 3627 5247
rect 4693 5233 4707 5247
rect 4833 5233 4847 5247
rect 5273 5233 5287 5247
rect 5733 5233 5747 5247
rect 5993 5233 6007 5247
rect 3133 5173 3147 5187
rect 3293 5173 3307 5187
rect 3593 5173 3607 5187
rect 4933 5174 4947 5188
rect 1113 5153 1127 5167
rect 1413 5153 1427 5167
rect 1573 5153 1587 5167
rect 2513 5153 2527 5167
rect 653 5133 667 5147
rect 793 5053 807 5067
rect 973 5053 987 5067
rect 1254 5133 1268 5147
rect 1253 5093 1267 5107
rect 1133 5053 1147 5067
rect 1113 5013 1127 5027
rect 1573 5033 1587 5047
rect 2473 5033 2487 5047
rect 3113 5133 3127 5147
rect 2653 5053 2667 5067
rect 3093 5053 3107 5067
rect 2633 5013 2647 5027
rect 3092 5013 3106 5027
rect 2473 4993 2487 5007
rect 2513 4993 2527 5007
rect 3273 5153 3287 5167
rect 3133 5013 3147 5027
rect 3313 5153 3327 5167
rect 3313 5033 3327 5047
rect 3293 5013 3307 5027
rect 4353 5133 4367 5147
rect 3733 5093 3747 5107
rect 3733 5013 3747 5027
rect 3273 4993 3287 5007
rect 3593 4993 3607 5007
rect 4493 5113 4507 5127
rect 5513 5173 5527 5187
rect 5393 5133 5407 5147
rect 4493 4993 4507 5007
rect 4933 4993 4947 5007
rect 5673 5153 5687 5167
rect 6053 5153 6067 5167
rect 5973 5133 5987 5147
rect 5673 5073 5687 5087
rect 6053 5093 6067 5107
rect 5953 5053 5967 5067
rect 5514 5033 5528 5047
rect 653 4973 667 4987
rect 813 4973 827 4987
rect 973 4973 987 4987
rect 1133 4973 1147 4987
rect 1393 4973 1407 4987
rect 3113 4973 3127 4987
rect 4353 4973 4367 4987
rect 5393 4973 5407 4987
rect 1653 4913 1667 4927
rect 2513 4913 2527 4927
rect 4193 4913 4207 4927
rect 4633 4913 4647 4927
rect 4772 4913 4786 4927
rect 5213 4913 5227 4927
rect 5353 4913 5367 4927
rect 5913 4913 5927 4927
rect 6033 4913 6047 4927
rect 453 4873 467 4887
rect 593 4853 607 4867
rect 1213 4813 1227 4827
rect 2092 4893 2106 4907
rect 1953 4853 1967 4867
rect 2093 4853 2107 4867
rect 1633 4773 1647 4787
rect 593 4733 607 4747
rect 1212 4733 1226 4747
rect 2533 4893 2547 4907
rect 3553 4893 3567 4907
rect 4034 4893 4048 4907
rect 2213 4833 2227 4847
rect 2513 4833 2527 4847
rect 2673 4853 2687 4867
rect 2833 4853 2847 4867
rect 3533 4853 3547 4867
rect 2533 4753 2547 4767
rect 2673 4753 2687 4767
rect 3273 4753 3287 4767
rect 2833 4733 2847 4747
rect 3893 4853 3907 4867
rect 3553 4733 3567 4747
rect 4233 4893 4247 4907
rect 4333 4893 4347 4907
rect 4233 4853 4247 4867
rect 4193 4753 4207 4767
rect 5093 4853 5107 4867
rect 4773 4813 4787 4827
rect 5073 4793 5087 4807
rect 4633 4753 4647 4767
rect 4033 4733 4047 4747
rect 4353 4733 4367 4747
rect 5233 4833 5247 4847
rect 5212 4753 5226 4767
rect 5234 4753 5248 4767
rect 5893 4873 5907 4887
rect 5913 4833 5927 4847
rect 6053 4893 6067 4907
rect 6032 4813 6046 4827
rect 6033 4773 6047 4787
rect 5893 4733 5907 4747
rect 6054 4733 6068 4747
rect 453 4713 467 4727
rect 1953 4713 1967 4727
rect 2213 4713 2227 4727
rect 3273 4713 3287 4727
rect 3533 4713 3547 4727
rect 3893 4713 3907 4727
rect 5072 4713 5086 4727
rect 5094 4713 5108 4727
rect 5353 4713 5367 4727
rect 6032 4713 6046 4727
rect 2292 4653 2306 4667
rect 2553 4653 2567 4667
rect 612 4633 626 4647
rect 1233 4633 1247 4647
rect 2113 4633 2127 4647
rect 2252 4633 2266 4647
rect 1073 4573 1087 4587
rect 1073 4513 1087 4527
rect 593 4473 607 4487
rect 1553 4613 1567 4627
rect 1673 4613 1687 4627
rect 1553 4573 1567 4587
rect 1553 4473 1567 4487
rect 1993 4513 2007 4527
rect 2273 4593 2287 4607
rect 2413 4613 2427 4627
rect 2293 4513 2307 4527
rect 2692 4633 2706 4647
rect 2714 4633 2728 4647
rect 2553 4473 2567 4487
rect 3513 4653 3527 4667
rect 3673 4653 3687 4667
rect 3833 4653 3847 4667
rect 4253 4653 4267 4667
rect 4372 4653 4386 4667
rect 4413 4653 4427 4667
rect 4813 4653 4827 4667
rect 5013 4653 5027 4667
rect 5153 4653 5167 4667
rect 5313 4653 5327 4667
rect 5613 4653 5627 4667
rect 6033 4653 6047 4667
rect 2734 4613 2748 4627
rect 2993 4613 3007 4627
rect 2853 4593 2867 4607
rect 2873 4573 2887 4587
rect 2853 4553 2867 4567
rect 2753 4513 2767 4527
rect 2873 4493 2887 4507
rect 3493 4533 3507 4547
rect 3514 4493 3528 4507
rect 3993 4613 4007 4627
rect 3833 4513 3847 4527
rect 3492 4473 3506 4487
rect 3673 4473 3687 4487
rect 4093 4593 4107 4607
rect 4093 4487 4107 4501
rect 4373 4493 4387 4507
rect 4413 4473 4427 4487
rect 4873 4633 4887 4647
rect 4853 4553 4867 4567
rect 5013 4533 5027 4547
rect 4893 4513 4907 4527
rect 5773 4633 5787 4647
rect 5913 4633 5927 4647
rect 5613 4513 5627 4527
rect 5934 4573 5948 4587
rect 5933 4533 5947 4547
rect 5773 4473 5787 4487
rect 5913 4473 5927 4487
rect 1233 4453 1247 4467
rect 1673 4453 1687 4467
rect 1993 4453 2007 4467
rect 2092 4453 2106 4467
rect 2313 4453 2327 4467
rect 2413 4453 2427 4467
rect 2713 4453 2727 4467
rect 2753 4453 2767 4467
rect 2993 4453 3007 4467
rect 3994 4453 4008 4467
rect 4253 4453 4267 4467
rect 4833 4453 4847 4467
rect 4893 4453 4907 4467
rect 5134 4453 5148 4467
rect 5313 4453 5327 4467
rect 6053 4453 6067 4467
rect 1573 4393 1587 4407
rect 1734 4393 1748 4407
rect 1927 4393 1941 4407
rect 2173 4393 2187 4407
rect 2953 4393 2967 4407
rect 3874 4393 3888 4407
rect 4933 4393 4947 4407
rect 5713 4393 5727 4407
rect 333 4373 347 4387
rect 193 4293 207 4307
rect 1573 4293 1587 4307
rect 1193 4273 1207 4287
rect 333 4233 347 4247
rect 1193 4233 1207 4247
rect 1873 4373 1887 4387
rect 2194 4373 2208 4387
rect 3214 4373 3228 4387
rect 1913 4333 1927 4347
rect 2733 4333 2747 4347
rect 2953 4333 2967 4347
rect 1873 4293 1887 4307
rect 2193 4293 2207 4307
rect 4793 4353 4807 4367
rect 3913 4333 3927 4347
rect 2773 4233 2787 4247
rect 3213 4233 3227 4247
rect 3873 4233 3887 4247
rect 3913 4233 3927 4247
rect 5133 4353 5147 4367
rect 4953 4293 4967 4307
rect 4933 4253 4947 4267
rect 4973 4233 4987 4247
rect 5273 4333 5287 4347
rect 5273 4253 5287 4267
rect 5733 4333 5747 4347
rect 5733 4233 5747 4247
rect 192 4193 206 4207
rect 1733 4193 1747 4207
rect 2173 4193 2187 4207
rect 2732 4193 2746 4207
rect 2754 4193 2768 4207
rect 4793 4193 4807 4207
rect 5133 4193 5147 4207
rect 5713 4193 5727 4207
rect 1552 4133 1566 4147
rect 2313 4133 2327 4147
rect 2493 4133 2507 4147
rect 3053 4133 3067 4147
rect 5272 4133 5286 4147
rect 5294 4133 5308 4147
rect 5913 4133 5927 4147
rect 493 4113 507 4127
rect 473 4013 487 4027
rect 853 4073 867 4087
rect 514 3993 528 4007
rect 853 3993 867 4007
rect 473 3953 487 3967
rect 2172 4093 2186 4107
rect 2313 4073 2327 4087
rect 3793 4093 3807 4107
rect 4233 4093 4247 4107
rect 2493 3953 2507 3967
rect 3053 3953 3067 3967
rect 5273 4073 5287 4087
rect 5273 3993 5287 4007
rect 5593 4113 5607 4127
rect 5453 4093 5467 4107
rect 5293 3953 5307 3967
rect 5453 3953 5467 3967
rect 5773 4093 5787 4107
rect 5772 3993 5786 4007
rect 1553 3933 1567 3947
rect 2173 3933 2187 3947
rect 3793 3933 3807 3947
rect 4233 3933 4247 3947
rect 5273 3933 5287 3947
rect 5593 3933 5607 3947
rect 5913 3933 5927 3947
rect 12 3873 26 3887
rect 613 3873 627 3887
rect 4173 3873 4187 3887
rect 4812 3873 4826 3887
rect 4834 3873 4848 3887
rect 13 3833 27 3847
rect 313 3813 327 3827
rect 313 3713 327 3727
rect 2533 3853 2547 3867
rect 3753 3853 3767 3867
rect 814 3813 828 3827
rect 1333 3813 1347 3827
rect 2373 3813 2387 3827
rect 774 3753 788 3767
rect 772 3693 786 3707
rect 1093 3753 1107 3767
rect 1333 3693 1347 3707
rect 2673 3813 2687 3827
rect 3412 3813 3426 3827
rect 2533 3713 2547 3727
rect 3113 3753 3127 3767
rect 2673 3693 2687 3707
rect 4173 3833 4187 3847
rect 3873 3813 3887 3827
rect 3853 3753 3867 3767
rect 3753 3713 3767 3727
rect 3873 3733 3887 3747
rect 5214 3853 5228 3867
rect 4833 3833 4847 3847
rect 4813 3713 4827 3727
rect 613 3673 627 3687
rect 793 3673 807 3687
rect 1093 3673 1107 3687
rect 2373 3673 2387 3687
rect 3114 3673 3128 3687
rect 3413 3673 3427 3687
rect 3854 3673 3868 3687
rect 5213 3673 5227 3687
rect 1273 3613 1287 3627
rect 3053 3613 3067 3627
rect 3353 3613 3367 3627
rect 4273 3613 4287 3627
rect 4433 3613 4447 3627
rect 5353 3613 5367 3627
rect 293 3593 307 3607
rect 573 3573 587 3587
rect 1273 3533 1287 3547
rect 573 3473 587 3487
rect 2413 3473 2427 3487
rect 573 3433 587 3447
rect 4273 3453 4287 3467
rect 4433 3453 4447 3467
rect 3353 3433 3367 3447
rect 5953 3553 5967 3567
rect 5953 3433 5967 3447
rect 293 3413 307 3427
rect 2414 3413 2428 3427
rect 3054 3413 3068 3427
rect 5353 3413 5367 3427
rect 353 3353 367 3367
rect 633 3353 647 3367
rect 873 3353 887 3367
rect 2633 3353 2647 3367
rect 3073 3353 3087 3367
rect 3233 3353 3247 3367
rect 3813 3353 3827 3367
rect 5473 3353 5487 3367
rect 5613 3353 5627 3367
rect 5893 3353 5907 3367
rect 873 3293 887 3307
rect 2633 3293 2647 3307
rect 3053 3233 3067 3247
rect 633 3193 647 3207
rect 3254 3293 3268 3307
rect 3073 3193 3087 3207
rect 3233 3193 3247 3207
rect 4113 3293 4127 3307
rect 4694 3293 4708 3307
rect 3813 3233 3827 3247
rect 4113 3193 4127 3207
rect 4693 3193 4707 3207
rect 3053 3173 3067 3187
rect 3253 3173 3267 3187
rect 5752 3293 5766 3307
rect 5893 3293 5907 3307
rect 5753 3193 5767 3207
rect 5613 3173 5627 3187
rect 333 3153 347 3167
rect 5473 3153 5487 3167
rect 5353 3093 5367 3107
rect 2573 3073 2587 3087
rect 2873 3073 2887 3087
rect 213 3033 227 3047
rect 213 2953 227 2967
rect 3173 3053 3187 3067
rect 5333 3013 5347 3027
rect 3172 2953 3186 2967
rect 2573 2913 2587 2927
rect 2874 2913 2888 2927
rect 5332 2913 5346 2927
rect 5953 2953 5967 2967
rect 5354 2893 5368 2907
rect 5953 2893 5967 2907
rect 293 2813 307 2827
rect 1773 2793 1787 2807
rect 2073 2793 2087 2807
rect 293 2673 307 2687
rect 1653 2673 1667 2687
rect 1773 2653 1787 2667
rect 3373 2773 3387 2787
rect 4733 2773 4747 2787
rect 4873 2773 4887 2787
rect 5433 2773 5447 2787
rect 4733 2693 4747 2707
rect 3373 2653 3387 2667
rect 1653 2633 1667 2647
rect 2073 2633 2087 2647
rect 4873 2633 4887 2647
rect 5433 2633 5447 2647
rect 1233 2573 1247 2587
rect 1533 2573 1547 2587
rect 3473 2573 3487 2587
rect 5513 2573 5527 2587
rect 1213 2493 1227 2507
rect 1353 2533 1367 2547
rect 1233 2453 1247 2467
rect 1212 2433 1226 2447
rect 2113 2533 2127 2547
rect 1953 2493 1967 2507
rect 4273 2513 4287 2527
rect 4613 2513 4627 2527
rect 3473 2473 3487 2487
rect 2113 2433 2127 2447
rect 4273 2393 4287 2407
rect 4613 2393 4627 2407
rect 1353 2373 1367 2387
rect 1553 2373 1567 2387
rect 1953 2373 1967 2387
rect 5513 2373 5527 2387
rect 4093 2313 4107 2327
rect 553 2273 567 2287
rect 5193 2293 5207 2307
rect 3373 2253 3387 2267
rect 4093 2253 4107 2267
rect 5933 2253 5947 2267
rect 5193 2233 5207 2247
rect 3373 2173 3387 2187
rect 553 2153 567 2167
rect 5933 2113 5947 2127
rect 1413 2033 1427 2047
rect 1413 1853 1427 1867
rect 193 1793 207 1807
rect 3433 1793 3447 1807
rect 4773 1793 4787 1807
rect 3033 1753 3047 1767
rect 1613 1733 1627 1747
rect 1313 1673 1327 1687
rect 2993 1693 3007 1707
rect 193 1633 207 1647
rect 1314 1633 1328 1647
rect 1613 1633 1627 1647
rect 3413 1713 3427 1727
rect 3413 1653 3427 1667
rect 4533 1693 4547 1707
rect 3034 1613 3048 1627
rect 3433 1613 3447 1627
rect 5353 1773 5367 1787
rect 5653 1753 5667 1767
rect 4773 1633 4787 1647
rect 5353 1633 5367 1647
rect 5653 1633 5667 1647
rect 4753 1613 4767 1627
rect 4793 1613 4807 1627
rect 2993 1593 3007 1607
rect 4533 1593 4547 1607
rect 2953 1533 2967 1547
rect 5893 1533 5907 1547
rect 2813 1513 2827 1527
rect 473 1493 487 1507
rect 2633 1473 2647 1487
rect 473 1433 487 1447
rect 2813 1373 2827 1387
rect 4593 1433 4607 1447
rect 2953 1353 2967 1367
rect 2633 1333 2647 1347
rect 4593 1333 4607 1347
rect 5893 1333 5907 1347
rect 2133 1273 2147 1287
rect 2453 1273 2467 1287
rect 2853 1273 2867 1287
rect 593 1213 607 1227
rect 2433 1173 2447 1187
rect 2433 1093 2447 1107
rect 593 1073 607 1087
rect 2133 1074 2147 1088
rect 5213 1253 5227 1267
rect 2853 1213 2867 1227
rect 3373 1213 3387 1227
rect 4154 1173 4168 1187
rect 5213 1113 5227 1127
rect 3373 1093 3387 1107
rect 4153 1093 4167 1107
rect 2453 1073 2467 1087
rect 313 1013 327 1027
rect 833 1013 847 1027
rect 633 993 647 1007
rect 334 973 348 987
rect 493 973 507 987
rect 313 873 327 887
rect 493 873 507 887
rect 333 833 347 847
rect 3113 993 3127 1007
rect 2933 973 2947 987
rect 2913 953 2927 967
rect 833 913 847 927
rect 2933 913 2947 927
rect 3253 973 3267 987
rect 3112 873 3126 887
rect 2913 833 2927 847
rect 5233 953 5247 967
rect 5233 873 5247 887
rect 633 813 647 827
rect 3253 813 3267 827
rect 654 753 668 767
rect 1593 753 1607 767
rect 2533 753 2547 767
rect 3113 753 3127 767
rect 4032 753 4046 767
rect 4313 753 4327 767
rect 793 693 807 707
rect 1293 653 1307 667
rect 793 593 807 607
rect 1593 633 1607 647
rect 2933 733 2947 747
rect 2933 633 2947 647
rect 2552 593 2566 607
rect 2532 573 2546 587
rect 3633 733 3647 747
rect 3273 713 3287 727
rect 3094 573 3108 587
rect 4333 733 4347 747
rect 4813 733 4827 747
rect 4313 593 4327 607
rect 4353 633 4367 647
rect 4033 573 4047 587
rect 4332 573 4346 587
rect 5913 633 5927 647
rect 4813 593 4827 607
rect 653 553 667 567
rect 1293 553 1307 567
rect 2554 553 2568 567
rect 3272 553 3286 567
rect 3633 553 3647 567
rect 4353 553 4367 567
rect 5913 553 5927 567
rect 613 493 627 507
rect 1033 473 1047 487
rect 773 413 787 427
rect 613 313 627 327
rect 3493 453 3507 467
rect 2573 433 2587 447
rect 1713 413 1727 427
rect 1033 353 1047 367
rect 2733 413 2747 427
rect 5633 433 5647 447
rect 3493 393 3507 407
rect 1713 313 1727 327
rect 2573 313 2587 327
rect 2733 313 2747 327
rect 5633 313 5647 327
rect 773 293 787 307
rect 153 233 167 247
rect 2953 233 2967 247
rect 5112 233 5126 247
rect 2113 193 2127 207
rect 1793 173 1807 187
rect 2953 113 2967 127
rect 2113 73 2127 87
rect 153 33 167 47
rect 1793 33 1807 47
rect 5113 33 5127 47
<< metal2 >>
rect 1107 5996 1313 6003
rect 1467 5996 3523 6003
rect 147 5976 213 5983
rect 227 5976 833 5983
rect 907 5976 1133 5983
rect 1147 5976 1293 5983
rect 2307 5976 2653 5983
rect 2767 5976 2893 5983
rect 2947 5976 3073 5983
rect 3087 5976 3213 5983
rect 3327 5976 3493 5983
rect 3516 5983 3523 5996
rect 3687 5996 4133 6003
rect 4147 5996 4603 6003
rect 3516 5976 3713 5983
rect 3767 5976 3833 5983
rect 3847 5976 4293 5983
rect 4307 5976 4393 5983
rect 4596 5983 4603 5996
rect 4627 5996 5173 6003
rect 5267 5996 5513 6003
rect 4596 5976 4913 5983
rect 4967 5976 5213 5983
rect 5307 5976 5353 5983
rect 447 5956 513 5963
rect 527 5956 1673 5963
rect 1947 5956 2013 5963
rect 2027 5956 4093 5963
rect 4107 5956 4323 5963
rect 467 5936 613 5943
rect 627 5936 1233 5943
rect 1627 5936 1873 5943
rect 2207 5936 2253 5943
rect 2567 5936 2613 5943
rect 2847 5936 3173 5943
rect 3187 5936 3433 5943
rect 3607 5936 3673 5943
rect 4316 5943 4323 5956
rect 4847 5956 5113 5963
rect 5127 5956 5252 5963
rect 5288 5956 5333 5963
rect 5347 5956 5373 5963
rect 5447 5956 5473 5963
rect 4316 5936 4653 5943
rect 2753 5927 2767 5933
rect 2247 5916 2293 5923
rect 2687 5916 2753 5923
rect 3567 5916 3613 5923
rect 3493 5907 3507 5913
rect 4456 5907 4463 5936
rect 4747 5936 4793 5943
rect 4927 5936 4953 5943
rect 5407 5936 5553 5943
rect 5567 5936 5773 5943
rect 5127 5913 5133 5927
rect 5267 5916 5333 5923
rect 187 5896 253 5903
rect 306 5893 312 5907
rect 348 5896 413 5903
rect 567 5893 573 5907
rect 707 5896 753 5903
rect 847 5896 913 5903
rect 1347 5893 1353 5907
rect 1487 5896 1533 5903
rect 1687 5896 1753 5903
rect 2507 5896 2553 5903
rect 2667 5896 2713 5903
rect 3267 5896 3333 5903
rect 3427 5896 3453 5903
rect 3587 5896 3653 5903
rect 3707 5896 3793 5903
rect 3887 5896 3973 5903
rect 4067 5893 4073 5907
rect 5227 5896 5253 5903
rect 5507 5896 5573 5903
rect 5667 5896 5733 5903
rect 687 5876 713 5883
rect 867 5873 873 5887
rect 2547 5876 2573 5883
rect 1847 5856 1893 5863
rect 2067 5856 2113 5863
rect 2367 5856 2433 5863
rect 2687 5856 2773 5863
rect 3067 5853 3073 5867
rect 4107 5853 4113 5867
rect 4127 5856 4193 5863
rect 4407 5853 4413 5867
rect 4707 5856 4772 5863
rect 4808 5853 4813 5867
rect 5220 5863 5233 5867
rect 5207 5856 5233 5863
rect 5220 5853 5233 5856
rect 5967 5856 6073 5863
rect 4273 5847 4287 5853
rect 527 5836 553 5843
rect 687 5836 733 5843
rect 827 5836 893 5843
rect 960 5843 973 5847
rect 947 5836 973 5843
rect 960 5833 973 5836
rect 1067 5836 1133 5843
rect 1187 5836 1233 5843
rect 3607 5843 3620 5847
rect 3700 5843 3713 5847
rect 3607 5836 3633 5843
rect 3687 5836 3713 5843
rect 3607 5833 3620 5836
rect 3700 5833 3713 5836
rect 3866 5833 3873 5847
rect 4567 5833 4573 5847
rect 2553 5827 2567 5833
rect 3433 5827 3447 5833
rect 796 5816 853 5823
rect 527 5796 593 5803
rect 647 5796 673 5803
rect 796 5803 803 5816
rect 2727 5816 2793 5823
rect 2967 5816 3033 5823
rect 3107 5816 3233 5823
rect 3247 5816 3273 5823
rect 3673 5827 3687 5833
rect 4247 5816 4473 5823
rect 4996 5823 5003 5853
rect 5687 5836 5793 5843
rect 4747 5816 5003 5823
rect 5116 5816 5393 5823
rect 747 5796 803 5803
rect 867 5796 893 5803
rect 947 5796 1033 5803
rect 1047 5796 1533 5803
rect 1547 5796 1593 5803
rect 1687 5796 2313 5803
rect 2327 5796 3013 5803
rect 3027 5796 4073 5803
rect 5116 5807 5123 5816
rect 5407 5813 5412 5827
rect 5433 5813 5434 5820
rect 4147 5796 4193 5803
rect 4307 5796 4913 5803
rect 4927 5796 5113 5803
rect 5256 5796 5293 5803
rect 787 5776 973 5783
rect 987 5776 1313 5783
rect 1427 5776 1763 5783
rect 1756 5767 1763 5776
rect 1788 5776 1823 5783
rect 107 5756 233 5763
rect 307 5756 333 5763
rect 527 5753 532 5767
rect 568 5756 693 5763
rect 807 5756 953 5763
rect 967 5756 1153 5763
rect 1167 5756 1573 5763
rect 1587 5756 1743 5763
rect 127 5736 273 5743
rect 287 5736 693 5743
rect 1467 5736 1713 5743
rect 1736 5743 1743 5756
rect 1767 5756 1793 5763
rect 1816 5763 1823 5776
rect 2127 5776 2173 5783
rect 2187 5776 2333 5783
rect 2347 5776 2792 5783
rect 2828 5776 2993 5783
rect 3047 5776 3383 5783
rect 1816 5756 2433 5763
rect 2527 5756 2673 5763
rect 2727 5756 2863 5763
rect 1736 5736 2133 5743
rect 2647 5736 2753 5743
rect 2767 5736 2833 5743
rect 2856 5743 2863 5756
rect 2927 5756 3313 5763
rect 3376 5763 3383 5776
rect 3407 5776 3513 5783
rect 3527 5776 4073 5783
rect 4187 5776 4233 5783
rect 4287 5776 4533 5783
rect 4547 5776 4593 5783
rect 4667 5776 4732 5783
rect 4768 5776 4913 5783
rect 4987 5776 5153 5783
rect 5256 5783 5263 5796
rect 5433 5807 5447 5813
rect 5427 5800 5447 5807
rect 5427 5796 5444 5800
rect 5427 5793 5440 5796
rect 5527 5796 5633 5803
rect 5907 5796 5973 5803
rect 5167 5776 5263 5783
rect 5287 5786 5300 5787
rect 5287 5773 5293 5786
rect 5427 5776 5473 5783
rect 3376 5756 3572 5763
rect 3608 5756 3873 5763
rect 3887 5756 3943 5763
rect 2856 5736 2953 5743
rect 3007 5736 3123 5743
rect 1507 5716 1733 5723
rect 2007 5716 2073 5723
rect 2087 5716 2813 5723
rect 2887 5716 3093 5723
rect 3116 5723 3123 5736
rect 3596 5743 3603 5753
rect 3287 5736 3603 5743
rect 3936 5743 3943 5756
rect 3967 5756 4093 5763
rect 4107 5756 4233 5763
rect 4496 5756 4693 5763
rect 4496 5743 4503 5756
rect 4707 5756 5033 5763
rect 5266 5753 5267 5760
rect 5288 5756 5433 5763
rect 3647 5736 3823 5743
rect 3936 5736 4503 5743
rect 3116 5716 3273 5723
rect 3327 5716 3793 5723
rect 3816 5723 3823 5736
rect 4627 5736 4833 5743
rect 5253 5743 5267 5753
rect 5253 5740 5413 5743
rect 5256 5736 5413 5740
rect 3816 5716 3873 5723
rect 4007 5716 4293 5723
rect 4487 5716 4653 5723
rect 4716 5716 4852 5723
rect 927 5696 1013 5703
rect 1027 5696 1233 5703
rect 1247 5696 1673 5703
rect 1767 5696 1833 5703
rect 2447 5696 2653 5703
rect 2847 5696 2953 5703
rect 2967 5696 3133 5703
rect 3267 5696 3293 5703
rect 3347 5696 3673 5703
rect 3687 5694 3692 5707
rect 3680 5693 3692 5694
rect 3728 5696 3753 5703
rect 4347 5696 4573 5703
rect 4716 5703 4723 5716
rect 4888 5716 5333 5723
rect 5347 5720 5683 5723
rect 5347 5716 5687 5720
rect 5673 5707 5687 5716
rect 4587 5696 4723 5703
rect 4747 5696 4792 5703
rect 4828 5696 5053 5703
rect 5107 5696 5373 5703
rect 5467 5696 5553 5703
rect 1327 5676 1373 5683
rect 1507 5676 2253 5683
rect 2267 5676 2713 5683
rect 2727 5676 2873 5683
rect 2987 5676 3323 5683
rect 127 5656 233 5663
rect 447 5656 553 5663
rect 767 5656 1213 5663
rect 1227 5656 1253 5663
rect 1527 5656 2033 5663
rect 2427 5656 2553 5663
rect 2667 5656 3133 5663
rect 3316 5663 3323 5676
rect 3407 5676 3433 5683
rect 3447 5676 3673 5683
rect 3727 5673 3733 5687
rect 3827 5676 3953 5683
rect 4147 5676 4773 5683
rect 4947 5676 4972 5683
rect 5008 5676 5173 5683
rect 5247 5676 5273 5683
rect 5587 5676 5773 5683
rect 3316 5656 3633 5663
rect 3787 5656 3852 5663
rect 3888 5656 4213 5663
rect 1307 5636 1353 5643
rect 1687 5636 1783 5643
rect 647 5613 653 5627
rect 847 5616 893 5623
rect 1776 5607 1783 5636
rect 1807 5636 1943 5643
rect 1936 5607 1943 5636
rect 3007 5636 3063 5643
rect 2647 5613 2653 5627
rect 2940 5623 2953 5627
rect 2927 5616 2953 5623
rect 2940 5613 2953 5616
rect 2133 5607 2147 5613
rect 3056 5607 3063 5636
rect 4056 5627 4063 5656
rect 4227 5656 4373 5663
rect 4427 5656 4593 5663
rect 4667 5656 5293 5663
rect 5387 5656 5733 5663
rect 5747 5656 5813 5663
rect 5827 5656 5993 5663
rect 4736 5636 4793 5643
rect 3147 5616 3213 5623
rect 3587 5616 3633 5623
rect 3687 5616 3733 5623
rect 4027 5623 4040 5627
rect 4027 5616 4053 5623
rect 4027 5613 4040 5616
rect 1267 5596 1333 5603
rect 1387 5596 1473 5603
rect 2227 5596 2273 5603
rect 4147 5596 4213 5603
rect 4267 5593 4273 5607
rect 4287 5593 4293 5607
rect 4736 5587 4743 5636
rect 4816 5636 4913 5643
rect 4816 5607 4823 5636
rect 5800 5623 5813 5627
rect 5787 5616 5813 5623
rect 5800 5613 5813 5616
rect 5173 5607 5187 5613
rect 5187 5596 5253 5603
rect 5620 5603 5633 5607
rect 5507 5596 5593 5603
rect 5607 5596 5633 5603
rect 5620 5593 5633 5596
rect 4727 5576 4743 5587
rect 4727 5573 4740 5576
rect 5827 5574 5833 5587
rect 5827 5573 5840 5574
rect 307 5553 313 5567
rect 640 5563 653 5567
rect 627 5556 653 5563
rect 640 5553 653 5556
rect 707 5563 720 5567
rect 707 5556 733 5563
rect 707 5553 720 5556
rect 1167 5563 1180 5567
rect 1167 5556 1193 5563
rect 1167 5553 1180 5556
rect 1547 5556 1613 5563
rect 2367 5556 2413 5563
rect 2807 5556 2833 5563
rect 3387 5556 3473 5563
rect 3527 5556 3613 5563
rect 3707 5556 3753 5563
rect 3807 5556 3873 5563
rect 4607 5556 4673 5563
rect 5040 5563 5053 5567
rect 5027 5556 5053 5563
rect 5040 5553 5053 5556
rect 5327 5553 5333 5567
rect 5487 5556 5533 5563
rect 5840 5566 5860 5567
rect 5667 5556 5753 5563
rect 93 5547 107 5553
rect 413 5547 427 5553
rect 487 5536 513 5543
rect 187 5516 253 5523
rect 627 5516 773 5523
rect 787 5516 833 5523
rect 1036 5523 1043 5553
rect 1753 5523 1767 5533
rect 856 5516 1043 5523
rect 1556 5516 1767 5523
rect 507 5496 653 5503
rect 856 5503 863 5516
rect 667 5496 863 5503
rect 1007 5496 1173 5503
rect 1367 5496 1453 5503
rect 1467 5496 1533 5503
rect 47 5476 313 5483
rect 867 5476 1213 5483
rect 1227 5476 1373 5483
rect 1556 5483 1563 5516
rect 2187 5516 2213 5523
rect 2507 5516 2613 5523
rect 2736 5523 2743 5553
rect 3913 5547 3927 5553
rect 2787 5536 2853 5543
rect 3087 5536 3153 5543
rect 2627 5516 2743 5523
rect 3147 5516 3333 5523
rect 3507 5516 3552 5523
rect 3588 5516 3653 5523
rect 4036 5523 4043 5553
rect 4513 5547 4527 5553
rect 5847 5563 5860 5566
rect 5847 5556 5873 5563
rect 5847 5553 5860 5556
rect 5967 5556 6013 5563
rect 4747 5536 4793 5543
rect 4907 5536 4953 5543
rect 5216 5536 5273 5543
rect 4333 5527 4347 5533
rect 3887 5516 4203 5523
rect 1647 5496 1793 5503
rect 1807 5496 1953 5503
rect 1967 5496 2153 5503
rect 2207 5496 2573 5503
rect 2667 5496 2753 5503
rect 2847 5496 3033 5503
rect 3147 5496 3253 5503
rect 3387 5496 3853 5503
rect 4196 5503 4203 5516
rect 4227 5516 4333 5523
rect 4467 5516 4773 5523
rect 4927 5516 5092 5523
rect 5216 5523 5223 5536
rect 5627 5536 5713 5543
rect 6067 5533 6073 5547
rect 5116 5516 5223 5523
rect 4196 5496 4393 5503
rect 4687 5496 4713 5503
rect 4767 5496 4833 5503
rect 4847 5496 4892 5503
rect 5116 5507 5123 5516
rect 5247 5516 5433 5523
rect 5787 5516 5893 5523
rect 5907 5516 6013 5523
rect 4928 5496 4973 5503
rect 5047 5496 5113 5503
rect 1487 5476 1563 5483
rect 1607 5476 1813 5483
rect 1827 5476 1993 5483
rect 2047 5476 2973 5483
rect 3167 5476 3213 5483
rect 3307 5476 3533 5483
rect 3547 5476 3693 5483
rect 3767 5476 4653 5483
rect 4707 5476 4913 5483
rect 5233 5483 5247 5493
rect 4967 5480 5247 5483
rect 5256 5496 5373 5503
rect 4967 5476 5243 5480
rect 1307 5456 1753 5463
rect 1767 5456 2073 5463
rect 2287 5456 2473 5463
rect 2776 5456 2892 5463
rect 107 5436 193 5443
rect 327 5436 653 5443
rect 767 5436 793 5443
rect 807 5436 833 5443
rect 1107 5436 1413 5443
rect 1727 5433 1733 5447
rect 1887 5436 1913 5443
rect 1987 5436 2133 5443
rect 2147 5436 2353 5443
rect 2776 5443 2783 5456
rect 2928 5456 2993 5463
rect 3047 5460 3124 5463
rect 3047 5456 3127 5460
rect 3113 5447 3127 5456
rect 3207 5456 3333 5463
rect 3347 5456 3493 5463
rect 3607 5456 3733 5463
rect 5256 5467 5263 5496
rect 5467 5496 5493 5503
rect 5587 5496 5613 5503
rect 5667 5493 5673 5507
rect 6067 5493 6073 5507
rect 5447 5476 5693 5483
rect 3867 5456 4053 5463
rect 4067 5456 4413 5463
rect 4527 5456 5193 5463
rect 5247 5456 5263 5467
rect 5247 5453 5260 5456
rect 5347 5463 5360 5467
rect 5347 5460 5363 5463
rect 5347 5453 5367 5460
rect 5387 5456 5773 5463
rect 5967 5456 5993 5463
rect 2736 5436 2783 5443
rect 147 5416 413 5423
rect 487 5416 553 5423
rect 576 5416 673 5423
rect 576 5387 583 5416
rect 807 5416 1053 5423
rect 1207 5416 1513 5423
rect 2367 5416 2393 5423
rect 2736 5423 2743 5436
rect 2807 5436 3092 5443
rect 3113 5440 3114 5447
rect 3167 5436 3413 5443
rect 3467 5436 3553 5443
rect 3687 5436 3813 5443
rect 3827 5436 3853 5443
rect 4087 5436 4153 5443
rect 4167 5436 4373 5443
rect 4387 5436 4473 5443
rect 4707 5436 4733 5443
rect 4807 5436 4953 5443
rect 5196 5443 5203 5453
rect 5353 5447 5367 5453
rect 5196 5436 5313 5443
rect 5367 5436 5513 5443
rect 5527 5436 5712 5443
rect 5748 5436 5833 5443
rect 5947 5436 6013 5443
rect 2487 5416 2743 5423
rect 1387 5396 1413 5403
rect 2467 5396 2493 5403
rect 2676 5387 2683 5416
rect 2767 5416 2903 5423
rect 2896 5387 2903 5416
rect 2947 5416 3163 5423
rect 3013 5387 3027 5393
rect 3156 5387 3163 5416
rect 3187 5416 3293 5423
rect 3516 5416 3613 5423
rect 3227 5396 3293 5403
rect 3387 5396 3433 5403
rect 3516 5387 3523 5416
rect 3787 5416 3913 5423
rect 4027 5416 4072 5423
rect 4108 5416 4173 5423
rect 4327 5416 4393 5423
rect 4407 5416 4613 5423
rect 4667 5416 4833 5423
rect 5007 5416 5053 5423
rect 5067 5416 5493 5423
rect 5507 5416 5593 5423
rect 5927 5416 5993 5423
rect 4207 5396 4233 5403
rect 4527 5396 4553 5403
rect 4687 5393 4693 5407
rect 247 5383 260 5387
rect 247 5376 273 5383
rect 247 5373 260 5376
rect 327 5376 373 5383
rect 727 5373 733 5387
rect 927 5376 993 5383
rect 1047 5373 1053 5387
rect 1127 5376 1173 5383
rect 1276 5380 1313 5383
rect 1273 5376 1313 5380
rect 1273 5367 1287 5376
rect 1327 5373 1333 5387
rect 1747 5373 1753 5387
rect 1867 5376 1933 5383
rect 2187 5376 2233 5383
rect 2740 5383 2753 5387
rect 2727 5376 2753 5383
rect 2740 5373 2753 5376
rect 4027 5376 4073 5383
rect 4127 5373 4133 5387
rect 4287 5373 4293 5387
rect 4647 5376 4733 5383
rect 4907 5376 4993 5383
rect 5127 5376 5173 5383
rect 5187 5376 5213 5383
rect 5647 5376 5733 5383
rect 5980 5383 5993 5387
rect 5967 5376 5993 5383
rect 5980 5373 5993 5376
rect 3307 5333 3313 5347
rect 3587 5336 3653 5343
rect 3887 5336 3953 5343
rect 4247 5334 4253 5347
rect 4240 5333 4253 5334
rect 4640 5343 4653 5347
rect 4627 5336 4653 5343
rect 4640 5333 4653 5336
rect 5306 5333 5307 5340
rect 5987 5336 6033 5343
rect 1453 5327 1467 5333
rect 687 5316 753 5323
rect 847 5316 893 5323
rect 1107 5316 1153 5323
rect 1616 5303 1623 5333
rect 3353 5327 3367 5333
rect 1767 5313 1773 5327
rect 2507 5316 2553 5323
rect 2607 5316 2653 5323
rect 2747 5316 2833 5323
rect 2927 5316 2953 5323
rect 3113 5307 3127 5313
rect 1407 5296 1623 5303
rect 2787 5293 2793 5307
rect 3327 5296 3453 5303
rect 3696 5303 3703 5333
rect 3813 5327 3827 5333
rect 4247 5316 4313 5323
rect 4407 5316 4453 5323
rect 4687 5316 4713 5323
rect 5293 5327 5307 5333
rect 5793 5327 5807 5333
rect 5306 5320 5307 5327
rect 5328 5313 5333 5327
rect 5347 5316 5393 5323
rect 3567 5296 3703 5303
rect 4267 5303 4280 5307
rect 4267 5293 4283 5303
rect 4647 5296 4713 5303
rect 127 5276 153 5283
rect 387 5276 453 5283
rect 607 5276 793 5283
rect 1027 5276 1093 5283
rect 1327 5276 1433 5283
rect 1527 5276 1653 5283
rect 1667 5276 1713 5283
rect 1827 5276 1873 5283
rect 1967 5276 2113 5283
rect 2127 5276 2173 5283
rect 2267 5276 2313 5283
rect 2336 5276 2833 5283
rect 987 5256 1392 5263
rect 1428 5256 1453 5263
rect 2336 5263 2343 5276
rect 2887 5276 2913 5283
rect 2987 5276 3033 5283
rect 3047 5276 3253 5283
rect 3327 5276 3433 5283
rect 3687 5276 4253 5283
rect 4276 5283 4283 5293
rect 5287 5303 5300 5307
rect 5287 5293 5303 5303
rect 5387 5296 5443 5303
rect 4276 5276 4913 5283
rect 4967 5276 5193 5283
rect 5296 5283 5303 5293
rect 5296 5276 5353 5283
rect 5436 5283 5443 5296
rect 5436 5276 5573 5283
rect 5596 5276 5793 5283
rect 1587 5256 2343 5263
rect 2407 5256 2533 5263
rect 2547 5256 2712 5263
rect 2748 5253 2752 5267
rect 2788 5253 2793 5267
rect 2867 5256 2912 5263
rect 2948 5256 3133 5263
rect 3467 5256 3613 5263
rect 3627 5256 3773 5263
rect 3827 5256 4093 5263
rect 4247 5256 4333 5263
rect 4567 5256 4633 5263
rect 4647 5256 4673 5263
rect 5107 5256 5153 5263
rect 5167 5256 5323 5263
rect 193 5247 207 5253
rect 627 5236 673 5243
rect 1127 5233 1133 5247
rect 1227 5236 1332 5243
rect 1368 5236 1653 5243
rect 1807 5236 1832 5243
rect 1868 5236 1913 5243
rect 2007 5236 2273 5243
rect 2327 5236 2493 5243
rect 2516 5236 2553 5243
rect 687 5216 853 5223
rect 927 5216 1113 5223
rect 1207 5216 1393 5223
rect 1527 5216 1573 5223
rect 1916 5223 1923 5233
rect 1916 5216 2053 5223
rect 2307 5216 2393 5223
rect 2516 5223 2523 5236
rect 2707 5236 2773 5243
rect 2847 5236 2933 5243
rect 3007 5236 3193 5243
rect 3247 5236 3273 5243
rect 3287 5236 3373 5243
rect 3547 5236 3573 5243
rect 3627 5236 3673 5243
rect 3727 5236 3813 5243
rect 3827 5236 4473 5243
rect 4707 5236 4753 5243
rect 4847 5236 4893 5243
rect 4907 5236 5263 5243
rect 2447 5216 2523 5223
rect 2536 5216 2653 5223
rect 727 5196 793 5203
rect 1147 5196 1293 5203
rect 1347 5196 1413 5203
rect 2536 5203 2543 5216
rect 2667 5216 2953 5223
rect 3067 5216 3332 5223
rect 3368 5216 3933 5223
rect 4007 5216 4073 5223
rect 4127 5216 4193 5223
rect 4296 5216 4413 5223
rect 1567 5196 2543 5203
rect 2567 5196 2772 5203
rect 2808 5196 2903 5203
rect 2896 5187 2903 5196
rect 3056 5203 3063 5213
rect 4296 5203 4303 5216
rect 4487 5216 4693 5223
rect 4747 5216 4853 5223
rect 4927 5216 5033 5223
rect 5256 5223 5263 5236
rect 5287 5233 5293 5247
rect 5316 5243 5323 5256
rect 5596 5263 5603 5276
rect 5807 5276 5932 5283
rect 5968 5276 6013 5283
rect 5467 5256 5603 5263
rect 5316 5236 5733 5243
rect 5947 5236 5993 5243
rect 5256 5216 5893 5223
rect 3007 5196 3063 5203
rect 3576 5196 4303 5203
rect 4356 5196 4713 5203
rect 127 5176 253 5183
rect 267 5176 553 5183
rect 567 5176 1693 5183
rect 1887 5176 2093 5183
rect 2147 5176 2713 5183
rect 2907 5176 2932 5183
rect 2968 5176 3133 5183
rect 3147 5176 3293 5183
rect 3576 5183 3583 5196
rect 3307 5176 3583 5183
rect 4356 5183 4363 5196
rect 4847 5196 5133 5203
rect 5176 5196 5273 5203
rect 3607 5176 4363 5183
rect 4527 5176 4933 5183
rect 5176 5183 5183 5196
rect 5047 5176 5183 5183
rect 5207 5176 5513 5183
rect 5987 5176 6083 5183
rect 587 5156 723 5163
rect 716 5147 723 5156
rect 1107 5153 1113 5167
rect 1407 5153 1413 5167
rect 1467 5156 1573 5163
rect 1787 5156 1913 5163
rect 1927 5156 2073 5163
rect 2087 5156 2353 5163
rect 2376 5156 2432 5163
rect 667 5133 673 5147
rect 727 5136 833 5143
rect 847 5136 1153 5143
rect 1207 5136 1232 5143
rect 1268 5136 1293 5143
rect 1387 5136 1573 5143
rect 1587 5136 1713 5143
rect 1867 5136 1943 5143
rect 1936 5107 1943 5136
rect 2376 5143 2383 5156
rect 2468 5156 2513 5163
rect 2527 5156 2573 5163
rect 2687 5156 3273 5163
rect 3327 5156 3653 5163
rect 4087 5156 4273 5163
rect 4676 5156 4873 5163
rect 1967 5136 2383 5143
rect 2427 5136 2633 5143
rect 2747 5136 3073 5143
rect 3127 5136 3233 5143
rect 3327 5136 3352 5143
rect 3388 5136 3553 5143
rect 3687 5136 3733 5143
rect 3907 5136 4053 5143
rect 4107 5136 4273 5143
rect 4367 5136 4453 5143
rect 4676 5143 4683 5156
rect 4947 5156 5213 5163
rect 5687 5156 6053 5163
rect 6076 5163 6083 5176
rect 6076 5156 6123 5163
rect 4607 5136 4683 5143
rect 2987 5116 3013 5123
rect 3393 5116 3433 5123
rect 3393 5107 3407 5116
rect 4427 5116 4493 5123
rect 4636 5123 4643 5136
rect 4707 5136 4833 5143
rect 4947 5136 5013 5143
rect 5127 5136 5173 5143
rect 5247 5136 5293 5143
rect 5407 5136 5473 5143
rect 5987 5136 6033 5143
rect 4636 5116 4673 5123
rect 5527 5116 5693 5123
rect 5927 5116 6073 5123
rect 6116 5116 6123 5156
rect 107 5096 153 5103
rect 607 5096 673 5103
rect 1127 5096 1193 5103
rect 1247 5093 1253 5107
rect 1887 5093 1893 5107
rect 2107 5096 2193 5103
rect 3560 5103 3573 5107
rect 3547 5096 3573 5103
rect 3560 5093 3573 5096
rect 3647 5093 3653 5107
rect 3747 5103 3760 5107
rect 3747 5096 3773 5103
rect 3747 5093 3760 5096
rect 4307 5096 4353 5103
rect 4747 5096 4793 5103
rect 4967 5096 5033 5103
rect 5327 5096 5393 5103
rect 6067 5096 6103 5103
rect 793 5067 807 5073
rect 2507 5076 2533 5083
rect 4427 5076 4473 5083
rect 5607 5076 5673 5083
rect 5907 5076 5973 5083
rect 6027 5076 6073 5083
rect 6096 5083 6103 5096
rect 6096 5076 6123 5083
rect 973 5067 987 5073
rect 1107 5056 1133 5063
rect 2647 5054 2653 5067
rect 2640 5053 2653 5054
rect 3107 5053 3113 5067
rect 5967 5066 5980 5067
rect 5967 5053 5973 5066
rect 307 5036 393 5043
rect 507 5043 520 5047
rect 507 5036 533 5043
rect 507 5033 520 5036
rect 627 5036 693 5043
rect 747 5036 813 5043
rect 947 5036 1013 5043
rect 1127 5036 1173 5043
rect 1267 5036 1333 5043
rect 1427 5036 1493 5043
rect 1587 5036 1633 5043
rect 1980 5043 1993 5047
rect 1967 5036 1993 5043
rect 1980 5033 1993 5036
rect 2207 5036 2253 5043
rect 2487 5036 2553 5043
rect 2647 5036 2713 5043
rect 2927 5033 2933 5047
rect 3067 5033 3072 5047
rect 3108 5036 3153 5043
rect 3260 5043 3273 5047
rect 3247 5036 3273 5043
rect 3260 5033 3273 5036
rect 3327 5036 3373 5043
rect 3607 5043 3620 5047
rect 3607 5036 3633 5043
rect 3607 5033 3620 5036
rect 3847 5033 3852 5047
rect 3888 5036 3973 5043
rect 4027 5036 4093 5043
rect 4147 5036 4233 5043
rect 4667 5036 4753 5043
rect 5007 5033 5013 5047
rect 5067 5036 5133 5043
rect 5307 5036 5413 5043
rect 5480 5043 5492 5047
rect 5467 5036 5492 5043
rect 5480 5033 5492 5036
rect 5528 5043 5540 5047
rect 5528 5036 5553 5043
rect 5528 5033 5540 5036
rect 5760 5043 5773 5047
rect 5747 5036 5773 5043
rect 5760 5033 5773 5036
rect 893 5027 907 5033
rect 1013 5027 1027 5033
rect 2293 5027 2307 5033
rect 1087 5016 1113 5023
rect 2393 5027 2407 5033
rect 2627 5013 2633 5027
rect 2873 5023 2887 5033
rect 3413 5027 3427 5033
rect 4013 5027 4027 5033
rect 2787 5016 2887 5023
rect 3106 5013 3107 5020
rect 3128 5013 3133 5027
rect 3307 5013 3313 5027
rect 3707 5016 3733 5023
rect 4356 5016 4393 5023
rect 227 4996 293 5003
rect 407 4996 653 5003
rect 767 4996 873 5003
rect 1047 4996 1473 5003
rect 1667 4996 1713 5003
rect 1736 4996 2143 5003
rect 587 4976 653 4983
rect 727 4976 793 4983
rect 807 4973 813 4987
rect 987 4976 1053 4983
rect 1067 4976 1093 4983
rect 1147 4976 1193 4983
rect 1207 4976 1323 4983
rect 1316 4967 1323 4976
rect 1387 4973 1393 4987
rect 1736 4983 1743 4996
rect 2136 4987 2143 4996
rect 2387 4996 2473 5003
rect 3093 5003 3107 5013
rect 2527 5000 3107 5003
rect 2527 4996 3103 5000
rect 3207 4996 3233 5003
rect 3287 4996 3593 5003
rect 3647 4996 3793 5003
rect 3836 4996 3892 5003
rect 1616 4976 1743 4983
rect 127 4956 173 4963
rect 387 4956 553 4963
rect 567 4956 613 4963
rect 667 4956 893 4963
rect 1327 4956 1493 4963
rect 1616 4963 1623 4976
rect 1787 4976 2013 4983
rect 2147 4976 2313 4983
rect 2327 4976 2673 4983
rect 2727 4976 2753 4983
rect 2807 4976 2893 4983
rect 3027 4976 3113 4983
rect 3227 4976 3352 4983
rect 3388 4976 3653 4983
rect 3836 4983 3843 4996
rect 3928 4996 4113 5003
rect 4167 4996 4292 5003
rect 4356 5003 4363 5016
rect 4328 4996 4363 5003
rect 4507 4996 4533 5003
rect 4576 5007 4583 5033
rect 4896 5020 4903 5033
rect 4893 5007 4907 5020
rect 4576 4996 4593 5007
rect 4580 4993 4593 4996
rect 4616 4996 4853 5003
rect 3667 4976 3843 4983
rect 3867 4976 3973 4983
rect 4287 4976 4353 4983
rect 4447 4976 4533 4983
rect 4547 4976 4573 4983
rect 4616 4983 4623 4996
rect 5856 5003 5863 5033
rect 4947 4996 5863 5003
rect 4587 4976 4623 4983
rect 4807 4976 5033 4983
rect 5047 4976 5073 4983
rect 5147 4976 5193 4983
rect 5407 4976 5433 4983
rect 5487 4976 5673 4983
rect 5887 4976 5993 4983
rect 1507 4956 1623 4963
rect 1647 4956 2053 4963
rect 2116 4956 2513 4963
rect 107 4936 193 4943
rect 487 4936 593 4943
rect 847 4936 1113 4943
rect 1687 4936 1873 4943
rect 2116 4943 2123 4956
rect 2647 4956 2913 4963
rect 2967 4956 3433 4963
rect 3447 4956 3753 4963
rect 3767 4956 3793 4963
rect 3816 4956 4332 4963
rect 1947 4936 2123 4943
rect 2247 4936 2393 4943
rect 2587 4936 2872 4943
rect 2908 4936 3373 4943
rect 3816 4943 3823 4956
rect 4368 4956 4903 4963
rect 3427 4936 3823 4943
rect 3947 4936 4133 4943
rect 4527 4936 4792 4943
rect 4828 4936 4873 4943
rect 4896 4943 4903 4956
rect 4927 4956 5053 4963
rect 6033 4963 6047 4973
rect 5667 4960 6047 4963
rect 5667 4956 6043 4960
rect 4896 4936 4953 4943
rect 4967 4936 5153 4943
rect 5167 4936 5253 4943
rect 5336 4936 5393 4943
rect 27 4916 253 4923
rect 276 4920 413 4923
rect 273 4916 413 4920
rect 273 4907 287 4916
rect 547 4916 653 4923
rect 667 4916 1173 4923
rect 1287 4916 1312 4923
rect 1348 4916 1433 4923
rect 1667 4916 1713 4923
rect 1827 4916 2292 4923
rect 2328 4916 2513 4923
rect 2667 4916 2713 4923
rect 2867 4916 3143 4923
rect 67 4896 243 4903
rect 236 4867 243 4896
rect 327 4896 373 4903
rect 767 4896 843 4903
rect 467 4876 493 4883
rect 413 4867 427 4873
rect 836 4867 843 4896
rect 867 4896 1003 4903
rect 996 4867 1003 4896
rect 1067 4896 1193 4903
rect 1407 4896 1732 4903
rect 1768 4896 1863 4903
rect 1173 4867 1187 4873
rect 1856 4867 1863 4896
rect 1887 4896 1993 4903
rect 2007 4896 2092 4903
rect 2128 4896 2213 4903
rect 2227 4896 2503 4903
rect 2496 4883 2503 4896
rect 2547 4896 2953 4903
rect 3047 4896 3113 4903
rect 3136 4903 3143 4916
rect 3167 4916 3453 4923
rect 3467 4916 4193 4923
rect 4247 4916 4313 4923
rect 4387 4916 4633 4923
rect 4687 4916 4772 4923
rect 4808 4916 4832 4923
rect 4868 4916 4993 4923
rect 5336 4923 5343 4936
rect 5947 4936 6033 4943
rect 5227 4916 5343 4923
rect 5367 4916 5433 4923
rect 5927 4916 5953 4923
rect 6007 4916 6033 4923
rect 3136 4896 3233 4903
rect 3307 4896 3443 4903
rect 2496 4876 2573 4883
rect 2753 4867 2767 4873
rect 3436 4867 3443 4896
rect 3527 4896 3553 4903
rect 3567 4896 4012 4903
rect 4048 4893 4053 4907
rect 4247 4896 4333 4903
rect 4427 4896 4493 4903
rect 4567 4896 4713 4903
rect 4987 4896 5093 4903
rect 5147 4896 5353 4903
rect 5427 4896 5513 4903
rect 5687 4896 5733 4903
rect 5927 4896 6053 4903
rect 4347 4876 4373 4883
rect 5907 4876 5933 4883
rect 487 4856 553 4863
rect 607 4856 673 4863
rect 1467 4856 1553 4863
rect 1707 4853 1713 4867
rect 1967 4856 2013 4863
rect 2107 4856 2153 4863
rect 2507 4856 2593 4863
rect 2820 4863 2833 4867
rect 2687 4856 2753 4863
rect 2807 4856 2833 4863
rect 2820 4853 2833 4856
rect 2887 4853 2893 4867
rect 3267 4856 3313 4863
rect 3487 4856 3533 4863
rect 3647 4853 3653 4867
rect 3907 4856 3953 4863
rect 4047 4863 4060 4867
rect 4047 4856 4073 4863
rect 4047 4853 4060 4856
rect 4127 4856 4233 4863
rect 4287 4856 4353 4863
rect 4587 4856 4633 4863
rect 5027 4856 5093 4863
rect 5116 4856 5153 4863
rect 2207 4833 2213 4847
rect 2527 4833 2533 4847
rect 5116 4843 5123 4856
rect 5587 4856 5653 4863
rect 5807 4853 5813 4867
rect 5913 4847 5927 4853
rect 5067 4836 5123 4843
rect 5207 4836 5233 4843
rect 1227 4816 1293 4823
rect 3547 4816 3613 4823
rect 3687 4813 3693 4827
rect 3847 4816 3893 4823
rect 4787 4816 4853 4823
rect 5707 4816 5753 4823
rect 6027 4813 6032 4827
rect 6068 4816 6123 4823
rect 447 4796 533 4803
rect 1336 4796 1433 4803
rect 96 4763 103 4793
rect 813 4783 827 4793
rect 727 4776 827 4783
rect 1336 4783 1343 4796
rect 2327 4796 2373 4803
rect 2667 4796 2733 4803
rect 2827 4796 2913 4803
rect 1267 4776 1343 4783
rect 1647 4773 1653 4787
rect 2367 4776 2413 4783
rect 2467 4776 2493 4783
rect 3776 4783 3783 4813
rect 3987 4796 4053 4803
rect 4367 4803 4380 4807
rect 4367 4796 4393 4803
rect 4367 4793 4380 4796
rect 4607 4796 4653 4803
rect 5087 4796 5133 4803
rect 5547 4793 5553 4807
rect 5567 4796 5633 4803
rect 3536 4776 3783 4783
rect 96 4756 213 4763
rect 287 4756 353 4763
rect 447 4756 1423 4763
rect 247 4736 313 4743
rect 327 4736 593 4743
rect 827 4736 1153 4743
rect 1167 4736 1212 4743
rect 1248 4736 1393 4743
rect 1416 4743 1423 4756
rect 1547 4756 1812 4763
rect 1848 4756 2173 4763
rect 2187 4756 2313 4763
rect 2327 4756 2533 4763
rect 2627 4756 2673 4763
rect 2787 4756 2813 4763
rect 2927 4756 3113 4763
rect 3136 4756 3273 4763
rect 1416 4736 1733 4743
rect 1816 4743 1823 4753
rect 1816 4736 1933 4743
rect 2047 4736 2333 4743
rect 2356 4736 2833 4743
rect 387 4716 453 4723
rect 727 4716 1113 4723
rect 1416 4720 1773 4723
rect 1413 4716 1773 4720
rect 1413 4707 1427 4716
rect 1967 4716 2013 4723
rect 2147 4716 2213 4723
rect 2356 4723 2363 4736
rect 3136 4743 3143 4756
rect 3327 4756 3493 4763
rect 3536 4763 3543 4776
rect 4787 4776 4933 4783
rect 6047 4773 6053 4787
rect 3507 4756 3543 4763
rect 3687 4756 3793 4763
rect 3807 4756 4053 4763
rect 4107 4756 4193 4763
rect 4207 4756 4413 4763
rect 4567 4756 4633 4763
rect 4647 4756 4693 4763
rect 4707 4756 4833 4763
rect 4887 4756 5033 4763
rect 5096 4756 5212 4763
rect 3047 4736 3143 4743
rect 3167 4736 3273 4743
rect 3347 4736 3373 4743
rect 3507 4736 3553 4743
rect 3747 4736 3853 4743
rect 3867 4736 3933 4743
rect 4047 4736 4073 4743
rect 4187 4736 4253 4743
rect 4347 4733 4353 4747
rect 4487 4736 4593 4743
rect 4647 4736 4733 4743
rect 2267 4716 2363 4723
rect 2387 4716 2613 4723
rect 2627 4716 2833 4723
rect 2947 4716 3153 4723
rect 3167 4716 3193 4723
rect 3287 4716 3463 4723
rect 687 4696 933 4703
rect 1027 4696 1303 4703
rect 927 4676 1053 4683
rect 1127 4676 1253 4683
rect 1296 4683 1303 4696
rect 1587 4696 1693 4703
rect 1796 4696 1873 4703
rect 1296 4676 1593 4683
rect 1796 4683 1803 4696
rect 1967 4696 2033 4703
rect 2056 4696 2653 4703
rect 2056 4683 2063 4696
rect 2707 4696 2732 4703
rect 2768 4696 3073 4703
rect 3227 4696 3293 4703
rect 3367 4696 3433 4703
rect 3456 4703 3463 4716
rect 3487 4716 3533 4723
rect 3736 4723 3743 4733
rect 3647 4716 3743 4723
rect 3907 4716 3952 4723
rect 3988 4716 4132 4723
rect 4168 4716 4213 4723
rect 4476 4723 4483 4733
rect 4887 4736 4993 4743
rect 5096 4743 5103 4756
rect 5248 4756 5373 4763
rect 5527 4756 5793 4763
rect 5807 4756 5933 4763
rect 5067 4736 5103 4743
rect 5127 4736 5573 4743
rect 5647 4736 5893 4743
rect 6053 4733 6054 4740
rect 6053 4727 6067 4733
rect 4307 4716 4483 4723
rect 4507 4716 4713 4723
rect 4867 4716 4953 4723
rect 5047 4716 5072 4723
rect 5108 4716 5253 4723
rect 5327 4716 5353 4723
rect 5767 4716 6032 4723
rect 6053 4720 6054 4727
rect 3456 4696 3603 4703
rect 1647 4676 1803 4683
rect 1956 4676 2063 4683
rect 407 4656 753 4663
rect 867 4656 953 4663
rect 967 4656 1433 4663
rect 1956 4663 1963 4676
rect 2087 4676 2392 4683
rect 2428 4676 2593 4683
rect 2687 4676 3373 4683
rect 3387 4676 3533 4683
rect 3596 4683 3603 4696
rect 3627 4696 3793 4703
rect 3896 4696 4193 4703
rect 3896 4683 3903 4696
rect 4207 4696 4513 4703
rect 4587 4696 4912 4703
rect 4948 4696 5113 4703
rect 5136 4696 5233 4703
rect 3596 4676 3903 4683
rect 3927 4676 4553 4683
rect 4727 4676 4913 4683
rect 5136 4683 5143 4696
rect 5247 4696 5273 4703
rect 5347 4696 5433 4703
rect 5487 4696 5613 4703
rect 4927 4676 5143 4683
rect 5167 4676 5413 4683
rect 5507 4676 5853 4683
rect 5867 4676 5973 4683
rect 6067 4676 6103 4683
rect 1807 4656 1963 4663
rect 1987 4656 2053 4663
rect 2207 4656 2292 4663
rect 2328 4656 2413 4663
rect 2487 4656 2513 4663
rect 2567 4656 2933 4663
rect 2947 4656 3033 4663
rect 3056 4656 3313 4663
rect 127 4636 433 4643
rect 607 4633 612 4647
rect 648 4636 1172 4643
rect 1208 4636 1233 4643
rect 1287 4636 1373 4643
rect 1607 4636 1673 4643
rect 1787 4636 1853 4643
rect 1867 4636 2073 4643
rect 2127 4636 2252 4643
rect 2288 4636 2493 4643
rect 2547 4636 2692 4643
rect 2728 4633 2733 4647
rect 2747 4636 2863 4643
rect 96 4616 193 4623
rect 96 4587 103 4616
rect 207 4616 253 4623
rect 587 4616 793 4623
rect 807 4616 993 4623
rect 1167 4616 1333 4623
rect 1507 4616 1553 4623
rect 1687 4616 2373 4623
rect 2427 4616 2712 4623
rect 2856 4623 2863 4636
rect 3056 4643 3063 4656
rect 3336 4656 3472 4663
rect 2887 4636 3063 4643
rect 3336 4643 3343 4656
rect 3508 4653 3513 4667
rect 3567 4656 3673 4663
rect 3687 4653 3693 4667
rect 3747 4656 3833 4663
rect 3847 4656 4153 4663
rect 4267 4656 4293 4663
rect 4347 4656 4372 4663
rect 4408 4654 4413 4667
rect 4400 4653 4413 4654
rect 4827 4653 4833 4667
rect 5027 4656 5053 4663
rect 5107 4656 5153 4663
rect 5327 4656 5373 4663
rect 5627 4656 5753 4663
rect 5767 4656 5813 4663
rect 6047 4656 6073 4663
rect 5913 4647 5927 4653
rect 3087 4636 3343 4643
rect 3356 4636 3913 4643
rect 2748 4616 2843 4623
rect 2856 4616 2993 4623
rect 2836 4607 2843 4616
rect 3356 4623 3363 4636
rect 4027 4636 4173 4643
rect 4396 4636 4773 4643
rect 4396 4627 4403 4636
rect 4827 4636 4873 4643
rect 4967 4636 5033 4643
rect 5087 4636 5393 4643
rect 5787 4636 5873 4643
rect 6096 4643 6103 4676
rect 6076 4640 6103 4643
rect 6073 4636 6103 4640
rect 6073 4627 6087 4636
rect 3227 4616 3363 4623
rect 3427 4616 3473 4623
rect 3547 4616 3673 4623
rect 3767 4616 3993 4623
rect 4047 4616 4072 4623
rect 4093 4613 4094 4620
rect 4367 4616 4392 4623
rect 4428 4616 4873 4623
rect 4887 4616 4993 4623
rect 5067 4616 5203 4623
rect 4093 4607 4107 4613
rect 2107 4596 2153 4603
rect 2287 4593 2293 4607
rect 2627 4603 2640 4607
rect 2627 4593 2647 4603
rect 2836 4596 2853 4607
rect 2840 4593 2853 4596
rect 4547 4596 4613 4603
rect 4627 4596 4733 4603
rect 2633 4587 2647 4593
rect 2933 4587 2947 4593
rect 5196 4587 5203 4616
rect 5247 4616 5293 4623
rect 5907 4616 6033 4623
rect 5747 4596 5847 4603
rect 5833 4587 5847 4596
rect 547 4576 633 4583
rect 1087 4576 1153 4583
rect 1567 4583 1580 4587
rect 1567 4576 1593 4583
rect 1567 4573 1580 4576
rect 1767 4576 1813 4583
rect 2260 4583 2273 4587
rect 2247 4576 2273 4583
rect 2260 4573 2273 4576
rect 2400 4583 2413 4587
rect 2387 4576 2413 4583
rect 2400 4573 2413 4576
rect 2747 4576 2793 4583
rect 2887 4573 2893 4587
rect 3687 4583 3700 4587
rect 3687 4576 3713 4583
rect 3687 4573 3700 4576
rect 3767 4576 3833 4583
rect 4047 4576 4113 4583
rect 5948 4576 5993 4583
rect 993 4567 1007 4573
rect 1047 4556 1093 4563
rect 2847 4553 2853 4567
rect 4647 4556 4693 4563
rect 4867 4553 4873 4567
rect 1687 4536 1733 4543
rect 2267 4536 2313 4543
rect 3507 4536 3533 4543
rect 4987 4536 5013 4543
rect 5907 4536 5933 4543
rect 6027 4536 6053 4543
rect 307 4516 373 4523
rect 1067 4513 1073 4527
rect 1147 4523 1160 4527
rect 1147 4516 1173 4523
rect 1147 4513 1160 4516
rect 1287 4523 1300 4527
rect 1287 4516 1313 4523
rect 1287 4513 1300 4516
rect 1487 4516 1573 4523
rect 1927 4516 1993 4523
rect 2307 4516 2353 4523
rect 2407 4516 2493 4523
rect 2667 4516 2753 4523
rect 2867 4516 2913 4523
rect 2927 4516 3013 4523
rect 3147 4516 3213 4523
rect 3847 4513 3853 4527
rect 4407 4516 4473 4523
rect 4787 4516 4893 4523
rect 4947 4516 5033 4523
rect 5307 4516 5333 4523
rect 5387 4516 5473 4523
rect 5567 4516 5613 4523
rect 213 4507 227 4513
rect 267 4476 473 4483
rect 656 4483 663 4513
rect 656 4476 713 4483
rect 836 4483 843 4513
rect 2173 4507 2187 4513
rect 767 4476 843 4483
rect 1167 4476 1233 4483
rect 1307 4476 1353 4483
rect 1367 4476 1433 4483
rect 1567 4473 1573 4487
rect 1827 4476 2013 4483
rect 2216 4483 2223 4513
rect 2613 4507 2627 4513
rect 3093 4507 3107 4513
rect 3573 4507 3587 4513
rect 2547 4496 2573 4503
rect 2860 4506 2873 4507
rect 2867 4493 2873 4506
rect 2967 4496 3013 4503
rect 3513 4493 3514 4500
rect 3773 4507 3787 4513
rect 3933 4507 3947 4513
rect 4173 4507 4187 4513
rect 3513 4487 3527 4493
rect 4333 4507 4347 4513
rect 5073 4507 5087 4513
rect 4387 4506 4400 4507
rect 4387 4493 4393 4506
rect 5256 4487 5263 4513
rect 5693 4507 5707 4513
rect 5853 4507 5867 4513
rect 2067 4476 2223 4483
rect 2287 4476 2353 4483
rect 2527 4476 2553 4483
rect 2576 4476 2803 4483
rect 593 4467 607 4473
rect 1027 4456 1113 4463
rect 1127 4456 1223 4463
rect 927 4436 1173 4443
rect 1216 4443 1223 4456
rect 1247 4453 1253 4467
rect 1467 4456 1673 4463
rect 1687 4456 1713 4463
rect 2007 4456 2092 4463
rect 2128 4456 2233 4463
rect 2307 4453 2313 4467
rect 2336 4456 2413 4463
rect 1216 4436 1393 4443
rect 1507 4436 1623 4443
rect 1616 4427 1623 4436
rect 1667 4436 1913 4443
rect 2087 4436 2213 4443
rect 2336 4443 2343 4456
rect 2576 4463 2583 4476
rect 2487 4456 2583 4463
rect 2707 4453 2713 4467
rect 2767 4463 2780 4467
rect 2796 4463 2803 4476
rect 2847 4476 3253 4483
rect 3327 4476 3492 4483
rect 3513 4480 3514 4487
rect 3567 4476 3633 4483
rect 3687 4476 3793 4483
rect 3807 4476 4013 4483
rect 4067 4476 4093 4483
rect 4247 4476 4292 4483
rect 4328 4476 4413 4483
rect 4707 4476 5213 4483
rect 5267 4476 5513 4483
rect 5687 4476 5732 4483
rect 5768 4473 5773 4487
rect 5927 4476 5993 4483
rect 2767 4453 2783 4463
rect 2796 4456 2953 4463
rect 3007 4456 3233 4463
rect 3287 4456 3453 4463
rect 3467 4456 3563 4463
rect 2227 4436 2343 4443
rect 2447 4436 2572 4443
rect 2608 4436 2713 4443
rect 2776 4443 2783 4453
rect 2776 4436 3053 4443
rect 3207 4436 3333 4443
rect 3427 4436 3533 4443
rect 3556 4443 3563 4456
rect 3627 4456 3673 4463
rect 3747 4456 3972 4463
rect 3993 4453 3994 4460
rect 4047 4456 4153 4463
rect 4227 4456 4253 4463
rect 4387 4456 4453 4463
rect 4467 4456 4533 4463
rect 4667 4456 4733 4463
rect 4807 4456 4833 4463
rect 4907 4456 5023 4463
rect 3556 4436 3693 4443
rect 3993 4443 4007 4453
rect 3827 4440 4007 4443
rect 3827 4436 4003 4440
rect 4096 4436 4353 4443
rect 107 4416 373 4423
rect 587 4416 653 4423
rect 1087 4416 1193 4423
rect 1387 4416 1453 4423
rect 1627 4416 1863 4423
rect 56 4387 63 4413
rect 1573 4407 1587 4413
rect 87 4396 213 4403
rect 227 4396 253 4403
rect 447 4396 873 4403
rect 1147 4396 1213 4403
rect 1267 4396 1493 4403
rect 1507 4396 1533 4403
rect 1667 4396 1712 4403
rect 1748 4396 1833 4403
rect 1856 4403 1863 4416
rect 1907 4416 2012 4423
rect 2048 4416 2952 4423
rect 2988 4416 3153 4423
rect 3167 4416 3312 4423
rect 3336 4423 3343 4433
rect 4096 4423 4103 4436
rect 4436 4436 4493 4443
rect 3336 4416 4103 4423
rect 4436 4423 4443 4436
rect 4787 4436 4853 4443
rect 5016 4443 5023 4456
rect 5047 4456 5112 4463
rect 5148 4453 5152 4467
rect 5188 4456 5313 4463
rect 5327 4456 5393 4463
rect 5487 4456 5543 4463
rect 5016 4436 5493 4443
rect 5536 4443 5543 4456
rect 5567 4456 5853 4463
rect 6047 4453 6053 4467
rect 5536 4436 5592 4443
rect 5628 4436 5713 4443
rect 4127 4416 4443 4423
rect 4587 4416 4733 4423
rect 4847 4416 5073 4423
rect 5287 4416 5313 4423
rect 1856 4396 1903 4403
rect 147 4376 293 4383
rect 307 4376 333 4383
rect 647 4376 913 4383
rect 1407 4376 1593 4383
rect 1647 4376 1873 4383
rect 1896 4383 1903 4396
rect 1941 4396 2173 4403
rect 2347 4396 2493 4403
rect 2727 4396 2873 4403
rect 2967 4396 2992 4403
rect 3028 4396 3133 4403
rect 3307 4396 3453 4403
rect 3707 4396 3852 4403
rect 3888 4396 3953 4403
rect 3976 4396 4033 4403
rect 1896 4376 2172 4383
rect 2208 4376 2353 4383
rect 2747 4376 2813 4383
rect 2867 4376 3192 4383
rect 3228 4376 3393 4383
rect 3976 4383 3983 4396
rect 4187 4396 4253 4403
rect 4307 4396 4373 4403
rect 4507 4396 4573 4403
rect 4707 4396 4872 4403
rect 4908 4396 4933 4403
rect 5096 4396 5573 4403
rect 5096 4387 5103 4396
rect 5727 4396 5752 4403
rect 5788 4396 5873 4403
rect 3947 4376 3983 4383
rect 4007 4376 4093 4383
rect 4167 4376 4423 4383
rect 3047 4356 3093 4363
rect 3747 4356 3773 4363
rect 93 4347 107 4353
rect 873 4347 887 4353
rect 1973 4347 1987 4353
rect 4416 4347 4423 4376
rect 4907 4376 5093 4383
rect 5167 4376 5313 4383
rect 5467 4376 5493 4383
rect 5927 4376 5973 4383
rect 4747 4356 4793 4363
rect 5147 4366 5160 4367
rect 5147 4353 5153 4366
rect 5847 4356 5947 4363
rect 5933 4347 5947 4356
rect 320 4343 333 4347
rect 307 4336 333 4343
rect 320 4333 333 4336
rect 667 4333 673 4347
rect 727 4336 793 4343
rect 1296 4336 1333 4343
rect 1296 4327 1303 4336
rect 1347 4336 1373 4343
rect 1587 4336 1653 4343
rect 1867 4336 1913 4343
rect 2027 4336 2113 4343
rect 2287 4336 2373 4343
rect 2747 4336 2773 4343
rect 2867 4336 2953 4343
rect 3127 4333 3133 4347
rect 3927 4336 3973 4343
rect 4027 4336 4073 4343
rect 4887 4336 4953 4343
rect 5047 4336 5083 4343
rect 1287 4316 1303 4327
rect 1287 4313 1300 4316
rect 3187 4316 3213 4323
rect 5076 4323 5083 4336
rect 5107 4336 5193 4343
rect 5287 4336 5333 4343
rect 5467 4343 5480 4347
rect 5467 4336 5493 4343
rect 5467 4333 5480 4336
rect 5747 4343 5760 4347
rect 5747 4336 5773 4343
rect 5747 4333 5760 4336
rect 6000 4343 6013 4347
rect 5987 4336 6013 4343
rect 6000 4333 6013 4336
rect 5076 4316 5153 4323
rect 193 4307 207 4313
rect 487 4296 553 4303
rect 1247 4293 1253 4307
rect 1567 4293 1573 4307
rect 1767 4293 1773 4307
rect 1847 4296 1873 4303
rect 1887 4296 1913 4303
rect 2187 4293 2193 4307
rect 3847 4296 3913 4303
rect 4727 4293 4733 4307
rect 4967 4293 4973 4307
rect 327 4276 413 4283
rect 427 4276 513 4283
rect 1147 4276 1193 4283
rect 2847 4273 2853 4287
rect 567 4256 613 4263
rect 1027 4256 1053 4263
rect 1147 4256 1313 4263
rect 1787 4256 1913 4263
rect 2253 4263 2267 4273
rect 2167 4256 2267 4263
rect 2976 4263 2983 4293
rect 3207 4276 3273 4283
rect 4287 4273 4293 4287
rect 2927 4256 3033 4263
rect 4596 4263 4603 4293
rect 5653 4287 5667 4293
rect 5307 4273 5313 4287
rect 4476 4256 4603 4263
rect 4476 4247 4483 4256
rect 4627 4256 4833 4263
rect 4947 4256 4973 4263
rect 5247 4256 5273 4263
rect 5407 4256 5443 4263
rect 247 4236 333 4243
rect 767 4236 853 4243
rect 1207 4236 1233 4243
rect 1296 4236 1353 4243
rect 627 4216 893 4223
rect 1296 4223 1303 4236
rect 1527 4236 1713 4243
rect 1787 4236 1853 4243
rect 1976 4236 2093 4243
rect 1976 4227 1983 4236
rect 2767 4233 2773 4247
rect 3027 4236 3213 4243
rect 3367 4236 3393 4243
rect 3767 4236 3873 4243
rect 3927 4236 4133 4243
rect 4227 4236 4253 4243
rect 4367 4236 4393 4243
rect 4476 4243 4493 4247
rect 4447 4236 4493 4243
rect 4480 4233 4493 4236
rect 4687 4236 4973 4243
rect 4987 4233 4993 4247
rect 5276 4243 5283 4253
rect 5147 4236 5223 4243
rect 5276 4236 5393 4243
rect 1187 4216 1303 4223
rect 1327 4216 1973 4223
rect 2167 4216 2333 4223
rect 2387 4216 2493 4223
rect 2747 4216 2972 4223
rect 3008 4216 3053 4223
rect 3067 4216 3113 4223
rect 3247 4216 3303 4223
rect 127 4196 192 4203
rect 228 4196 1613 4203
rect 1747 4196 1933 4203
rect 2187 4196 2613 4203
rect 2687 4196 2732 4203
rect 2768 4193 2773 4207
rect 2947 4196 3273 4203
rect 3296 4203 3303 4216
rect 3827 4216 4573 4223
rect 5216 4223 5223 4236
rect 5436 4243 5443 4256
rect 5436 4236 5473 4243
rect 5607 4236 5733 4243
rect 5807 4236 5873 4243
rect 5887 4236 5913 4243
rect 4967 4216 5203 4223
rect 5216 4216 5493 4223
rect 3296 4196 3513 4203
rect 3807 4196 4313 4203
rect 4327 4196 4673 4203
rect 4807 4196 4933 4203
rect 5087 4196 5133 4203
rect 5196 4203 5203 4216
rect 5196 4196 5633 4203
rect 5700 4203 5713 4207
rect 5696 4193 5713 4203
rect 27 4176 73 4183
rect 147 4176 1033 4183
rect 1087 4176 1793 4183
rect 1927 4176 2153 4183
rect 2247 4176 2313 4183
rect 2367 4180 2443 4183
rect 2367 4176 2447 4180
rect 2433 4167 2447 4176
rect 2467 4176 2923 4183
rect 187 4156 333 4163
rect 707 4156 813 4163
rect 827 4156 1253 4163
rect 1336 4156 1513 4163
rect 47 4136 253 4143
rect 307 4136 673 4143
rect 687 4136 1153 4143
rect 1336 4143 1343 4156
rect 1707 4156 2412 4163
rect 2433 4160 2434 4167
rect 2507 4156 2793 4163
rect 2916 4163 2923 4176
rect 2967 4176 3352 4183
rect 3388 4176 3493 4183
rect 3547 4176 3573 4183
rect 3687 4176 3823 4183
rect 2916 4156 3432 4163
rect 3313 4147 3327 4156
rect 3468 4156 3793 4163
rect 3816 4163 3823 4176
rect 3867 4176 4073 4183
rect 4087 4176 4453 4183
rect 4467 4176 4653 4183
rect 4707 4176 4893 4183
rect 5227 4176 5463 4183
rect 5456 4167 5463 4176
rect 5696 4183 5703 4193
rect 5627 4176 5703 4183
rect 5727 4176 5873 4183
rect 3816 4156 4003 4163
rect 1247 4136 1343 4143
rect 1367 4136 1552 4143
rect 1588 4136 1773 4143
rect 1887 4136 2313 4143
rect 2336 4136 2493 4143
rect 27 4116 333 4123
rect 507 4116 613 4123
rect 867 4116 933 4123
rect 1387 4116 1533 4123
rect 1827 4116 2072 4123
rect 2108 4116 2233 4123
rect 2336 4123 2343 4136
rect 2587 4136 2773 4143
rect 2787 4136 3053 4143
rect 3387 4136 3473 4143
rect 3567 4136 3633 4143
rect 3996 4143 4003 4156
rect 4847 4156 5223 4163
rect 3996 4136 5133 4143
rect 5216 4143 5223 4156
rect 5467 4156 5513 4163
rect 5587 4156 5652 4163
rect 5688 4156 5733 4163
rect 5987 4156 6013 4163
rect 6087 4163 6100 4167
rect 6087 4154 6103 4163
rect 6080 4153 6103 4154
rect 5216 4136 5272 4143
rect 5308 4136 5413 4143
rect 5927 4136 5993 4143
rect 6047 4136 6073 4143
rect 5593 4127 5607 4133
rect 2307 4116 2343 4123
rect 2356 4116 2393 4123
rect -24 4096 213 4103
rect -24 4076 -17 4096
rect 907 4096 993 4103
rect 1247 4096 1413 4103
rect 1516 4096 1613 4103
rect 827 4076 853 4083
rect 973 4076 1013 4083
rect 973 4067 987 4076
rect 1516 4067 1523 4096
rect 1727 4096 2033 4103
rect 2147 4096 2172 4103
rect 2208 4096 2273 4103
rect 2356 4103 2363 4116
rect 2447 4116 2673 4123
rect 3247 4116 3333 4123
rect 3767 4116 3853 4123
rect 3967 4116 4433 4123
rect 4727 4116 4773 4123
rect 5127 4116 5153 4123
rect 5376 4116 5433 4123
rect 2287 4096 2363 4103
rect 2376 4096 2493 4103
rect 2376 4083 2383 4096
rect 2627 4096 2733 4103
rect 3047 4096 3093 4103
rect 3147 4096 3193 4103
rect 3747 4096 3793 4103
rect 4127 4096 4153 4103
rect 4247 4096 4373 4103
rect 4587 4096 5073 4103
rect 5376 4103 5383 4116
rect 5667 4116 5693 4123
rect 6096 4123 6103 4153
rect 6047 4116 6103 4123
rect 5136 4096 5383 4103
rect 5136 4087 5143 4096
rect 5407 4096 5453 4103
rect 5787 4096 5833 4103
rect 5847 4096 5993 4103
rect 2327 4076 2383 4083
rect 4667 4076 4767 4083
rect 4753 4067 4767 4076
rect 5127 4076 5143 4087
rect 5127 4073 5140 4076
rect 5287 4076 5333 4083
rect 347 4056 393 4063
rect 2727 4053 2733 4067
rect 5447 4056 5513 4063
rect 5887 4053 5893 4067
rect -24 4036 13 4043
rect 840 4043 853 4047
rect 827 4036 853 4043
rect 840 4033 853 4036
rect 1967 4033 1973 4047
rect 2887 4033 2893 4047
rect 473 4027 487 4033
rect 5907 4016 5933 4023
rect 5273 4007 5287 4013
rect 427 3996 492 4003
rect 528 4003 540 4007
rect 528 3996 553 4003
rect 528 3993 540 3996
rect 867 3996 953 4003
rect 1647 3996 1713 4003
rect 1787 3996 1873 4003
rect 2027 3996 2073 4003
rect 2320 4003 2333 4007
rect 2307 3996 2333 4003
rect 2320 3993 2333 3996
rect 2487 3996 2553 4003
rect 3167 3993 3173 4007
rect 3607 3996 3673 4003
rect 4227 3996 4293 4003
rect 4507 3996 4613 4003
rect 5067 3996 5133 4003
rect 5387 3993 5393 4007
rect 5560 4003 5573 4007
rect 5547 3996 5573 4003
rect 5560 3993 5573 3996
rect 5687 3996 5772 4003
rect 5808 3993 5813 4007
rect 233 3987 247 3993
rect 1353 3987 1367 3993
rect 127 3956 313 3963
rect 947 3956 973 3963
rect 1496 3963 1503 3993
rect 2253 3987 2267 3993
rect 1347 3956 1503 3963
rect 1667 3956 1793 3963
rect 2416 3963 2423 3993
rect 2047 3956 2423 3963
rect 2716 3963 2723 3993
rect 3833 3987 3847 3993
rect 4013 3987 4027 3993
rect 2507 3956 2723 3963
rect 3067 3956 3113 3963
rect 3307 3956 3353 3963
rect 3707 3956 3913 3963
rect 3927 3956 4053 3963
rect 4176 3963 4183 3993
rect 4067 3956 4183 3963
rect 4456 3963 4463 3993
rect 4773 3987 4787 3993
rect 4913 3987 4927 3993
rect 4327 3956 4463 3963
rect 4667 3956 4713 3963
rect 5047 3956 5083 3963
rect 473 3947 487 3953
rect 347 3936 373 3943
rect 1407 3936 1473 3943
rect 1567 3936 1893 3943
rect 2187 3936 2273 3943
rect 2287 3936 2433 3943
rect 2527 3936 2793 3943
rect 3747 3936 3793 3943
rect 3807 3936 3873 3943
rect 3947 3936 4233 3943
rect 4307 3936 4333 3943
rect 4427 3936 4953 3943
rect 5076 3943 5083 3956
rect 5147 3956 5193 3963
rect 5216 3963 5223 3993
rect 5267 3976 5293 3983
rect 5927 3976 5953 3983
rect 5216 3956 5243 3963
rect 5076 3936 5213 3943
rect 5236 3927 5243 3956
rect 5307 3956 5333 3963
rect 5467 3956 5493 3963
rect 5687 3956 5733 3963
rect 6016 3963 6023 3993
rect 5887 3956 6023 3963
rect 5267 3933 5273 3947
rect 5527 3936 5593 3943
rect 5927 3933 5933 3947
rect 307 3916 353 3923
rect 427 3916 1753 3923
rect 2127 3916 2333 3923
rect 2507 3916 3253 3923
rect 3727 3916 3993 3923
rect 4087 3916 4593 3923
rect 4847 3916 5053 3923
rect 5507 3916 5633 3923
rect 16 3900 73 3903
rect 13 3896 73 3900
rect 13 3887 27 3896
rect 287 3896 583 3903
rect 26 3880 27 3887
rect 48 3876 133 3883
rect 507 3876 553 3883
rect 576 3883 583 3896
rect 647 3896 673 3903
rect 687 3896 753 3903
rect 827 3896 933 3903
rect 947 3896 1033 3903
rect 1107 3896 1353 3903
rect 1547 3896 1813 3903
rect 2156 3896 2463 3903
rect 576 3876 613 3883
rect 636 3876 953 3883
rect 107 3856 393 3863
rect 447 3856 593 3863
rect 636 3863 643 3876
rect 967 3876 993 3883
rect 1007 3876 1173 3883
rect 1187 3876 1473 3883
rect 1667 3876 1713 3883
rect 2156 3883 2163 3896
rect 1727 3876 2163 3883
rect 2456 3887 2463 3896
rect 2607 3896 2713 3903
rect 2727 3896 2913 3903
rect 3227 3896 3593 3903
rect 3647 3896 4003 3903
rect 2187 3876 2313 3883
rect 2327 3876 2373 3883
rect 2467 3876 2753 3883
rect 3327 3876 3433 3883
rect 3547 3876 3713 3883
rect 3996 3883 4003 3896
rect 4027 3896 4793 3903
rect 5487 3896 5993 3903
rect 4796 3887 4803 3893
rect 3996 3876 4053 3883
rect 4167 3873 4173 3887
rect 4267 3876 4453 3883
rect 4627 3876 4783 3883
rect 4796 3876 4812 3887
rect 4776 3867 4783 3876
rect 4800 3873 4812 3876
rect 4848 3876 5253 3883
rect 5467 3876 5713 3883
rect 607 3856 643 3863
rect 1067 3856 1153 3863
rect 1167 3856 1493 3863
rect 1887 3856 2032 3863
rect 2068 3856 2113 3863
rect 2127 3856 2173 3863
rect 2347 3856 2473 3863
rect 2547 3856 2633 3863
rect 2867 3856 3073 3863
rect 3247 3856 3373 3863
rect 3707 3856 3753 3863
rect 3847 3856 3873 3863
rect 4147 3856 4213 3863
rect 4227 3856 4273 3863
rect 4367 3856 4752 3863
rect 4788 3856 4913 3863
rect 5167 3856 5192 3863
rect 5228 3856 5503 3863
rect 27 3833 33 3847
rect 4167 3833 4173 3847
rect 4827 3833 4833 3847
rect 4847 3833 4853 3847
rect 5367 3836 5467 3843
rect 1693 3827 1707 3833
rect 5453 3827 5467 3836
rect 5496 3827 5503 3856
rect 5756 3856 5953 3863
rect 5756 3827 5763 3856
rect 327 3816 413 3823
rect 467 3816 553 3823
rect 667 3813 673 3827
rect 727 3816 792 3823
rect 828 3813 833 3827
rect 987 3813 993 3827
rect 1347 3823 1360 3827
rect 1347 3816 1373 3823
rect 1347 3813 1360 3816
rect 1507 3823 1520 3827
rect 1507 3816 1533 3823
rect 1507 3813 1520 3816
rect 1767 3816 1833 3823
rect 1987 3813 1993 3827
rect 2247 3823 2260 3827
rect 2247 3816 2273 3823
rect 2247 3813 2260 3816
rect 2387 3816 2433 3823
rect 2627 3816 2673 3823
rect 2747 3816 2853 3823
rect 3067 3816 3112 3823
rect 3148 3816 3193 3823
rect 3287 3823 3300 3827
rect 3287 3816 3313 3823
rect 3287 3813 3300 3816
rect 3367 3816 3412 3823
rect 3448 3816 3493 3823
rect 3607 3816 3653 3823
rect 3887 3816 3933 3823
rect 3987 3816 4073 3823
rect 4187 3816 4253 3823
rect 4547 3813 4553 3827
rect 4667 3816 4713 3823
rect 4927 3813 4933 3827
rect 5207 3816 5293 3823
rect 5927 3816 5993 3823
rect -24 3776 13 3783
rect 4007 3776 4093 3783
rect 6047 3776 6123 3783
rect 747 3753 752 3767
rect 788 3756 853 3763
rect 967 3753 973 3767
rect 1027 3756 1093 3763
rect 1267 3756 1353 3763
rect 1487 3756 1553 3763
rect 1947 3756 2013 3763
rect 3127 3756 3173 3763
rect 3387 3756 3453 3763
rect 3727 3756 3773 3763
rect 3840 3763 3853 3767
rect 3827 3756 3853 3763
rect 3840 3753 3853 3756
rect 127 3716 213 3723
rect 267 3716 313 3723
rect 447 3716 493 3723
rect 696 3723 703 3753
rect 1013 3747 1027 3753
rect 507 3716 743 3723
rect 367 3696 533 3703
rect 547 3696 713 3703
rect 736 3703 743 3716
rect 767 3716 893 3723
rect 1147 3716 1293 3723
rect 1867 3716 2053 3723
rect 2156 3723 2163 3753
rect 3213 3743 3227 3753
rect 3213 3736 3313 3743
rect 3867 3733 3873 3747
rect 5036 3743 5043 3773
rect 5087 3756 5113 3763
rect 5127 3756 5173 3763
rect 5036 3736 5093 3743
rect 2067 3716 2273 3723
rect 2387 3716 2493 3723
rect 2507 3716 2533 3723
rect 2767 3716 2853 3723
rect 2867 3716 2913 3723
rect 3107 3716 3473 3723
rect 3527 3716 3753 3723
rect 3767 3716 3913 3723
rect 3927 3716 3993 3723
rect 4247 3716 4313 3723
rect 4747 3716 4813 3723
rect 4827 3716 4853 3723
rect 5616 3723 5623 3753
rect 5616 3716 5733 3723
rect 5896 3723 5903 3753
rect 5787 3716 5903 3723
rect 736 3696 772 3703
rect 808 3696 873 3703
rect 887 3696 1073 3703
rect 1207 3696 1273 3703
rect 1347 3696 1433 3703
rect 1607 3696 2193 3703
rect 2687 3696 3633 3703
rect 3807 3696 3933 3703
rect 3947 3696 4493 3703
rect 4627 3696 4713 3703
rect 4727 3696 4813 3703
rect 5247 3696 5633 3703
rect 5647 3696 5753 3703
rect 5767 3696 5833 3703
rect 487 3676 573 3683
rect 627 3676 753 3683
rect 807 3673 813 3687
rect 867 3676 973 3683
rect 1107 3676 1673 3683
rect 2247 3676 2293 3683
rect 2347 3676 2373 3683
rect 2387 3676 2453 3683
rect 2767 3676 2793 3683
rect 2807 3676 3092 3683
rect 3113 3673 3114 3680
rect 3367 3676 3413 3683
rect 3787 3676 3832 3683
rect 3868 3676 3953 3683
rect 4247 3676 4353 3683
rect 5047 3676 5213 3683
rect 5327 3676 5473 3683
rect 27 3656 543 3663
rect 227 3636 513 3643
rect 536 3643 543 3656
rect 907 3656 933 3663
rect 947 3656 1043 3663
rect 536 3636 1013 3643
rect 1036 3643 1043 3656
rect 1087 3656 1593 3663
rect 1887 3656 2153 3663
rect 2167 3656 2253 3663
rect 3113 3663 3127 3673
rect 3087 3660 3127 3663
rect 3087 3656 3123 3660
rect 3567 3656 3673 3663
rect 3687 3656 3853 3663
rect 4067 3656 4393 3663
rect 4967 3656 5913 3663
rect 1036 3636 1113 3643
rect 2276 3636 2713 3643
rect 27 3616 1273 3623
rect 2276 3623 2283 3636
rect 2807 3636 2953 3643
rect 3107 3636 3133 3643
rect 3147 3636 3193 3643
rect 3327 3636 3453 3643
rect 5167 3636 5233 3643
rect 5407 3636 5433 3643
rect 1287 3616 2283 3623
rect 2387 3616 2753 3623
rect 2916 3616 3053 3623
rect 187 3596 293 3603
rect 427 3596 693 3603
rect 707 3596 813 3603
rect 1467 3596 1793 3603
rect 1835 3600 2113 3603
rect 1833 3596 2113 3600
rect 1833 3587 1847 3596
rect 2207 3596 2593 3603
rect 2916 3603 2923 3616
rect 3147 3616 3233 3623
rect 3247 3616 3353 3623
rect 3367 3616 3593 3623
rect 3747 3616 3853 3623
rect 3867 3616 4063 3623
rect 4056 3607 4063 3616
rect 4287 3616 4433 3623
rect 4447 3616 4533 3623
rect 4847 3616 5053 3623
rect 5067 3616 5193 3623
rect 5367 3613 5373 3627
rect 2667 3596 2923 3603
rect 2967 3596 3093 3603
rect 3167 3596 3273 3603
rect 3287 3596 3393 3603
rect 3407 3596 3873 3603
rect 4067 3596 4173 3603
rect 4527 3596 4733 3603
rect 5167 3596 5443 3603
rect 247 3576 273 3583
rect 327 3576 473 3583
rect 487 3576 573 3583
rect 1347 3576 1393 3583
rect 1547 3576 1593 3583
rect 1707 3576 1753 3583
rect 1846 3580 1847 3587
rect 1868 3576 2133 3583
rect 2147 3576 2333 3583
rect 2847 3576 2993 3583
rect 3007 3576 3113 3583
rect 3127 3576 3593 3583
rect 3787 3576 3893 3583
rect 3907 3576 4553 3583
rect 4567 3576 4693 3583
rect 4707 3576 4943 3583
rect 4936 3567 4943 3576
rect 5436 3587 5443 3596
rect 5587 3596 5633 3603
rect 5887 3596 5913 3603
rect 4987 3576 5193 3583
rect 5207 3576 5313 3583
rect 5367 3576 5393 3583
rect 5447 3576 5533 3583
rect 5607 3576 5793 3583
rect 5807 3576 5873 3583
rect 6007 3576 6073 3583
rect 5953 3567 5967 3573
rect 193 3547 207 3553
rect 1147 3556 1207 3563
rect 693 3547 707 3553
rect 1193 3547 1207 3556
rect 2476 3556 2553 3563
rect -24 3536 13 3543
rect 147 3536 193 3543
rect 287 3536 373 3543
rect 1287 3536 1353 3543
rect 2476 3527 2483 3556
rect 3647 3556 3693 3563
rect 4947 3556 4973 3563
rect 3247 3543 3260 3547
rect 3247 3536 3273 3543
rect 3247 3533 3260 3536
rect 4067 3536 4153 3543
rect 4407 3536 4473 3543
rect 4860 3543 4873 3547
rect 4847 3536 4873 3543
rect 4860 3533 4873 3536
rect 5307 3536 5353 3543
rect 5587 3536 5673 3543
rect 5947 3536 6013 3543
rect 847 3513 853 3527
rect 2647 3513 2653 3527
rect 4300 3523 4313 3527
rect 4296 3513 4313 3523
rect 4296 3503 4303 3513
rect 4267 3496 4303 3503
rect 267 3476 333 3483
rect 407 3476 453 3483
rect 587 3476 633 3483
rect 1267 3476 1373 3483
rect 1607 3476 1633 3483
rect 1767 3476 1813 3483
rect 2327 3476 2413 3483
rect 2747 3483 2760 3487
rect 2747 3476 2773 3483
rect 2747 3473 2760 3476
rect 2887 3476 2933 3483
rect 3467 3476 3553 3483
rect 3687 3476 3733 3483
rect 3947 3476 3993 3483
rect 4087 3476 4173 3483
rect 4327 3473 4333 3487
rect 4487 3473 4493 3487
rect 4687 3476 4723 3483
rect 127 3436 573 3443
rect 676 3443 683 3473
rect 1213 3467 1227 3473
rect 867 3456 893 3463
rect 1673 3467 1687 3473
rect 676 3436 873 3443
rect 967 3436 1013 3443
rect 1107 3436 1953 3443
rect 1976 3443 1983 3473
rect 2173 3467 2187 3473
rect 1976 3436 2253 3443
rect 3096 3443 3103 3473
rect 3253 3467 3267 3473
rect 2967 3436 3313 3443
rect 3367 3436 3413 3443
rect 3596 3443 3603 3473
rect 4267 3453 4273 3467
rect 4407 3456 4433 3463
rect 4716 3463 4723 3476
rect 4747 3476 4813 3483
rect 5056 3476 5133 3483
rect 4716 3456 4753 3463
rect 5056 3463 5063 3476
rect 5467 3476 5553 3483
rect 5787 3476 5853 3483
rect 5027 3456 5063 3463
rect 5693 3467 5707 3473
rect 5893 3467 5907 3473
rect 3596 3436 3953 3443
rect 4007 3436 4533 3443
rect 4547 3436 4933 3443
rect 5427 3436 5513 3443
rect 5627 3436 5653 3443
rect 5953 3427 5967 3433
rect 287 3413 293 3427
rect 1127 3416 1173 3423
rect 1187 3416 1453 3423
rect 1807 3416 2043 3423
rect 347 3396 1593 3403
rect 1636 3396 1993 3403
rect 547 3376 733 3383
rect 867 3376 1213 3383
rect 1636 3383 1643 3396
rect 2036 3403 2043 3416
rect 2067 3416 2173 3423
rect 2187 3416 2392 3423
rect 2428 3416 2793 3423
rect 2807 3416 3032 3423
rect 3068 3416 4433 3423
rect 4807 3416 4833 3423
rect 5107 3416 5213 3423
rect 5367 3413 5373 3427
rect 5887 3416 5953 3423
rect 2036 3396 2113 3403
rect 2127 3396 2373 3403
rect 2527 3396 2873 3403
rect 2987 3396 3353 3403
rect 3707 3396 4073 3403
rect 5187 3396 5413 3403
rect 1347 3376 1643 3383
rect 1687 3376 2293 3383
rect 2507 3376 3133 3383
rect 3147 3376 3373 3383
rect 3567 3376 3633 3383
rect 4947 3376 4993 3383
rect 5087 3376 5253 3383
rect 6047 3376 6073 3383
rect 287 3356 353 3363
rect 647 3356 693 3363
rect 847 3356 873 3363
rect 2607 3356 2633 3363
rect 2887 3356 3073 3363
rect 3207 3356 3233 3363
rect 3587 3356 3813 3363
rect 4067 3356 4313 3363
rect 4367 3356 4393 3363
rect 4847 3356 5143 3363
rect 5136 3347 5143 3356
rect 5487 3353 5493 3367
rect 5627 3356 5893 3363
rect 6007 3356 6033 3363
rect 67 3336 133 3343
rect 147 3336 253 3343
rect 367 3336 393 3343
rect 747 3336 853 3343
rect 1387 3336 1433 3343
rect 2347 3336 2393 3343
rect 2847 3336 3253 3343
rect 3267 3336 3493 3343
rect 3507 3336 3773 3343
rect 3967 3336 4173 3343
rect 5067 3336 5093 3343
rect 5147 3336 5553 3343
rect 5707 3336 5853 3343
rect 5867 3336 5973 3343
rect 733 3327 747 3333
rect 4827 3316 4853 3323
rect 87 3293 93 3307
rect 567 3296 633 3303
rect 887 3296 973 3303
rect 1647 3296 1693 3303
rect 1896 3296 1933 3303
rect 2447 3296 2513 3303
rect 2647 3296 2693 3303
rect 2920 3303 2933 3307
rect 2747 3296 2853 3303
rect 2907 3296 2933 3303
rect 2920 3293 2933 3296
rect 3187 3296 3232 3303
rect 3268 3303 3280 3307
rect 3268 3296 3293 3303
rect 3268 3293 3280 3296
rect 3387 3296 3453 3303
rect 3767 3296 3873 3303
rect 3927 3296 3973 3303
rect 4067 3296 4113 3303
rect 4207 3296 4273 3303
rect 4407 3296 4473 3303
rect 4627 3296 4672 3303
rect 4708 3296 4753 3303
rect 4987 3296 5053 3303
rect 5247 3296 5313 3303
rect 5487 3303 5500 3307
rect 5487 3296 5513 3303
rect 5487 3293 5500 3296
rect 5567 3296 5653 3303
rect 5707 3296 5752 3303
rect 5788 3303 5800 3307
rect 5788 3296 5813 3303
rect 5788 3293 5800 3296
rect 5907 3296 5973 3303
rect 767 3253 773 3267
rect 1027 3256 1073 3263
rect 1160 3263 1173 3267
rect 1147 3256 1173 3263
rect 1160 3253 1173 3256
rect 2167 3256 2233 3263
rect 2600 3263 2613 3267
rect 2587 3256 2613 3263
rect 2600 3253 2613 3256
rect 4287 3256 4333 3263
rect 4867 3256 4913 3263
rect 5407 3256 5493 3263
rect 713 3247 727 3253
rect 2053 3247 2067 3253
rect 587 3236 643 3243
rect 413 3227 427 3233
rect 536 3203 543 3233
rect 636 3223 643 3236
rect 3040 3243 3053 3247
rect 3027 3236 3053 3243
rect 3040 3233 3053 3236
rect 3407 3236 3433 3243
rect 3567 3236 3613 3243
rect 3627 3236 3693 3243
rect 3827 3236 3893 3243
rect 636 3216 673 3223
rect 307 3196 633 3203
rect 787 3196 813 3203
rect 1396 3203 1403 3233
rect 4907 3216 4973 3223
rect 1247 3196 1403 3203
rect 1767 3196 1813 3203
rect 1887 3196 1913 3203
rect 2307 3196 2413 3203
rect 2727 3196 2793 3203
rect 2807 3196 2833 3203
rect 2887 3196 3033 3203
rect 3087 3196 3113 3203
rect 3247 3196 3473 3203
rect 3647 3196 3733 3203
rect 4127 3196 4213 3203
rect 4227 3196 4373 3203
rect 4387 3196 4553 3203
rect 4647 3196 4693 3203
rect 4787 3196 5073 3203
rect 5427 3196 5573 3203
rect 5587 3196 5713 3203
rect 5767 3196 5833 3203
rect 127 3176 273 3183
rect 287 3176 413 3183
rect 647 3176 953 3183
rect 2267 3176 2373 3183
rect 2387 3176 2693 3183
rect 2876 3183 2883 3193
rect 2767 3176 2883 3183
rect 3067 3176 3152 3183
rect 3188 3176 3253 3183
rect 4607 3176 4893 3183
rect 5547 3176 5613 3183
rect 347 3153 353 3167
rect 727 3156 1393 3163
rect 1407 3156 1873 3163
rect 1927 3156 2073 3163
rect 2747 3156 2853 3163
rect 4507 3156 4633 3163
rect 5487 3156 5573 3163
rect 47 3136 153 3143
rect 167 3136 233 3143
rect 247 3136 673 3143
rect 1287 3136 1653 3143
rect 1947 3136 2153 3143
rect 2167 3136 2473 3143
rect 2707 3136 2813 3143
rect 2827 3136 3093 3143
rect 4187 3136 4353 3143
rect 5227 3136 5393 3143
rect 1247 3116 2413 3123
rect 2476 3123 2483 3133
rect 2476 3116 2953 3123
rect 4247 3116 4273 3123
rect 5447 3116 5513 3123
rect 1087 3096 1293 3103
rect 1567 3096 1813 3103
rect 1887 3096 2333 3103
rect 2347 3096 2913 3103
rect 3147 3096 3213 3103
rect 3967 3096 4273 3103
rect 4287 3096 4693 3103
rect 5267 3096 5353 3103
rect 5407 3096 5453 3103
rect 5507 3096 5653 3103
rect 5667 3096 5833 3103
rect 1027 3076 1153 3083
rect 1387 3076 1433 3083
rect 1627 3076 1733 3083
rect 1747 3076 2133 3083
rect 2407 3076 2433 3083
rect 2527 3076 2573 3083
rect 2627 3076 2793 3083
rect 2807 3076 2873 3083
rect 3067 3076 3493 3083
rect 3687 3076 3813 3083
rect 3827 3076 4153 3083
rect 4447 3076 4633 3083
rect 4647 3076 4853 3083
rect 5027 3076 5473 3083
rect 5647 3076 5733 3083
rect 127 3056 183 3063
rect 176 3043 183 3056
rect 227 3056 793 3063
rect 807 3056 2673 3063
rect 2687 3056 2753 3063
rect 2947 3056 3133 3063
rect 3187 3056 3393 3063
rect 3867 3056 3933 3063
rect 3947 3056 4893 3063
rect 4907 3056 4973 3063
rect 4987 3056 5693 3063
rect 5707 3056 5773 3063
rect 5947 3056 6013 3063
rect 176 3036 213 3043
rect 1827 3036 1983 3043
rect 1976 3027 1983 3036
rect 5207 3043 5220 3047
rect 5207 3033 5223 3043
rect 1007 3016 1073 3023
rect 1987 3016 2013 3023
rect 2107 3016 2153 3023
rect 2447 3016 2513 3023
rect 2527 3016 2593 3023
rect 3267 3016 3313 3023
rect 4067 3016 4133 3023
rect 4727 3013 4733 3027
rect 5216 3023 5223 3033
rect 5320 3023 5333 3027
rect 5216 3016 5293 3023
rect 5307 3016 5333 3023
rect 5320 3013 5333 3016
rect 5527 3016 5573 3023
rect 5727 3016 5773 3023
rect 1527 2996 1593 3003
rect 1827 2996 1913 3003
rect 5227 2996 5253 3003
rect 5347 2996 5393 3003
rect 5887 2996 5933 3003
rect 227 2956 273 2963
rect 327 2956 433 2963
rect 587 2956 673 2963
rect 2147 2963 2160 2967
rect 2147 2956 2173 2963
rect 2147 2953 2160 2956
rect 2267 2956 2373 2963
rect 2667 2953 2673 2967
rect 2987 2956 3053 2963
rect 3127 2956 3172 2963
rect 3208 2963 3220 2967
rect 3208 2956 3233 2963
rect 3208 2953 3220 2956
rect 3327 2956 3373 2963
rect 3387 2956 3473 2963
rect 3567 2956 3653 2963
rect 3747 2956 3793 2963
rect 4167 2956 4253 2963
rect 4467 2956 4513 2963
rect 4607 2953 4613 2967
rect 4787 2956 4833 2963
rect 5127 2963 5140 2967
rect 5127 2956 5153 2963
rect 5127 2953 5140 2956
rect 5327 2956 5413 2963
rect 5967 2963 5980 2967
rect 5967 2956 5993 2963
rect 5967 2953 5980 2956
rect 1273 2947 1287 2953
rect 920 2943 933 2947
rect 796 2936 853 2943
rect 907 2936 933 2943
rect 127 2916 173 2923
rect 267 2916 463 2923
rect 456 2907 463 2916
rect 547 2916 713 2923
rect 796 2923 803 2936
rect 920 2933 933 2936
rect 767 2916 803 2923
rect 1107 2916 1333 2923
rect 1347 2916 1473 2923
rect 1756 2923 1763 2953
rect 2073 2947 2087 2953
rect 2773 2947 2787 2953
rect 1567 2916 1763 2923
rect 2127 2916 2213 2923
rect 2587 2916 2852 2923
rect 2888 2916 2933 2923
rect 3696 2923 3703 2953
rect 3487 2916 3703 2923
rect 3836 2923 3843 2953
rect 3993 2947 4007 2953
rect 3767 2916 3843 2923
rect 3867 2916 4113 2923
rect 4996 2923 5003 2953
rect 4127 2916 5003 2923
rect 5346 2913 5347 2920
rect 5407 2916 5553 2923
rect 5696 2923 5703 2953
rect 5567 2916 5953 2923
rect 167 2896 453 2903
rect 467 2896 593 2903
rect 607 2896 733 2903
rect 1096 2903 1103 2913
rect 747 2896 1103 2903
rect 1247 2896 1313 2903
rect 5333 2907 5347 2913
rect 1607 2896 1713 2903
rect 1767 2896 2253 2903
rect 2427 2896 2613 2903
rect 3667 2896 4033 2903
rect 4247 2896 4293 2903
rect 4367 2896 4413 2903
rect 4587 2896 4863 2903
rect 1327 2876 1553 2883
rect 1647 2876 2233 2883
rect 4207 2876 4313 2883
rect 4387 2876 4553 2883
rect 4856 2883 4863 2896
rect 4887 2896 5013 2903
rect 5346 2900 5347 2907
rect 5353 2893 5354 2900
rect 5967 2893 5973 2907
rect 4856 2876 5133 2883
rect 5147 2876 5223 2883
rect 67 2856 273 2863
rect 427 2856 573 2863
rect 927 2856 953 2863
rect 1087 2856 1133 2863
rect 1447 2856 1493 2863
rect 1687 2856 1833 2863
rect 2867 2856 3253 2863
rect 3787 2856 4033 2863
rect 4047 2856 4853 2863
rect 4867 2856 5153 2863
rect 5216 2863 5223 2876
rect 5353 2883 5367 2893
rect 5327 2880 5367 2883
rect 5327 2876 5363 2880
rect 5216 2856 5733 2863
rect 1747 2836 1883 2843
rect 307 2816 373 2823
rect 747 2816 773 2823
rect 913 2807 927 2813
rect 1876 2807 1883 2836
rect 2027 2836 2653 2843
rect 2727 2836 3193 2843
rect 3207 2836 3233 2843
rect 3547 2836 4513 2843
rect 4527 2836 4653 2843
rect 4707 2836 4773 2843
rect 5227 2836 5633 2843
rect 5847 2836 5893 2843
rect 5907 2836 5933 2843
rect 2033 2807 2047 2813
rect 2167 2816 2373 2823
rect 2387 2816 2513 2823
rect 3087 2816 3423 2823
rect 2073 2807 2087 2813
rect 827 2796 873 2803
rect 1787 2796 1833 2803
rect 1967 2803 1980 2807
rect 1967 2796 1993 2803
rect 1967 2793 1980 2796
rect 3416 2787 3423 2816
rect 3447 2816 4003 2823
rect 3996 2807 4003 2816
rect 4267 2816 4393 2823
rect 3947 2796 3993 2803
rect 4733 2787 4747 2793
rect 687 2776 773 2783
rect 1667 2776 1713 2783
rect 2307 2776 2413 2783
rect 2487 2776 2533 2783
rect 2847 2776 2893 2783
rect 3287 2776 3373 2783
rect 3527 2776 3573 2783
rect 3667 2776 3753 2783
rect 3807 2776 3873 2783
rect 4180 2783 4193 2787
rect 4167 2776 4193 2783
rect 4180 2773 4193 2776
rect 4287 2776 4333 2783
rect 4827 2776 4873 2783
rect 5387 2776 5433 2783
rect -24 2703 -17 2743
rect 527 2733 533 2747
rect 1947 2736 2013 2743
rect 2027 2736 2073 2743
rect 2287 2736 2353 2743
rect 2707 2736 2773 2743
rect 3020 2743 3033 2747
rect 3007 2736 3033 2743
rect 3020 2733 3033 2736
rect 4687 2736 4733 2743
rect 5120 2743 5132 2747
rect 5107 2736 5132 2743
rect 5120 2733 5132 2736
rect 5168 2736 5233 2743
rect 5447 2736 5513 2743
rect 5567 2736 5653 2743
rect 5907 2736 5953 2743
rect 93 2727 107 2733
rect 893 2727 907 2733
rect -24 2696 33 2703
rect 1387 2696 1433 2703
rect 1856 2703 1863 2733
rect 2107 2723 2120 2727
rect 2107 2716 2133 2723
rect 2107 2713 2120 2716
rect 1856 2696 1993 2703
rect 3116 2703 3123 2733
rect 3987 2723 4000 2727
rect 3987 2716 4013 2723
rect 4147 2716 4213 2723
rect 3987 2713 4000 2716
rect 4427 2716 4493 2723
rect 4967 2716 5053 2723
rect 3007 2696 3123 2703
rect 307 2676 333 2683
rect 1667 2676 2473 2683
rect 2996 2683 3003 2693
rect 2867 2676 3393 2683
rect 3407 2676 3473 2683
rect 3487 2676 3633 2683
rect 3647 2676 3733 2683
rect 3747 2676 3893 2683
rect 4536 2683 4543 2713
rect 4747 2696 4773 2703
rect 5796 2703 5803 2733
rect 5647 2696 5803 2703
rect 5867 2696 5973 2703
rect 4536 2676 4693 2683
rect 4867 2676 4893 2683
rect 5267 2676 5513 2683
rect 5527 2676 5893 2683
rect 1647 2656 1773 2663
rect 2247 2656 3153 2663
rect 3387 2656 4153 2663
rect 4167 2656 4653 2663
rect 4667 2656 4833 2663
rect 4987 2656 5293 2663
rect 407 2636 593 2643
rect 1027 2636 1653 2643
rect 2087 2636 2153 2643
rect 2227 2636 2753 2643
rect 2767 2636 2953 2643
rect 3607 2636 3793 2643
rect 3867 2636 3973 2643
rect 3996 2636 4593 2643
rect 1087 2616 1313 2623
rect 1667 2616 1733 2623
rect 2567 2616 2693 2623
rect 3127 2616 3153 2623
rect 3996 2623 4003 2636
rect 4867 2633 4873 2647
rect 5407 2636 5433 2643
rect 3167 2616 4003 2623
rect 4907 2616 5433 2623
rect 1136 2596 1433 2603
rect 1136 2587 1143 2596
rect 1847 2596 2273 2603
rect 2667 2596 2753 2603
rect 2767 2596 3033 2603
rect 5367 2596 5573 2603
rect 287 2576 453 2583
rect 467 2576 1133 2583
rect 1207 2576 1233 2583
rect 1547 2576 2893 2583
rect 3187 2576 3473 2583
rect 5527 2576 5633 2583
rect 4307 2556 4353 2563
rect 4367 2556 4573 2563
rect 727 2536 873 2543
rect 1287 2536 1353 2543
rect 1847 2536 1873 2543
rect 2127 2536 2353 2543
rect 3047 2536 3073 2543
rect 4347 2536 4393 2543
rect 4747 2536 4813 2543
rect 5147 2536 5253 2543
rect 5307 2536 5433 2543
rect 1507 2516 1533 2523
rect 1547 2516 1653 2523
rect 3467 2516 3653 2523
rect 4247 2516 4273 2523
rect 4507 2516 4613 2523
rect 5007 2516 5053 2523
rect 5147 2516 5263 2523
rect 1227 2493 1233 2507
rect 1967 2496 2013 2503
rect 2067 2496 2113 2503
rect 4587 2496 4653 2503
rect 333 2487 347 2493
rect 5256 2487 5263 2516
rect 147 2473 153 2487
rect 807 2476 873 2483
rect 887 2476 933 2483
rect 1060 2483 1073 2487
rect 1047 2476 1073 2483
rect 1060 2473 1073 2476
rect 1607 2476 1713 2483
rect 1767 2476 1833 2483
rect 2487 2476 2573 2483
rect 3487 2476 3553 2483
rect 4447 2476 4533 2483
rect 5487 2476 5553 2483
rect 1807 2456 1853 2463
rect 1233 2447 1247 2453
rect 1167 2436 1212 2443
rect 1233 2440 1234 2447
rect 1320 2443 1333 2447
rect 1307 2436 1333 2443
rect 1320 2433 1333 2436
rect 1387 2436 1453 2443
rect 2047 2436 2113 2443
rect 2547 2436 2593 2443
rect 3207 2433 3213 2447
rect 3727 2436 3813 2443
rect 4727 2433 4733 2447
rect 4900 2443 4913 2447
rect 4887 2436 4913 2443
rect 4900 2433 4913 2436
rect 5427 2436 5533 2443
rect 5607 2436 5653 2443
rect 5747 2433 5753 2447
rect 693 2427 707 2433
rect 1640 2423 1653 2427
rect 1536 2416 1573 2423
rect 1627 2416 1653 2423
rect 747 2396 793 2403
rect 947 2396 993 2403
rect 1007 2396 1113 2403
rect 1536 2403 1543 2416
rect 1640 2413 1653 2416
rect 1507 2396 1543 2403
rect 1896 2403 1903 2433
rect 2173 2427 2187 2433
rect 2333 2427 2347 2433
rect 3013 2427 3027 2433
rect 2447 2413 2453 2427
rect 3487 2416 3533 2423
rect 1827 2396 2313 2403
rect 3187 2396 3233 2403
rect 3827 2396 3853 2403
rect 4376 2403 4383 2433
rect 4287 2396 4383 2403
rect 4627 2396 4673 2403
rect 5327 2396 5473 2403
rect 5547 2396 5592 2403
rect 5628 2396 5713 2403
rect 767 2376 973 2383
rect 987 2376 1183 2383
rect 1176 2367 1183 2376
rect 1307 2376 1353 2383
rect 1547 2373 1553 2387
rect 1787 2376 1953 2383
rect 4447 2376 4633 2383
rect 4647 2376 4773 2383
rect 5507 2373 5513 2387
rect 187 2356 213 2363
rect 227 2356 273 2363
rect 467 2356 593 2363
rect 1187 2356 1373 2363
rect 1487 2356 1633 2363
rect 1987 2356 2233 2363
rect 2387 2356 2493 2363
rect 2507 2356 2753 2363
rect 2847 2356 3173 2363
rect 3227 2356 3313 2363
rect 3387 2356 3513 2363
rect 3847 2356 4013 2363
rect 4027 2356 4253 2363
rect 4927 2356 5713 2363
rect 1327 2336 1393 2343
rect 1447 2336 1813 2343
rect 2607 2336 2873 2343
rect 2887 2336 2953 2343
rect 3087 2336 3133 2343
rect 5553 2347 5567 2356
rect 5787 2356 5813 2363
rect 3267 2336 3353 2343
rect 3416 2336 3573 2343
rect 3416 2327 3423 2336
rect 3927 2336 3973 2343
rect 4587 2336 5233 2343
rect 456 2316 573 2323
rect 456 2287 463 2316
rect 1467 2316 1593 2323
rect 2287 2316 2313 2323
rect 2767 2316 2913 2323
rect 3267 2316 3413 2323
rect 4067 2316 4093 2323
rect 4227 2316 4313 2323
rect 5767 2316 5813 2323
rect 593 2287 607 2293
rect 716 2296 753 2303
rect 507 2276 553 2283
rect 716 2283 723 2296
rect 1407 2296 1633 2303
rect 1767 2296 1973 2303
rect 2127 2296 2193 2303
rect 2207 2296 2243 2303
rect 647 2276 723 2283
rect 987 2276 1073 2283
rect 2236 2267 2243 2296
rect 2847 2296 2893 2303
rect 4527 2296 4573 2303
rect 5087 2296 5193 2303
rect 5376 2296 5413 2303
rect 2287 2276 2333 2283
rect 2707 2273 2713 2287
rect 3987 2283 4000 2287
rect 3987 2276 4013 2283
rect 3987 2273 4000 2276
rect 4267 2273 4273 2287
rect 5376 2283 5383 2296
rect 5747 2296 5873 2303
rect 5927 2296 5953 2303
rect 5347 2276 5383 2283
rect 5853 2267 5867 2273
rect 47 2263 60 2267
rect 47 2256 73 2263
rect 47 2253 60 2256
rect 1427 2256 1473 2263
rect 1827 2256 1913 2263
rect 2827 2263 2840 2267
rect 2827 2256 2853 2263
rect 2827 2253 2840 2256
rect 3307 2256 3373 2263
rect 4107 2256 4153 2263
rect 4487 2256 4553 2263
rect 5127 2263 5140 2267
rect 5127 2256 5153 2263
rect 5167 2256 5253 2263
rect 5127 2253 5140 2256
rect 5587 2256 5633 2263
rect 5947 2256 5993 2263
rect 6007 2253 6013 2267
rect 5207 2236 5273 2243
rect 500 2223 513 2227
rect 387 2216 473 2223
rect 487 2216 513 2223
rect 500 2213 513 2216
rect 587 2223 600 2227
rect 587 2216 613 2223
rect 587 2213 600 2216
rect 1267 2216 1313 2223
rect 1807 2213 1813 2227
rect 2067 2213 2073 2227
rect 2127 2216 2193 2223
rect 2367 2213 2373 2227
rect 2747 2216 2813 2223
rect 3327 2216 3433 2223
rect 3807 2213 3813 2227
rect 4287 2213 4293 2227
rect 4807 2213 4813 2227
rect 4947 2216 4993 2223
rect 5340 2223 5353 2227
rect 5327 2216 5353 2223
rect 5340 2213 5353 2216
rect 4033 2207 4047 2213
rect 4613 2207 4627 2213
rect 107 2193 113 2207
rect 347 2193 353 2207
rect 1507 2196 1583 2203
rect 213 2187 227 2193
rect 1576 2187 1583 2196
rect 1707 2196 1753 2203
rect 3187 2196 3233 2203
rect 4200 2203 4213 2207
rect 4187 2196 4213 2203
rect 4200 2193 4213 2196
rect 4467 2196 4513 2203
rect 5187 2193 5193 2207
rect 5707 2196 5793 2203
rect 5927 2196 5993 2203
rect 1576 2176 1593 2187
rect 1580 2173 1593 2176
rect 3387 2176 3473 2183
rect 3567 2176 3613 2183
rect 567 2156 733 2163
rect 1487 2156 1573 2163
rect 1587 2156 1813 2163
rect 1827 2156 1893 2163
rect 1947 2156 2273 2163
rect 3227 2156 3253 2163
rect 4427 2156 4753 2163
rect 5176 2163 5183 2193
rect 5176 2156 5353 2163
rect 5407 2156 5433 2163
rect 5887 2156 5973 2163
rect 4667 2136 4793 2143
rect 747 2116 1133 2123
rect 1207 2116 1233 2123
rect 2087 2116 2133 2123
rect 2147 2116 3253 2123
rect 3407 2116 4833 2123
rect 5007 2116 5193 2123
rect 5887 2116 5933 2123
rect 987 2096 1213 2103
rect 1427 2096 1533 2103
rect 3127 2096 3493 2103
rect 3747 2096 4173 2103
rect 4187 2096 4233 2103
rect 4247 2096 4733 2103
rect 4747 2096 4873 2103
rect 4887 2096 4933 2103
rect 4947 2096 5473 2103
rect 5487 2096 5773 2103
rect 5787 2096 5813 2103
rect 527 2076 673 2083
rect 1107 2076 1553 2083
rect 1627 2076 2113 2083
rect 2647 2076 3153 2083
rect 3167 2076 3853 2083
rect 4327 2076 5753 2083
rect 247 2056 433 2063
rect 447 2056 693 2063
rect 1167 2056 1333 2063
rect 1347 2056 1473 2063
rect 2287 2056 2713 2063
rect 2967 2056 3313 2063
rect 3327 2056 3353 2063
rect 3367 2056 3573 2063
rect 3587 2056 3693 2063
rect 4827 2056 5233 2063
rect 5447 2056 5513 2063
rect 5527 2056 5953 2063
rect 207 2036 853 2043
rect 1327 2036 1413 2043
rect 2347 2036 2493 2043
rect 307 2016 563 2023
rect 556 1987 563 2016
rect 1307 2016 1373 2023
rect 2387 2016 2453 2023
rect 5287 2016 5393 2023
rect 1227 1996 1313 2003
rect 1787 1996 1833 2003
rect 1907 1996 1993 2003
rect 3707 1996 3823 2003
rect 1267 1976 1333 1983
rect 3007 1976 3073 1983
rect 3816 1967 3823 1996
rect 4627 1996 4673 2003
rect 4387 1976 4453 1983
rect 1680 1963 1693 1967
rect 1667 1956 1693 1963
rect 1680 1953 1693 1956
rect 2127 1956 2173 1963
rect 3607 1963 3620 1967
rect 3607 1956 3633 1963
rect 3607 1953 3620 1956
rect 5427 1953 5433 1967
rect 5827 1956 5913 1963
rect 207 1923 220 1927
rect 207 1916 233 1923
rect 207 1913 220 1916
rect 327 1916 413 1923
rect 507 1916 573 1923
rect 600 1923 613 1927
rect 587 1916 613 1923
rect 600 1913 613 1916
rect 707 1916 793 1923
rect 847 1916 913 1923
rect 1247 1916 1313 1923
rect 1507 1916 1553 1923
rect 1987 1923 2000 1927
rect 1987 1916 2013 1923
rect 1987 1913 2000 1916
rect 3087 1913 3093 1927
rect 4107 1916 4153 1923
rect 4447 1923 4460 1927
rect 4447 1916 4473 1923
rect 4447 1913 4460 1916
rect 4827 1923 4840 1927
rect 4827 1916 4853 1923
rect 4827 1913 4840 1916
rect 1353 1907 1367 1913
rect 2473 1907 2487 1913
rect 147 1893 153 1907
rect 307 1896 353 1903
rect 1547 1896 1633 1903
rect 1907 1903 1920 1907
rect 1907 1893 1923 1903
rect 2107 1896 2353 1903
rect 2367 1896 2393 1903
rect 3133 1907 3147 1913
rect 3433 1907 3447 1913
rect 3847 1896 3953 1903
rect 767 1876 953 1883
rect 967 1876 1013 1883
rect 1916 1883 1923 1893
rect 1916 1876 2373 1883
rect 3027 1876 3113 1883
rect 5207 1876 5253 1883
rect 1407 1853 1413 1867
rect 1627 1856 1673 1863
rect 1927 1856 2113 1863
rect 2127 1856 2513 1863
rect 3467 1856 3493 1863
rect 5367 1856 5393 1863
rect 387 1836 973 1843
rect 987 1836 1233 1843
rect 1256 1836 1353 1843
rect 156 1816 533 1823
rect 156 1807 163 1816
rect 927 1816 993 1823
rect 1256 1823 1263 1836
rect 1787 1836 1953 1843
rect 2287 1836 2433 1843
rect 2447 1836 2603 1843
rect 1167 1816 1263 1823
rect 1347 1816 1913 1823
rect 2067 1816 2133 1823
rect 2487 1816 2573 1823
rect 2596 1823 2603 1836
rect 2627 1836 2773 1843
rect 3227 1836 3273 1843
rect 3367 1836 3473 1843
rect 3536 1836 4053 1843
rect 2596 1816 2893 1823
rect 3536 1823 3543 1836
rect 4387 1836 4873 1843
rect 4967 1836 5113 1843
rect 5627 1836 5653 1843
rect 5667 1836 5793 1843
rect 2907 1816 3543 1823
rect 3556 1816 3593 1823
rect 167 1796 193 1803
rect 587 1796 653 1803
rect 1687 1796 1733 1803
rect 1847 1796 1893 1803
rect 2567 1796 2873 1803
rect 2947 1796 2993 1803
rect 3387 1796 3433 1803
rect 3556 1803 3563 1816
rect 3647 1816 3893 1823
rect 4127 1816 4433 1823
rect 5307 1816 5493 1823
rect 5507 1816 5973 1823
rect 3487 1796 3563 1803
rect 4047 1796 4153 1803
rect 4207 1796 4273 1803
rect 4287 1796 4353 1803
rect 4487 1796 4773 1803
rect 5747 1796 5913 1803
rect 93 1767 107 1773
rect 536 1776 613 1783
rect 147 1756 213 1763
rect 536 1763 543 1776
rect 1167 1776 1333 1783
rect 1547 1776 1873 1783
rect 2607 1776 2633 1783
rect 3156 1776 3193 1783
rect 753 1767 767 1773
rect 487 1756 543 1763
rect 807 1756 873 1763
rect 2987 1756 3033 1763
rect 3156 1763 3163 1776
rect 3207 1776 3513 1783
rect 4467 1776 4673 1783
rect 4716 1776 4993 1783
rect 3127 1756 3163 1763
rect 2553 1747 2567 1753
rect 3893 1747 3907 1753
rect 4553 1747 4567 1753
rect 4716 1747 4723 1776
rect 5307 1776 5353 1783
rect 5467 1776 5533 1783
rect 5667 1763 5680 1767
rect 5667 1756 5693 1763
rect 5667 1753 5680 1756
rect 5807 1763 5820 1767
rect 5807 1756 5833 1763
rect 5807 1753 5820 1756
rect 1327 1736 1393 1743
rect 1487 1736 1553 1743
rect 1627 1736 1673 1743
rect 1827 1733 1833 1747
rect 2147 1736 2233 1743
rect 2407 1736 2513 1743
rect 3427 1736 3473 1743
rect 3947 1736 4033 1743
rect 4547 1733 4553 1747
rect 4787 1736 4873 1743
rect 5027 1736 5093 1743
rect 5167 1736 5213 1743
rect 3407 1713 3413 1727
rect 140 1703 153 1707
rect 127 1696 153 1703
rect 140 1693 153 1696
rect 687 1696 773 1703
rect 2887 1696 2953 1703
rect 3007 1696 3093 1703
rect 3527 1693 3533 1707
rect 4147 1703 4160 1707
rect 4147 1696 4173 1703
rect 4147 1693 4160 1696
rect 4467 1696 4533 1703
rect 5727 1696 5773 1703
rect 5827 1703 5840 1707
rect 5827 1696 5853 1703
rect 6027 1696 6123 1703
rect 5827 1693 5840 1696
rect 1073 1687 1087 1693
rect 1307 1673 1313 1687
rect 1440 1683 1453 1687
rect 1427 1676 1453 1683
rect 1440 1673 1453 1676
rect 1600 1683 1613 1687
rect 1587 1676 1613 1683
rect 1600 1673 1613 1676
rect 2647 1676 2693 1683
rect 3227 1676 3293 1683
rect 4587 1673 4593 1687
rect 4607 1676 4653 1683
rect 4907 1676 4953 1683
rect 5187 1676 5233 1683
rect 5527 1676 5593 1683
rect 1147 1656 1243 1663
rect 207 1636 233 1643
rect 547 1636 593 1643
rect 1236 1643 1243 1656
rect 1236 1636 1292 1643
rect 1328 1636 1613 1643
rect 1816 1643 1823 1673
rect 2373 1667 2387 1673
rect 2287 1656 2313 1663
rect 2416 1647 2423 1673
rect 3427 1656 3533 1663
rect 1707 1636 1893 1643
rect 2407 1643 2423 1647
rect 2407 1636 2613 1643
rect 2407 1633 2420 1636
rect 2787 1636 3293 1643
rect 3387 1636 3433 1643
rect 4016 1643 4023 1673
rect 3787 1636 4503 1643
rect 1207 1616 1313 1623
rect 1747 1616 1833 1623
rect 2267 1616 2293 1623
rect 2307 1616 2573 1623
rect 2596 1616 2733 1623
rect 827 1596 1333 1603
rect 1767 1596 1853 1603
rect 1867 1596 1953 1603
rect 2047 1596 2133 1603
rect 2596 1603 2603 1616
rect 2847 1616 3012 1623
rect 3048 1616 3213 1623
rect 3447 1613 3453 1627
rect 3847 1616 4313 1623
rect 4496 1623 4503 1636
rect 4767 1633 4773 1647
rect 5227 1636 5313 1643
rect 5367 1636 5493 1643
rect 5607 1636 5653 1643
rect 4496 1616 4753 1623
rect 4807 1616 4993 1623
rect 5107 1616 5433 1623
rect 2187 1596 2603 1603
rect 2647 1596 2813 1603
rect 2867 1596 2993 1603
rect 3016 1603 3023 1613
rect 3016 1596 3073 1603
rect 3247 1596 3863 1603
rect 3233 1587 3247 1593
rect 207 1576 473 1583
rect 647 1576 1473 1583
rect 1927 1576 2053 1583
rect 3227 1580 3247 1587
rect 3227 1576 3243 1580
rect 3227 1573 3240 1576
rect 3267 1576 3833 1583
rect 3856 1583 3863 1596
rect 3887 1596 4053 1603
rect 4067 1596 4493 1603
rect 4547 1596 4743 1603
rect 3856 1576 4413 1583
rect 4736 1583 4743 1596
rect 5047 1596 5173 1603
rect 4736 1576 5233 1583
rect 5247 1576 5353 1583
rect 447 1556 893 1563
rect 907 1556 1253 1563
rect 1827 1556 2213 1563
rect 2236 1556 2773 1563
rect 587 1536 673 1543
rect 747 1536 933 1543
rect 1287 1536 1553 1543
rect 1687 1536 2093 1543
rect 2236 1543 2243 1556
rect 3016 1556 3173 1563
rect 2107 1536 2243 1543
rect 2427 1536 2663 1543
rect 287 1516 373 1523
rect 1787 1516 1873 1523
rect 2007 1516 2173 1523
rect 2656 1523 2663 1536
rect 2827 1536 2873 1543
rect 3016 1543 3023 1556
rect 3196 1556 3373 1563
rect 2967 1536 3023 1543
rect 3196 1543 3203 1556
rect 3747 1556 4093 1563
rect 4107 1556 4593 1563
rect 5356 1563 5363 1573
rect 5356 1556 5613 1563
rect 3047 1536 3203 1543
rect 3307 1536 3493 1543
rect 3507 1536 4452 1543
rect 4488 1536 4693 1543
rect 4707 1536 4813 1543
rect 4827 1536 4853 1543
rect 4867 1536 4953 1543
rect 5087 1536 5733 1543
rect 5787 1536 5893 1543
rect 2656 1516 2813 1523
rect 3427 1516 3653 1523
rect 4427 1516 4773 1523
rect 5047 1516 5093 1523
rect 107 1496 253 1503
rect 267 1496 473 1503
rect 1667 1496 2113 1503
rect 2240 1503 2253 1507
rect 2127 1496 2253 1503
rect 2236 1493 2253 1496
rect 2327 1496 2353 1503
rect 2747 1496 2872 1503
rect 2908 1496 2993 1503
rect 3007 1496 3093 1503
rect 3547 1496 3593 1503
rect 4227 1496 4663 1503
rect 347 1476 433 1483
rect 847 1476 893 1483
rect 1767 1483 1780 1487
rect 1767 1473 1787 1483
rect 1907 1476 2033 1483
rect 1773 1467 1787 1473
rect 2236 1467 2243 1493
rect 4656 1487 4663 1496
rect 5016 1496 5133 1503
rect 2607 1476 2633 1483
rect 3347 1476 3513 1483
rect 4447 1476 4533 1483
rect 4667 1476 4693 1483
rect 5016 1467 5023 1496
rect 5967 1496 5993 1503
rect 1387 1456 1453 1463
rect 2380 1463 2393 1467
rect 2367 1456 2393 1463
rect 2380 1453 2393 1456
rect 4107 1456 4173 1463
rect 5160 1463 5173 1467
rect 5147 1456 5173 1463
rect 5160 1453 5173 1456
rect 733 1447 747 1453
rect 2873 1447 2887 1453
rect 5733 1447 5747 1453
rect 427 1436 463 1443
rect 456 1423 463 1436
rect 487 1436 553 1443
rect 3387 1443 3400 1447
rect 3387 1436 3413 1443
rect 3387 1433 3400 1436
rect 4547 1436 4593 1443
rect 4667 1433 4673 1447
rect 5507 1436 5553 1443
rect 456 1416 513 1423
rect 127 1396 213 1403
rect 987 1396 1073 1403
rect 1567 1396 1633 1403
rect 1807 1396 1893 1403
rect 2067 1403 2080 1407
rect 2067 1396 2093 1403
rect 2067 1393 2080 1396
rect 2187 1396 2253 1403
rect 2407 1393 2413 1407
rect 2627 1396 2713 1403
rect 2947 1396 3013 1403
rect 3587 1396 3673 1403
rect 4287 1396 4393 1403
rect 5140 1403 5153 1407
rect 4887 1396 4993 1403
rect 5127 1396 5153 1403
rect 5140 1393 5153 1396
rect 5907 1396 5973 1403
rect 253 1387 267 1393
rect 307 1356 333 1363
rect 907 1356 1053 1363
rect 1476 1363 1483 1393
rect 2333 1387 2347 1393
rect 2607 1376 2673 1383
rect 2827 1383 2840 1387
rect 2827 1376 2853 1383
rect 2827 1373 2840 1376
rect 1476 1356 1613 1363
rect 2147 1356 2213 1363
rect 3056 1363 3063 1393
rect 3347 1376 3393 1383
rect 2967 1356 3063 1363
rect 3727 1356 3773 1363
rect 4236 1363 4243 1393
rect 4833 1387 4847 1393
rect 4476 1376 4513 1383
rect 4027 1356 4243 1363
rect 4476 1363 4483 1376
rect 4607 1376 4653 1383
rect 5627 1376 5673 1383
rect 4447 1356 4483 1363
rect 1367 1336 1393 1343
rect 1527 1336 1733 1343
rect 1927 1336 1953 1343
rect 2647 1336 2923 1343
rect 667 1316 893 1323
rect 1107 1316 1153 1323
rect 1167 1316 1373 1323
rect 1647 1316 2273 1323
rect 2287 1316 2653 1323
rect 2767 1316 2893 1323
rect 107 1296 133 1303
rect 627 1296 753 1303
rect 927 1296 1253 1303
rect 1507 1296 1773 1303
rect 1787 1296 2373 1303
rect 2387 1296 2633 1303
rect 2916 1303 2923 1336
rect 3607 1336 3753 1343
rect 4436 1343 4443 1353
rect 4087 1336 4443 1343
rect 4547 1336 4593 1343
rect 4847 1336 5183 1343
rect 3127 1316 3173 1323
rect 3187 1316 3623 1323
rect 3116 1303 3123 1313
rect 2916 1296 3123 1303
rect 3167 1296 3593 1303
rect 3616 1303 3623 1316
rect 3667 1316 3873 1323
rect 4076 1323 4083 1333
rect 3987 1316 4083 1323
rect 5107 1316 5153 1323
rect 5176 1323 5183 1336
rect 5907 1336 6013 1343
rect 5176 1316 5313 1323
rect 5687 1316 5893 1323
rect 3616 1296 3693 1303
rect 5287 1296 5513 1303
rect 5827 1300 5903 1303
rect 5827 1296 5907 1300
rect 5893 1287 5907 1296
rect 167 1276 193 1283
rect 687 1276 933 1283
rect 1327 1276 1433 1283
rect 2147 1276 2173 1283
rect 2227 1276 2453 1283
rect 2867 1276 2893 1283
rect 3027 1276 3053 1283
rect 3067 1276 3273 1283
rect 3287 1276 3413 1283
rect 3847 1276 4133 1283
rect 4147 1276 4293 1283
rect 4307 1276 4393 1283
rect 4587 1276 4653 1283
rect 4707 1276 4813 1283
rect 5027 1276 5473 1283
rect 327 1256 353 1263
rect 1187 1256 1303 1263
rect 627 1233 633 1247
rect 1296 1227 1303 1256
rect 1707 1256 1813 1263
rect 1827 1256 1893 1263
rect 2147 1256 2243 1263
rect 2236 1227 2243 1256
rect 2367 1256 2493 1263
rect 2747 1256 2853 1263
rect 2927 1256 3093 1263
rect 4267 1256 4453 1263
rect 4816 1256 4853 1263
rect 4816 1243 4823 1256
rect 5087 1256 5133 1263
rect 5187 1256 5213 1263
rect 5256 1247 5263 1276
rect 5487 1276 5853 1283
rect 5447 1256 5553 1263
rect 4747 1236 4823 1243
rect 5516 1243 5523 1256
rect 5947 1256 6013 1263
rect 5453 1236 5523 1243
rect 5453 1227 5467 1236
rect 267 1216 333 1223
rect 527 1216 593 1223
rect 920 1223 933 1227
rect 907 1216 933 1223
rect 920 1213 933 1216
rect 1607 1216 1713 1223
rect 2307 1216 2373 1223
rect 2787 1216 2853 1223
rect 3067 1216 3093 1223
rect 3327 1216 3363 1223
rect 3356 1203 3363 1216
rect 3387 1216 3433 1223
rect 3927 1213 3933 1227
rect 4447 1216 4493 1223
rect 5367 1216 5413 1223
rect 5627 1216 5673 1223
rect 3356 1196 3393 1203
rect 107 1173 113 1187
rect 647 1173 653 1187
rect 1387 1176 1433 1183
rect 1587 1176 1633 1183
rect 1787 1176 1833 1183
rect 2447 1176 2513 1183
rect 4127 1173 4132 1187
rect 4168 1176 4233 1183
rect 4467 1176 4553 1183
rect 4567 1176 4673 1183
rect 4727 1173 4733 1187
rect 5227 1176 5273 1183
rect 5807 1183 5820 1187
rect 5807 1176 5833 1183
rect 5807 1173 5820 1176
rect 4873 1167 4887 1173
rect 287 1156 393 1163
rect 907 1153 913 1167
rect 2887 1163 2900 1167
rect 2887 1156 2913 1163
rect 2887 1153 2900 1156
rect 3360 1163 3373 1167
rect 3347 1156 3373 1163
rect 3360 1153 3373 1156
rect 4007 1156 4073 1163
rect 5327 1156 5433 1163
rect 5527 1156 5573 1163
rect 5947 1153 5953 1167
rect 2353 1147 2367 1153
rect 127 1136 153 1143
rect 167 1136 213 1143
rect 3813 1147 3827 1153
rect 4507 1136 4813 1143
rect 347 1116 533 1123
rect 1287 1116 1733 1123
rect 1747 1116 1773 1123
rect 2127 1116 2243 1123
rect 467 1096 613 1103
rect 1296 1096 1433 1103
rect 1296 1083 1303 1096
rect 2236 1103 2243 1116
rect 2667 1116 3033 1123
rect 3047 1116 3253 1123
rect 3967 1116 4013 1123
rect 4087 1116 4373 1123
rect 5127 1116 5213 1123
rect 5696 1123 5703 1153
rect 5567 1116 5703 1123
rect 2236 1096 2433 1103
rect 3387 1096 3473 1103
rect 3947 1096 3973 1103
rect 3987 1096 4153 1103
rect 4347 1096 4413 1103
rect 607 1076 1303 1083
rect 2087 1076 2133 1083
rect 2467 1076 3213 1083
rect 3387 1076 3513 1083
rect 3887 1076 4913 1083
rect 5007 1076 5153 1083
rect 5167 1076 5393 1083
rect 5447 1076 5533 1083
rect 627 1056 1153 1063
rect 1167 1056 1373 1063
rect 1527 1056 1783 1063
rect 1776 1047 1783 1056
rect 1847 1056 2132 1063
rect 2168 1056 2193 1063
rect 2207 1056 2373 1063
rect 2727 1056 2793 1063
rect 3376 1063 3383 1073
rect 2807 1056 3383 1063
rect 3487 1056 3633 1063
rect 4587 1056 5233 1063
rect 107 1036 203 1043
rect 127 1016 153 1023
rect 196 1003 203 1036
rect 267 1036 533 1043
rect 787 1036 1073 1043
rect 1087 1036 1233 1043
rect 1247 1036 1273 1043
rect 1327 1036 1593 1043
rect 1787 1036 2013 1043
rect 2027 1036 2112 1043
rect 2148 1036 2313 1043
rect 2407 1036 2493 1043
rect 2507 1036 3153 1043
rect 3307 1036 3353 1043
rect 4287 1036 4513 1043
rect 227 1016 273 1023
rect 327 1016 493 1023
rect 847 1016 1913 1023
rect 1967 1016 2033 1023
rect 2267 1016 2353 1023
rect 2947 1016 3173 1023
rect 3267 1016 3773 1023
rect 3787 1016 4053 1023
rect 4327 1016 4703 1023
rect 633 1007 647 1013
rect 4696 1007 4703 1016
rect 4847 1016 4873 1023
rect 196 996 233 1003
rect 2307 996 2333 1003
rect 2687 996 2733 1003
rect 3127 996 3433 1003
rect 3487 996 3513 1003
rect 3647 996 4013 1003
rect 4707 996 4753 1003
rect 4767 996 4993 1003
rect 167 976 273 983
rect 287 976 312 983
rect 348 976 373 983
rect 507 976 693 983
rect 1187 976 1253 983
rect 2227 976 2433 983
rect 2447 976 2753 983
rect 2947 976 2973 983
rect 3207 976 3253 983
rect 3407 976 3593 983
rect 3607 976 3893 983
rect 4887 976 4953 983
rect 4967 976 5173 983
rect 5187 976 5293 983
rect 647 956 883 963
rect 507 943 520 947
rect 507 936 533 943
rect 507 933 520 936
rect 876 927 883 956
rect 2647 956 2772 963
rect 2808 956 2833 963
rect 2847 956 2913 963
rect 5207 956 5233 963
rect 2367 936 2473 943
rect 2547 936 2593 943
rect 4007 943 4020 947
rect 4007 936 4033 943
rect 4007 933 4020 936
rect 4367 933 4373 947
rect 4747 936 4793 943
rect 5060 943 5073 947
rect 5047 936 5073 943
rect 5060 933 5073 936
rect 5507 936 5573 943
rect 5707 936 5773 943
rect 4693 927 4707 933
rect 767 916 833 923
rect 947 916 1033 923
rect 2087 916 2133 923
rect 2707 923 2720 927
rect 2707 916 2733 923
rect 2707 913 2720 916
rect 2787 916 2853 923
rect 2867 916 2933 923
rect 3327 916 3393 923
rect 6047 896 6073 903
rect 267 876 313 883
rect 447 876 493 883
rect 607 876 673 883
rect 1467 876 1523 883
rect 93 867 107 873
rect 1516 867 1523 876
rect 3047 876 3112 883
rect 3148 883 3160 887
rect 3148 876 3173 883
rect 3148 873 3160 876
rect 3480 883 3492 887
rect 3467 876 3492 883
rect 3480 873 3492 876
rect 3528 876 3613 883
rect 3927 876 4013 883
rect 4227 876 4333 883
rect 4747 873 4753 887
rect 5027 876 5113 883
rect 5380 883 5393 887
rect 5247 876 5313 883
rect 5367 876 5393 883
rect 5380 873 5393 876
rect 5547 876 5633 883
rect 5927 873 5933 887
rect 5947 876 6053 883
rect 327 856 373 863
rect 847 853 853 867
rect 1067 853 1073 867
rect 1516 856 1533 867
rect 1520 853 1533 856
rect 267 836 333 843
rect 407 836 553 843
rect 607 836 653 843
rect 1187 836 1253 843
rect 2427 836 2473 843
rect 2927 836 2993 843
rect 3407 836 3693 843
rect 3756 843 3763 873
rect 3756 836 4133 843
rect 4176 843 4183 873
rect 4853 867 4867 873
rect 4176 836 4273 843
rect 5156 843 5163 873
rect 5156 836 5213 843
rect 5476 843 5483 873
rect 5447 836 5483 843
rect 5587 836 5753 843
rect 5767 836 5953 843
rect 147 816 173 823
rect 187 816 233 823
rect 467 816 613 823
rect 627 813 633 827
rect 1027 816 1193 823
rect 2487 816 2653 823
rect 2707 816 2833 823
rect 2887 816 3013 823
rect 3327 816 3353 823
rect 3507 816 4383 823
rect 107 796 313 803
rect 907 796 933 803
rect 1087 796 1133 803
rect 1427 796 1643 803
rect 1636 787 1643 796
rect 1967 796 2013 803
rect 2627 796 2973 803
rect 3253 803 3267 813
rect 2987 796 3913 803
rect 4376 803 4383 816
rect 5347 816 5473 823
rect 4376 796 4593 803
rect 4647 796 5653 803
rect 5667 796 5893 803
rect 307 776 493 783
rect 567 780 663 783
rect 567 776 667 780
rect 653 767 667 776
rect 707 776 773 783
rect 987 776 1153 783
rect 1207 776 1293 783
rect 1487 776 1533 783
rect 1647 776 1833 783
rect 1927 776 3253 783
rect 3376 776 3453 783
rect 207 756 253 763
rect 427 756 632 763
rect 653 760 654 767
rect 1407 756 1453 763
rect 1607 756 1713 763
rect 1727 756 1973 763
rect 2027 756 2253 763
rect 2547 756 2573 763
rect 2667 756 2733 763
rect 2747 756 2793 763
rect 3107 753 3113 767
rect 3376 763 3383 776
rect 3787 780 4042 783
rect 3787 776 4047 780
rect 4033 767 4047 776
rect 4336 776 4373 783
rect 4336 767 4343 776
rect 4827 776 5593 783
rect 5607 776 5693 783
rect 3207 756 3383 763
rect 3707 756 3753 763
rect 4046 760 4047 767
rect 4068 756 4113 763
rect 4327 756 4343 767
rect 4327 753 4340 756
rect 4367 756 4473 763
rect 4607 756 4693 763
rect 5767 756 5793 763
rect 576 736 653 743
rect 576 707 583 736
rect 1527 736 1633 743
rect 1676 736 1913 743
rect 1267 716 1353 723
rect 1533 707 1547 713
rect 1676 707 1683 736
rect 2067 736 2233 743
rect 2347 736 2373 743
rect 2647 736 2673 743
rect 2947 736 3013 743
rect 3027 736 3233 743
rect 3247 736 3333 743
rect 3647 736 3673 743
rect 4187 736 4293 743
rect 4347 736 4373 743
rect 4827 736 4853 743
rect 4927 736 4993 743
rect 3287 713 3293 727
rect 307 696 373 703
rect 807 696 853 703
rect 1727 696 1813 703
rect 2587 693 2593 707
rect 2647 696 2693 703
rect 3187 693 3192 707
rect 3228 696 3333 703
rect 3587 696 3633 703
rect 3727 696 3773 703
rect 3887 696 3913 703
rect 4287 696 4333 703
rect 4427 696 4473 703
rect 4787 696 4873 703
rect 5327 696 5393 703
rect 5487 696 5533 703
rect 5787 696 5853 703
rect 147 656 193 663
rect 447 656 493 663
rect 947 656 993 663
rect 1307 656 1373 663
rect 2087 656 2133 663
rect 2147 653 2153 667
rect 2207 656 2293 663
rect 2767 656 2833 663
rect 3047 656 3113 663
rect 4107 656 4173 663
rect 4307 656 4353 663
rect 4587 656 4633 663
rect 4747 656 4813 663
rect 5027 653 5033 667
rect 5967 663 5980 667
rect 5967 656 5993 663
rect 5967 653 5980 656
rect 1993 647 2007 653
rect 5713 647 5727 653
rect 727 636 793 643
rect 1580 643 1593 647
rect 1567 636 1593 643
rect 1580 633 1593 636
rect 2467 636 2573 643
rect 2887 636 2933 643
rect 4167 636 4213 643
rect 4267 636 4353 643
rect 5927 633 5933 647
rect 87 616 173 623
rect 716 603 723 633
rect 1793 627 1807 633
rect 3353 627 3367 633
rect 1967 616 2233 623
rect 3467 616 3513 623
rect 3647 616 3673 623
rect 5927 616 5973 623
rect 607 596 723 603
rect 807 596 953 603
rect 1367 596 1653 603
rect 1847 596 2073 603
rect 2547 593 2552 607
rect 2588 596 2613 603
rect 2867 596 3253 603
rect 4327 596 4393 603
rect 4827 596 4853 603
rect 4907 596 4953 603
rect 4967 596 5013 603
rect 387 576 673 583
rect 687 576 873 583
rect 2546 573 2547 580
rect 2907 576 2932 583
rect 2968 576 3072 583
rect 3108 576 3153 583
rect 4047 576 4113 583
rect 4247 576 4332 583
rect 4368 576 4553 583
rect 4567 576 4673 583
rect 2533 567 2547 573
rect 427 556 573 563
rect 647 553 653 567
rect 747 556 1013 563
rect 1027 556 1293 563
rect 2546 560 2547 567
rect 2568 553 2573 567
rect 2587 556 3272 563
rect 3308 556 3333 563
rect 3627 553 3633 567
rect 3647 556 3713 563
rect 4236 563 4243 573
rect 3727 556 4243 563
rect 4367 556 4433 563
rect 4547 556 4773 563
rect 5027 556 5833 563
rect 5907 553 5913 567
rect 127 536 213 543
rect 1047 536 1253 543
rect 1267 536 1493 543
rect 1507 536 1573 543
rect 1587 536 1873 543
rect 2047 536 2153 543
rect 2307 536 2473 543
rect 2487 536 4753 543
rect 4807 536 4833 543
rect 5287 536 5633 543
rect 216 523 223 533
rect 216 516 413 523
rect 2007 516 3183 523
rect 287 496 613 503
rect 627 496 693 503
rect 867 496 932 503
rect 968 496 1073 503
rect 1487 496 1553 503
rect 1807 496 2053 503
rect 3176 503 3183 516
rect 3207 516 3753 523
rect 3767 516 4013 523
rect 4527 516 4573 523
rect 2207 496 3163 503
rect 3176 496 3843 503
rect 107 476 333 483
rect 1047 476 1233 483
rect 3156 483 3163 496
rect 3156 476 3673 483
rect 3836 483 3843 496
rect 3867 496 3953 503
rect 3967 496 4153 503
rect 4267 496 5093 503
rect 3836 476 3893 483
rect 4027 476 4433 483
rect 5247 476 5313 483
rect 5707 476 5773 483
rect 227 456 433 463
rect 507 456 693 463
rect 707 456 993 463
rect 1007 456 1093 463
rect 1167 456 1393 463
rect 2627 456 2773 463
rect 3167 456 3493 463
rect 4047 456 4373 463
rect 4767 456 5013 463
rect 5307 456 5393 463
rect 5487 456 5533 463
rect 5627 456 5753 463
rect 5907 456 5933 463
rect 2573 447 2587 453
rect 347 436 373 443
rect 2167 436 2293 443
rect 4447 436 4473 443
rect 5607 436 5633 443
rect 553 427 567 433
rect 787 416 833 423
rect 1727 416 1773 423
rect 2667 416 2733 423
rect 3247 416 3333 423
rect 3467 413 3473 427
rect 5387 413 5393 427
rect 5987 423 6000 427
rect 5987 416 6013 423
rect 5987 413 6000 416
rect 433 407 447 413
rect 2193 407 2207 413
rect 127 396 193 403
rect 647 403 660 407
rect 647 396 673 403
rect 647 393 660 396
rect 1147 396 1193 403
rect 2527 396 2573 403
rect 2827 393 2833 407
rect 2887 393 2893 407
rect 3107 396 3153 403
rect 3507 396 3593 403
rect 3767 393 3773 407
rect 4167 396 4233 403
rect 4827 396 4893 403
rect 5067 396 5133 403
rect 267 356 333 363
rect 767 356 853 363
rect 987 356 1033 363
rect 1280 363 1293 367
rect 1267 356 1293 363
rect 1280 353 1293 356
rect 1427 356 1473 363
rect 1727 356 1793 363
rect 2067 356 2133 363
rect 2727 356 2753 363
rect 3087 353 3093 367
rect 3367 353 3373 367
rect 3487 353 3493 367
rect 4667 356 4713 363
rect 5167 363 5180 367
rect 5167 356 5193 363
rect 5167 353 5180 356
rect 5307 356 5353 363
rect 2673 347 2687 353
rect 1467 336 1493 343
rect 1567 336 1613 343
rect 4547 336 4593 343
rect 3573 327 3587 333
rect 1707 313 1713 327
rect 1727 316 1853 323
rect 2347 316 2473 323
rect 2587 316 2633 323
rect 2647 316 2693 323
rect 2747 313 2753 327
rect 2807 316 2873 323
rect 3267 316 3503 323
rect 613 307 627 313
rect 687 296 773 303
rect 796 296 1033 303
rect 796 283 803 296
rect 1567 296 1613 303
rect 1947 296 1993 303
rect 2187 296 2233 303
rect 2307 296 2853 303
rect 3147 296 3473 303
rect 3496 303 3503 316
rect 4687 316 4813 323
rect 5147 316 5193 323
rect 5207 316 5233 323
rect 5247 316 5313 323
rect 5736 323 5743 353
rect 5873 347 5887 353
rect 5647 316 5743 323
rect 5807 316 5993 323
rect 3496 296 3753 303
rect 4927 296 5393 303
rect 507 276 803 283
rect 1027 276 1093 283
rect 1227 276 2213 283
rect 2547 276 2713 283
rect 2767 276 3113 283
rect 3127 276 3333 283
rect 3687 276 4072 283
rect 4108 276 4633 283
rect 5887 276 5953 283
rect 307 256 1363 263
rect 167 236 233 243
rect 687 236 793 243
rect 1356 243 1363 256
rect 1387 256 1453 263
rect 1467 256 1813 263
rect 1827 256 1893 263
rect 1907 256 2373 263
rect 2527 256 2633 263
rect 2687 256 3053 263
rect 3107 256 3613 263
rect 3627 256 3693 263
rect 3707 256 3833 263
rect 3847 256 3933 263
rect 3947 256 4213 263
rect 4227 256 4873 263
rect 4887 256 4913 263
rect 4927 256 5073 263
rect 5115 260 5153 263
rect 5113 256 5153 260
rect 5113 247 5127 256
rect 5327 256 5913 263
rect 1356 236 1533 243
rect 1787 236 2213 243
rect 2267 236 2453 243
rect 2927 236 2953 243
rect 3747 236 4293 243
rect 5126 240 5127 247
rect 5148 236 5173 243
rect 5567 236 5613 243
rect 116 216 293 223
rect 116 187 123 216
rect 636 216 913 223
rect 233 187 247 193
rect 636 187 643 216
rect 2456 223 2463 233
rect 2456 216 2593 223
rect 3587 216 3773 223
rect 3787 216 4053 223
rect 4067 216 4213 223
rect 4267 216 4583 223
rect 2107 193 2113 207
rect 2687 196 2733 203
rect 3227 196 3253 203
rect 4293 187 4307 193
rect 4576 187 4583 216
rect 4807 216 4873 223
rect 5167 216 5233 223
rect 5327 196 5373 203
rect 5567 196 5613 203
rect 967 176 1013 183
rect 1267 176 1333 183
rect 1507 173 1513 187
rect 1807 176 1873 183
rect 2407 176 2473 183
rect 2527 173 2533 187
rect 2907 173 2913 187
rect 3347 176 3393 183
rect 3607 176 3693 183
rect 3827 176 3893 183
rect 4407 183 4420 187
rect 4407 176 4433 183
rect 4407 173 4420 176
rect 4647 176 4713 183
rect 4907 176 4943 183
rect 4936 163 4943 176
rect 4967 176 5033 183
rect 5147 183 5160 187
rect 5147 176 5173 183
rect 5147 173 5160 176
rect 5467 183 5480 187
rect 5467 176 5493 183
rect 5467 173 5480 176
rect 5707 176 5773 183
rect 4936 156 4993 163
rect 827 136 893 143
rect 4467 133 4473 147
rect 4607 133 4613 147
rect 4747 133 4753 147
rect 2033 127 2047 133
rect 107 116 173 123
rect 667 116 713 123
rect 1247 116 1313 123
rect 1787 116 1853 123
rect 2233 127 2247 133
rect 3073 127 3087 133
rect 2440 123 2453 127
rect 2427 116 2453 123
rect 2440 113 2453 116
rect 2940 123 2953 127
rect 2927 116 2953 123
rect 2940 113 2953 116
rect 1647 96 1693 103
rect 907 76 933 83
rect 1307 76 1473 83
rect 1856 83 1863 113
rect 2007 96 2273 103
rect 3787 96 3833 103
rect 4336 103 4343 133
rect 5807 116 5853 123
rect 4336 96 4773 103
rect 5687 96 5753 103
rect 5936 103 5943 133
rect 5847 96 5943 103
rect 5987 96 6033 103
rect 1856 76 2113 83
rect 2427 76 2553 83
rect 2827 76 3033 83
rect 3367 76 4153 83
rect 4207 76 4953 83
rect 5067 76 5233 83
rect 2087 56 2173 63
rect 3427 56 3713 63
rect 3927 56 5153 63
rect 167 36 203 43
rect 196 23 203 36
rect 267 36 333 43
rect 987 36 1253 43
rect 1527 36 1793 43
rect 2247 36 3293 43
rect 3347 36 3373 43
rect 3487 36 3573 43
rect 5127 36 5373 43
rect 196 16 433 23
rect 2047 16 3413 23
rect 3467 16 3493 23
<< m3contact >>
rect 1093 5993 1107 6007
rect 1313 5993 1327 6007
rect 1453 5993 1467 6007
rect 133 5973 147 5987
rect 213 5973 227 5987
rect 833 5973 847 5987
rect 893 5973 907 5987
rect 1133 5973 1147 5987
rect 1293 5973 1307 5987
rect 2293 5973 2307 5987
rect 2653 5973 2667 5987
rect 2753 5973 2767 5987
rect 2893 5973 2907 5987
rect 2933 5973 2947 5987
rect 3073 5973 3087 5987
rect 3213 5973 3227 5987
rect 3313 5973 3327 5987
rect 3493 5973 3507 5987
rect 3673 5993 3687 6007
rect 4133 5993 4147 6007
rect 3713 5973 3727 5987
rect 3753 5973 3767 5987
rect 3833 5973 3847 5987
rect 4293 5973 4307 5987
rect 4393 5973 4407 5987
rect 4613 5993 4627 6007
rect 5173 5993 5187 6007
rect 5253 5993 5267 6007
rect 5513 5993 5527 6007
rect 4913 5973 4927 5987
rect 4953 5973 4967 5987
rect 5213 5973 5227 5987
rect 5293 5973 5307 5987
rect 5353 5973 5367 5987
rect 433 5953 447 5967
rect 1673 5953 1687 5967
rect 1933 5953 1947 5967
rect 2013 5953 2027 5967
rect 4093 5953 4107 5967
rect 453 5933 467 5947
rect 613 5933 627 5947
rect 1233 5933 1247 5947
rect 1613 5933 1627 5947
rect 1873 5933 1887 5947
rect 2193 5933 2207 5947
rect 2253 5933 2267 5947
rect 2553 5933 2567 5947
rect 2613 5933 2627 5947
rect 2753 5933 2767 5947
rect 2833 5933 2847 5947
rect 3173 5933 3187 5947
rect 3673 5933 3687 5947
rect 4833 5953 4847 5967
rect 5252 5953 5266 5967
rect 5333 5953 5347 5967
rect 5373 5953 5387 5967
rect 5473 5953 5487 5967
rect 2233 5913 2247 5927
rect 2293 5913 2307 5927
rect 2793 5913 2807 5927
rect 3493 5913 3507 5927
rect 3553 5913 3567 5927
rect 3613 5913 3627 5927
rect 4253 5913 4267 5927
rect 4293 5913 4307 5927
rect 4653 5933 4667 5947
rect 4793 5933 4807 5947
rect 4953 5933 4967 5947
rect 5393 5933 5407 5947
rect 5553 5933 5567 5947
rect 5773 5933 5787 5947
rect 4973 5913 4987 5927
rect 5013 5913 5027 5927
rect 5133 5913 5147 5927
rect 5253 5913 5267 5927
rect 5373 5913 5387 5927
rect 93 5893 107 5907
rect 133 5893 147 5907
rect 173 5893 187 5907
rect 253 5893 267 5907
rect 334 5893 348 5907
rect 453 5893 467 5907
rect 613 5893 627 5907
rect 793 5893 807 5907
rect 833 5893 847 5907
rect 953 5893 967 5907
rect 1033 5893 1047 5907
rect 1153 5893 1167 5907
rect 1293 5893 1307 5907
rect 1353 5893 1367 5907
rect 1533 5893 1547 5907
rect 1573 5893 1587 5907
rect 1613 5893 1627 5907
rect 1673 5893 1687 5907
rect 1933 5893 1947 5907
rect 2013 5893 2027 5907
rect 2193 5893 2207 5907
rect 2333 5893 2347 5907
rect 2613 5893 2627 5907
rect 2653 5893 2667 5907
rect 2893 5893 2907 5907
rect 3013 5893 3027 5907
rect 3193 5893 3207 5907
rect 3253 5893 3267 5907
rect 3373 5893 3387 5907
rect 3413 5893 3427 5907
rect 3453 5893 3467 5907
rect 3533 5893 3547 5907
rect 3573 5893 3587 5907
rect 3693 5893 3707 5907
rect 3833 5893 3847 5907
rect 3873 5893 3887 5907
rect 4053 5893 4067 5907
rect 4073 5893 4087 5907
rect 4573 5893 4587 5907
rect 4653 5893 4667 5907
rect 4833 5893 4847 5907
rect 5173 5893 5187 5907
rect 5213 5893 5227 5907
rect 5573 5893 5587 5907
rect 5613 5893 5627 5907
rect 5733 5893 5747 5907
rect 5773 5893 5787 5907
rect 5913 5893 5927 5907
rect 713 5873 727 5887
rect 873 5873 887 5887
rect 2533 5873 2547 5887
rect 2573 5873 2587 5887
rect 1833 5853 1847 5867
rect 2113 5853 2127 5867
rect 2293 5853 2307 5867
rect 2433 5853 2447 5867
rect 2673 5853 2687 5867
rect 3073 5853 3087 5867
rect 3173 5853 3187 5867
rect 3233 5853 3247 5867
rect 4093 5853 4107 5867
rect 4193 5853 4207 5867
rect 4233 5853 4247 5867
rect 4313 5853 4327 5867
rect 4393 5853 4407 5867
rect 4772 5853 4786 5867
rect 4794 5853 4808 5867
rect 4873 5853 4887 5867
rect 4953 5853 4967 5867
rect 5033 5853 5047 5867
rect 5133 5853 5147 5867
rect 5193 5853 5207 5867
rect 5233 5853 5247 5867
rect 5313 5853 5327 5867
rect 5353 5853 5367 5867
rect 5393 5853 5407 5867
rect 6073 5853 6087 5867
rect 113 5833 127 5847
rect 153 5833 167 5847
rect 233 5833 247 5847
rect 273 5833 287 5847
rect 433 5833 447 5847
rect 473 5833 487 5847
rect 513 5833 527 5847
rect 553 5833 567 5847
rect 593 5833 607 5847
rect 633 5833 647 5847
rect 673 5833 687 5847
rect 733 5833 747 5847
rect 773 5833 787 5847
rect 813 5833 827 5847
rect 893 5833 907 5847
rect 973 5833 987 5847
rect 1133 5833 1147 5847
rect 1233 5833 1247 5847
rect 1273 5833 1287 5847
rect 1313 5833 1327 5847
rect 1453 5833 1467 5847
rect 1493 5833 1507 5847
rect 1593 5833 1607 5847
rect 1633 5833 1647 5847
rect 1733 5833 1747 5847
rect 1773 5833 1787 5847
rect 2173 5833 2187 5847
rect 2213 5833 2227 5847
rect 2473 5833 2487 5847
rect 2513 5833 2527 5847
rect 2593 5833 2607 5847
rect 2633 5833 2647 5847
rect 2873 5833 2887 5847
rect 2913 5833 2927 5847
rect 3353 5833 3367 5847
rect 3393 5833 3407 5847
rect 3513 5833 3527 5847
rect 3553 5833 3567 5847
rect 3713 5833 3727 5847
rect 3813 5833 3827 5847
rect 3953 5833 3967 5847
rect 3993 5833 4007 5847
rect 4273 5833 4287 5847
rect 4573 5833 4587 5847
rect 593 5793 607 5807
rect 633 5793 647 5807
rect 733 5793 747 5807
rect 853 5813 867 5827
rect 2553 5813 2567 5827
rect 2713 5813 2727 5827
rect 2793 5813 2807 5827
rect 2953 5813 2967 5827
rect 3033 5813 3047 5827
rect 3093 5813 3107 5827
rect 3233 5813 3247 5827
rect 3273 5813 3287 5827
rect 3433 5813 3447 5827
rect 3673 5813 3687 5827
rect 4233 5813 4247 5827
rect 4473 5813 4487 5827
rect 4733 5813 4747 5827
rect 5473 5833 5487 5847
rect 5513 5833 5527 5847
rect 5633 5833 5647 5847
rect 5893 5833 5907 5847
rect 893 5793 907 5807
rect 933 5793 947 5807
rect 1033 5793 1047 5807
rect 1533 5793 1547 5807
rect 1593 5793 1607 5807
rect 1673 5793 1687 5807
rect 2313 5793 2327 5807
rect 3013 5793 3027 5807
rect 4073 5794 4087 5808
rect 5393 5813 5407 5827
rect 5434 5813 5448 5827
rect 4133 5793 4147 5807
rect 4193 5793 4207 5807
rect 4293 5793 4307 5807
rect 4913 5793 4927 5807
rect 5113 5793 5127 5807
rect 773 5773 787 5787
rect 973 5773 987 5787
rect 1313 5773 1327 5787
rect 1413 5773 1427 5787
rect 1774 5773 1788 5787
rect 93 5753 107 5767
rect 233 5753 247 5767
rect 293 5753 307 5767
rect 513 5753 527 5767
rect 554 5753 568 5767
rect 793 5753 807 5767
rect 953 5753 967 5767
rect 1153 5753 1167 5767
rect 1573 5753 1587 5767
rect 113 5733 127 5747
rect 273 5733 287 5747
rect 693 5733 707 5747
rect 1453 5733 1467 5747
rect 1713 5733 1727 5747
rect 1753 5753 1767 5767
rect 1793 5753 1807 5767
rect 2113 5773 2127 5787
rect 2173 5773 2187 5787
rect 2333 5773 2347 5787
rect 2792 5773 2806 5787
rect 2814 5773 2828 5787
rect 2993 5773 3007 5787
rect 3033 5773 3047 5787
rect 2433 5753 2447 5767
rect 2513 5753 2527 5767
rect 2133 5733 2147 5747
rect 2633 5733 2647 5747
rect 2753 5733 2767 5747
rect 2833 5733 2847 5747
rect 2913 5753 2927 5767
rect 3313 5753 3327 5767
rect 3393 5773 3407 5787
rect 3513 5773 3527 5787
rect 4073 5772 4087 5786
rect 4173 5773 4187 5787
rect 4233 5774 4247 5788
rect 4273 5773 4287 5787
rect 4533 5773 4547 5787
rect 4593 5773 4607 5787
rect 4653 5773 4667 5787
rect 4754 5773 4768 5787
rect 4973 5773 4987 5787
rect 5153 5773 5167 5787
rect 5293 5794 5307 5808
rect 5413 5793 5427 5807
rect 5513 5793 5527 5807
rect 5633 5793 5647 5807
rect 5893 5793 5907 5807
rect 5973 5793 5987 5807
rect 5293 5772 5307 5786
rect 5473 5773 5487 5787
rect 3594 5753 3608 5767
rect 2953 5733 2967 5747
rect 2993 5733 3007 5747
rect 1493 5713 1507 5727
rect 1733 5713 1747 5727
rect 1993 5713 2007 5727
rect 2073 5713 2087 5727
rect 2813 5713 2827 5727
rect 2873 5713 2887 5727
rect 3093 5713 3107 5727
rect 3273 5734 3287 5748
rect 3633 5733 3647 5747
rect 3953 5753 3967 5767
rect 4093 5753 4107 5767
rect 4233 5752 4247 5766
rect 4693 5753 4707 5767
rect 5033 5753 5047 5767
rect 5274 5753 5288 5767
rect 3273 5712 3287 5726
rect 3313 5713 3327 5727
rect 3793 5713 3807 5727
rect 4613 5733 4627 5747
rect 4833 5733 4847 5747
rect 5413 5733 5427 5747
rect 3873 5713 3887 5727
rect 3993 5713 4007 5727
rect 4293 5713 4307 5727
rect 4473 5713 4487 5727
rect 4653 5713 4667 5727
rect 913 5693 927 5707
rect 1013 5693 1027 5707
rect 1233 5693 1247 5707
rect 1753 5693 1767 5707
rect 1833 5693 1847 5707
rect 2433 5693 2447 5707
rect 2833 5693 2847 5707
rect 3133 5693 3147 5707
rect 3293 5693 3307 5707
rect 3333 5693 3347 5707
rect 3673 5694 3687 5708
rect 3714 5693 3728 5707
rect 3753 5693 3767 5707
rect 4573 5693 4587 5707
rect 4852 5713 4866 5727
rect 4874 5713 4888 5727
rect 5333 5713 5347 5727
rect 4792 5693 4806 5707
rect 4814 5693 4828 5707
rect 5093 5693 5107 5707
rect 5373 5693 5387 5707
rect 5453 5693 5467 5707
rect 5553 5693 5567 5707
rect 1313 5673 1327 5687
rect 1493 5673 1507 5687
rect 2253 5673 2267 5687
rect 2713 5673 2727 5687
rect 2873 5673 2887 5687
rect 2973 5673 2987 5687
rect 113 5653 127 5667
rect 233 5653 247 5667
rect 433 5653 447 5667
rect 553 5653 567 5667
rect 753 5653 767 5667
rect 1213 5653 1227 5667
rect 1253 5653 1267 5667
rect 1513 5653 1527 5667
rect 2033 5653 2047 5667
rect 2413 5653 2427 5667
rect 2553 5653 2567 5667
rect 3393 5673 3407 5687
rect 3433 5673 3447 5687
rect 3673 5672 3687 5686
rect 3733 5673 3747 5687
rect 3813 5673 3827 5687
rect 3953 5673 3967 5687
rect 4133 5673 4147 5687
rect 4773 5673 4787 5687
rect 4933 5673 4947 5687
rect 4972 5673 4986 5687
rect 4994 5673 5008 5687
rect 5173 5673 5187 5687
rect 5273 5673 5287 5687
rect 5573 5673 5587 5687
rect 5773 5673 5787 5687
rect 3633 5653 3647 5667
rect 3773 5653 3787 5667
rect 3852 5653 3866 5667
rect 3874 5653 3888 5667
rect 1293 5633 1307 5647
rect 1353 5633 1367 5647
rect 113 5613 127 5627
rect 153 5613 167 5627
rect 233 5613 247 5627
rect 273 5613 287 5627
rect 433 5613 447 5627
rect 473 5613 487 5627
rect 553 5613 567 5627
rect 593 5613 607 5627
rect 633 5613 647 5627
rect 753 5613 767 5627
rect 793 5613 807 5627
rect 1013 5613 1027 5627
rect 1053 5613 1067 5627
rect 1173 5613 1187 5627
rect 1213 5613 1227 5627
rect 1593 5613 1607 5627
rect 1633 5613 1647 5627
rect 1793 5633 1807 5647
rect 2993 5633 3007 5647
rect 2133 5613 2147 5627
rect 2433 5613 2447 5627
rect 2473 5613 2487 5627
rect 2593 5613 2607 5627
rect 2633 5613 2647 5627
rect 2713 5613 2727 5627
rect 2753 5613 2767 5627
rect 2873 5613 2887 5627
rect 4213 5653 4227 5667
rect 4373 5653 4387 5667
rect 4413 5653 4427 5667
rect 4593 5653 4607 5667
rect 4653 5653 4667 5667
rect 5293 5653 5307 5667
rect 5733 5653 5747 5667
rect 5813 5653 5827 5667
rect 5993 5653 6007 5667
rect 3133 5613 3147 5627
rect 3213 5613 3227 5627
rect 3313 5613 3327 5627
rect 3353 5613 3367 5627
rect 3493 5613 3507 5627
rect 3533 5613 3547 5627
rect 3673 5613 3687 5627
rect 3773 5613 3787 5627
rect 3893 5613 3907 5627
rect 3933 5613 3947 5627
rect 4013 5613 4027 5627
rect 4093 5613 4107 5627
rect 4393 5613 4407 5627
rect 4493 5613 4507 5627
rect 4533 5613 4547 5627
rect 4653 5613 4667 5627
rect 4693 5613 4707 5627
rect 1253 5593 1267 5607
rect 1733 5593 1747 5607
rect 1813 5593 1827 5607
rect 1993 5593 2007 5607
rect 2093 5593 2107 5607
rect 2173 5593 2187 5607
rect 2213 5593 2227 5607
rect 3013 5593 3027 5607
rect 3093 5593 3107 5607
rect 4133 5593 4147 5607
rect 4253 5593 4267 5607
rect 4293 5593 4307 5607
rect 4793 5633 4807 5647
rect 4953 5613 4967 5627
rect 4993 5613 5007 5627
rect 5173 5613 5187 5627
rect 5293 5613 5307 5627
rect 5333 5613 5347 5627
rect 5413 5613 5427 5627
rect 5453 5613 5467 5627
rect 5733 5613 5747 5627
rect 5773 5613 5787 5627
rect 5853 5613 5867 5627
rect 5893 5613 5907 5627
rect 5993 5613 6007 5627
rect 6033 5613 6047 5627
rect 4773 5593 4787 5607
rect 4853 5593 4867 5607
rect 5113 5593 5127 5607
rect 5253 5593 5267 5607
rect 5493 5593 5507 5607
rect 5633 5593 5647 5607
rect 4713 5573 4727 5587
rect 5833 5574 5847 5588
rect 133 5553 147 5567
rect 253 5553 267 5567
rect 313 5553 327 5567
rect 453 5553 467 5567
rect 573 5553 587 5567
rect 653 5553 667 5567
rect 693 5553 707 5567
rect 773 5553 787 5567
rect 913 5553 927 5567
rect 993 5553 1007 5567
rect 1153 5553 1167 5567
rect 1233 5553 1247 5567
rect 1533 5553 1547 5567
rect 1953 5553 1967 5567
rect 2313 5553 2327 5567
rect 2353 5553 2367 5567
rect 2453 5553 2467 5567
rect 2573 5553 2587 5567
rect 2613 5553 2627 5567
rect 2793 5553 2807 5567
rect 2893 5553 2907 5567
rect 2933 5553 2947 5567
rect 3193 5553 3207 5567
rect 3333 5553 3347 5567
rect 3373 5553 3387 5567
rect 3613 5553 3627 5567
rect 3653 5553 3667 5567
rect 3693 5553 3707 5567
rect 3793 5553 3807 5567
rect 3873 5553 3887 5567
rect 4073 5553 4087 5567
rect 4233 5553 4247 5567
rect 4373 5553 4387 5567
rect 4553 5553 4567 5567
rect 4593 5553 4607 5567
rect 4973 5553 4987 5567
rect 5153 5553 5167 5567
rect 5333 5553 5347 5567
rect 5433 5553 5447 5567
rect 5533 5553 5547 5567
rect 5653 5553 5667 5567
rect 93 5533 107 5547
rect 413 5533 427 5547
rect 473 5533 487 5547
rect 513 5533 527 5547
rect 173 5513 187 5527
rect 253 5513 267 5527
rect 613 5513 627 5527
rect 773 5513 787 5527
rect 1313 5533 1327 5547
rect 1353 5533 1367 5547
rect 1453 5533 1467 5547
rect 1493 5533 1507 5547
rect 1753 5533 1767 5547
rect 1793 5533 1807 5547
rect 2113 5533 2127 5547
rect 2153 5533 2167 5547
rect 493 5493 507 5507
rect 993 5493 1007 5507
rect 1173 5493 1187 5507
rect 1353 5493 1367 5507
rect 1453 5493 1467 5507
rect 1533 5493 1547 5507
rect 33 5473 47 5487
rect 313 5473 327 5487
rect 853 5473 867 5487
rect 1213 5473 1227 5487
rect 1373 5473 1387 5487
rect 1473 5473 1487 5487
rect 2173 5513 2187 5527
rect 2213 5513 2227 5527
rect 2493 5513 2507 5527
rect 2613 5513 2627 5527
rect 2773 5533 2787 5547
rect 2853 5533 2867 5547
rect 3033 5533 3047 5547
rect 3073 5533 3087 5547
rect 3153 5533 3167 5547
rect 3913 5533 3927 5547
rect 3333 5513 3347 5527
rect 3493 5513 3507 5527
rect 3574 5513 3588 5527
rect 3653 5513 3667 5527
rect 3873 5513 3887 5527
rect 5833 5552 5847 5566
rect 5953 5553 5967 5567
rect 4513 5533 4527 5547
rect 4833 5533 4847 5547
rect 4953 5533 4967 5547
rect 1633 5493 1647 5507
rect 1793 5493 1807 5507
rect 1953 5493 1967 5507
rect 2153 5493 2167 5507
rect 2193 5493 2207 5507
rect 2573 5493 2587 5507
rect 2653 5493 2667 5507
rect 2753 5493 2767 5507
rect 3033 5493 3047 5507
rect 3133 5493 3147 5507
rect 3373 5493 3387 5507
rect 3853 5493 3867 5507
rect 4213 5513 4227 5527
rect 4333 5513 4347 5527
rect 4453 5513 4467 5527
rect 4773 5513 4787 5527
rect 5092 5513 5106 5527
rect 5273 5533 5287 5547
rect 5573 5533 5587 5547
rect 5613 5533 5627 5547
rect 5713 5533 5727 5547
rect 6073 5533 6087 5547
rect 4393 5493 4407 5507
rect 4673 5493 4687 5507
rect 4713 5493 4727 5507
rect 4753 5493 4767 5507
rect 4833 5493 4847 5507
rect 4914 5494 4928 5508
rect 5233 5513 5247 5527
rect 5433 5513 5447 5527
rect 5773 5513 5787 5527
rect 5893 5513 5907 5527
rect 6013 5513 6027 5527
rect 4973 5493 4987 5507
rect 5033 5493 5047 5507
rect 5113 5493 5127 5507
rect 1593 5473 1607 5487
rect 1813 5473 1827 5487
rect 1993 5473 2007 5487
rect 2033 5473 2047 5487
rect 2973 5473 2987 5487
rect 3153 5473 3167 5487
rect 3213 5473 3227 5487
rect 3293 5473 3307 5487
rect 3533 5473 3547 5487
rect 3693 5473 3707 5487
rect 3753 5473 3767 5487
rect 4653 5473 4667 5487
rect 4693 5473 4707 5487
rect 4913 5472 4927 5486
rect 4953 5473 4967 5487
rect 1293 5453 1307 5467
rect 1753 5453 1767 5467
rect 2073 5453 2087 5467
rect 2273 5453 2287 5467
rect 2473 5453 2487 5467
rect 93 5433 107 5447
rect 313 5433 327 5447
rect 653 5433 667 5447
rect 753 5433 767 5447
rect 793 5434 807 5448
rect 1413 5433 1427 5447
rect 1733 5433 1747 5447
rect 1873 5433 1887 5447
rect 1913 5433 1927 5447
rect 1973 5433 1987 5447
rect 2133 5433 2147 5447
rect 2353 5434 2367 5448
rect 2892 5453 2906 5467
rect 2914 5453 2928 5467
rect 2993 5453 3007 5467
rect 3033 5453 3047 5467
rect 3193 5453 3207 5467
rect 3333 5453 3347 5467
rect 3493 5453 3507 5467
rect 3593 5453 3607 5467
rect 3733 5453 3747 5467
rect 3853 5454 3867 5468
rect 5453 5493 5467 5507
rect 5493 5493 5507 5507
rect 5573 5493 5587 5507
rect 5613 5493 5627 5507
rect 5673 5493 5687 5507
rect 6073 5493 6087 5507
rect 5433 5473 5447 5487
rect 5693 5473 5707 5487
rect 4053 5453 4067 5467
rect 4413 5453 4427 5467
rect 4513 5453 4527 5467
rect 5193 5453 5207 5467
rect 5233 5453 5247 5467
rect 5333 5453 5347 5467
rect 5373 5453 5387 5467
rect 5773 5453 5787 5467
rect 5953 5453 5967 5467
rect 5993 5453 6007 5467
rect 133 5413 147 5427
rect 413 5413 427 5427
rect 473 5413 487 5427
rect 553 5413 567 5427
rect 793 5412 807 5426
rect 1053 5413 1067 5427
rect 1193 5413 1207 5427
rect 1513 5413 1527 5427
rect 2353 5412 2367 5426
rect 2393 5413 2407 5427
rect 2473 5413 2487 5427
rect 3092 5433 3106 5447
rect 3153 5433 3167 5447
rect 3413 5433 3427 5447
rect 3453 5433 3467 5447
rect 3553 5433 3567 5447
rect 3673 5433 3687 5447
rect 3813 5433 3827 5447
rect 3853 5432 3867 5446
rect 4153 5433 4167 5447
rect 4373 5433 4387 5447
rect 4473 5433 4487 5447
rect 4733 5433 4747 5447
rect 4793 5433 4807 5447
rect 5313 5433 5327 5447
rect 5353 5433 5367 5447
rect 5513 5433 5527 5447
rect 5712 5433 5726 5447
rect 5833 5433 5847 5447
rect 5933 5433 5947 5447
rect 1373 5393 1387 5407
rect 2453 5393 2467 5407
rect 2493 5393 2507 5407
rect 2753 5413 2767 5427
rect 3013 5393 3027 5407
rect 3173 5413 3187 5427
rect 3293 5414 3307 5428
rect 3213 5393 3227 5407
rect 3293 5392 3307 5406
rect 3333 5393 3347 5407
rect 3373 5393 3387 5407
rect 3773 5413 3787 5427
rect 3913 5413 3927 5427
rect 4013 5413 4027 5427
rect 4072 5413 4086 5427
rect 4173 5413 4187 5427
rect 4313 5413 4327 5427
rect 4613 5413 4627 5427
rect 4653 5413 4667 5427
rect 4993 5413 5007 5427
rect 5053 5413 5067 5427
rect 5493 5413 5507 5427
rect 5593 5413 5607 5427
rect 5913 5413 5927 5427
rect 5993 5413 6007 5427
rect 3673 5393 3687 5407
rect 3713 5393 3727 5407
rect 4193 5393 4207 5407
rect 4513 5393 4527 5407
rect 4553 5393 4567 5407
rect 4693 5393 4707 5407
rect 5773 5393 5787 5407
rect 5813 5393 5827 5407
rect 93 5373 107 5387
rect 133 5373 147 5387
rect 233 5373 247 5387
rect 313 5373 327 5387
rect 373 5373 387 5387
rect 433 5373 447 5387
rect 473 5373 487 5387
rect 613 5373 627 5387
rect 713 5373 727 5387
rect 773 5373 787 5387
rect 913 5373 927 5387
rect 993 5373 1007 5387
rect 1053 5373 1067 5387
rect 1213 5373 1227 5387
rect 1313 5373 1327 5387
rect 1473 5373 1487 5387
rect 1653 5373 1667 5387
rect 1733 5373 1747 5387
rect 1793 5373 1807 5387
rect 1973 5373 1987 5387
rect 2093 5373 2107 5387
rect 2133 5373 2147 5387
rect 2173 5373 2187 5387
rect 2273 5373 2287 5387
rect 2393 5373 2407 5387
rect 2433 5373 2447 5387
rect 2573 5373 2587 5387
rect 2853 5373 2867 5387
rect 3053 5373 3067 5387
rect 3193 5373 3207 5387
rect 3553 5373 3567 5387
rect 3853 5373 3867 5387
rect 4113 5373 4127 5387
rect 4173 5373 4187 5387
rect 4273 5373 4287 5387
rect 4333 5373 4347 5387
rect 4473 5373 4487 5387
rect 4593 5373 4607 5387
rect 4633 5373 4647 5387
rect 4773 5373 4787 5387
rect 4993 5373 5007 5387
rect 5033 5373 5047 5387
rect 5073 5373 5087 5387
rect 5113 5373 5127 5387
rect 5173 5373 5187 5387
rect 5353 5373 5367 5387
rect 5433 5373 5447 5387
rect 5473 5373 5487 5387
rect 5593 5373 5607 5387
rect 5733 5373 5747 5387
rect 5913 5373 5927 5387
rect 1273 5353 1287 5367
rect 1513 5333 1527 5347
rect 3293 5333 3307 5347
rect 3313 5333 3327 5347
rect 3393 5333 3407 5347
rect 3573 5333 3587 5347
rect 3653 5333 3667 5347
rect 3733 5333 3747 5347
rect 3953 5333 3967 5347
rect 4233 5334 4247 5348
rect 4553 5333 4567 5347
rect 4653 5333 4667 5347
rect 5292 5333 5306 5347
rect 5973 5333 5987 5347
rect 6033 5333 6047 5347
rect 113 5313 127 5327
rect 153 5313 167 5327
rect 253 5313 267 5327
rect 293 5313 307 5327
rect 413 5313 427 5327
rect 453 5313 467 5327
rect 593 5313 607 5327
rect 633 5313 647 5327
rect 673 5313 687 5327
rect 753 5313 767 5327
rect 793 5313 807 5327
rect 1013 5313 1027 5327
rect 1053 5313 1067 5327
rect 1193 5313 1207 5327
rect 1313 5313 1327 5327
rect 1353 5313 1367 5327
rect 1453 5313 1467 5327
rect 1393 5293 1407 5307
rect 1753 5313 1767 5327
rect 1813 5313 1827 5327
rect 1913 5313 1927 5327
rect 1953 5313 1967 5327
rect 2073 5313 2087 5327
rect 2113 5313 2127 5327
rect 2253 5313 2267 5327
rect 2293 5313 2307 5327
rect 2413 5313 2427 5327
rect 2453 5313 2467 5327
rect 2493 5313 2507 5327
rect 2553 5313 2567 5327
rect 2593 5313 2607 5327
rect 2693 5313 2707 5327
rect 2733 5313 2747 5327
rect 2873 5313 2887 5327
rect 2953 5313 2967 5327
rect 2993 5313 3007 5327
rect 3033 5313 3047 5327
rect 3173 5313 3187 5327
rect 3213 5313 3227 5327
rect 3353 5313 3367 5327
rect 3493 5313 3507 5327
rect 3533 5313 3547 5327
rect 2793 5293 2807 5307
rect 3113 5293 3127 5307
rect 3313 5294 3327 5308
rect 3553 5293 3567 5307
rect 3813 5313 3827 5327
rect 3993 5313 4007 5327
rect 4033 5313 4047 5327
rect 4153 5313 4167 5327
rect 4193 5313 4207 5327
rect 4233 5312 4247 5326
rect 4313 5313 4327 5327
rect 4353 5313 4367 5327
rect 4673 5313 4687 5327
rect 4713 5314 4727 5328
rect 4753 5313 4767 5327
rect 4793 5313 4807 5327
rect 4873 5313 4887 5327
rect 4913 5313 4927 5327
rect 5053 5313 5067 5327
rect 5093 5313 5107 5327
rect 5193 5313 5207 5327
rect 5233 5313 5247 5327
rect 5314 5313 5328 5327
rect 5393 5313 5407 5327
rect 5453 5313 5467 5327
rect 5493 5313 5507 5327
rect 5613 5313 5627 5327
rect 5653 5313 5667 5327
rect 5793 5313 5807 5327
rect 5893 5313 5907 5327
rect 5933 5313 5947 5327
rect 4633 5293 4647 5307
rect 113 5273 127 5287
rect 153 5273 167 5287
rect 373 5273 387 5287
rect 453 5273 467 5287
rect 593 5273 607 5287
rect 793 5273 807 5287
rect 1013 5273 1027 5287
rect 1313 5273 1327 5287
rect 1433 5273 1447 5287
rect 1513 5273 1527 5287
rect 1653 5273 1667 5287
rect 1813 5273 1827 5287
rect 1873 5273 1887 5287
rect 1953 5273 1967 5287
rect 2113 5273 2127 5287
rect 2173 5273 2187 5287
rect 2253 5273 2267 5287
rect 973 5253 987 5267
rect 1392 5253 1406 5267
rect 1453 5253 1467 5267
rect 1573 5253 1587 5267
rect 2833 5273 2847 5287
rect 2873 5273 2887 5287
rect 2913 5273 2927 5287
rect 2973 5273 2987 5287
rect 3033 5273 3047 5287
rect 3253 5273 3267 5287
rect 3313 5272 3327 5286
rect 3673 5273 3687 5287
rect 4253 5273 4267 5287
rect 4713 5292 4727 5306
rect 5273 5293 5287 5307
rect 5373 5293 5387 5307
rect 4913 5273 4927 5287
rect 5193 5273 5207 5287
rect 5353 5273 5367 5287
rect 5573 5273 5587 5287
rect 2393 5253 2407 5267
rect 2533 5253 2547 5267
rect 2712 5253 2726 5267
rect 2734 5253 2748 5267
rect 2774 5253 2788 5267
rect 2853 5253 2867 5267
rect 2934 5253 2948 5267
rect 3133 5253 3147 5267
rect 3613 5253 3627 5267
rect 3773 5253 3787 5267
rect 3813 5254 3827 5268
rect 4333 5253 4347 5267
rect 4553 5253 4567 5267
rect 4633 5253 4647 5267
rect 5093 5253 5107 5267
rect 5153 5253 5167 5267
rect 193 5233 207 5247
rect 613 5233 627 5247
rect 1133 5233 1147 5247
rect 1213 5233 1227 5247
rect 1332 5233 1346 5247
rect 1354 5233 1368 5247
rect 1653 5233 1667 5247
rect 1793 5233 1807 5247
rect 1854 5233 1868 5247
rect 1913 5233 1927 5247
rect 1993 5233 2007 5247
rect 2273 5233 2287 5247
rect 2493 5233 2507 5247
rect 673 5213 687 5227
rect 853 5213 867 5227
rect 913 5213 927 5227
rect 1113 5213 1127 5227
rect 1193 5213 1207 5227
rect 1393 5213 1407 5227
rect 1513 5213 1527 5227
rect 1573 5213 1587 5227
rect 2053 5213 2067 5227
rect 2293 5213 2307 5227
rect 2393 5213 2407 5227
rect 2433 5213 2447 5227
rect 2553 5233 2567 5247
rect 2693 5233 2707 5247
rect 2833 5233 2847 5247
rect 2993 5233 3007 5247
rect 3193 5233 3207 5247
rect 3233 5233 3247 5247
rect 3273 5233 3287 5247
rect 3373 5233 3387 5247
rect 3533 5233 3547 5247
rect 3573 5233 3587 5247
rect 3673 5233 3687 5247
rect 3713 5233 3727 5247
rect 3813 5232 3827 5246
rect 4473 5234 4487 5248
rect 4753 5233 4767 5247
rect 4893 5233 4907 5247
rect 713 5193 727 5207
rect 793 5193 807 5207
rect 1133 5193 1147 5207
rect 1293 5193 1307 5207
rect 1333 5193 1347 5207
rect 1413 5193 1427 5207
rect 1553 5193 1567 5207
rect 2653 5213 2667 5227
rect 2953 5213 2967 5227
rect 3053 5213 3067 5227
rect 3332 5213 3346 5227
rect 3354 5213 3368 5227
rect 3933 5213 3947 5227
rect 3993 5213 4007 5227
rect 4073 5213 4087 5227
rect 4113 5213 4127 5227
rect 4193 5213 4207 5227
rect 2553 5193 2567 5207
rect 2772 5193 2786 5207
rect 2794 5193 2808 5207
rect 2993 5193 3007 5207
rect 4413 5213 4427 5227
rect 4473 5212 4487 5226
rect 4693 5213 4707 5227
rect 4733 5213 4747 5227
rect 4853 5213 4867 5227
rect 4913 5213 4927 5227
rect 5033 5213 5047 5227
rect 5293 5233 5307 5247
rect 5453 5253 5467 5267
rect 5793 5273 5807 5287
rect 5932 5273 5946 5287
rect 5954 5273 5968 5287
rect 5933 5233 5947 5247
rect 5893 5213 5907 5227
rect 113 5173 127 5187
rect 253 5173 267 5187
rect 553 5173 567 5187
rect 1693 5173 1707 5187
rect 1873 5173 1887 5187
rect 2093 5173 2107 5187
rect 2133 5173 2147 5187
rect 2713 5173 2727 5187
rect 2893 5173 2907 5187
rect 2932 5173 2946 5187
rect 2954 5173 2968 5187
rect 4713 5193 4727 5207
rect 4833 5193 4847 5207
rect 5133 5193 5147 5207
rect 4513 5173 4527 5187
rect 5033 5173 5047 5187
rect 5273 5193 5287 5207
rect 5193 5173 5207 5187
rect 5973 5173 5987 5187
rect 573 5153 587 5167
rect 1093 5153 1107 5167
rect 1393 5153 1407 5167
rect 1453 5153 1467 5167
rect 1773 5153 1787 5167
rect 1913 5153 1927 5167
rect 2073 5153 2087 5167
rect 2353 5153 2367 5167
rect 673 5133 687 5147
rect 713 5133 727 5147
rect 833 5133 847 5147
rect 1153 5133 1167 5147
rect 1193 5133 1207 5147
rect 1232 5133 1246 5147
rect 1293 5133 1307 5147
rect 1373 5133 1387 5147
rect 1573 5133 1587 5147
rect 1713 5133 1727 5147
rect 1853 5133 1867 5147
rect 1953 5133 1967 5147
rect 2432 5153 2446 5167
rect 2454 5153 2468 5167
rect 2573 5153 2587 5167
rect 2673 5153 2687 5167
rect 3653 5153 3667 5167
rect 4073 5153 4087 5167
rect 4273 5154 4287 5168
rect 2413 5133 2427 5147
rect 2633 5133 2647 5147
rect 2733 5133 2747 5147
rect 3073 5133 3087 5147
rect 3233 5133 3247 5147
rect 3313 5133 3327 5147
rect 3352 5133 3366 5147
rect 3374 5133 3388 5147
rect 3553 5133 3567 5147
rect 3673 5133 3687 5147
rect 3733 5133 3747 5147
rect 3893 5133 3907 5147
rect 4053 5133 4067 5147
rect 4093 5133 4107 5147
rect 4273 5132 4287 5146
rect 4453 5133 4467 5147
rect 4593 5133 4607 5147
rect 4873 5153 4887 5167
rect 4933 5154 4947 5168
rect 5213 5153 5227 5167
rect 2973 5113 2987 5127
rect 3013 5113 3027 5127
rect 3433 5113 3447 5127
rect 4413 5113 4427 5127
rect 4693 5133 4707 5147
rect 4833 5133 4847 5147
rect 4933 5132 4947 5146
rect 5013 5133 5027 5147
rect 5113 5133 5127 5147
rect 5173 5133 5187 5147
rect 5233 5133 5247 5147
rect 5293 5133 5307 5147
rect 5473 5133 5487 5147
rect 6033 5133 6047 5147
rect 4673 5113 4687 5127
rect 5513 5113 5527 5127
rect 5693 5113 5707 5127
rect 5913 5113 5927 5127
rect 6073 5113 6087 5127
rect 153 5093 167 5107
rect 193 5093 207 5107
rect 233 5093 247 5107
rect 373 5093 387 5107
rect 413 5093 427 5107
rect 553 5093 567 5107
rect 593 5093 607 5107
rect 673 5093 687 5107
rect 713 5093 727 5107
rect 753 5093 767 5107
rect 833 5093 847 5107
rect 873 5093 887 5107
rect 1033 5093 1047 5107
rect 1073 5093 1087 5107
rect 1113 5093 1127 5107
rect 1193 5093 1207 5107
rect 1313 5093 1327 5107
rect 1353 5093 1367 5107
rect 1473 5093 1487 5107
rect 1513 5093 1527 5107
rect 1653 5093 1667 5107
rect 1773 5093 1787 5107
rect 1813 5093 1827 5107
rect 1873 5093 1887 5107
rect 2053 5093 2067 5107
rect 2093 5093 2107 5107
rect 2193 5093 2207 5107
rect 2233 5093 2247 5107
rect 2273 5093 2287 5107
rect 2413 5093 2427 5107
rect 2453 5093 2467 5107
rect 2573 5093 2587 5107
rect 2613 5093 2627 5107
rect 2733 5093 2747 5107
rect 2773 5093 2787 5107
rect 2853 5093 2867 5107
rect 2893 5093 2907 5107
rect 3033 5093 3047 5107
rect 3073 5093 3087 5107
rect 3173 5093 3187 5107
rect 3213 5093 3227 5107
rect 3353 5093 3367 5107
rect 3533 5093 3547 5107
rect 3573 5093 3587 5107
rect 3633 5093 3647 5107
rect 3653 5093 3667 5107
rect 3693 5093 3707 5107
rect 3773 5093 3787 5107
rect 3813 5093 3827 5107
rect 3953 5093 3967 5107
rect 3993 5093 4007 5107
rect 4113 5093 4127 5107
rect 4153 5093 4167 5107
rect 4253 5093 4267 5107
rect 4293 5093 4307 5107
rect 4353 5093 4367 5107
rect 4553 5093 4567 5107
rect 4593 5093 4607 5107
rect 4793 5093 4807 5107
rect 4833 5093 4847 5107
rect 4873 5093 4887 5107
rect 4953 5093 4967 5107
rect 5033 5093 5047 5107
rect 5113 5093 5127 5107
rect 5153 5093 5167 5107
rect 5273 5093 5287 5107
rect 5313 5093 5327 5107
rect 5393 5093 5407 5107
rect 5433 5093 5447 5107
rect 5473 5093 5487 5107
rect 5713 5093 5727 5107
rect 5753 5093 5767 5107
rect 793 5073 807 5087
rect 973 5073 987 5087
rect 2493 5073 2507 5087
rect 2533 5073 2547 5087
rect 4473 5073 4487 5087
rect 5973 5074 5987 5088
rect 6073 5073 6087 5087
rect 1093 5053 1107 5067
rect 2633 5054 2647 5068
rect 3113 5053 3127 5067
rect 5973 5052 5987 5066
rect 113 5033 127 5047
rect 213 5033 227 5047
rect 253 5033 267 5047
rect 293 5033 307 5047
rect 433 5033 447 5047
rect 493 5033 507 5047
rect 573 5033 587 5047
rect 613 5033 627 5047
rect 733 5033 747 5047
rect 813 5033 827 5047
rect 853 5033 867 5047
rect 933 5033 947 5047
rect 1053 5033 1067 5047
rect 1113 5033 1127 5047
rect 1213 5033 1227 5047
rect 1253 5033 1267 5047
rect 1413 5033 1427 5047
rect 1533 5033 1547 5047
rect 1633 5033 1647 5047
rect 1753 5033 1767 5047
rect 1793 5033 1807 5047
rect 1913 5033 1927 5047
rect 1993 5033 2007 5047
rect 2073 5033 2087 5047
rect 2113 5033 2127 5047
rect 2193 5033 2207 5047
rect 2433 5033 2447 5047
rect 2593 5033 2607 5047
rect 2633 5033 2647 5047
rect 2753 5033 2767 5047
rect 2873 5033 2887 5047
rect 2933 5033 2947 5047
rect 3013 5033 3027 5047
rect 3072 5033 3086 5047
rect 3094 5033 3108 5047
rect 3153 5033 3167 5047
rect 3193 5033 3207 5047
rect 3273 5033 3287 5047
rect 3513 5033 3527 5047
rect 3593 5033 3607 5047
rect 3673 5033 3687 5047
rect 3793 5033 3807 5047
rect 3852 5033 3866 5047
rect 3874 5033 3888 5047
rect 4093 5033 4107 5047
rect 4233 5033 4247 5047
rect 4273 5033 4287 5047
rect 4313 5033 4327 5047
rect 4533 5033 4547 5047
rect 4613 5033 4627 5047
rect 4653 5033 4667 5047
rect 4753 5033 4767 5047
rect 4853 5033 4867 5047
rect 4993 5033 5007 5047
rect 5053 5033 5067 5047
rect 5253 5033 5267 5047
rect 5413 5033 5427 5047
rect 5492 5033 5506 5047
rect 5693 5033 5707 5047
rect 5773 5033 5787 5047
rect 893 5013 907 5027
rect 1013 5013 1027 5027
rect 1073 5013 1087 5027
rect 2293 5013 2307 5027
rect 2393 5013 2407 5027
rect 2613 5013 2627 5027
rect 2773 5013 2787 5027
rect 3114 5013 3128 5027
rect 3313 5013 3327 5027
rect 3413 5013 3427 5027
rect 3693 5013 3707 5027
rect 4013 5013 4027 5027
rect 213 4993 227 5007
rect 293 4993 307 5007
rect 393 4993 407 5007
rect 653 4993 667 5007
rect 753 4993 767 5007
rect 873 4993 887 5007
rect 1033 4993 1047 5007
rect 1473 4993 1487 5007
rect 1653 4993 1667 5007
rect 1713 4993 1727 5007
rect 573 4973 587 4987
rect 713 4973 727 4987
rect 793 4973 807 4987
rect 1053 4973 1067 4987
rect 1093 4973 1107 4987
rect 1193 4973 1207 4987
rect 1373 4973 1387 4987
rect 2373 4993 2387 5007
rect 3193 4993 3207 5007
rect 3233 4993 3247 5007
rect 3633 4993 3647 5007
rect 3793 4993 3807 5007
rect 113 4953 127 4967
rect 173 4953 187 4967
rect 373 4953 387 4967
rect 553 4953 567 4967
rect 613 4953 627 4967
rect 653 4953 667 4967
rect 893 4953 907 4967
rect 1313 4953 1327 4967
rect 1493 4953 1507 4967
rect 1773 4973 1787 4987
rect 2013 4973 2027 4987
rect 2133 4973 2147 4987
rect 2313 4973 2327 4987
rect 2673 4973 2687 4987
rect 2713 4973 2727 4987
rect 2753 4973 2767 4987
rect 2793 4973 2807 4987
rect 2893 4973 2907 4987
rect 3013 4973 3027 4987
rect 3213 4973 3227 4987
rect 3352 4973 3366 4987
rect 3374 4973 3388 4987
rect 3653 4973 3667 4987
rect 3892 4993 3906 5007
rect 3914 4993 3928 5007
rect 4113 4993 4127 5007
rect 4153 4993 4167 5007
rect 4292 4993 4306 5007
rect 4314 4993 4328 5007
rect 4393 5013 4407 5027
rect 4433 5013 4447 5027
rect 4533 4994 4547 5008
rect 4593 4993 4607 5007
rect 3853 4973 3867 4987
rect 3973 4973 3987 4987
rect 4273 4973 4287 4987
rect 4433 4973 4447 4987
rect 4533 4972 4547 4986
rect 4573 4973 4587 4987
rect 4853 4993 4867 5007
rect 4893 4993 4907 5007
rect 5993 5013 6007 5027
rect 6033 5013 6047 5027
rect 4793 4973 4807 4987
rect 5033 4973 5047 4987
rect 5073 4973 5087 4987
rect 5133 4973 5147 4987
rect 5193 4973 5207 4987
rect 5433 4973 5447 4987
rect 5473 4973 5487 4987
rect 5673 4973 5687 4987
rect 5873 4973 5887 4987
rect 5993 4973 6007 4987
rect 6033 4973 6047 4987
rect 1633 4953 1647 4967
rect 2053 4953 2067 4967
rect 93 4933 107 4947
rect 193 4933 207 4947
rect 473 4933 487 4947
rect 593 4933 607 4947
rect 833 4933 847 4947
rect 1113 4933 1127 4947
rect 1673 4933 1687 4947
rect 1873 4933 1887 4947
rect 1933 4933 1947 4947
rect 2513 4953 2527 4967
rect 2633 4953 2647 4967
rect 2913 4953 2927 4967
rect 2953 4953 2967 4967
rect 3433 4953 3447 4967
rect 3753 4953 3767 4967
rect 3793 4953 3807 4967
rect 2233 4933 2247 4947
rect 2393 4933 2407 4947
rect 2573 4933 2587 4947
rect 2872 4933 2886 4947
rect 2894 4933 2908 4947
rect 3373 4933 3387 4947
rect 3413 4933 3427 4947
rect 4332 4953 4346 4967
rect 4354 4953 4368 4967
rect 3933 4933 3947 4947
rect 4133 4933 4147 4947
rect 4513 4933 4527 4947
rect 4792 4934 4806 4948
rect 4814 4933 4828 4947
rect 4873 4933 4887 4947
rect 4913 4953 4927 4967
rect 5053 4953 5067 4967
rect 5653 4953 5667 4967
rect 4953 4933 4967 4947
rect 5153 4933 5167 4947
rect 5253 4933 5267 4947
rect 13 4913 27 4927
rect 253 4913 267 4927
rect 413 4913 427 4927
rect 533 4913 547 4927
rect 653 4913 667 4927
rect 1173 4913 1187 4927
rect 1273 4913 1287 4927
rect 1312 4913 1326 4927
rect 1334 4913 1348 4927
rect 1433 4913 1447 4927
rect 1713 4913 1727 4927
rect 1813 4913 1827 4927
rect 2292 4913 2306 4927
rect 2314 4913 2328 4927
rect 2653 4913 2667 4927
rect 2713 4913 2727 4927
rect 2853 4913 2867 4927
rect 53 4893 67 4907
rect 273 4893 287 4907
rect 313 4893 327 4907
rect 373 4893 387 4907
rect 753 4893 767 4907
rect 413 4873 427 4887
rect 493 4873 507 4887
rect 853 4893 867 4907
rect 1053 4893 1067 4907
rect 1193 4893 1207 4907
rect 1393 4893 1407 4907
rect 1732 4893 1746 4907
rect 1754 4893 1768 4907
rect 1173 4873 1187 4887
rect 1273 4873 1287 4887
rect 1313 4873 1327 4887
rect 1873 4893 1887 4907
rect 1993 4893 2007 4907
rect 2114 4893 2128 4907
rect 2213 4893 2227 4907
rect 2953 4893 2967 4907
rect 3033 4893 3047 4907
rect 3113 4893 3127 4907
rect 3153 4913 3167 4927
rect 3453 4913 3467 4927
rect 4233 4913 4247 4927
rect 4313 4913 4327 4927
rect 4373 4913 4387 4927
rect 4673 4913 4687 4927
rect 4794 4912 4808 4926
rect 4832 4913 4846 4927
rect 4854 4913 4868 4927
rect 4993 4913 5007 4927
rect 5393 4933 5407 4947
rect 5933 4933 5947 4947
rect 6033 4933 6047 4947
rect 5433 4913 5447 4927
rect 5953 4913 5967 4927
rect 5993 4913 6007 4927
rect 3233 4893 3247 4907
rect 3293 4893 3307 4907
rect 2573 4873 2587 4887
rect 2753 4873 2767 4887
rect 3513 4893 3527 4907
rect 4012 4893 4026 4907
rect 4053 4893 4067 4907
rect 4413 4893 4427 4907
rect 4493 4893 4507 4907
rect 4553 4893 4567 4907
rect 4713 4893 4727 4907
rect 4973 4893 4987 4907
rect 5093 4893 5107 4907
rect 5133 4893 5147 4907
rect 5353 4893 5367 4907
rect 5413 4893 5427 4907
rect 5513 4893 5527 4907
rect 5673 4893 5687 4907
rect 5733 4893 5747 4907
rect 5913 4893 5927 4907
rect 4333 4873 4347 4887
rect 4373 4873 4387 4887
rect 4833 4873 4847 4887
rect 4873 4873 4887 4887
rect 5933 4873 5947 4887
rect 113 4853 127 4867
rect 193 4853 207 4867
rect 373 4853 387 4867
rect 473 4853 487 4867
rect 553 4853 567 4867
rect 713 4853 727 4867
rect 793 4853 807 4867
rect 953 4853 967 4867
rect 1133 4853 1147 4867
rect 1413 4853 1427 4867
rect 1453 4853 1467 4867
rect 1693 4853 1707 4867
rect 1753 4853 1767 4867
rect 2053 4853 2067 4867
rect 2293 4853 2307 4867
rect 2453 4853 2467 4867
rect 2493 4853 2507 4867
rect 2593 4853 2607 4867
rect 2633 4853 2647 4867
rect 2873 4853 2887 4867
rect 3033 4853 3047 4867
rect 3133 4853 3147 4867
rect 3173 4853 3187 4867
rect 3253 4853 3267 4867
rect 3653 4853 3667 4867
rect 3793 4853 3807 4867
rect 3993 4853 4007 4867
rect 4033 4853 4047 4867
rect 4073 4853 4087 4867
rect 4353 4853 4367 4867
rect 4413 4853 4427 4867
rect 4453 4853 4467 4867
rect 4633 4853 4647 4867
rect 4673 4853 4687 4867
rect 4713 4853 4727 4867
rect 4973 4853 4987 4867
rect 2193 4833 2207 4847
rect 2533 4833 2547 4847
rect 5053 4833 5067 4847
rect 5293 4853 5307 4867
rect 5433 4853 5447 4867
rect 5533 4853 5547 4867
rect 5573 4853 5587 4867
rect 5793 4853 5807 4867
rect 5913 4853 5927 4867
rect 5953 4853 5967 4867
rect 5993 4853 6007 4867
rect 5193 4833 5207 4847
rect 2413 4813 2427 4827
rect 2473 4813 2487 4827
rect 3533 4813 3547 4827
rect 3693 4813 3707 4827
rect 3833 4813 3847 4827
rect 3893 4813 3907 4827
rect 5753 4813 5767 4827
rect 6013 4813 6027 4827
rect 6054 4813 6068 4827
rect 213 4793 227 4807
rect 253 4793 267 4807
rect 353 4793 367 4807
rect 393 4793 407 4807
rect 433 4793 447 4807
rect 653 4793 667 4807
rect 693 4793 707 4807
rect 813 4793 827 4807
rect 853 4793 867 4807
rect 973 4793 987 4807
rect 1013 4793 1027 4807
rect 1113 4793 1127 4807
rect 1153 4793 1167 4807
rect 713 4773 727 4787
rect 1253 4773 1267 4787
rect 1533 4793 1547 4807
rect 1573 4793 1587 4807
rect 1693 4793 1707 4807
rect 1733 4793 1747 4807
rect 1833 4793 1847 4807
rect 1873 4793 1887 4807
rect 1993 4793 2007 4807
rect 2033 4793 2047 4807
rect 2133 4793 2147 4807
rect 2173 4793 2187 4807
rect 2273 4793 2287 4807
rect 2313 4793 2327 4807
rect 2373 4793 2387 4807
rect 2573 4793 2587 4807
rect 2613 4793 2627 4807
rect 2653 4793 2667 4807
rect 2773 4793 2787 4807
rect 2813 4793 2827 4807
rect 3013 4793 3027 4807
rect 3153 4793 3167 4807
rect 3193 4793 3207 4807
rect 3293 4793 3307 4807
rect 3333 4793 3347 4807
rect 3453 4793 3467 4807
rect 3493 4793 3507 4807
rect 1653 4773 1667 4787
rect 2353 4773 2367 4787
rect 2413 4773 2427 4787
rect 2453 4773 2467 4787
rect 2493 4773 2507 4787
rect 3933 4793 3947 4807
rect 3973 4793 3987 4807
rect 4053 4793 4067 4807
rect 4093 4793 4107 4807
rect 4133 4793 4147 4807
rect 4253 4793 4267 4807
rect 4293 4793 4307 4807
rect 4353 4793 4367 4807
rect 4433 4793 4447 4807
rect 4553 4793 4567 4807
rect 4593 4793 4607 4807
rect 4653 4793 4667 4807
rect 4693 4793 4707 4807
rect 4733 4793 4747 4807
rect 4993 4793 5007 4807
rect 5033 4793 5047 4807
rect 5133 4793 5147 4807
rect 5173 4793 5187 4807
rect 5273 4793 5287 4807
rect 5313 4793 5327 4807
rect 5453 4793 5467 4807
rect 5533 4793 5547 4807
rect 5633 4793 5647 4807
rect 5793 4793 5807 4807
rect 5833 4793 5847 4807
rect 5933 4793 5947 4807
rect 5973 4793 5987 4807
rect 213 4753 227 4767
rect 273 4753 287 4767
rect 353 4753 367 4767
rect 433 4753 447 4767
rect 233 4733 247 4747
rect 313 4733 327 4747
rect 813 4733 827 4747
rect 1153 4733 1167 4747
rect 1234 4733 1248 4747
rect 1393 4733 1407 4747
rect 1533 4753 1547 4767
rect 1812 4753 1826 4767
rect 1834 4753 1848 4767
rect 2173 4753 2187 4767
rect 2313 4753 2327 4767
rect 2613 4753 2627 4767
rect 2773 4753 2787 4767
rect 2813 4753 2827 4767
rect 2913 4753 2927 4767
rect 3113 4753 3127 4767
rect 1733 4733 1747 4747
rect 1933 4733 1947 4747
rect 2033 4733 2047 4747
rect 2333 4733 2347 4747
rect 373 4713 387 4727
rect 713 4713 727 4727
rect 1113 4713 1127 4727
rect 1773 4713 1787 4727
rect 2013 4713 2027 4727
rect 2133 4713 2147 4727
rect 2253 4713 2267 4727
rect 3033 4733 3047 4747
rect 3313 4753 3327 4767
rect 3493 4754 3507 4768
rect 4773 4773 4787 4787
rect 4933 4773 4947 4787
rect 6053 4773 6067 4787
rect 3673 4753 3687 4767
rect 3793 4753 3807 4767
rect 4053 4753 4067 4767
rect 4093 4753 4107 4767
rect 4413 4753 4427 4767
rect 4553 4753 4567 4767
rect 4693 4753 4707 4767
rect 4833 4753 4847 4767
rect 4873 4754 4887 4768
rect 5033 4753 5047 4767
rect 3153 4734 3167 4748
rect 3273 4733 3287 4747
rect 3333 4733 3347 4747
rect 3373 4733 3387 4747
rect 3493 4732 3507 4746
rect 3733 4733 3747 4747
rect 3853 4733 3867 4747
rect 3933 4733 3947 4747
rect 4073 4733 4087 4747
rect 4173 4733 4187 4747
rect 4253 4733 4267 4747
rect 4333 4733 4347 4747
rect 4473 4733 4487 4747
rect 4593 4733 4607 4747
rect 4633 4733 4647 4747
rect 4733 4733 4747 4747
rect 2373 4713 2387 4727
rect 2613 4713 2627 4727
rect 2833 4713 2847 4727
rect 2933 4713 2947 4727
rect 3153 4712 3167 4726
rect 3193 4713 3207 4727
rect 673 4693 687 4707
rect 933 4693 947 4707
rect 1013 4693 1027 4707
rect 913 4673 927 4687
rect 1053 4673 1067 4687
rect 1113 4673 1127 4687
rect 1253 4673 1267 4687
rect 1413 4693 1427 4707
rect 1573 4693 1587 4707
rect 1693 4693 1707 4707
rect 1593 4673 1607 4687
rect 1633 4673 1647 4687
rect 1873 4693 1887 4707
rect 1953 4693 1967 4707
rect 2033 4693 2047 4707
rect 2653 4693 2667 4707
rect 2693 4693 2707 4707
rect 2732 4693 2746 4707
rect 2754 4693 2768 4707
rect 3073 4693 3087 4707
rect 3213 4693 3227 4707
rect 3293 4693 3307 4707
rect 3353 4693 3367 4707
rect 3433 4693 3447 4707
rect 3473 4713 3487 4727
rect 3633 4713 3647 4727
rect 3952 4713 3966 4727
rect 3974 4713 3988 4727
rect 4132 4713 4146 4727
rect 4154 4713 4168 4727
rect 4213 4713 4227 4727
rect 4293 4713 4307 4727
rect 4873 4732 4887 4746
rect 4993 4733 5007 4747
rect 5053 4733 5067 4747
rect 5373 4753 5387 4767
rect 5513 4753 5527 4767
rect 5793 4753 5807 4767
rect 5933 4753 5947 4767
rect 5113 4733 5127 4747
rect 5573 4733 5587 4747
rect 5633 4733 5647 4747
rect 4493 4713 4507 4727
rect 4713 4713 4727 4727
rect 4853 4713 4867 4727
rect 4953 4713 4967 4727
rect 5033 4713 5047 4727
rect 5253 4713 5267 4727
rect 5313 4713 5327 4727
rect 5753 4713 5767 4727
rect 6054 4713 6068 4727
rect 393 4653 407 4667
rect 753 4653 767 4667
rect 853 4653 867 4667
rect 953 4653 967 4667
rect 1433 4653 1447 4667
rect 1793 4653 1807 4667
rect 2073 4673 2087 4687
rect 2392 4673 2406 4687
rect 2414 4674 2428 4688
rect 2593 4673 2607 4687
rect 2673 4673 2687 4687
rect 3373 4673 3387 4687
rect 3533 4673 3547 4687
rect 3613 4693 3627 4707
rect 3793 4693 3807 4707
rect 4193 4693 4207 4707
rect 4513 4693 4527 4707
rect 4573 4693 4587 4707
rect 4912 4694 4926 4708
rect 4934 4693 4948 4707
rect 5113 4693 5127 4707
rect 3913 4673 3927 4687
rect 4553 4673 4567 4687
rect 4713 4673 4727 4687
rect 4913 4672 4927 4686
rect 5233 4693 5247 4707
rect 5273 4693 5287 4707
rect 5333 4693 5347 4707
rect 5433 4693 5447 4707
rect 5473 4693 5487 4707
rect 5613 4693 5627 4707
rect 5153 4673 5167 4687
rect 5413 4673 5427 4687
rect 5493 4673 5507 4687
rect 5853 4673 5867 4687
rect 5973 4673 5987 4687
rect 6053 4673 6067 4687
rect 1973 4653 1987 4667
rect 2053 4653 2067 4667
rect 2193 4653 2207 4667
rect 2314 4653 2328 4667
rect 2413 4652 2427 4666
rect 2473 4653 2487 4667
rect 2513 4653 2527 4667
rect 2933 4653 2947 4667
rect 3033 4653 3047 4667
rect 113 4633 127 4647
rect 433 4633 447 4647
rect 593 4633 607 4647
rect 634 4633 648 4647
rect 1172 4633 1186 4647
rect 1194 4633 1208 4647
rect 1273 4633 1287 4647
rect 1373 4633 1387 4647
rect 1593 4633 1607 4647
rect 1673 4633 1687 4647
rect 1773 4633 1787 4647
rect 1853 4633 1867 4647
rect 2073 4633 2087 4647
rect 2274 4633 2288 4647
rect 2493 4633 2507 4647
rect 2533 4633 2547 4647
rect 2733 4633 2747 4647
rect 193 4613 207 4627
rect 253 4613 267 4627
rect 573 4613 587 4627
rect 793 4613 807 4627
rect 993 4613 1007 4627
rect 1153 4613 1167 4627
rect 1333 4613 1347 4627
rect 1493 4613 1507 4627
rect 2373 4613 2387 4627
rect 2712 4613 2726 4627
rect 2873 4633 2887 4647
rect 3313 4653 3327 4667
rect 3073 4633 3087 4647
rect 3472 4653 3486 4667
rect 3494 4653 3508 4667
rect 3553 4653 3567 4667
rect 3693 4653 3707 4667
rect 3733 4653 3747 4667
rect 4153 4653 4167 4667
rect 4293 4653 4307 4667
rect 4333 4653 4347 4667
rect 4394 4654 4408 4668
rect 4833 4653 4847 4667
rect 5053 4653 5067 4667
rect 5093 4653 5107 4667
rect 5373 4653 5387 4667
rect 5753 4653 5767 4667
rect 5813 4653 5827 4667
rect 5913 4653 5927 4667
rect 6073 4653 6087 4667
rect 3213 4613 3227 4627
rect 3913 4633 3927 4647
rect 4013 4633 4027 4647
rect 4173 4633 4187 4647
rect 4773 4633 4787 4647
rect 4813 4633 4827 4647
rect 4953 4633 4967 4647
rect 5033 4633 5047 4647
rect 5073 4633 5087 4647
rect 5393 4633 5407 4647
rect 5873 4633 5887 4647
rect 3413 4613 3427 4627
rect 3473 4613 3487 4627
rect 3533 4613 3547 4627
rect 3673 4613 3687 4627
rect 3753 4613 3767 4627
rect 4033 4613 4047 4627
rect 4072 4613 4086 4627
rect 4094 4613 4108 4627
rect 4353 4613 4367 4627
rect 4392 4613 4406 4627
rect 4414 4613 4428 4627
rect 4873 4613 4887 4627
rect 4993 4613 5007 4627
rect 5053 4613 5067 4627
rect 2093 4593 2107 4607
rect 2153 4593 2167 4607
rect 2293 4593 2307 4607
rect 2613 4593 2627 4607
rect 2933 4593 2947 4607
rect 4533 4593 4547 4607
rect 4613 4593 4627 4607
rect 4733 4593 4747 4607
rect 5233 4613 5247 4627
rect 5293 4613 5307 4627
rect 5893 4613 5907 4627
rect 6033 4613 6047 4627
rect 6073 4613 6087 4627
rect 5733 4593 5747 4607
rect 233 4573 247 4587
rect 273 4573 287 4587
rect 393 4573 407 4587
rect 433 4573 447 4587
rect 633 4573 647 4587
rect 673 4573 687 4587
rect 713 4573 727 4587
rect 813 4573 827 4587
rect 853 4573 867 4587
rect 993 4573 1007 4587
rect 1153 4573 1167 4587
rect 1193 4573 1207 4587
rect 1293 4573 1307 4587
rect 1333 4573 1347 4587
rect 1453 4573 1467 4587
rect 1493 4573 1507 4587
rect 1633 4573 1647 4587
rect 1813 4573 1827 4587
rect 1853 4573 1867 4587
rect 1893 4573 1907 4587
rect 2013 4573 2027 4587
rect 2053 4573 2067 4587
rect 2193 4573 2207 4587
rect 2233 4573 2247 4587
rect 2273 4573 2287 4587
rect 2333 4573 2347 4587
rect 2413 4573 2427 4587
rect 2473 4573 2487 4587
rect 2513 4573 2527 4587
rect 2673 4573 2687 4587
rect 2733 4573 2747 4587
rect 3033 4573 3047 4587
rect 3073 4573 3087 4587
rect 3233 4573 3247 4587
rect 3353 4573 3367 4587
rect 3473 4573 3487 4587
rect 3593 4573 3607 4587
rect 3633 4573 3647 4587
rect 3673 4573 3687 4587
rect 3713 4573 3727 4587
rect 3753 4573 3767 4587
rect 3833 4573 3847 4587
rect 3873 4573 3887 4587
rect 3913 4573 3927 4587
rect 4033 4573 4047 4587
rect 4113 4573 4127 4587
rect 4153 4573 4167 4587
rect 4193 4573 4207 4587
rect 4313 4573 4327 4587
rect 4353 4573 4367 4587
rect 4453 4573 4467 4587
rect 4493 4573 4507 4587
rect 4753 4573 4767 4587
rect 4793 4573 4807 4587
rect 4913 4573 4927 4587
rect 4953 4573 4967 4587
rect 5053 4573 5067 4587
rect 5093 4573 5107 4587
rect 5193 4573 5207 4587
rect 5233 4573 5247 4587
rect 5353 4573 5367 4587
rect 5393 4573 5407 4587
rect 5493 4573 5507 4587
rect 5533 4573 5547 4587
rect 5673 4573 5687 4587
rect 5713 4573 5727 4587
rect 5833 4573 5847 4587
rect 5873 4573 5887 4587
rect 953 4553 967 4567
rect 1033 4553 1047 4567
rect 1093 4553 1107 4567
rect 2833 4553 2847 4567
rect 4693 4553 4707 4567
rect 4873 4553 4887 4567
rect 1673 4533 1687 4547
rect 1733 4533 1747 4547
rect 2253 4533 2267 4547
rect 2313 4533 2327 4547
rect 3533 4533 3547 4547
rect 4973 4533 4987 4547
rect 5893 4533 5907 4547
rect 6013 4533 6027 4547
rect 6053 4533 6067 4547
rect 113 4513 127 4527
rect 253 4513 267 4527
rect 293 4513 307 4527
rect 413 4513 427 4527
rect 553 4513 567 4527
rect 693 4513 707 4527
rect 793 4513 807 4527
rect 1053 4513 1067 4527
rect 1133 4513 1147 4527
rect 1273 4513 1287 4527
rect 1353 4513 1367 4527
rect 1433 4513 1447 4527
rect 1573 4513 1587 4527
rect 1613 4513 1627 4527
rect 1773 4513 1787 4527
rect 1873 4513 1887 4527
rect 2033 4513 2047 4527
rect 2073 4513 2087 4527
rect 2393 4513 2407 4527
rect 2813 4513 2827 4527
rect 2853 4514 2867 4528
rect 3013 4514 3027 4528
rect 3053 4513 3067 4527
rect 3133 4513 3147 4527
rect 3213 4513 3227 4527
rect 3333 4513 3347 4527
rect 3453 4513 3467 4527
rect 3613 4513 3627 4527
rect 3733 4513 3747 4527
rect 3853 4513 3867 4527
rect 3893 4513 3907 4527
rect 4053 4513 4067 4527
rect 4293 4513 4307 4527
rect 4393 4514 4407 4528
rect 4733 4513 4747 4527
rect 5033 4513 5047 4527
rect 5113 4513 5127 4527
rect 5213 4513 5227 4527
rect 5293 4513 5307 4527
rect 5333 4513 5347 4527
rect 5473 4513 5487 4527
rect 5513 4513 5527 4527
rect 5733 4513 5747 4527
rect 5813 4513 5827 4527
rect 5973 4513 5987 4527
rect 213 4493 227 4507
rect 253 4473 267 4487
rect 473 4473 487 4487
rect 713 4473 727 4487
rect 753 4473 767 4487
rect 973 4493 987 4507
rect 1013 4493 1027 4507
rect 2173 4493 2187 4507
rect 1153 4473 1167 4487
rect 1233 4473 1247 4487
rect 1293 4473 1307 4487
rect 1353 4473 1367 4487
rect 1433 4473 1447 4487
rect 1573 4473 1587 4487
rect 1813 4473 1827 4487
rect 2013 4473 2027 4487
rect 2053 4473 2067 4487
rect 2533 4493 2547 4507
rect 2573 4493 2587 4507
rect 2613 4493 2627 4507
rect 2853 4492 2867 4506
rect 2953 4493 2967 4507
rect 3013 4492 3027 4506
rect 3093 4493 3107 4507
rect 3573 4493 3587 4507
rect 3773 4493 3787 4507
rect 3933 4493 3947 4507
rect 4173 4493 4187 4507
rect 4333 4493 4347 4507
rect 4393 4492 4407 4506
rect 4613 4493 4627 4507
rect 4653 4493 4667 4507
rect 5073 4493 5087 4507
rect 5693 4493 5707 4507
rect 5853 4493 5867 4507
rect 2273 4473 2287 4487
rect 2353 4473 2367 4487
rect 2513 4473 2527 4487
rect 593 4453 607 4467
rect 1013 4453 1027 4467
rect 1113 4453 1127 4467
rect 913 4433 927 4447
rect 1173 4433 1187 4447
rect 1253 4453 1267 4467
rect 1453 4453 1467 4467
rect 1713 4453 1727 4467
rect 2114 4453 2128 4467
rect 2233 4453 2247 4467
rect 2293 4453 2307 4467
rect 1393 4433 1407 4447
rect 1493 4433 1507 4447
rect 1653 4433 1667 4447
rect 1913 4433 1927 4447
rect 2073 4433 2087 4447
rect 2213 4433 2227 4447
rect 2473 4453 2487 4467
rect 2693 4453 2707 4467
rect 2833 4473 2847 4487
rect 3253 4473 3267 4487
rect 3313 4473 3327 4487
rect 3514 4473 3528 4487
rect 3553 4473 3567 4487
rect 3633 4473 3647 4487
rect 3793 4473 3807 4487
rect 4013 4473 4027 4487
rect 4053 4473 4067 4487
rect 4093 4473 4107 4487
rect 4233 4473 4247 4487
rect 4292 4473 4306 4487
rect 4314 4473 4328 4487
rect 4693 4473 4707 4487
rect 5213 4473 5227 4487
rect 5253 4473 5267 4487
rect 5513 4473 5527 4487
rect 5673 4473 5687 4487
rect 5732 4473 5746 4487
rect 5754 4473 5768 4487
rect 5993 4473 6007 4487
rect 2953 4453 2967 4467
rect 3233 4453 3247 4467
rect 3273 4453 3287 4467
rect 3453 4453 3467 4467
rect 2433 4433 2447 4447
rect 2572 4433 2586 4447
rect 2594 4433 2608 4447
rect 2713 4433 2727 4447
rect 3053 4433 3067 4447
rect 3193 4433 3207 4447
rect 3333 4433 3347 4447
rect 3413 4433 3427 4447
rect 3533 4433 3547 4447
rect 3613 4453 3627 4467
rect 3673 4453 3687 4467
rect 3733 4453 3747 4467
rect 3972 4453 3986 4467
rect 4033 4453 4047 4467
rect 4153 4453 4167 4467
rect 4213 4453 4227 4467
rect 4373 4453 4387 4467
rect 4453 4453 4467 4467
rect 4533 4453 4547 4467
rect 4653 4453 4667 4467
rect 4733 4453 4747 4467
rect 4793 4453 4807 4467
rect 3693 4433 3707 4447
rect 3813 4433 3827 4447
rect 53 4413 67 4427
rect 93 4413 107 4427
rect 373 4413 387 4427
rect 573 4413 587 4427
rect 653 4413 667 4427
rect 1073 4413 1087 4427
rect 1193 4413 1207 4427
rect 1373 4413 1387 4427
rect 1453 4413 1467 4427
rect 1573 4413 1587 4427
rect 1613 4413 1627 4427
rect 73 4393 87 4407
rect 213 4393 227 4407
rect 253 4393 267 4407
rect 433 4393 447 4407
rect 873 4393 887 4407
rect 1133 4393 1147 4407
rect 1213 4393 1227 4407
rect 1253 4393 1267 4407
rect 1493 4393 1507 4407
rect 1533 4393 1547 4407
rect 1653 4393 1667 4407
rect 1712 4393 1726 4407
rect 1833 4393 1847 4407
rect 1893 4413 1907 4427
rect 2012 4413 2026 4427
rect 2034 4413 2048 4427
rect 2952 4413 2966 4427
rect 2974 4413 2988 4427
rect 3153 4413 3167 4427
rect 3312 4413 3326 4427
rect 4353 4433 4367 4447
rect 4113 4413 4127 4427
rect 4493 4433 4507 4447
rect 4773 4433 4787 4447
rect 4853 4433 4867 4447
rect 5033 4453 5047 4467
rect 5112 4453 5126 4467
rect 5152 4453 5166 4467
rect 5174 4453 5188 4467
rect 5393 4453 5407 4467
rect 5473 4453 5487 4467
rect 5493 4433 5507 4447
rect 5553 4453 5567 4467
rect 5853 4453 5867 4467
rect 6033 4453 6047 4467
rect 5592 4433 5606 4447
rect 5614 4433 5628 4447
rect 5713 4433 5727 4447
rect 4573 4414 4587 4428
rect 4733 4413 4747 4427
rect 4833 4413 4847 4427
rect 5073 4413 5087 4427
rect 5273 4413 5287 4427
rect 5313 4413 5327 4427
rect 53 4373 67 4387
rect 133 4373 147 4387
rect 293 4373 307 4387
rect 633 4373 647 4387
rect 913 4373 927 4387
rect 1393 4373 1407 4387
rect 1593 4373 1607 4387
rect 1633 4373 1647 4387
rect 1913 4393 1927 4407
rect 2333 4393 2347 4407
rect 2493 4393 2507 4407
rect 2713 4393 2727 4407
rect 2873 4393 2887 4407
rect 2992 4393 3006 4407
rect 3014 4393 3028 4407
rect 3133 4393 3147 4407
rect 3293 4393 3307 4407
rect 3453 4393 3467 4407
rect 3693 4393 3707 4407
rect 3852 4393 3866 4407
rect 3953 4393 3967 4407
rect 2172 4373 2186 4387
rect 2353 4373 2367 4387
rect 2733 4373 2747 4387
rect 2813 4373 2827 4387
rect 2853 4373 2867 4387
rect 3192 4373 3206 4387
rect 3393 4373 3407 4387
rect 3933 4373 3947 4387
rect 4033 4393 4047 4407
rect 4173 4393 4187 4407
rect 4253 4393 4267 4407
rect 4293 4393 4307 4407
rect 4373 4393 4387 4407
rect 4493 4393 4507 4407
rect 4573 4392 4587 4406
rect 4693 4393 4707 4407
rect 4872 4393 4886 4407
rect 4894 4394 4908 4408
rect 5573 4393 5587 4407
rect 5752 4393 5766 4407
rect 5774 4393 5788 4407
rect 5873 4393 5887 4407
rect 3993 4373 4007 4387
rect 4093 4373 4107 4387
rect 4153 4373 4167 4387
rect 93 4353 107 4367
rect 533 4353 547 4367
rect 573 4353 587 4367
rect 873 4353 887 4367
rect 1213 4353 1227 4367
rect 1253 4353 1267 4367
rect 1973 4353 1987 4367
rect 3033 4353 3047 4367
rect 3093 4353 3107 4367
rect 3733 4353 3747 4367
rect 3773 4353 3787 4367
rect 4893 4372 4907 4386
rect 5093 4373 5107 4387
rect 5153 4374 5167 4388
rect 5313 4373 5327 4387
rect 5453 4373 5467 4387
rect 5493 4373 5507 4387
rect 5913 4373 5927 4387
rect 5973 4373 5987 4387
rect 4693 4353 4707 4367
rect 4733 4353 4747 4367
rect 5153 4352 5167 4366
rect 5833 4353 5847 4367
rect 133 4333 147 4347
rect 253 4333 267 4347
rect 333 4333 347 4347
rect 433 4333 447 4347
rect 653 4333 667 4347
rect 713 4333 727 4347
rect 793 4333 807 4347
rect 833 4333 847 4347
rect 1113 4333 1127 4347
rect 1333 4333 1347 4347
rect 1533 4333 1547 4347
rect 1573 4333 1587 4347
rect 1693 4333 1707 4347
rect 1813 4333 1827 4347
rect 1853 4333 1867 4347
rect 2013 4333 2027 4347
rect 2153 4333 2167 4347
rect 2233 4333 2247 4347
rect 2373 4333 2387 4347
rect 2433 4333 2447 4347
rect 2473 4333 2487 4347
rect 2693 4333 2707 4347
rect 2773 4333 2787 4347
rect 2813 4333 2827 4347
rect 2993 4333 3007 4347
rect 3113 4333 3127 4347
rect 3293 4333 3307 4347
rect 3413 4333 3427 4347
rect 3453 4333 3467 4347
rect 3673 4333 3687 4347
rect 3813 4333 3827 4347
rect 4073 4333 4087 4347
rect 4113 4333 4127 4347
rect 4153 4333 4167 4347
rect 4253 4333 4267 4347
rect 4373 4333 4387 4347
rect 4573 4333 4587 4347
rect 4833 4333 4847 4347
rect 4953 4333 4967 4347
rect 4993 4333 5007 4347
rect 193 4313 207 4327
rect 1273 4313 1287 4327
rect 3173 4313 3187 4327
rect 3213 4313 3227 4327
rect 5093 4333 5107 4347
rect 5233 4333 5247 4347
rect 5453 4333 5467 4347
rect 5613 4333 5627 4347
rect 5813 4333 5827 4347
rect 5933 4333 5947 4347
rect 6013 4333 6027 4347
rect 5153 4313 5167 4327
rect 473 4293 487 4307
rect 933 4293 947 4307
rect 993 4293 1007 4307
rect 1253 4293 1267 4307
rect 1553 4293 1567 4307
rect 1753 4293 1767 4307
rect 1773 4293 1787 4307
rect 1913 4293 1927 4307
rect 2173 4293 2187 4307
rect 2513 4293 2527 4307
rect 2573 4293 2587 4307
rect 3033 4293 3047 4307
rect 3493 4293 3507 4307
rect 3553 4293 3567 4307
rect 3773 4293 3787 4307
rect 3913 4293 3927 4307
rect 4533 4293 4547 4307
rect 4733 4293 4747 4307
rect 4973 4293 4987 4307
rect 113 4273 127 4287
rect 153 4273 167 4287
rect 233 4273 247 4287
rect 273 4273 287 4287
rect 313 4273 327 4287
rect 513 4273 527 4287
rect 693 4273 707 4287
rect 733 4273 747 4287
rect 813 4273 827 4287
rect 853 4273 867 4287
rect 1133 4274 1147 4288
rect 1353 4273 1367 4287
rect 1393 4273 1407 4287
rect 1513 4273 1527 4287
rect 1633 4273 1647 4287
rect 1673 4273 1687 4287
rect 1953 4273 1967 4287
rect 1993 4273 2007 4287
rect 2093 4273 2107 4287
rect 2133 4273 2147 4287
rect 2253 4273 2267 4287
rect 2293 4273 2307 4287
rect 2413 4273 2427 4287
rect 2453 4273 2467 4287
rect 2793 4273 2807 4287
rect 2833 4273 2847 4287
rect 2853 4273 2867 4287
rect 553 4253 567 4267
rect 613 4253 627 4267
rect 1013 4253 1027 4267
rect 1053 4253 1067 4267
rect 1133 4252 1147 4266
rect 1313 4253 1327 4267
rect 1773 4254 1787 4268
rect 1913 4253 1927 4267
rect 2153 4253 2167 4267
rect 2913 4253 2927 4267
rect 3113 4273 3127 4287
rect 3153 4273 3167 4287
rect 3193 4273 3207 4287
rect 3393 4273 3407 4287
rect 3433 4273 3447 4287
rect 3953 4273 3967 4287
rect 3993 4273 4007 4287
rect 4133 4273 4147 4287
rect 4173 4273 4187 4287
rect 4293 4273 4307 4287
rect 4393 4273 4407 4287
rect 4433 4273 4447 4287
rect 3033 4253 3047 4267
rect 4853 4273 4867 4287
rect 4893 4273 4907 4287
rect 5013 4273 5027 4287
rect 5053 4273 5067 4287
rect 5173 4273 5187 4287
rect 5213 4273 5227 4287
rect 5293 4273 5307 4287
rect 5313 4273 5327 4287
rect 5353 4273 5367 4287
rect 5473 4273 5487 4287
rect 5513 4273 5527 4287
rect 5593 4273 5607 4287
rect 5653 4273 5667 4287
rect 5793 4273 5807 4287
rect 5833 4273 5847 4287
rect 5913 4273 5927 4287
rect 5953 4273 5967 4287
rect 4613 4253 4627 4267
rect 4833 4253 4847 4267
rect 4973 4253 4987 4267
rect 5233 4253 5247 4267
rect 5393 4254 5407 4268
rect 233 4233 247 4247
rect 753 4233 767 4247
rect 853 4233 867 4247
rect 1233 4233 1247 4247
rect 613 4213 627 4227
rect 893 4213 907 4227
rect 1173 4213 1187 4227
rect 1353 4233 1367 4247
rect 1513 4233 1527 4247
rect 1713 4233 1727 4247
rect 1773 4232 1787 4246
rect 1853 4233 1867 4247
rect 2093 4233 2107 4247
rect 2753 4233 2767 4247
rect 3013 4233 3027 4247
rect 3353 4233 3367 4247
rect 3393 4233 3407 4247
rect 3753 4233 3767 4247
rect 4133 4233 4147 4247
rect 4213 4233 4227 4247
rect 4253 4233 4267 4247
rect 4353 4233 4367 4247
rect 4393 4233 4407 4247
rect 4433 4233 4447 4247
rect 4493 4233 4507 4247
rect 4673 4233 4687 4247
rect 4993 4233 5007 4247
rect 5133 4233 5147 4247
rect 1313 4213 1327 4227
rect 1973 4213 1987 4227
rect 2153 4213 2167 4227
rect 2333 4213 2347 4227
rect 2373 4213 2387 4227
rect 2493 4213 2507 4227
rect 2733 4213 2747 4227
rect 2972 4213 2986 4227
rect 2994 4213 3008 4227
rect 3053 4213 3067 4227
rect 3113 4213 3127 4227
rect 3233 4213 3247 4227
rect 113 4193 127 4207
rect 214 4193 228 4207
rect 1613 4193 1627 4207
rect 1933 4193 1947 4207
rect 2613 4193 2627 4207
rect 2673 4193 2687 4207
rect 2773 4193 2787 4207
rect 2933 4193 2947 4207
rect 3273 4193 3287 4207
rect 3813 4213 3827 4227
rect 4573 4213 4587 4227
rect 4953 4213 4967 4227
rect 5393 4232 5407 4246
rect 5473 4233 5487 4247
rect 5593 4233 5607 4247
rect 5793 4233 5807 4247
rect 5873 4233 5887 4247
rect 5913 4233 5927 4247
rect 3513 4193 3527 4207
rect 3793 4193 3807 4207
rect 4313 4193 4327 4207
rect 4673 4193 4687 4207
rect 4933 4193 4947 4207
rect 5073 4193 5087 4207
rect 5493 4213 5507 4227
rect 5633 4193 5647 4207
rect 13 4173 27 4187
rect 73 4173 87 4187
rect 133 4173 147 4187
rect 1033 4173 1047 4187
rect 1073 4173 1087 4187
rect 1793 4173 1807 4187
rect 1913 4173 1927 4187
rect 2153 4173 2167 4187
rect 2233 4173 2247 4187
rect 2313 4173 2327 4187
rect 2353 4173 2367 4187
rect 2453 4173 2467 4187
rect 173 4153 187 4167
rect 333 4153 347 4167
rect 693 4153 707 4167
rect 813 4153 827 4167
rect 1253 4153 1267 4167
rect 33 4133 47 4147
rect 253 4133 267 4147
rect 293 4133 307 4147
rect 673 4133 687 4147
rect 1153 4133 1167 4147
rect 1233 4133 1247 4147
rect 1513 4153 1527 4167
rect 1693 4153 1707 4167
rect 2412 4153 2426 4167
rect 2434 4153 2448 4167
rect 2493 4153 2507 4167
rect 2793 4153 2807 4167
rect 2953 4173 2967 4187
rect 3352 4173 3366 4187
rect 3374 4173 3388 4187
rect 3493 4173 3507 4187
rect 3533 4173 3547 4187
rect 3573 4173 3587 4187
rect 3673 4173 3687 4187
rect 3432 4153 3446 4167
rect 3454 4153 3468 4167
rect 3793 4153 3807 4167
rect 3853 4173 3867 4187
rect 4073 4173 4087 4187
rect 4453 4173 4467 4187
rect 4653 4173 4667 4187
rect 4693 4173 4707 4187
rect 4893 4173 4907 4187
rect 5213 4173 5227 4187
rect 5613 4173 5627 4187
rect 5713 4173 5727 4187
rect 5873 4173 5887 4187
rect 1353 4133 1367 4147
rect 1574 4133 1588 4147
rect 1773 4133 1787 4147
rect 1873 4133 1887 4147
rect 13 4113 27 4127
rect 333 4113 347 4127
rect 613 4113 627 4127
rect 853 4113 867 4127
rect 933 4113 947 4127
rect 1373 4113 1387 4127
rect 1533 4113 1547 4127
rect 1813 4113 1827 4127
rect 2072 4113 2086 4127
rect 2094 4113 2108 4127
rect 2233 4113 2247 4127
rect 2293 4113 2307 4127
rect 2573 4133 2587 4147
rect 2773 4133 2787 4147
rect 3313 4133 3327 4147
rect 3373 4133 3387 4147
rect 3473 4133 3487 4147
rect 3553 4133 3567 4147
rect 3633 4133 3647 4147
rect 4833 4153 4847 4167
rect 5133 4133 5147 4147
rect 5453 4153 5467 4167
rect 5513 4153 5527 4167
rect 5573 4153 5587 4167
rect 5652 4153 5666 4167
rect 5674 4153 5688 4167
rect 5733 4153 5747 4167
rect 5973 4153 5987 4167
rect 6013 4153 6027 4167
rect 6073 4154 6087 4168
rect 5413 4133 5427 4147
rect 5593 4133 5607 4147
rect 5993 4133 6007 4147
rect 6033 4134 6047 4148
rect 6073 4132 6087 4146
rect 213 4093 227 4107
rect 893 4093 907 4107
rect 993 4093 1007 4107
rect 1233 4093 1247 4107
rect 1413 4093 1427 4107
rect 813 4073 827 4087
rect 1013 4073 1027 4087
rect 1613 4093 1627 4107
rect 1713 4093 1727 4107
rect 2033 4093 2047 4107
rect 2133 4093 2147 4107
rect 2194 4093 2208 4107
rect 2273 4093 2287 4107
rect 2393 4113 2407 4127
rect 2433 4113 2447 4127
rect 2673 4113 2687 4127
rect 3233 4113 3247 4127
rect 3333 4113 3347 4127
rect 3753 4113 3767 4127
rect 3853 4113 3867 4127
rect 3953 4113 3967 4127
rect 4433 4113 4447 4127
rect 4713 4113 4727 4127
rect 4773 4113 4787 4127
rect 5113 4113 5127 4127
rect 5153 4113 5167 4127
rect 2493 4093 2507 4107
rect 2613 4093 2627 4107
rect 2733 4093 2747 4107
rect 3033 4093 3047 4107
rect 3093 4093 3107 4107
rect 3133 4093 3147 4107
rect 3193 4093 3207 4107
rect 3733 4093 3747 4107
rect 4113 4093 4127 4107
rect 4153 4093 4167 4107
rect 4373 4093 4387 4107
rect 4573 4093 4587 4107
rect 5073 4093 5087 4107
rect 5433 4113 5447 4127
rect 5653 4113 5667 4127
rect 5693 4113 5707 4127
rect 6033 4112 6047 4126
rect 5393 4093 5407 4107
rect 5833 4093 5847 4107
rect 5993 4093 6007 4107
rect 4653 4073 4667 4087
rect 5113 4073 5127 4087
rect 5333 4073 5347 4087
rect 93 4053 107 4067
rect 133 4053 147 4067
rect 253 4053 267 4067
rect 293 4053 307 4067
rect 333 4053 347 4067
rect 393 4053 407 4067
rect 433 4053 447 4067
rect 533 4053 547 4067
rect 573 4053 587 4067
rect 933 4053 947 4067
rect 1333 4053 1347 4067
rect 1373 4053 1387 4067
rect 1473 4053 1487 4067
rect 1613 4053 1627 4067
rect 1653 4053 1667 4067
rect 1753 4053 1767 4067
rect 1793 4053 1807 4067
rect 2093 4053 2107 4067
rect 2133 4053 2147 4067
rect 2233 4053 2247 4067
rect 2273 4053 2287 4067
rect 2393 4053 2407 4067
rect 2433 4053 2447 4067
rect 2573 4053 2587 4067
rect 2613 4053 2627 4067
rect 2713 4053 2727 4067
rect 2773 4053 2787 4067
rect 3093 4053 3107 4067
rect 3133 4053 3147 4067
rect 3273 4053 3287 4067
rect 3313 4053 3327 4067
rect 3693 4053 3707 4067
rect 3733 4053 3747 4067
rect 3853 4053 3867 4067
rect 3893 4053 3907 4067
rect 3993 4053 4007 4067
rect 4033 4053 4047 4067
rect 4153 4053 4167 4067
rect 4193 4053 4207 4067
rect 4313 4053 4327 4067
rect 4353 4053 4367 4067
rect 4433 4053 4447 4067
rect 4473 4053 4487 4067
rect 4593 4053 4607 4067
rect 4633 4053 4647 4067
rect 4753 4053 4767 4067
rect 4793 4053 4807 4067
rect 4893 4053 4907 4067
rect 4933 4053 4947 4067
rect 5033 4053 5047 4067
rect 5073 4053 5087 4067
rect 5193 4053 5207 4067
rect 5233 4053 5247 4067
rect 5353 4053 5367 4067
rect 5393 4053 5407 4067
rect 5433 4053 5447 4067
rect 5513 4053 5527 4067
rect 5553 4053 5567 4067
rect 5653 4053 5667 4067
rect 5693 4053 5707 4067
rect 5833 4053 5847 4067
rect 5873 4053 5887 4067
rect 5893 4053 5907 4067
rect 5953 4053 5967 4067
rect 5993 4053 6007 4067
rect 13 4033 27 4047
rect 473 4033 487 4047
rect 753 4033 767 4047
rect 813 4033 827 4047
rect 853 4033 867 4047
rect 1033 4033 1047 4047
rect 1093 4033 1107 4047
rect 1893 4033 1907 4047
rect 1973 4033 1987 4047
rect 2813 4033 2827 4047
rect 2893 4033 2907 4047
rect 3373 4033 3387 4047
rect 3433 4033 3447 4047
rect 5273 4013 5287 4027
rect 5893 4013 5907 4027
rect 5933 4013 5947 4027
rect 113 3993 127 4007
rect 273 3993 287 4007
rect 492 3993 506 4007
rect 593 3993 607 4007
rect 633 3993 647 4007
rect 993 3993 1007 4007
rect 1213 3993 1227 4007
rect 1393 3993 1407 4007
rect 1713 3993 1727 4007
rect 1873 3993 1887 4007
rect 1933 3993 1947 4007
rect 2013 3993 2027 4007
rect 2113 3993 2127 4007
rect 2293 3993 2307 4007
rect 2333 3993 2347 4007
rect 2373 3993 2387 4007
rect 2473 3993 2487 4007
rect 2593 3993 2607 4007
rect 2753 3993 2767 4007
rect 2993 3993 3007 4007
rect 3113 3993 3127 4007
rect 3173 3993 3187 4007
rect 3293 3993 3307 4007
rect 3333 3993 3347 4007
rect 3553 3993 3567 4007
rect 3593 3993 3607 4007
rect 3713 3993 3727 4007
rect 3873 3993 3887 4007
rect 4053 3993 4067 4007
rect 4213 3993 4227 4007
rect 4333 3993 4347 4007
rect 4493 3993 4507 4007
rect 4653 3993 4667 4007
rect 4733 3993 4747 4007
rect 5053 3993 5067 4007
rect 5133 3993 5147 4007
rect 5173 3993 5187 4007
rect 5333 3993 5347 4007
rect 5393 3993 5407 4007
rect 5493 3993 5507 4007
rect 5573 3993 5587 4007
rect 5794 3993 5808 4007
rect 5853 3993 5867 4007
rect 5973 3993 5987 4007
rect 233 3973 247 3987
rect 1353 3973 1367 3987
rect 113 3953 127 3967
rect 313 3953 327 3967
rect 933 3953 947 3967
rect 973 3953 987 3967
rect 1333 3953 1347 3967
rect 2253 3973 2267 3987
rect 1653 3953 1667 3967
rect 1793 3953 1807 3967
rect 2033 3953 2047 3967
rect 3833 3973 3847 3987
rect 4013 3973 4027 3987
rect 3113 3953 3127 3967
rect 3293 3953 3307 3967
rect 3353 3953 3367 3967
rect 3693 3953 3707 3967
rect 3913 3953 3927 3967
rect 4053 3953 4067 3967
rect 4313 3953 4327 3967
rect 4773 3973 4787 3987
rect 4913 3973 4927 3987
rect 4653 3953 4667 3967
rect 4713 3953 4727 3967
rect 5033 3953 5047 3967
rect 333 3933 347 3947
rect 373 3933 387 3947
rect 473 3933 487 3947
rect 1393 3933 1407 3947
rect 1473 3933 1487 3947
rect 1893 3933 1907 3947
rect 2273 3933 2287 3947
rect 2433 3933 2447 3947
rect 2513 3933 2527 3947
rect 2793 3933 2807 3947
rect 3733 3933 3747 3947
rect 3873 3933 3887 3947
rect 3933 3933 3947 3947
rect 4293 3933 4307 3947
rect 4333 3933 4347 3947
rect 4413 3933 4427 3947
rect 4953 3933 4967 3947
rect 5133 3953 5147 3967
rect 5193 3953 5207 3967
rect 5253 3973 5267 3987
rect 5293 3973 5307 3987
rect 5913 3973 5927 3987
rect 5953 3973 5967 3987
rect 5213 3933 5227 3947
rect 5333 3953 5347 3967
rect 5493 3953 5507 3967
rect 5673 3953 5687 3967
rect 5733 3953 5747 3967
rect 5873 3953 5887 3967
rect 5253 3933 5267 3947
rect 5513 3933 5527 3947
rect 5933 3933 5947 3947
rect 293 3913 307 3927
rect 353 3913 367 3927
rect 413 3913 427 3927
rect 1753 3913 1767 3927
rect 2113 3913 2127 3927
rect 2333 3913 2347 3927
rect 2493 3913 2507 3927
rect 3253 3913 3267 3927
rect 3713 3913 3727 3927
rect 3993 3913 4007 3927
rect 4073 3913 4087 3927
rect 4593 3913 4607 3927
rect 4833 3913 4847 3927
rect 5053 3913 5067 3927
rect 5233 3913 5247 3927
rect 5493 3913 5507 3927
rect 5633 3913 5647 3927
rect 73 3893 87 3907
rect 273 3893 287 3907
rect 34 3873 48 3887
rect 133 3873 147 3887
rect 493 3873 507 3887
rect 553 3873 567 3887
rect 633 3893 647 3907
rect 673 3893 687 3907
rect 753 3893 767 3907
rect 813 3893 827 3907
rect 933 3893 947 3907
rect 1033 3893 1047 3907
rect 1093 3893 1107 3907
rect 1353 3893 1367 3907
rect 1533 3893 1547 3907
rect 1813 3893 1827 3907
rect 93 3853 107 3867
rect 393 3853 407 3867
rect 433 3853 447 3867
rect 593 3853 607 3867
rect 953 3873 967 3887
rect 993 3873 1007 3887
rect 1173 3873 1187 3887
rect 1473 3873 1487 3887
rect 1653 3873 1667 3887
rect 1713 3873 1727 3887
rect 2173 3874 2187 3888
rect 2593 3893 2607 3907
rect 2713 3893 2727 3907
rect 2913 3893 2927 3907
rect 3213 3893 3227 3907
rect 3593 3893 3607 3907
rect 3633 3893 3647 3907
rect 2313 3873 2327 3887
rect 2373 3873 2387 3887
rect 2453 3873 2467 3887
rect 2753 3873 2767 3887
rect 3313 3873 3327 3887
rect 3433 3873 3447 3887
rect 3533 3873 3547 3887
rect 3713 3873 3727 3887
rect 4013 3893 4027 3907
rect 4793 3893 4807 3907
rect 5473 3893 5487 3907
rect 5993 3893 6007 3907
rect 4053 3873 4067 3887
rect 4153 3873 4167 3887
rect 4253 3873 4267 3887
rect 4453 3873 4467 3887
rect 4613 3873 4627 3887
rect 5253 3873 5267 3887
rect 5453 3873 5467 3887
rect 5713 3873 5727 3887
rect 1053 3853 1067 3867
rect 1153 3853 1167 3867
rect 1493 3853 1507 3867
rect 1873 3853 1887 3867
rect 2032 3853 2046 3867
rect 2054 3853 2068 3867
rect 2113 3853 2127 3867
rect 2173 3852 2187 3866
rect 2333 3853 2347 3867
rect 2473 3853 2487 3867
rect 2633 3853 2647 3867
rect 2853 3853 2867 3867
rect 3073 3853 3087 3867
rect 3233 3853 3247 3867
rect 3373 3853 3387 3867
rect 3693 3853 3707 3867
rect 3833 3853 3847 3867
rect 3873 3853 3887 3867
rect 4133 3853 4147 3867
rect 4213 3853 4227 3867
rect 4273 3853 4287 3867
rect 4353 3853 4367 3867
rect 4752 3853 4766 3867
rect 4774 3853 4788 3867
rect 4913 3853 4927 3867
rect 5153 3853 5167 3867
rect 5192 3853 5206 3867
rect 33 3833 47 3847
rect 1693 3833 1707 3847
rect 4153 3833 4167 3847
rect 4813 3833 4827 3847
rect 4853 3833 4867 3847
rect 5013 3833 5027 3847
rect 5053 3833 5067 3847
rect 5353 3833 5367 3847
rect 5953 3853 5967 3867
rect 113 3813 127 3827
rect 233 3813 247 3827
rect 273 3813 287 3827
rect 453 3813 467 3827
rect 653 3813 667 3827
rect 713 3813 727 3827
rect 792 3813 806 3827
rect 873 3813 887 3827
rect 973 3813 987 3827
rect 1153 3813 1167 3827
rect 1233 3813 1247 3827
rect 1413 3813 1427 3827
rect 1493 3813 1507 3827
rect 1573 3813 1587 3827
rect 1753 3813 1767 3827
rect 1873 3813 1887 3827
rect 1973 3813 1987 3827
rect 2033 3813 2047 3827
rect 2173 3813 2187 3827
rect 2233 3813 2247 3827
rect 2313 3813 2327 3827
rect 2473 3813 2487 3827
rect 2853 3813 2867 3827
rect 2893 3813 2907 3827
rect 2933 3813 2947 3827
rect 3112 3813 3126 3827
rect 3134 3813 3148 3827
rect 3233 3813 3247 3827
rect 3273 3813 3287 3827
rect 3313 3813 3327 3827
rect 3434 3813 3448 3827
rect 3533 3813 3547 3827
rect 3593 3813 3607 3827
rect 3693 3813 3707 3827
rect 3833 3813 3847 3827
rect 3933 3813 3947 3827
rect 4073 3813 4087 3827
rect 4113 3813 4127 3827
rect 4173 3813 4187 3827
rect 4413 3813 4427 3827
rect 4453 3813 4467 3827
rect 4533 3813 4547 3827
rect 4593 3813 4607 3827
rect 4653 3813 4667 3827
rect 4753 3813 4767 3827
rect 4873 3813 4887 3827
rect 4933 3813 4947 3827
rect 5153 3813 5167 3827
rect 5193 3813 5207 3827
rect 5333 3813 5347 3827
rect 5453 3813 5467 3827
rect 5633 3813 5647 3827
rect 5793 3813 5807 3827
rect 5873 3813 5887 3827
rect 5913 3813 5927 3827
rect 13 3773 27 3787
rect 3993 3773 4007 3787
rect 4153 3773 4167 3787
rect 93 3753 107 3767
rect 133 3753 147 3767
rect 213 3753 227 3767
rect 253 3753 267 3767
rect 393 3753 407 3767
rect 433 3753 447 3767
rect 533 3753 547 3767
rect 573 3753 587 3767
rect 752 3753 766 3767
rect 893 3753 907 3767
rect 953 3753 967 3767
rect 973 3753 987 3767
rect 1133 3753 1147 3767
rect 1353 3753 1367 3767
rect 1393 3753 1407 3767
rect 1433 3753 1447 3767
rect 1473 3753 1487 3767
rect 1553 3753 1567 3767
rect 1593 3753 1607 3767
rect 1673 3753 1687 3767
rect 1713 3753 1727 3767
rect 1853 3753 1867 3767
rect 1893 3753 1907 3767
rect 1933 3753 1947 3767
rect 2013 3753 2027 3767
rect 2053 3753 2067 3767
rect 2293 3753 2307 3767
rect 2333 3753 2347 3767
rect 2453 3753 2467 3767
rect 2493 3753 2507 3767
rect 2593 3753 2607 3767
rect 2633 3753 2647 3767
rect 2713 3753 2727 3767
rect 2753 3753 2767 3767
rect 2873 3753 2887 3767
rect 2913 3753 2927 3767
rect 3033 3753 3047 3767
rect 3073 3753 3087 3767
rect 3173 3753 3187 3767
rect 3213 3753 3227 3767
rect 3333 3753 3347 3767
rect 3373 3753 3387 3767
rect 3453 3753 3467 3767
rect 3513 3753 3527 3767
rect 3553 3753 3567 3767
rect 3673 3753 3687 3767
rect 3713 3753 3727 3767
rect 3773 3753 3787 3767
rect 3913 3753 3927 3767
rect 3953 3753 3967 3767
rect 4233 3753 4247 3767
rect 4273 3753 4287 3767
rect 4393 3753 4407 3767
rect 4433 3753 4447 3767
rect 4573 3753 4587 3767
rect 4613 3753 4627 3767
rect 4733 3753 4747 3767
rect 4773 3753 4787 3767
rect 4853 3753 4867 3767
rect 4893 3753 4907 3767
rect 113 3713 127 3727
rect 213 3713 227 3727
rect 253 3713 267 3727
rect 433 3713 447 3727
rect 493 3713 507 3727
rect 1013 3733 1027 3747
rect 353 3693 367 3707
rect 533 3693 547 3707
rect 713 3693 727 3707
rect 753 3713 767 3727
rect 893 3713 907 3727
rect 1133 3713 1147 3727
rect 1293 3713 1307 3727
rect 1853 3713 1867 3727
rect 2053 3713 2067 3727
rect 3313 3733 3327 3747
rect 3853 3733 3867 3747
rect 5073 3753 5087 3767
rect 5113 3753 5127 3767
rect 5313 3753 5327 3767
rect 5353 3753 5367 3767
rect 5433 3753 5447 3767
rect 5473 3753 5487 3767
rect 5733 3753 5747 3767
rect 5773 3753 5787 3767
rect 5093 3733 5107 3747
rect 2273 3713 2287 3727
rect 2373 3713 2387 3727
rect 2493 3713 2507 3727
rect 2753 3713 2767 3727
rect 2853 3713 2867 3727
rect 2913 3713 2927 3727
rect 3093 3713 3107 3727
rect 3473 3713 3487 3727
rect 3513 3713 3527 3727
rect 3913 3713 3927 3727
rect 3993 3713 4007 3727
rect 4233 3713 4247 3727
rect 4313 3713 4327 3727
rect 4733 3713 4747 3727
rect 4853 3713 4867 3727
rect 5733 3713 5747 3727
rect 5773 3713 5787 3727
rect 794 3693 808 3707
rect 873 3693 887 3707
rect 1073 3693 1087 3707
rect 1193 3693 1207 3707
rect 1273 3693 1287 3707
rect 1433 3693 1447 3707
rect 1593 3693 1607 3707
rect 2193 3693 2207 3707
rect 3633 3693 3647 3707
rect 3793 3693 3807 3707
rect 3933 3693 3947 3707
rect 4493 3693 4507 3707
rect 4613 3693 4627 3707
rect 4713 3693 4727 3707
rect 4813 3693 4827 3707
rect 5233 3693 5247 3707
rect 5633 3693 5647 3707
rect 5753 3693 5767 3707
rect 5833 3693 5847 3707
rect 473 3673 487 3687
rect 573 3673 587 3687
rect 753 3673 767 3687
rect 813 3673 827 3687
rect 853 3673 867 3687
rect 973 3673 987 3687
rect 1673 3673 1687 3687
rect 2233 3673 2247 3687
rect 2293 3673 2307 3687
rect 2333 3673 2347 3687
rect 2453 3673 2467 3687
rect 2753 3673 2767 3687
rect 2793 3673 2807 3687
rect 3092 3673 3106 3687
rect 3353 3673 3367 3687
rect 3773 3673 3787 3687
rect 3832 3673 3846 3687
rect 3953 3673 3967 3687
rect 4233 3673 4247 3687
rect 4353 3673 4367 3687
rect 5033 3673 5047 3687
rect 5313 3673 5327 3687
rect 5473 3673 5487 3687
rect 13 3653 27 3667
rect 213 3633 227 3647
rect 513 3633 527 3647
rect 893 3653 907 3667
rect 933 3653 947 3667
rect 1013 3633 1027 3647
rect 1073 3653 1087 3667
rect 1593 3653 1607 3667
rect 1873 3653 1887 3667
rect 2153 3653 2167 3667
rect 2253 3653 2267 3667
rect 3073 3653 3087 3667
rect 3553 3653 3567 3667
rect 3673 3653 3687 3667
rect 3853 3653 3867 3667
rect 4053 3653 4067 3667
rect 4393 3653 4407 3667
rect 4953 3653 4967 3667
rect 5913 3653 5927 3667
rect 1113 3633 1127 3647
rect 13 3613 27 3627
rect 2713 3633 2727 3647
rect 2793 3633 2807 3647
rect 2953 3633 2967 3647
rect 3093 3633 3107 3647
rect 3133 3634 3147 3648
rect 3193 3633 3207 3647
rect 3313 3633 3327 3647
rect 3453 3633 3467 3647
rect 5153 3633 5167 3647
rect 5233 3633 5247 3647
rect 5393 3633 5407 3647
rect 5433 3633 5447 3647
rect 2373 3613 2387 3627
rect 2753 3613 2767 3627
rect 173 3593 187 3607
rect 413 3593 427 3607
rect 693 3593 707 3607
rect 813 3593 827 3607
rect 1453 3593 1467 3607
rect 1793 3593 1807 3607
rect 2113 3593 2127 3607
rect 2193 3593 2207 3607
rect 2593 3593 2607 3607
rect 2653 3593 2667 3607
rect 3133 3612 3147 3626
rect 3233 3613 3247 3627
rect 3593 3613 3607 3627
rect 3733 3613 3747 3627
rect 3853 3613 3867 3627
rect 4533 3613 4547 3627
rect 4833 3613 4847 3627
rect 5053 3613 5067 3627
rect 5193 3613 5207 3627
rect 5373 3613 5387 3627
rect 2953 3593 2967 3607
rect 3093 3593 3107 3607
rect 3153 3593 3167 3607
rect 3273 3593 3287 3607
rect 3393 3593 3407 3607
rect 3873 3593 3887 3607
rect 4053 3593 4067 3607
rect 4173 3593 4187 3607
rect 4513 3593 4527 3607
rect 4733 3593 4747 3607
rect 5153 3593 5167 3607
rect 233 3573 247 3587
rect 273 3573 287 3587
rect 313 3573 327 3587
rect 473 3573 487 3587
rect 1333 3573 1347 3587
rect 1393 3573 1407 3587
rect 1533 3573 1547 3587
rect 1593 3573 1607 3587
rect 1693 3573 1707 3587
rect 1753 3573 1767 3587
rect 1832 3573 1846 3587
rect 1854 3573 1868 3587
rect 2133 3573 2147 3587
rect 2333 3573 2347 3587
rect 2833 3573 2847 3587
rect 2993 3573 3007 3587
rect 3113 3573 3127 3587
rect 3593 3573 3607 3587
rect 3773 3573 3787 3587
rect 3893 3573 3907 3587
rect 4553 3573 4567 3587
rect 4693 3573 4707 3587
rect 4973 3574 4987 3588
rect 5573 3593 5587 3607
rect 5633 3593 5647 3607
rect 5873 3594 5887 3608
rect 5913 3593 5927 3607
rect 5193 3573 5207 3587
rect 5313 3573 5327 3587
rect 5353 3573 5367 3587
rect 5393 3573 5407 3587
rect 5433 3573 5447 3587
rect 5533 3573 5547 3587
rect 5593 3573 5607 3587
rect 5793 3573 5807 3587
rect 5873 3572 5887 3586
rect 5953 3573 5967 3587
rect 5993 3573 6007 3587
rect 6073 3573 6087 3587
rect 193 3553 207 3567
rect 693 3553 707 3567
rect 1133 3553 1147 3567
rect 13 3533 27 3547
rect 93 3533 107 3547
rect 133 3533 147 3547
rect 233 3533 247 3547
rect 273 3533 287 3547
rect 473 3533 487 3547
rect 513 3533 527 3547
rect 653 3533 667 3547
rect 1233 3533 1247 3547
rect 1393 3533 1407 3547
rect 1493 3533 1507 3547
rect 1533 3533 1547 3547
rect 1653 3533 1667 3547
rect 1693 3533 1707 3547
rect 1833 3533 1847 3547
rect 1873 3533 1887 3547
rect 1993 3533 2007 3547
rect 2033 3533 2047 3547
rect 2113 3533 2127 3547
rect 2153 3533 2167 3547
rect 2293 3533 2307 3547
rect 2333 3533 2347 3547
rect 2553 3553 2567 3567
rect 3633 3553 3647 3567
rect 3693 3553 3707 3567
rect 4933 3553 4947 3567
rect 4973 3552 4987 3566
rect 2793 3533 2807 3547
rect 2833 3533 2847 3547
rect 2953 3533 2967 3547
rect 2993 3533 3007 3547
rect 3113 3533 3127 3547
rect 3153 3533 3167 3547
rect 3233 3533 3247 3547
rect 3313 3533 3327 3547
rect 3393 3533 3407 3547
rect 3433 3533 3447 3547
rect 3573 3533 3587 3547
rect 3613 3533 3627 3547
rect 3753 3533 3767 3547
rect 3793 3533 3807 3547
rect 3873 3533 3887 3547
rect 3913 3533 3927 3547
rect 4153 3533 4167 3547
rect 4193 3533 4207 3547
rect 4233 3533 4247 3547
rect 4353 3533 4367 3547
rect 4393 3533 4407 3547
rect 4473 3533 4487 3547
rect 4513 3533 4527 3547
rect 4553 3533 4567 3547
rect 4653 3533 4667 3547
rect 4693 3533 4707 3547
rect 4793 3533 4807 3547
rect 4833 3533 4847 3547
rect 4873 3533 4887 3547
rect 5153 3533 5167 3547
rect 5193 3533 5207 3547
rect 5353 3533 5367 3547
rect 5393 3533 5407 3547
rect 5433 3533 5447 3547
rect 5673 3533 5687 3547
rect 5713 3533 5727 3547
rect 5753 3533 5767 3547
rect 5833 3533 5847 3547
rect 5873 3533 5887 3547
rect 5933 3533 5947 3547
rect 853 3513 867 3527
rect 893 3513 907 3527
rect 953 3513 967 3527
rect 2433 3513 2447 3527
rect 2513 3513 2527 3527
rect 2653 3513 2667 3527
rect 4313 3513 4327 3527
rect 4953 3513 4967 3527
rect 4993 3513 5007 3527
rect 5033 3513 5047 3527
rect 4253 3493 4267 3507
rect 113 3473 127 3487
rect 213 3473 227 3487
rect 333 3473 347 3487
rect 393 3473 407 3487
rect 453 3473 467 3487
rect 493 3473 507 3487
rect 533 3473 547 3487
rect 793 3473 807 3487
rect 1073 3473 1087 3487
rect 1173 3473 1187 3487
rect 1253 3473 1267 3487
rect 1513 3473 1527 3487
rect 1553 3473 1567 3487
rect 1593 3473 1607 3487
rect 1633 3473 1647 3487
rect 1713 3473 1727 3487
rect 1753 3473 1767 3487
rect 1853 3473 1867 3487
rect 2013 3473 2027 3487
rect 2133 3473 2147 3487
rect 2273 3473 2287 3487
rect 2673 3473 2687 3487
rect 2733 3473 2747 3487
rect 2813 3473 2827 3487
rect 2873 3473 2887 3487
rect 2973 3473 2987 3487
rect 3133 3473 3147 3487
rect 3293 3473 3307 3487
rect 3413 3473 3427 3487
rect 3553 3473 3567 3487
rect 3633 3473 3647 3487
rect 3673 3473 3687 3487
rect 3773 3473 3787 3487
rect 3893 3473 3907 3487
rect 3993 3473 4007 3487
rect 4033 3473 4047 3487
rect 4073 3473 4087 3487
rect 4213 3473 4227 3487
rect 4313 3473 4327 3487
rect 4373 3473 4387 3487
rect 4473 3473 4487 3487
rect 4533 3473 4547 3487
rect 4633 3473 4647 3487
rect 113 3433 127 3447
rect 853 3453 867 3467
rect 893 3453 907 3467
rect 1213 3453 1227 3467
rect 1673 3453 1687 3467
rect 873 3433 887 3447
rect 953 3433 967 3447
rect 1013 3433 1027 3447
rect 1093 3433 1107 3447
rect 1953 3433 1967 3447
rect 2173 3453 2187 3467
rect 2453 3453 2467 3467
rect 2493 3453 2507 3467
rect 2253 3433 2267 3447
rect 2953 3433 2967 3447
rect 3253 3453 3267 3467
rect 3313 3433 3327 3447
rect 3413 3433 3427 3447
rect 4253 3453 4267 3467
rect 4393 3453 4407 3467
rect 4733 3473 4747 3487
rect 4753 3453 4767 3467
rect 4973 3453 4987 3467
rect 5173 3473 5187 3487
rect 5313 3473 5327 3487
rect 5413 3473 5427 3487
rect 5553 3473 5567 3487
rect 5593 3473 5607 3487
rect 5733 3473 5747 3487
rect 5773 3473 5787 3487
rect 5853 3473 5867 3487
rect 5993 3473 6007 3487
rect 5693 3453 5707 3467
rect 5893 3453 5907 3467
rect 3953 3433 3967 3447
rect 3993 3433 4007 3447
rect 4533 3433 4547 3447
rect 4933 3433 4947 3447
rect 5413 3433 5427 3447
rect 5513 3433 5527 3447
rect 5613 3433 5627 3447
rect 5653 3433 5667 3447
rect 273 3413 287 3427
rect 1113 3413 1127 3427
rect 1173 3413 1187 3427
rect 1453 3413 1467 3427
rect 1793 3413 1807 3427
rect 333 3393 347 3407
rect 1593 3393 1607 3407
rect 533 3373 547 3387
rect 733 3373 747 3387
rect 853 3373 867 3387
rect 1213 3373 1227 3387
rect 1333 3373 1347 3387
rect 1993 3393 2007 3407
rect 2053 3413 2067 3427
rect 2173 3413 2187 3427
rect 2392 3413 2406 3427
rect 2793 3413 2807 3427
rect 3032 3413 3046 3427
rect 4433 3413 4447 3427
rect 4793 3413 4807 3427
rect 4833 3413 4847 3427
rect 5093 3413 5107 3427
rect 5213 3413 5227 3427
rect 5373 3413 5387 3427
rect 5873 3413 5887 3427
rect 5953 3413 5967 3427
rect 2113 3393 2127 3407
rect 2373 3393 2387 3407
rect 2513 3393 2527 3407
rect 2873 3393 2887 3407
rect 2973 3393 2987 3407
rect 3353 3393 3367 3407
rect 3693 3393 3707 3407
rect 4073 3393 4087 3407
rect 5173 3393 5187 3407
rect 5413 3393 5427 3407
rect 1673 3373 1687 3387
rect 2293 3373 2307 3387
rect 2493 3373 2507 3387
rect 3133 3373 3147 3387
rect 3373 3373 3387 3387
rect 3553 3373 3567 3387
rect 3633 3373 3647 3387
rect 4933 3373 4947 3387
rect 4993 3373 5007 3387
rect 5073 3373 5087 3387
rect 5253 3373 5267 3387
rect 6033 3374 6047 3388
rect 6073 3373 6087 3387
rect 273 3353 287 3367
rect 693 3353 707 3367
rect 833 3353 847 3367
rect 2593 3353 2607 3367
rect 2873 3353 2887 3367
rect 3193 3353 3207 3367
rect 3573 3353 3587 3367
rect 4053 3353 4067 3367
rect 4313 3353 4327 3367
rect 4353 3353 4367 3367
rect 4393 3353 4407 3367
rect 4833 3353 4847 3367
rect 5493 3353 5507 3367
rect 5993 3353 6007 3367
rect 6033 3352 6047 3366
rect 53 3333 67 3347
rect 133 3333 147 3347
rect 253 3333 267 3347
rect 353 3333 367 3347
rect 393 3333 407 3347
rect 733 3333 747 3347
rect 853 3333 867 3347
rect 1373 3333 1387 3347
rect 1433 3333 1447 3347
rect 2333 3333 2347 3347
rect 2393 3333 2407 3347
rect 2833 3333 2847 3347
rect 3253 3333 3267 3347
rect 3493 3333 3507 3347
rect 3773 3333 3787 3347
rect 3953 3333 3967 3347
rect 4173 3333 4187 3347
rect 5053 3333 5067 3347
rect 5093 3333 5107 3347
rect 5133 3333 5147 3347
rect 5553 3333 5567 3347
rect 5693 3333 5707 3347
rect 5853 3333 5867 3347
rect 5973 3333 5987 3347
rect 693 3313 707 3327
rect 2553 3313 2567 3327
rect 2593 3313 2607 3327
rect 4313 3313 4327 3327
rect 4353 3313 4367 3327
rect 4813 3313 4827 3327
rect 4853 3313 4867 3327
rect 4893 3313 4907 3327
rect 4933 3313 4947 3327
rect 73 3293 87 3307
rect 133 3293 147 3307
rect 253 3293 267 3307
rect 293 3293 307 3307
rect 393 3293 407 3307
rect 633 3293 647 3307
rect 833 3293 847 3307
rect 1413 3293 1427 3307
rect 1693 3293 1707 3307
rect 1733 3293 1747 3307
rect 2253 3293 2267 3307
rect 2393 3293 2407 3307
rect 2513 3293 2527 3307
rect 2733 3293 2747 3307
rect 2933 3293 2947 3307
rect 3033 3293 3047 3307
rect 3133 3293 3147 3307
rect 3232 3293 3246 3307
rect 3333 3293 3347 3307
rect 3373 3293 3387 3307
rect 3493 3293 3507 3307
rect 3593 3293 3607 3307
rect 3713 3293 3727 3307
rect 3873 3293 3887 3307
rect 3913 3293 3927 3307
rect 3973 3293 3987 3307
rect 4013 3293 4027 3307
rect 4273 3293 4287 3307
rect 4393 3293 4407 3307
rect 4573 3293 4587 3307
rect 4672 3293 4686 3307
rect 4793 3293 4807 3307
rect 4973 3293 4987 3307
rect 5093 3293 5107 3307
rect 5313 3293 5327 3307
rect 5373 3293 5387 3307
rect 5473 3293 5487 3307
rect 5553 3293 5567 3307
rect 5653 3293 5667 3307
rect 5774 3293 5788 3307
rect 5853 3293 5867 3307
rect 673 3253 687 3267
rect 753 3253 767 3267
rect 773 3253 787 3267
rect 1073 3253 1087 3267
rect 1173 3253 1187 3267
rect 1273 3253 1287 3267
rect 1453 3253 1467 3267
rect 1513 3253 1527 3267
rect 2113 3253 2127 3267
rect 2153 3253 2167 3267
rect 2293 3253 2307 3267
rect 2613 3253 2627 3267
rect 4273 3253 4287 3267
rect 4853 3253 4867 3267
rect 5333 3253 5347 3267
rect 5493 3253 5507 3267
rect 113 3233 127 3247
rect 153 3233 167 3247
rect 233 3233 247 3247
rect 273 3233 287 3247
rect 413 3213 427 3227
rect 293 3193 307 3207
rect 713 3233 727 3247
rect 813 3233 827 3247
rect 853 3233 867 3247
rect 953 3233 967 3247
rect 1753 3233 1767 3247
rect 1873 3233 1887 3247
rect 2053 3233 2067 3247
rect 2373 3233 2387 3247
rect 2413 3233 2427 3247
rect 2713 3233 2727 3247
rect 2753 3233 2767 3247
rect 2833 3233 2847 3247
rect 2873 3233 2887 3247
rect 3113 3233 3127 3247
rect 3153 3233 3167 3247
rect 3313 3233 3327 3247
rect 3353 3233 3367 3247
rect 3393 3233 3407 3247
rect 3433 3233 3447 3247
rect 3473 3233 3487 3247
rect 3513 3233 3527 3247
rect 3553 3233 3567 3247
rect 3693 3233 3707 3247
rect 3733 3233 3747 3247
rect 3773 3233 3787 3247
rect 3993 3233 4007 3247
rect 4033 3233 4047 3247
rect 4173 3233 4187 3247
rect 4213 3233 4227 3247
rect 4453 3233 4467 3247
rect 4493 3233 4507 3247
rect 4593 3233 4607 3247
rect 4633 3233 4647 3247
rect 4773 3233 4787 3247
rect 4813 3233 4827 3247
rect 5073 3233 5087 3247
rect 5113 3233 5127 3247
rect 5213 3233 5227 3247
rect 5253 3233 5267 3247
rect 5533 3233 5547 3247
rect 5573 3233 5587 3247
rect 5673 3233 5687 3247
rect 5713 3233 5727 3247
rect 5833 3233 5847 3247
rect 5873 3233 5887 3247
rect 5953 3233 5967 3247
rect 5993 3233 6007 3247
rect 673 3213 687 3227
rect 773 3193 787 3207
rect 813 3193 827 3207
rect 1233 3193 1247 3207
rect 4893 3213 4907 3227
rect 4973 3213 4987 3227
rect 1753 3193 1767 3207
rect 1813 3193 1827 3207
rect 1873 3193 1887 3207
rect 1913 3193 1927 3207
rect 2293 3193 2307 3207
rect 2413 3193 2427 3207
rect 2713 3193 2727 3207
rect 2793 3193 2807 3207
rect 2833 3193 2847 3207
rect 2873 3193 2887 3207
rect 3033 3193 3047 3207
rect 3113 3193 3127 3207
rect 3473 3193 3487 3207
rect 3633 3193 3647 3207
rect 3733 3193 3747 3207
rect 4213 3193 4227 3207
rect 4373 3193 4387 3207
rect 4553 3193 4567 3207
rect 4633 3193 4647 3207
rect 4773 3193 4787 3207
rect 5073 3193 5087 3207
rect 5413 3193 5427 3207
rect 5573 3193 5587 3207
rect 5713 3193 5727 3207
rect 5833 3193 5847 3207
rect 113 3173 127 3187
rect 273 3173 287 3187
rect 413 3173 427 3187
rect 633 3173 647 3187
rect 953 3173 967 3187
rect 2253 3173 2267 3187
rect 2373 3173 2387 3187
rect 2693 3173 2707 3187
rect 2753 3173 2767 3187
rect 3152 3173 3166 3187
rect 3174 3173 3188 3187
rect 4593 3173 4607 3187
rect 4893 3173 4907 3187
rect 5533 3173 5547 3187
rect 353 3153 367 3167
rect 713 3153 727 3167
rect 1393 3153 1407 3167
rect 1873 3153 1887 3167
rect 1913 3153 1927 3167
rect 2073 3153 2087 3167
rect 2733 3153 2747 3167
rect 2853 3153 2867 3167
rect 4493 3153 4507 3167
rect 4633 3153 4647 3167
rect 5573 3153 5587 3167
rect 33 3133 47 3147
rect 153 3133 167 3147
rect 233 3133 247 3147
rect 673 3133 687 3147
rect 1273 3133 1287 3147
rect 1653 3133 1667 3147
rect 1933 3133 1947 3147
rect 2153 3133 2167 3147
rect 2473 3133 2487 3147
rect 2693 3133 2707 3147
rect 2813 3133 2827 3147
rect 3093 3133 3107 3147
rect 4173 3133 4187 3147
rect 4353 3133 4367 3147
rect 5213 3133 5227 3147
rect 5393 3133 5407 3147
rect 1233 3113 1247 3127
rect 2413 3113 2427 3127
rect 2953 3113 2967 3127
rect 4233 3113 4247 3127
rect 4273 3114 4287 3128
rect 5433 3113 5447 3127
rect 5513 3113 5527 3127
rect 1073 3093 1087 3107
rect 1293 3093 1307 3107
rect 1553 3093 1567 3107
rect 1813 3093 1827 3107
rect 1873 3093 1887 3107
rect 2333 3093 2347 3107
rect 2913 3093 2927 3107
rect 3133 3093 3147 3107
rect 3213 3093 3227 3107
rect 3953 3093 3967 3107
rect 4273 3092 4287 3106
rect 4693 3093 4707 3107
rect 5253 3093 5267 3107
rect 5393 3093 5407 3107
rect 5453 3093 5467 3107
rect 5493 3093 5507 3107
rect 5653 3093 5667 3107
rect 5833 3093 5847 3107
rect 1013 3073 1027 3087
rect 1153 3073 1167 3087
rect 1373 3073 1387 3087
rect 1433 3073 1447 3087
rect 1613 3073 1627 3087
rect 1733 3073 1747 3087
rect 2133 3073 2147 3087
rect 2393 3073 2407 3087
rect 2433 3073 2447 3087
rect 2513 3073 2527 3087
rect 2613 3073 2627 3087
rect 2793 3073 2807 3087
rect 3053 3073 3067 3087
rect 3493 3073 3507 3087
rect 3673 3073 3687 3087
rect 3813 3073 3827 3087
rect 4153 3073 4167 3087
rect 4433 3073 4447 3087
rect 4633 3073 4647 3087
rect 4853 3073 4867 3087
rect 5013 3073 5027 3087
rect 5473 3073 5487 3087
rect 5633 3073 5647 3087
rect 5733 3073 5747 3087
rect 113 3053 127 3067
rect 213 3053 227 3067
rect 793 3053 807 3067
rect 2673 3053 2687 3067
rect 2753 3053 2767 3067
rect 2933 3053 2947 3067
rect 3133 3053 3147 3067
rect 3393 3053 3407 3067
rect 3853 3053 3867 3067
rect 3933 3053 3947 3067
rect 4893 3053 4907 3067
rect 4973 3053 4987 3067
rect 5693 3053 5707 3067
rect 5773 3053 5787 3067
rect 5933 3053 5947 3067
rect 6013 3053 6027 3067
rect 1813 3033 1827 3047
rect 5193 3033 5207 3047
rect 113 3013 127 3027
rect 153 3013 167 3027
rect 253 3013 267 3027
rect 293 3013 307 3027
rect 413 3013 427 3027
rect 453 3013 467 3027
rect 553 3013 567 3027
rect 593 3013 607 3027
rect 693 3013 707 3027
rect 733 3013 747 3027
rect 993 3013 1007 3027
rect 1073 3013 1087 3027
rect 1113 3013 1127 3027
rect 1153 3013 1167 3027
rect 1293 3013 1307 3027
rect 1333 3013 1347 3027
rect 1433 3013 1447 3027
rect 1473 3013 1487 3027
rect 1733 3013 1747 3027
rect 1773 3013 1787 3027
rect 1973 3013 1987 3027
rect 2013 3013 2027 3027
rect 2053 3013 2067 3027
rect 2093 3013 2107 3027
rect 2153 3013 2167 3027
rect 2193 3013 2207 3027
rect 2233 3013 2247 3027
rect 2353 3013 2367 3027
rect 2393 3013 2407 3027
rect 2433 3013 2447 3027
rect 2593 3013 2607 3027
rect 2633 3013 2647 3027
rect 2673 3013 2687 3027
rect 2793 3013 2807 3027
rect 2833 3013 2847 3027
rect 2913 3013 2927 3027
rect 2953 3013 2967 3027
rect 3093 3013 3107 3027
rect 3133 3013 3147 3027
rect 3213 3013 3227 3027
rect 3253 3013 3267 3027
rect 3313 3013 3327 3027
rect 3353 3013 3367 3027
rect 3393 3013 3407 3027
rect 3493 3013 3507 3027
rect 3533 3013 3547 3027
rect 3673 3013 3687 3027
rect 3713 3013 3727 3027
rect 3813 3013 3827 3027
rect 3853 3013 3867 3027
rect 3973 3013 3987 3027
rect 4013 3013 4027 3027
rect 4053 3013 4067 3027
rect 4273 3013 4287 3027
rect 4313 3013 4327 3027
rect 4393 3013 4407 3027
rect 4433 3013 4447 3027
rect 4733 3013 4747 3027
rect 4853 3013 4867 3027
rect 4893 3013 4907 3027
rect 4973 3013 4987 3027
rect 5013 3013 5027 3027
rect 5133 3013 5147 3027
rect 5173 3013 5187 3027
rect 5433 3013 5447 3027
rect 5473 3013 5487 3027
rect 5513 3013 5527 3027
rect 5673 3013 5687 3027
rect 5713 3013 5727 3027
rect 5773 3013 5787 3027
rect 5813 3013 5827 3027
rect 5973 3013 5987 3027
rect 6013 3013 6027 3027
rect 873 2993 887 3007
rect 1513 2993 1527 3007
rect 1813 2993 1827 3007
rect 4573 2993 4587 3007
rect 5213 2993 5227 3007
rect 5253 2993 5267 3007
rect 5333 2993 5347 3007
rect 5393 2993 5407 3007
rect 5933 2993 5947 3007
rect 93 2953 107 2967
rect 133 2953 147 2967
rect 173 2953 187 2967
rect 313 2953 327 2967
rect 673 2953 687 2967
rect 713 2953 727 2967
rect 753 2953 767 2967
rect 973 2953 987 2967
rect 1093 2953 1107 2967
rect 1133 2953 1147 2967
rect 1313 2953 1327 2967
rect 1453 2953 1467 2967
rect 1493 2953 1507 2967
rect 1633 2953 1647 2967
rect 1713 2953 1727 2967
rect 1793 2953 1807 2967
rect 2133 2953 2147 2967
rect 2173 2953 2187 2967
rect 2213 2953 2227 2967
rect 2253 2953 2267 2967
rect 2413 2953 2427 2967
rect 2493 2953 2507 2967
rect 2613 2953 2627 2967
rect 2673 2953 2687 2967
rect 2813 2953 2827 2967
rect 2933 2953 2947 2967
rect 3053 2953 3067 2967
rect 3194 2953 3208 2967
rect 3313 2953 3327 2967
rect 3473 2953 3487 2967
rect 3513 2953 3527 2967
rect 3653 2953 3667 2967
rect 3733 2953 3747 2967
rect 3793 2953 3807 2967
rect 3953 2953 3967 2967
rect 4113 2953 4127 2967
rect 4153 2953 4167 2967
rect 4293 2953 4307 2967
rect 4413 2953 4427 2967
rect 4513 2953 4527 2967
rect 4593 2953 4607 2967
rect 4693 2953 4707 2967
rect 4773 2953 4787 2967
rect 4873 2953 4887 2967
rect 5113 2953 5127 2967
rect 5193 2953 5207 2967
rect 5273 2953 5287 2967
rect 5313 2953 5327 2967
rect 5453 2953 5467 2967
rect 5553 2953 5567 2967
rect 5833 2953 5847 2967
rect 113 2913 127 2927
rect 173 2913 187 2927
rect 253 2913 267 2927
rect 533 2913 547 2927
rect 713 2913 727 2927
rect 753 2913 767 2927
rect 933 2933 947 2947
rect 1273 2933 1287 2947
rect 1093 2913 1107 2927
rect 1333 2913 1347 2927
rect 1473 2913 1487 2927
rect 1553 2913 1567 2927
rect 1893 2933 1907 2947
rect 1933 2933 1947 2947
rect 2073 2933 2087 2947
rect 2773 2933 2787 2947
rect 2113 2913 2127 2927
rect 2213 2913 2227 2927
rect 2852 2913 2866 2927
rect 2933 2913 2947 2927
rect 3473 2913 3487 2927
rect 3753 2913 3767 2927
rect 3993 2933 4007 2947
rect 3853 2913 3867 2927
rect 4113 2913 4127 2927
rect 5393 2913 5407 2927
rect 5553 2913 5567 2927
rect 5953 2913 5967 2927
rect 153 2893 167 2907
rect 453 2893 467 2907
rect 593 2893 607 2907
rect 733 2893 747 2907
rect 1233 2893 1247 2907
rect 1313 2894 1327 2908
rect 1593 2893 1607 2907
rect 1713 2893 1727 2907
rect 1753 2893 1767 2907
rect 2253 2893 2267 2907
rect 2413 2893 2427 2907
rect 2613 2893 2627 2907
rect 3653 2893 3667 2907
rect 4033 2893 4047 2907
rect 4233 2893 4247 2907
rect 4293 2893 4307 2907
rect 4353 2893 4367 2907
rect 4413 2893 4427 2907
rect 4573 2893 4587 2907
rect 1313 2872 1327 2886
rect 1553 2873 1567 2887
rect 1633 2873 1647 2887
rect 2233 2873 2247 2887
rect 4193 2873 4207 2887
rect 4313 2873 4327 2887
rect 4373 2873 4387 2887
rect 4553 2873 4567 2887
rect 4873 2893 4887 2907
rect 5013 2893 5027 2907
rect 5332 2893 5346 2907
rect 5973 2893 5987 2907
rect 5133 2873 5147 2887
rect 53 2853 67 2867
rect 273 2853 287 2867
rect 413 2853 427 2867
rect 573 2853 587 2867
rect 913 2853 927 2867
rect 953 2853 967 2867
rect 1073 2853 1087 2867
rect 1133 2853 1147 2867
rect 1433 2853 1447 2867
rect 1493 2853 1507 2867
rect 1673 2853 1687 2867
rect 1833 2853 1847 2867
rect 2853 2853 2867 2867
rect 3253 2853 3267 2867
rect 3773 2853 3787 2867
rect 4033 2853 4047 2867
rect 4853 2853 4867 2867
rect 5153 2853 5167 2867
rect 5313 2873 5327 2887
rect 5733 2853 5747 2867
rect 1733 2833 1747 2847
rect 373 2813 387 2827
rect 733 2813 747 2827
rect 773 2813 787 2827
rect 913 2813 927 2827
rect 2013 2833 2027 2847
rect 2653 2833 2667 2847
rect 2713 2833 2727 2847
rect 3193 2833 3207 2847
rect 3233 2833 3247 2847
rect 3533 2833 3547 2847
rect 4513 2833 4527 2847
rect 4653 2833 4667 2847
rect 4693 2833 4707 2847
rect 4773 2833 4787 2847
rect 5213 2833 5227 2847
rect 5633 2833 5647 2847
rect 5833 2833 5847 2847
rect 5893 2833 5907 2847
rect 5933 2833 5947 2847
rect 2033 2813 2047 2827
rect 2073 2813 2087 2827
rect 2153 2813 2167 2827
rect 2373 2813 2387 2827
rect 2513 2813 2527 2827
rect 3073 2813 3087 2827
rect 813 2793 827 2807
rect 1953 2793 1967 2807
rect 2673 2793 2687 2807
rect 2713 2793 2727 2807
rect 3433 2813 3447 2827
rect 4253 2813 4267 2827
rect 4393 2813 4407 2827
rect 3933 2793 3947 2807
rect 3993 2793 4007 2807
rect 4653 2793 4667 2807
rect 4693 2793 4707 2807
rect 4733 2793 4747 2807
rect 5073 2793 5087 2807
rect 5113 2793 5127 2807
rect 5213 2793 5227 2807
rect 5253 2793 5267 2807
rect 5493 2793 5507 2807
rect 5533 2793 5547 2807
rect 5633 2793 5647 2807
rect 5673 2793 5687 2807
rect 5933 2793 5947 2807
rect 5973 2793 5987 2807
rect 213 2773 227 2787
rect 333 2773 347 2787
rect 373 2773 387 2787
rect 413 2773 427 2787
rect 633 2773 647 2787
rect 673 2773 687 2787
rect 773 2773 787 2787
rect 953 2773 967 2787
rect 1193 2773 1207 2787
rect 1613 2773 1627 2787
rect 1653 2773 1667 2787
rect 1713 2773 1727 2787
rect 2113 2773 2127 2787
rect 2233 2773 2247 2787
rect 2293 2773 2307 2787
rect 2473 2773 2487 2787
rect 2793 2773 2807 2787
rect 2893 2773 2907 2787
rect 2953 2773 2967 2787
rect 3153 2773 3167 2787
rect 3233 2773 3247 2787
rect 3453 2773 3467 2787
rect 3513 2773 3527 2787
rect 3613 2773 3627 2787
rect 3653 2773 3667 2787
rect 3793 2773 3807 2787
rect 3913 2773 3927 2787
rect 4033 2773 4047 2787
rect 4153 2773 4167 2787
rect 4193 2773 4207 2787
rect 4233 2773 4247 2787
rect 4333 2773 4347 2787
rect 4393 2773 4407 2787
rect 4553 2773 4567 2787
rect 4773 2773 4787 2787
rect 4973 2773 4987 2787
rect 5333 2773 5347 2787
rect 5813 2773 5827 2787
rect 33 2733 47 2747
rect 453 2733 467 2747
rect 533 2733 547 2747
rect 1073 2733 1087 2747
rect 1133 2733 1147 2747
rect 1313 2733 1327 2747
rect 1373 2733 1387 2747
rect 1433 2733 1447 2747
rect 1493 2733 1507 2747
rect 1933 2733 1947 2747
rect 2073 2733 2087 2747
rect 2353 2733 2367 2747
rect 2773 2733 2787 2747
rect 3033 2733 3047 2747
rect 4733 2733 4747 2747
rect 5132 2733 5146 2747
rect 5154 2733 5168 2747
rect 5433 2733 5447 2747
rect 5553 2733 5567 2747
rect 5853 2733 5867 2747
rect 5893 2733 5907 2747
rect 93 2713 107 2727
rect 353 2713 367 2727
rect 393 2713 407 2727
rect 753 2713 767 2727
rect 893 2713 907 2727
rect 1733 2713 1747 2727
rect 33 2693 47 2707
rect 1373 2693 1387 2707
rect 1433 2693 1447 2707
rect 2093 2713 2107 2727
rect 2393 2713 2407 2727
rect 2433 2713 2447 2727
rect 2513 2713 2527 2727
rect 2553 2713 2567 2727
rect 2813 2713 2827 2727
rect 2853 2713 2867 2727
rect 1993 2693 2007 2707
rect 2993 2693 3007 2707
rect 3253 2713 3267 2727
rect 3293 2713 3307 2727
rect 3433 2713 3447 2727
rect 3473 2713 3487 2727
rect 3593 2713 3607 2727
rect 3633 2713 3647 2727
rect 3733 2713 3747 2727
rect 3773 2713 3787 2727
rect 3893 2713 3907 2727
rect 3933 2713 3947 2727
rect 3973 2713 3987 2727
rect 4213 2713 4227 2727
rect 4253 2713 4267 2727
rect 4293 2713 4307 2727
rect 4493 2713 4507 2727
rect 4793 2713 4807 2727
rect 4833 2713 4847 2727
rect 5053 2713 5067 2727
rect 5353 2713 5367 2727
rect 5393 2713 5407 2727
rect 333 2673 347 2687
rect 2473 2673 2487 2687
rect 2853 2673 2867 2687
rect 3393 2673 3407 2687
rect 3473 2673 3487 2687
rect 3633 2673 3647 2687
rect 3733 2673 3747 2687
rect 3893 2673 3907 2687
rect 4773 2693 4787 2707
rect 5633 2693 5647 2707
rect 5853 2693 5867 2707
rect 5973 2693 5987 2707
rect 4693 2673 4707 2687
rect 4853 2673 4867 2687
rect 4893 2673 4907 2687
rect 5253 2673 5267 2687
rect 5513 2673 5527 2687
rect 5893 2673 5907 2687
rect 1633 2653 1647 2667
rect 2233 2653 2247 2667
rect 3153 2653 3167 2667
rect 4153 2653 4167 2667
rect 4653 2653 4667 2667
rect 4833 2653 4847 2667
rect 4973 2653 4987 2667
rect 5293 2653 5307 2667
rect 393 2633 407 2647
rect 593 2633 607 2647
rect 1013 2633 1027 2647
rect 2153 2633 2167 2647
rect 2213 2633 2227 2647
rect 2753 2633 2767 2647
rect 2953 2633 2967 2647
rect 3593 2633 3607 2647
rect 3793 2633 3807 2647
rect 3853 2633 3867 2647
rect 3973 2633 3987 2647
rect 1073 2613 1087 2627
rect 1313 2613 1327 2627
rect 1653 2613 1667 2627
rect 1733 2613 1747 2627
rect 2553 2613 2567 2627
rect 2693 2613 2707 2627
rect 3113 2613 3127 2627
rect 3153 2613 3167 2627
rect 4593 2633 4607 2647
rect 4853 2633 4867 2647
rect 5393 2633 5407 2647
rect 4893 2613 4907 2627
rect 5433 2613 5447 2627
rect 1433 2593 1447 2607
rect 1833 2593 1847 2607
rect 2273 2593 2287 2607
rect 2653 2593 2667 2607
rect 2753 2593 2767 2607
rect 3033 2593 3047 2607
rect 5353 2593 5367 2607
rect 5573 2593 5587 2607
rect 273 2573 287 2587
rect 453 2573 467 2587
rect 1133 2573 1147 2587
rect 1193 2573 1207 2587
rect 2893 2573 2907 2587
rect 3173 2573 3187 2587
rect 5633 2573 5647 2587
rect 4293 2553 4307 2567
rect 4353 2553 4367 2567
rect 4573 2553 4587 2567
rect 713 2533 727 2547
rect 873 2533 887 2547
rect 1273 2533 1287 2547
rect 1833 2533 1847 2547
rect 1873 2533 1887 2547
rect 2353 2533 2367 2547
rect 3033 2533 3047 2547
rect 3073 2533 3087 2547
rect 4333 2533 4347 2547
rect 4393 2533 4407 2547
rect 4733 2533 4747 2547
rect 4813 2533 4827 2547
rect 5133 2534 5147 2548
rect 5253 2533 5267 2547
rect 5293 2533 5307 2547
rect 5433 2533 5447 2547
rect 1493 2513 1507 2527
rect 1533 2513 1547 2527
rect 1653 2513 1667 2527
rect 3453 2513 3467 2527
rect 3653 2513 3667 2527
rect 4233 2513 4247 2527
rect 4493 2513 4507 2527
rect 4993 2513 5007 2527
rect 5053 2513 5067 2527
rect 5133 2512 5147 2526
rect 333 2493 347 2507
rect 573 2493 587 2507
rect 713 2493 727 2507
rect 753 2493 767 2507
rect 973 2493 987 2507
rect 1133 2493 1147 2507
rect 1173 2493 1187 2507
rect 1233 2493 1247 2507
rect 1273 2493 1287 2507
rect 1313 2493 1327 2507
rect 1433 2493 1447 2507
rect 1473 2493 1487 2507
rect 1873 2493 1887 2507
rect 1913 2493 1927 2507
rect 2013 2493 2027 2507
rect 2053 2493 2067 2507
rect 2113 2493 2127 2507
rect 2153 2493 2167 2507
rect 2193 2493 2207 2507
rect 2313 2493 2327 2507
rect 2353 2493 2367 2507
rect 2613 2493 2627 2507
rect 2653 2493 2667 2507
rect 2993 2493 3007 2507
rect 3033 2493 3047 2507
rect 3133 2493 3147 2507
rect 3173 2493 3187 2507
rect 3693 2493 3707 2507
rect 3733 2493 3747 2507
rect 3833 2493 3847 2507
rect 3873 2493 3887 2507
rect 3993 2493 4007 2507
rect 4353 2493 4367 2507
rect 4393 2493 4407 2507
rect 4573 2493 4587 2507
rect 4653 2493 4667 2507
rect 4693 2493 4707 2507
rect 4813 2493 4827 2507
rect 4853 2493 4867 2507
rect 5393 2493 5407 2507
rect 5433 2493 5447 2507
rect 5613 2493 5627 2507
rect 5713 2493 5727 2507
rect 5753 2493 5767 2507
rect 133 2473 147 2487
rect 213 2473 227 2487
rect 273 2473 287 2487
rect 793 2473 807 2487
rect 933 2473 947 2487
rect 1073 2473 1087 2487
rect 1713 2473 1727 2487
rect 1833 2473 1847 2487
rect 2573 2473 2587 2487
rect 2813 2473 2827 2487
rect 2873 2473 2887 2487
rect 3253 2473 3267 2487
rect 3313 2473 3327 2487
rect 4173 2473 4187 2487
rect 4233 2473 4247 2487
rect 4433 2473 4447 2487
rect 4933 2473 4947 2487
rect 4993 2473 5007 2487
rect 5213 2473 5227 2487
rect 5293 2473 5307 2487
rect 5473 2473 5487 2487
rect 5813 2473 5827 2487
rect 5873 2473 5887 2487
rect 1793 2453 1807 2467
rect 1853 2453 1867 2467
rect 33 2433 47 2447
rect 453 2433 467 2447
rect 593 2433 607 2447
rect 733 2433 747 2447
rect 993 2433 1007 2447
rect 1234 2433 1248 2447
rect 1333 2433 1347 2447
rect 1373 2433 1387 2447
rect 1493 2433 1507 2447
rect 1993 2433 2007 2447
rect 2533 2433 2547 2447
rect 2633 2433 2647 2447
rect 2693 2433 2707 2447
rect 2973 2433 2987 2447
rect 3153 2433 3167 2447
rect 3213 2433 3227 2447
rect 3433 2433 3447 2447
rect 3813 2433 3827 2447
rect 3853 2433 3867 2447
rect 3893 2433 3907 2447
rect 3973 2433 3987 2447
rect 4053 2433 4067 2447
rect 4333 2433 4347 2447
rect 4413 2433 4427 2447
rect 4673 2433 4687 2447
rect 4733 2433 4747 2447
rect 4833 2433 4847 2447
rect 4913 2433 4927 2447
rect 5113 2433 5127 2447
rect 5533 2433 5547 2447
rect 5593 2433 5607 2447
rect 5653 2433 5667 2447
rect 5693 2433 5707 2447
rect 5753 2433 5767 2447
rect 5993 2433 6007 2447
rect 693 2413 707 2427
rect 853 2413 867 2427
rect 893 2413 907 2427
rect 733 2393 747 2407
rect 793 2393 807 2407
rect 933 2393 947 2407
rect 993 2393 1007 2407
rect 1113 2393 1127 2407
rect 1493 2393 1507 2407
rect 1653 2413 1667 2427
rect 1733 2413 1747 2427
rect 1773 2413 1787 2427
rect 1813 2393 1827 2407
rect 2173 2413 2187 2427
rect 2333 2413 2347 2427
rect 2433 2413 2447 2427
rect 2493 2413 2507 2427
rect 3013 2413 3027 2427
rect 3473 2413 3487 2427
rect 3573 2413 3587 2427
rect 2313 2393 2327 2407
rect 3173 2393 3187 2407
rect 3233 2393 3247 2407
rect 3813 2393 3827 2407
rect 3853 2393 3867 2407
rect 4513 2413 4527 2427
rect 4553 2413 4567 2427
rect 5233 2413 5247 2427
rect 5273 2413 5287 2427
rect 4673 2393 4687 2407
rect 5313 2393 5327 2407
rect 5473 2393 5487 2407
rect 5533 2393 5547 2407
rect 5592 2393 5606 2407
rect 5614 2393 5628 2407
rect 5713 2393 5727 2407
rect 753 2373 767 2387
rect 973 2373 987 2387
rect 1293 2373 1307 2387
rect 1533 2373 1547 2387
rect 1773 2373 1787 2387
rect 4433 2373 4447 2387
rect 4633 2373 4647 2387
rect 4773 2373 4787 2387
rect 5493 2373 5507 2387
rect 173 2353 187 2367
rect 213 2353 227 2367
rect 273 2353 287 2367
rect 453 2353 467 2367
rect 593 2353 607 2367
rect 1173 2353 1187 2367
rect 1373 2353 1387 2367
rect 1473 2353 1487 2367
rect 1633 2353 1647 2367
rect 1973 2353 1987 2367
rect 2233 2353 2247 2367
rect 2373 2353 2387 2367
rect 2493 2353 2507 2367
rect 2753 2353 2767 2367
rect 2833 2353 2847 2367
rect 3173 2353 3187 2367
rect 3213 2353 3227 2367
rect 3313 2353 3327 2367
rect 3373 2353 3387 2367
rect 3513 2353 3527 2367
rect 3833 2353 3847 2367
rect 4013 2353 4027 2367
rect 4253 2353 4267 2367
rect 4913 2353 4927 2367
rect 1313 2333 1327 2347
rect 1393 2333 1407 2347
rect 1433 2333 1447 2347
rect 1813 2333 1827 2347
rect 2593 2333 2607 2347
rect 2873 2333 2887 2347
rect 2953 2333 2967 2347
rect 3073 2333 3087 2347
rect 3133 2333 3147 2347
rect 3253 2334 3267 2348
rect 5713 2353 5727 2367
rect 5773 2353 5787 2367
rect 5813 2353 5827 2367
rect 3353 2333 3367 2347
rect 3573 2333 3587 2347
rect 3913 2333 3927 2347
rect 3973 2333 3987 2347
rect 4573 2333 4587 2347
rect 5233 2333 5247 2347
rect 5553 2333 5567 2347
rect 573 2313 587 2327
rect 1453 2313 1467 2327
rect 1593 2313 1607 2327
rect 2273 2313 2287 2327
rect 2313 2313 2327 2327
rect 2753 2313 2767 2327
rect 2913 2313 2927 2327
rect 3253 2312 3267 2326
rect 3413 2313 3427 2327
rect 4053 2313 4067 2327
rect 4213 2313 4227 2327
rect 4313 2313 4327 2327
rect 5753 2313 5767 2327
rect 5813 2313 5827 2327
rect 593 2293 607 2307
rect 753 2293 767 2307
rect 1393 2293 1407 2307
rect 1633 2293 1647 2307
rect 1753 2293 1767 2307
rect 1973 2293 1987 2307
rect 2113 2293 2127 2307
rect 2193 2293 2207 2307
rect 973 2273 987 2287
rect 1073 2273 1087 2287
rect 2833 2293 2847 2307
rect 2893 2293 2907 2307
rect 4513 2293 4527 2307
rect 4573 2293 4587 2307
rect 5073 2293 5087 2307
rect 2273 2273 2287 2287
rect 2373 2273 2387 2287
rect 2693 2273 2707 2287
rect 2753 2273 2767 2287
rect 3413 2273 3427 2287
rect 3453 2273 3467 2287
rect 3973 2273 3987 2287
rect 4053 2273 4067 2287
rect 4253 2273 4267 2287
rect 4313 2273 4327 2287
rect 4593 2273 4607 2287
rect 4633 2273 4647 2287
rect 5293 2273 5307 2287
rect 5333 2273 5347 2287
rect 5413 2293 5427 2307
rect 5733 2293 5747 2307
rect 5873 2293 5887 2307
rect 5913 2293 5927 2307
rect 5953 2293 5967 2307
rect 5853 2273 5867 2287
rect 33 2253 47 2267
rect 73 2253 87 2267
rect 233 2253 247 2267
rect 353 2253 367 2267
rect 753 2253 767 2267
rect 793 2253 807 2267
rect 1113 2253 1127 2267
rect 1153 2253 1167 2267
rect 1373 2253 1387 2267
rect 1413 2253 1427 2267
rect 1473 2253 1487 2267
rect 1593 2253 1607 2267
rect 1633 2253 1647 2267
rect 1753 2253 1767 2267
rect 1813 2253 1827 2267
rect 2093 2253 2107 2267
rect 2413 2253 2427 2267
rect 2813 2253 2827 2267
rect 2893 2253 2907 2267
rect 3133 2253 3147 2267
rect 3253 2253 3267 2267
rect 3493 2253 3507 2267
rect 3913 2253 3927 2267
rect 4433 2253 4447 2267
rect 4553 2253 4567 2267
rect 4773 2253 4787 2267
rect 5053 2253 5067 2267
rect 5113 2253 5127 2267
rect 5253 2253 5267 2267
rect 5413 2253 5427 2267
rect 5633 2253 5647 2267
rect 5673 2253 5687 2267
rect 5813 2253 5827 2267
rect 5893 2253 5907 2267
rect 5993 2253 6007 2267
rect 5273 2233 5287 2247
rect 373 2213 387 2227
rect 513 2213 527 2227
rect 573 2213 587 2227
rect 913 2213 927 2227
rect 973 2213 987 2227
rect 1193 2213 1207 2227
rect 1313 2213 1327 2227
rect 1813 2213 1827 2227
rect 2073 2213 2087 2227
rect 2113 2213 2127 2227
rect 2373 2213 2387 2227
rect 2533 2213 2547 2227
rect 2593 2213 2607 2227
rect 2813 2213 2827 2227
rect 2953 2213 2967 2227
rect 3013 2213 3027 2227
rect 3313 2213 3327 2227
rect 3613 2213 3627 2227
rect 3673 2213 3687 2227
rect 3733 2213 3747 2227
rect 3813 2213 3827 2227
rect 4273 2213 4287 2227
rect 4573 2213 4587 2227
rect 4653 2213 4667 2227
rect 4793 2213 4807 2227
rect 4873 2213 4887 2227
rect 4993 2213 5007 2227
rect 5353 2213 5367 2227
rect 93 2193 107 2207
rect 113 2193 127 2207
rect 353 2193 367 2207
rect 733 2193 747 2207
rect 1093 2193 1107 2207
rect 1133 2193 1147 2207
rect 1493 2193 1507 2207
rect 213 2173 227 2187
rect 1613 2193 1627 2207
rect 1653 2193 1667 2207
rect 1693 2193 1707 2207
rect 1753 2193 1767 2207
rect 1893 2193 1907 2207
rect 1933 2193 1947 2207
rect 2873 2193 2887 2207
rect 2913 2193 2927 2207
rect 3173 2193 3187 2207
rect 3233 2193 3247 2207
rect 3273 2193 3287 2207
rect 4033 2193 4047 2207
rect 4213 2193 4227 2207
rect 4413 2193 4427 2207
rect 4453 2193 4467 2207
rect 4513 2193 4527 2207
rect 4613 2193 4627 2207
rect 4753 2193 4767 2207
rect 5193 2193 5207 2207
rect 5433 2193 5447 2207
rect 5553 2193 5567 2207
rect 5593 2193 5607 2207
rect 5793 2193 5807 2207
rect 5833 2193 5847 2207
rect 5873 2193 5887 2207
rect 5913 2193 5927 2207
rect 1593 2173 1607 2187
rect 3473 2173 3487 2187
rect 3553 2173 3567 2187
rect 3613 2173 3627 2187
rect 733 2153 747 2167
rect 1473 2153 1487 2167
rect 1573 2153 1587 2167
rect 1813 2153 1827 2167
rect 1893 2153 1907 2167
rect 1933 2153 1947 2167
rect 2273 2153 2287 2167
rect 3213 2153 3227 2167
rect 3253 2153 3267 2167
rect 4413 2153 4427 2167
rect 4753 2153 4767 2167
rect 5353 2153 5367 2167
rect 5393 2153 5407 2167
rect 5433 2153 5447 2167
rect 5873 2153 5887 2167
rect 5973 2153 5987 2167
rect 4653 2133 4667 2147
rect 4793 2133 4807 2147
rect 733 2113 747 2127
rect 1133 2113 1147 2127
rect 1193 2113 1207 2127
rect 1233 2113 1247 2127
rect 2073 2113 2087 2127
rect 2133 2113 2147 2127
rect 3253 2113 3267 2127
rect 3393 2113 3407 2127
rect 4833 2113 4847 2127
rect 4993 2113 5007 2127
rect 5193 2113 5207 2127
rect 5873 2113 5887 2127
rect 973 2093 987 2107
rect 1213 2093 1227 2107
rect 1413 2093 1427 2107
rect 1533 2093 1547 2107
rect 3113 2093 3127 2107
rect 3493 2093 3507 2107
rect 3733 2093 3747 2107
rect 4173 2093 4187 2107
rect 4233 2093 4247 2107
rect 4733 2093 4747 2107
rect 4873 2093 4887 2107
rect 4933 2093 4947 2107
rect 5473 2093 5487 2107
rect 5773 2093 5787 2107
rect 5813 2093 5827 2107
rect 513 2073 527 2087
rect 673 2073 687 2087
rect 1093 2073 1107 2087
rect 1553 2073 1567 2087
rect 1613 2073 1627 2087
rect 2113 2073 2127 2087
rect 2633 2073 2647 2087
rect 3153 2073 3167 2087
rect 3853 2073 3867 2087
rect 4313 2073 4327 2087
rect 5753 2073 5767 2087
rect 233 2053 247 2067
rect 433 2053 447 2067
rect 693 2053 707 2067
rect 1153 2053 1167 2067
rect 1333 2053 1347 2067
rect 1473 2053 1487 2067
rect 2273 2053 2287 2067
rect 2713 2053 2727 2067
rect 2953 2053 2967 2067
rect 3313 2053 3327 2067
rect 3353 2053 3367 2067
rect 3573 2053 3587 2067
rect 3693 2053 3707 2067
rect 4813 2053 4827 2067
rect 5233 2053 5247 2067
rect 5433 2053 5447 2067
rect 5513 2053 5527 2067
rect 5953 2053 5967 2067
rect 193 2033 207 2047
rect 853 2033 867 2047
rect 1313 2033 1327 2047
rect 2333 2033 2347 2047
rect 2493 2033 2507 2047
rect 293 2013 307 2027
rect 1293 2013 1307 2027
rect 1373 2013 1387 2027
rect 2373 2013 2387 2027
rect 2453 2013 2467 2027
rect 5273 2013 5287 2027
rect 5393 2013 5407 2027
rect 1213 1993 1227 2007
rect 1313 1993 1327 2007
rect 1773 1993 1787 2007
rect 1833 1993 1847 2007
rect 1893 1993 1907 2007
rect 1993 1993 2007 2007
rect 3693 1993 3707 2007
rect 253 1973 267 1987
rect 293 1973 307 1987
rect 393 1973 407 1987
rect 433 1973 447 1987
rect 673 1973 687 1987
rect 713 1973 727 1987
rect 813 1973 827 1987
rect 853 1973 867 1987
rect 973 1973 987 1987
rect 1253 1973 1267 1987
rect 1333 1973 1347 1987
rect 1373 1973 1387 1987
rect 1473 1973 1487 1987
rect 1513 1973 1527 1987
rect 2033 1973 2047 1987
rect 2073 1973 2087 1987
rect 2413 1973 2427 1987
rect 2453 1973 2467 1987
rect 2993 1973 3007 1987
rect 3413 1973 3427 1987
rect 3453 1973 3467 1987
rect 4613 1993 4627 2007
rect 4673 1993 4687 2007
rect 4073 1973 4087 1987
rect 4113 1973 4127 1987
rect 4373 1973 4387 1987
rect 4493 1973 4507 1987
rect 4833 1973 4847 1987
rect 4873 1973 4887 1987
rect 5233 1973 5247 1987
rect 5273 1973 5287 1987
rect 113 1953 127 1967
rect 1153 1953 1167 1967
rect 1213 1953 1227 1967
rect 1693 1953 1707 1967
rect 1833 1953 1847 1967
rect 1893 1953 1907 1967
rect 2113 1953 2127 1967
rect 2313 1953 2327 1967
rect 2533 1953 2547 1967
rect 2593 1953 2607 1967
rect 2893 1953 2907 1967
rect 2953 1953 2967 1967
rect 3253 1953 3267 1967
rect 3313 1953 3327 1967
rect 3593 1953 3607 1967
rect 3693 1953 3707 1967
rect 3953 1953 3967 1967
rect 4173 1953 4187 1967
rect 4233 1953 4247 1967
rect 4673 1953 4687 1967
rect 4733 1953 4747 1967
rect 4933 1953 4947 1967
rect 4993 1953 5007 1967
rect 5433 1953 5447 1967
rect 5473 1953 5487 1967
rect 5533 1953 5547 1967
rect 5773 1953 5787 1967
rect 5813 1953 5827 1967
rect 193 1913 207 1927
rect 273 1913 287 1927
rect 313 1913 327 1927
rect 453 1913 467 1927
rect 493 1913 507 1927
rect 573 1913 587 1927
rect 613 1913 627 1927
rect 653 1913 667 1927
rect 793 1913 807 1927
rect 913 1913 927 1927
rect 953 1913 967 1927
rect 1033 1913 1047 1927
rect 1233 1913 1247 1927
rect 1553 1913 1567 1927
rect 1713 1913 1727 1927
rect 1973 1913 1987 1927
rect 2053 1913 2067 1927
rect 2433 1913 2447 1927
rect 2713 1913 2727 1927
rect 2773 1913 2787 1927
rect 3073 1913 3087 1927
rect 3513 1913 3527 1927
rect 4053 1913 4067 1927
rect 4153 1913 4167 1927
rect 4353 1913 4367 1927
rect 4433 1913 4447 1927
rect 4553 1913 4567 1927
rect 4813 1913 4827 1927
rect 5113 1913 5127 1927
rect 5253 1913 5267 1927
rect 5293 1913 5307 1927
rect 5653 1913 5667 1927
rect 93 1893 107 1907
rect 153 1893 167 1907
rect 293 1893 307 1907
rect 353 1893 367 1907
rect 1353 1893 1367 1907
rect 1533 1893 1547 1907
rect 1633 1893 1647 1907
rect 1673 1893 1687 1907
rect 1893 1893 1907 1907
rect 2093 1893 2107 1907
rect 2353 1893 2367 1907
rect 2393 1893 2407 1907
rect 2473 1893 2487 1907
rect 3133 1893 3147 1907
rect 3433 1893 3447 1907
rect 3833 1893 3847 1907
rect 3953 1893 3967 1907
rect 5393 1893 5407 1907
rect 5433 1893 5447 1907
rect 753 1873 767 1887
rect 953 1873 967 1887
rect 1013 1873 1027 1887
rect 2373 1873 2387 1887
rect 3013 1873 3027 1887
rect 3113 1873 3127 1887
rect 5193 1873 5207 1887
rect 5253 1873 5267 1887
rect 1393 1853 1407 1867
rect 1613 1853 1627 1867
rect 1673 1853 1687 1867
rect 1913 1853 1927 1867
rect 2113 1853 2127 1867
rect 2513 1853 2527 1867
rect 3453 1853 3467 1867
rect 3493 1853 3507 1867
rect 5353 1853 5367 1867
rect 5393 1853 5407 1867
rect 373 1833 387 1847
rect 973 1833 987 1847
rect 1233 1833 1247 1847
rect 533 1813 547 1827
rect 913 1813 927 1827
rect 993 1813 1007 1827
rect 1153 1813 1167 1827
rect 1353 1833 1367 1847
rect 1773 1833 1787 1847
rect 1953 1833 1967 1847
rect 2273 1833 2287 1847
rect 2433 1833 2447 1847
rect 1333 1813 1347 1827
rect 1913 1813 1927 1827
rect 2053 1813 2067 1827
rect 2133 1813 2147 1827
rect 2473 1813 2487 1827
rect 2573 1813 2587 1827
rect 2613 1833 2627 1847
rect 2773 1833 2787 1847
rect 3213 1833 3227 1847
rect 3273 1833 3287 1847
rect 3353 1833 3367 1847
rect 3473 1833 3487 1847
rect 2893 1813 2907 1827
rect 4053 1833 4067 1847
rect 4373 1833 4387 1847
rect 4873 1833 4887 1847
rect 4953 1833 4967 1847
rect 5113 1833 5127 1847
rect 5613 1833 5627 1847
rect 5653 1833 5667 1847
rect 5793 1833 5807 1847
rect 153 1793 167 1807
rect 573 1793 587 1807
rect 653 1793 667 1807
rect 1673 1793 1687 1807
rect 1733 1793 1747 1807
rect 1833 1793 1847 1807
rect 1893 1793 1907 1807
rect 2553 1793 2567 1807
rect 2873 1793 2887 1807
rect 2933 1793 2947 1807
rect 2993 1793 3007 1807
rect 3373 1793 3387 1807
rect 3473 1793 3487 1807
rect 3593 1813 3607 1827
rect 3633 1813 3647 1827
rect 3893 1813 3907 1827
rect 4113 1813 4127 1827
rect 4433 1813 4447 1827
rect 5293 1813 5307 1827
rect 5493 1813 5507 1827
rect 5973 1813 5987 1827
rect 4033 1793 4047 1807
rect 4153 1793 4167 1807
rect 4193 1793 4207 1807
rect 4273 1793 4287 1807
rect 4353 1793 4367 1807
rect 4473 1793 4487 1807
rect 5733 1793 5747 1807
rect 5913 1793 5927 1807
rect 93 1773 107 1787
rect 213 1753 227 1767
rect 473 1753 487 1767
rect 613 1773 627 1787
rect 753 1773 767 1787
rect 1153 1773 1167 1787
rect 1333 1773 1347 1787
rect 1533 1773 1547 1787
rect 1873 1773 1887 1787
rect 2593 1773 2607 1787
rect 2633 1773 2647 1787
rect 873 1753 887 1767
rect 2553 1753 2567 1767
rect 2933 1753 2947 1767
rect 3073 1753 3087 1767
rect 3193 1773 3207 1787
rect 3513 1773 3527 1787
rect 4453 1773 4467 1787
rect 4673 1773 4687 1787
rect 3893 1753 3907 1767
rect 4153 1753 4167 1767
rect 4193 1753 4207 1767
rect 4553 1753 4567 1767
rect 4993 1773 5007 1787
rect 5293 1773 5307 1787
rect 5453 1773 5467 1787
rect 5533 1773 5547 1787
rect 5733 1753 5747 1767
rect 5793 1753 5807 1767
rect 5873 1753 5887 1767
rect 253 1733 267 1747
rect 293 1733 307 1747
rect 573 1733 587 1747
rect 613 1733 627 1747
rect 913 1733 927 1747
rect 953 1733 967 1747
rect 1233 1733 1247 1747
rect 1273 1733 1287 1747
rect 1313 1733 1327 1747
rect 1473 1733 1487 1747
rect 1813 1733 1827 1747
rect 1873 1733 1887 1747
rect 1913 1733 1927 1747
rect 2133 1733 2147 1747
rect 2273 1733 2287 1747
rect 2353 1733 2367 1747
rect 2513 1733 2527 1747
rect 2593 1733 2607 1747
rect 2673 1733 2687 1747
rect 2813 1733 2827 1747
rect 3193 1733 3207 1747
rect 3313 1733 3327 1747
rect 3353 1733 3367 1747
rect 3413 1733 3427 1747
rect 3473 1733 3487 1747
rect 3753 1733 3767 1747
rect 3853 1733 3867 1747
rect 3933 1733 3947 1747
rect 4533 1733 4547 1747
rect 4673 1733 4687 1747
rect 4773 1733 4787 1747
rect 5093 1733 5107 1747
rect 5213 1733 5227 1747
rect 5253 1733 5267 1747
rect 5293 1733 5307 1747
rect 5453 1733 5467 1747
rect 5493 1733 5507 1747
rect 5613 1733 5627 1747
rect 5973 1733 5987 1747
rect 3393 1713 3407 1727
rect 153 1693 167 1707
rect 413 1693 427 1707
rect 473 1693 487 1707
rect 673 1693 687 1707
rect 1133 1693 1147 1707
rect 2033 1693 2047 1707
rect 2093 1693 2107 1707
rect 2873 1693 2887 1707
rect 3533 1693 3547 1707
rect 3573 1693 3587 1707
rect 3633 1693 3647 1707
rect 4133 1693 4147 1707
rect 4313 1693 4327 1707
rect 5773 1693 5787 1707
rect 5813 1693 5827 1707
rect 233 1673 247 1687
rect 593 1673 607 1687
rect 633 1673 647 1687
rect 893 1673 907 1687
rect 1073 1673 1087 1687
rect 1253 1673 1267 1687
rect 1453 1673 1467 1687
rect 1533 1673 1547 1687
rect 1573 1673 1587 1687
rect 1613 1673 1627 1687
rect 1653 1673 1667 1687
rect 1693 1673 1707 1687
rect 1853 1673 1867 1687
rect 2213 1673 2227 1687
rect 2253 1673 2267 1687
rect 2533 1673 2547 1687
rect 2573 1673 2587 1687
rect 2633 1673 2647 1687
rect 2833 1673 2847 1687
rect 3213 1673 3227 1687
rect 3293 1673 3307 1687
rect 3333 1673 3347 1687
rect 3373 1673 3387 1687
rect 3873 1673 3887 1687
rect 3913 1673 3927 1687
rect 4053 1673 4067 1687
rect 4593 1673 4607 1687
rect 4653 1673 4667 1687
rect 4693 1673 4707 1687
rect 4733 1673 4747 1687
rect 4853 1673 4867 1687
rect 4953 1673 4967 1687
rect 4993 1673 5007 1687
rect 5033 1673 5047 1687
rect 5133 1673 5147 1687
rect 5173 1673 5187 1687
rect 5233 1673 5247 1687
rect 5273 1673 5287 1687
rect 5313 1673 5327 1687
rect 5433 1673 5447 1687
rect 5473 1673 5487 1687
rect 5513 1673 5527 1687
rect 5593 1673 5607 1687
rect 1133 1653 1147 1667
rect 233 1633 247 1647
rect 533 1633 547 1647
rect 593 1633 607 1647
rect 1292 1633 1306 1647
rect 1693 1633 1707 1647
rect 2273 1653 2287 1667
rect 2313 1653 2327 1667
rect 2373 1653 2387 1667
rect 3533 1653 3547 1667
rect 1893 1633 1907 1647
rect 2393 1633 2407 1647
rect 2613 1633 2627 1647
rect 2773 1633 2787 1647
rect 3293 1633 3307 1647
rect 3373 1633 3387 1647
rect 3433 1633 3447 1647
rect 3773 1633 3787 1647
rect 1193 1613 1207 1627
rect 1313 1613 1327 1627
rect 1733 1613 1747 1627
rect 1833 1613 1847 1627
rect 2253 1613 2267 1627
rect 2293 1613 2307 1627
rect 2573 1613 2587 1627
rect 813 1593 827 1607
rect 1333 1593 1347 1607
rect 1753 1593 1767 1607
rect 1853 1593 1867 1607
rect 1953 1593 1967 1607
rect 2033 1593 2047 1607
rect 2133 1593 2147 1607
rect 2173 1593 2187 1607
rect 2733 1613 2747 1627
rect 2833 1613 2847 1627
rect 3012 1613 3026 1627
rect 3213 1613 3227 1627
rect 3453 1613 3467 1627
rect 3833 1613 3847 1627
rect 4313 1613 4327 1627
rect 4753 1633 4767 1647
rect 5213 1633 5227 1647
rect 5313 1633 5327 1647
rect 5493 1633 5507 1647
rect 5593 1633 5607 1647
rect 4993 1613 5007 1627
rect 5093 1613 5107 1627
rect 5433 1613 5447 1627
rect 2633 1593 2647 1607
rect 2813 1593 2827 1607
rect 2853 1593 2867 1607
rect 3073 1593 3087 1607
rect 3233 1593 3247 1607
rect 193 1573 207 1587
rect 473 1573 487 1587
rect 633 1573 647 1587
rect 1473 1573 1487 1587
rect 1913 1573 1927 1587
rect 2053 1573 2067 1587
rect 3213 1573 3227 1587
rect 3253 1573 3267 1587
rect 3833 1573 3847 1587
rect 3873 1593 3887 1607
rect 4053 1593 4067 1607
rect 4493 1593 4507 1607
rect 4413 1573 4427 1587
rect 5033 1593 5047 1607
rect 5173 1593 5187 1607
rect 5233 1573 5247 1587
rect 5353 1573 5367 1587
rect 433 1553 447 1567
rect 893 1553 907 1567
rect 1253 1553 1267 1567
rect 1813 1553 1827 1567
rect 2213 1553 2227 1567
rect 573 1533 587 1547
rect 673 1533 687 1547
rect 733 1533 747 1547
rect 933 1533 947 1547
rect 1273 1533 1287 1547
rect 1553 1533 1567 1547
rect 1673 1533 1687 1547
rect 2093 1533 2107 1547
rect 2773 1553 2787 1567
rect 2413 1533 2427 1547
rect 273 1513 287 1527
rect 373 1513 387 1527
rect 1773 1513 1787 1527
rect 1873 1513 1887 1527
rect 1993 1513 2007 1527
rect 2173 1513 2187 1527
rect 2813 1533 2827 1547
rect 2873 1533 2887 1547
rect 3173 1553 3187 1567
rect 3033 1533 3047 1547
rect 3373 1553 3387 1567
rect 3733 1553 3747 1567
rect 4093 1553 4107 1567
rect 4593 1553 4607 1567
rect 5613 1553 5627 1567
rect 3293 1533 3307 1547
rect 3493 1533 3507 1547
rect 4452 1533 4466 1547
rect 4474 1533 4488 1547
rect 4693 1533 4707 1547
rect 4813 1533 4827 1547
rect 4853 1533 4867 1547
rect 4953 1533 4967 1547
rect 5073 1533 5087 1547
rect 5733 1533 5747 1547
rect 5773 1533 5787 1547
rect 3413 1513 3427 1527
rect 3653 1513 3667 1527
rect 4413 1513 4427 1527
rect 4773 1513 4787 1527
rect 5033 1513 5047 1527
rect 5093 1513 5107 1527
rect 93 1493 107 1507
rect 253 1493 267 1507
rect 1653 1493 1667 1507
rect 2113 1493 2127 1507
rect 2253 1493 2267 1507
rect 2313 1493 2327 1507
rect 2353 1493 2367 1507
rect 2733 1493 2747 1507
rect 2872 1493 2886 1507
rect 2894 1493 2908 1507
rect 2993 1493 3007 1507
rect 3093 1493 3107 1507
rect 3533 1493 3547 1507
rect 3593 1493 3607 1507
rect 4213 1493 4227 1507
rect 333 1473 347 1487
rect 433 1473 447 1487
rect 833 1473 847 1487
rect 893 1473 907 1487
rect 1753 1473 1767 1487
rect 1893 1473 1907 1487
rect 2033 1473 2047 1487
rect 2593 1473 2607 1487
rect 3333 1473 3347 1487
rect 3513 1473 3527 1487
rect 4433 1473 4447 1487
rect 4533 1473 4547 1487
rect 4653 1473 4667 1487
rect 4693 1473 4707 1487
rect 5133 1493 5147 1507
rect 5953 1493 5967 1507
rect 5993 1493 6007 1507
rect 93 1453 107 1467
rect 133 1453 147 1467
rect 233 1453 247 1467
rect 273 1453 287 1467
rect 733 1453 747 1467
rect 913 1453 927 1467
rect 953 1453 967 1467
rect 1053 1453 1067 1467
rect 1093 1453 1107 1467
rect 1373 1453 1387 1467
rect 1493 1453 1507 1467
rect 1613 1453 1627 1467
rect 1653 1453 1667 1467
rect 1773 1453 1787 1467
rect 1813 1453 1827 1467
rect 2073 1453 2087 1467
rect 2113 1453 2127 1467
rect 2313 1453 2327 1467
rect 2393 1453 2407 1467
rect 2733 1453 2747 1467
rect 2773 1453 2787 1467
rect 2873 1453 2887 1467
rect 2993 1453 3007 1467
rect 3033 1453 3047 1467
rect 3553 1453 3567 1467
rect 3593 1453 3607 1467
rect 3693 1453 3707 1467
rect 3733 1453 3747 1467
rect 4093 1453 4107 1467
rect 4173 1453 4187 1467
rect 4213 1453 4227 1467
rect 4253 1453 4267 1467
rect 4373 1453 4387 1467
rect 4413 1453 4427 1467
rect 4813 1453 4827 1467
rect 4853 1453 4867 1467
rect 4973 1453 4987 1467
rect 5093 1453 5107 1467
rect 5133 1453 5147 1467
rect 5173 1453 5187 1467
rect 5733 1453 5747 1467
rect 5993 1453 6007 1467
rect 6033 1453 6047 1467
rect 793 1433 807 1447
rect 1273 1433 1287 1447
rect 1333 1433 1347 1447
rect 1953 1433 1967 1447
rect 2533 1433 2547 1447
rect 2593 1433 2607 1447
rect 3113 1433 3127 1447
rect 3173 1433 3187 1447
rect 3373 1433 3387 1447
rect 3793 1433 3807 1447
rect 3853 1433 3867 1447
rect 4653 1433 4667 1447
rect 5313 1433 5327 1447
rect 5373 1433 5387 1447
rect 5493 1433 5507 1447
rect 5613 1433 5627 1447
rect 5673 1433 5687 1447
rect 513 1413 527 1427
rect 213 1393 227 1407
rect 293 1393 307 1407
rect 613 1393 627 1407
rect 893 1393 907 1407
rect 933 1393 947 1407
rect 973 1393 987 1407
rect 1153 1393 1167 1407
rect 1513 1393 1527 1407
rect 1553 1393 1567 1407
rect 1673 1393 1687 1407
rect 1753 1393 1767 1407
rect 1893 1393 1907 1407
rect 2053 1393 2067 1407
rect 2133 1393 2147 1407
rect 2173 1393 2187 1407
rect 2393 1393 2407 1407
rect 2413 1393 2427 1407
rect 2613 1393 2627 1407
rect 2753 1393 2767 1407
rect 2933 1393 2947 1407
rect 3013 1393 3027 1407
rect 3293 1393 3307 1407
rect 3673 1393 3687 1407
rect 3713 1393 3727 1407
rect 3753 1393 3767 1407
rect 3973 1393 3987 1407
rect 4073 1393 4087 1407
rect 4193 1393 4207 1407
rect 4273 1393 4287 1407
rect 4433 1393 4447 1407
rect 4793 1393 4807 1407
rect 4873 1393 4887 1407
rect 5153 1393 5167 1407
rect 5193 1393 5207 1407
rect 5433 1393 5447 1407
rect 5853 1393 5867 1407
rect 5893 1393 5907 1407
rect 6013 1393 6027 1407
rect 253 1373 267 1387
rect 393 1373 407 1387
rect 433 1373 447 1387
rect 533 1373 547 1387
rect 573 1373 587 1387
rect 293 1353 307 1367
rect 333 1353 347 1367
rect 893 1353 907 1367
rect 1053 1353 1067 1367
rect 1933 1373 1947 1387
rect 1973 1373 1987 1387
rect 2333 1373 2347 1387
rect 2593 1373 2607 1387
rect 2673 1373 2687 1387
rect 2893 1373 2907 1387
rect 1613 1353 1627 1367
rect 2133 1353 2147 1367
rect 2213 1353 2227 1367
rect 3333 1373 3347 1387
rect 3433 1373 3447 1387
rect 3713 1353 3727 1367
rect 3773 1353 3787 1367
rect 4013 1353 4027 1367
rect 4433 1353 4447 1367
rect 4553 1373 4567 1387
rect 4593 1373 4607 1387
rect 4693 1373 4707 1387
rect 4833 1373 4847 1387
rect 5613 1373 5627 1387
rect 5673 1373 5687 1387
rect 1353 1333 1367 1347
rect 1393 1333 1407 1347
rect 1513 1333 1527 1347
rect 1733 1333 1747 1347
rect 1913 1333 1927 1347
rect 1953 1333 1967 1347
rect 653 1313 667 1327
rect 893 1313 907 1327
rect 1093 1313 1107 1327
rect 1153 1313 1167 1327
rect 1373 1313 1387 1327
rect 1633 1313 1647 1327
rect 2273 1313 2287 1327
rect 2653 1313 2667 1327
rect 2753 1313 2767 1327
rect 2893 1313 2907 1327
rect 93 1293 107 1307
rect 133 1293 147 1307
rect 613 1293 627 1307
rect 753 1293 767 1307
rect 913 1293 927 1307
rect 1253 1293 1267 1307
rect 1493 1293 1507 1307
rect 1773 1293 1787 1307
rect 2373 1293 2387 1307
rect 2633 1293 2647 1307
rect 3593 1333 3607 1347
rect 3753 1333 3767 1347
rect 4073 1333 4087 1347
rect 4533 1333 4547 1347
rect 4833 1333 4847 1347
rect 3113 1313 3127 1327
rect 3173 1313 3187 1327
rect 3153 1293 3167 1307
rect 3593 1293 3607 1307
rect 3653 1313 3667 1327
rect 3873 1313 3887 1327
rect 3973 1313 3987 1327
rect 5093 1313 5107 1327
rect 5153 1313 5167 1327
rect 6013 1333 6027 1347
rect 5313 1313 5327 1327
rect 5673 1313 5687 1327
rect 5893 1313 5907 1327
rect 3693 1293 3707 1307
rect 5273 1293 5287 1307
rect 5513 1293 5527 1307
rect 5813 1293 5827 1307
rect 153 1273 167 1287
rect 193 1273 207 1287
rect 673 1273 687 1287
rect 933 1273 947 1287
rect 1313 1273 1327 1287
rect 1433 1273 1447 1287
rect 2173 1273 2187 1287
rect 2213 1273 2227 1287
rect 2893 1273 2907 1287
rect 3013 1273 3027 1287
rect 3053 1273 3067 1287
rect 3273 1273 3287 1287
rect 3413 1273 3427 1287
rect 3833 1273 3847 1287
rect 4133 1273 4147 1287
rect 4293 1273 4307 1287
rect 4393 1273 4407 1287
rect 4573 1273 4587 1287
rect 4653 1273 4667 1287
rect 4693 1273 4707 1287
rect 4813 1273 4827 1287
rect 5013 1273 5027 1287
rect 313 1253 327 1267
rect 353 1253 367 1267
rect 1173 1253 1187 1267
rect 93 1233 107 1247
rect 133 1233 147 1247
rect 613 1233 627 1247
rect 673 1233 687 1247
rect 1693 1253 1707 1267
rect 1813 1253 1827 1267
rect 1893 1253 1907 1267
rect 2133 1253 2147 1267
rect 2353 1253 2367 1267
rect 2493 1253 2507 1267
rect 2733 1253 2747 1267
rect 2853 1253 2867 1267
rect 2913 1253 2927 1267
rect 3093 1253 3107 1267
rect 4253 1253 4267 1267
rect 4453 1253 4467 1267
rect 4093 1233 4107 1247
rect 4133 1233 4147 1247
rect 4533 1233 4547 1247
rect 4573 1233 4587 1247
rect 4693 1233 4707 1247
rect 4733 1233 4747 1247
rect 4853 1253 4867 1267
rect 5073 1253 5087 1267
rect 5133 1253 5147 1267
rect 5173 1253 5187 1267
rect 5473 1273 5487 1287
rect 5853 1273 5867 1287
rect 5893 1273 5907 1287
rect 5433 1253 5447 1267
rect 5293 1233 5307 1247
rect 5553 1253 5567 1267
rect 5933 1253 5947 1267
rect 6013 1253 6027 1267
rect 5813 1233 5827 1247
rect 5853 1233 5867 1247
rect 213 1213 227 1227
rect 333 1213 347 1227
rect 373 1213 387 1227
rect 773 1213 787 1227
rect 933 1213 947 1227
rect 973 1213 987 1227
rect 1253 1213 1267 1227
rect 1593 1213 1607 1227
rect 1873 1213 1887 1227
rect 1913 1213 1927 1227
rect 2193 1213 2207 1227
rect 2293 1213 2307 1227
rect 2893 1213 2907 1227
rect 3053 1213 3067 1227
rect 3093 1213 3107 1227
rect 3513 1213 3527 1227
rect 3833 1213 3847 1227
rect 3913 1213 3927 1227
rect 3973 1213 3987 1227
rect 4253 1213 4267 1227
rect 4393 1213 4407 1227
rect 4493 1213 4507 1227
rect 4853 1213 4867 1227
rect 5013 1213 5027 1227
rect 5133 1213 5147 1227
rect 5173 1213 5187 1227
rect 5353 1213 5367 1227
rect 5553 1213 5567 1227
rect 5613 1213 5627 1227
rect 5673 1213 5687 1227
rect 5973 1213 5987 1227
rect 3393 1193 3407 1207
rect 93 1173 107 1187
rect 633 1173 647 1187
rect 1093 1173 1107 1187
rect 1153 1173 1167 1187
rect 1373 1173 1387 1187
rect 1633 1173 1647 1187
rect 1773 1173 1787 1187
rect 2033 1173 2047 1187
rect 2093 1173 2107 1187
rect 2653 1173 2667 1187
rect 3033 1173 3047 1187
rect 3173 1173 3187 1187
rect 3633 1173 3647 1187
rect 3693 1173 3707 1187
rect 4132 1173 4146 1187
rect 4293 1173 4307 1187
rect 4453 1173 4467 1187
rect 4673 1173 4687 1187
rect 4733 1173 4747 1187
rect 4813 1173 4827 1187
rect 5213 1173 5227 1187
rect 5793 1173 5807 1187
rect 233 1153 247 1167
rect 493 1153 507 1167
rect 533 1153 547 1167
rect 793 1153 807 1167
rect 893 1153 907 1167
rect 913 1153 927 1167
rect 1273 1153 1287 1167
rect 1313 1153 1327 1167
rect 1693 1153 1707 1167
rect 1733 1153 1747 1167
rect 2213 1153 2227 1167
rect 2253 1153 2267 1167
rect 2393 1153 2407 1167
rect 2753 1153 2767 1167
rect 2793 1153 2807 1167
rect 2873 1153 2887 1167
rect 3293 1153 3307 1167
rect 3373 1153 3387 1167
rect 3413 1153 3427 1167
rect 3453 1153 3467 1167
rect 3953 1153 3967 1167
rect 3993 1153 4007 1167
rect 4073 1153 4087 1167
rect 4373 1153 4387 1167
rect 4413 1153 4427 1167
rect 4873 1153 4887 1167
rect 4993 1153 5007 1167
rect 5113 1153 5127 1167
rect 5153 1153 5167 1167
rect 5313 1153 5327 1167
rect 5433 1153 5447 1167
rect 5473 1153 5487 1167
rect 5513 1153 5527 1167
rect 5573 1153 5587 1167
rect 5933 1153 5947 1167
rect 113 1133 127 1147
rect 153 1133 167 1147
rect 213 1133 227 1147
rect 2353 1133 2367 1147
rect 3813 1133 3827 1147
rect 4493 1133 4507 1147
rect 4813 1133 4827 1147
rect 333 1113 347 1127
rect 533 1113 547 1127
rect 1273 1113 1287 1127
rect 1733 1113 1747 1127
rect 1773 1113 1787 1127
rect 2113 1113 2127 1127
rect 453 1093 467 1107
rect 613 1093 627 1107
rect 1433 1093 1447 1107
rect 2653 1113 2667 1127
rect 3033 1113 3047 1127
rect 3253 1113 3267 1127
rect 3953 1113 3967 1127
rect 4013 1113 4027 1127
rect 4073 1113 4087 1127
rect 4373 1113 4387 1127
rect 5113 1113 5127 1127
rect 5553 1113 5567 1127
rect 3473 1093 3487 1107
rect 3933 1093 3947 1107
rect 3973 1093 3987 1107
rect 4333 1093 4347 1107
rect 4413 1093 4427 1107
rect 2073 1073 2087 1087
rect 3213 1073 3227 1087
rect 3373 1073 3387 1087
rect 3513 1073 3527 1087
rect 3873 1073 3887 1087
rect 4913 1073 4927 1087
rect 4993 1073 5007 1087
rect 5153 1073 5167 1087
rect 5393 1073 5407 1087
rect 5433 1073 5447 1087
rect 5533 1073 5547 1087
rect 613 1053 627 1067
rect 1153 1053 1167 1067
rect 1373 1053 1387 1067
rect 1513 1053 1527 1067
rect 1833 1053 1847 1067
rect 2132 1054 2146 1068
rect 2154 1053 2168 1067
rect 2193 1053 2207 1067
rect 2373 1053 2387 1067
rect 2713 1053 2727 1067
rect 2793 1053 2807 1067
rect 3473 1053 3487 1067
rect 3633 1053 3647 1067
rect 4573 1053 4587 1067
rect 5233 1053 5247 1067
rect 93 1033 107 1047
rect 113 1013 127 1027
rect 153 1013 167 1027
rect 253 1033 267 1047
rect 533 1033 547 1047
rect 773 1033 787 1047
rect 1073 1033 1087 1047
rect 1233 1033 1247 1047
rect 1273 1033 1287 1047
rect 1313 1033 1327 1047
rect 1593 1033 1607 1047
rect 1773 1033 1787 1047
rect 2013 1033 2027 1047
rect 2112 1033 2126 1047
rect 2134 1032 2148 1046
rect 2313 1033 2327 1047
rect 2393 1033 2407 1047
rect 2493 1033 2507 1047
rect 3153 1033 3167 1047
rect 3293 1033 3307 1047
rect 3353 1033 3367 1047
rect 4273 1033 4287 1047
rect 4513 1033 4527 1047
rect 213 1013 227 1027
rect 273 1013 287 1027
rect 493 1013 507 1027
rect 633 1013 647 1027
rect 1913 1013 1927 1027
rect 1953 1013 1967 1027
rect 2033 1013 2047 1027
rect 2253 1013 2267 1027
rect 2353 1013 2367 1027
rect 2933 1013 2947 1027
rect 3173 1013 3187 1027
rect 3253 1013 3267 1027
rect 3773 1013 3787 1027
rect 4053 1013 4067 1027
rect 4313 1013 4327 1027
rect 4833 1013 4847 1027
rect 4873 1013 4887 1027
rect 233 993 247 1007
rect 2293 993 2307 1007
rect 2333 993 2347 1007
rect 2673 993 2687 1007
rect 2733 993 2747 1007
rect 3433 993 3447 1007
rect 3473 993 3487 1007
rect 3513 993 3527 1007
rect 3633 993 3647 1007
rect 4013 993 4027 1007
rect 4693 993 4707 1007
rect 4753 993 4767 1007
rect 4993 993 5007 1007
rect 153 973 167 987
rect 273 973 287 987
rect 312 973 326 987
rect 373 973 387 987
rect 693 973 707 987
rect 1173 973 1187 987
rect 1253 973 1267 987
rect 2213 973 2227 987
rect 2433 973 2447 987
rect 2753 973 2767 987
rect 2973 973 2987 987
rect 3193 973 3207 987
rect 3393 973 3407 987
rect 3593 973 3607 987
rect 3893 973 3907 987
rect 4873 973 4887 987
rect 4953 973 4967 987
rect 5173 973 5187 987
rect 5293 973 5307 987
rect 633 953 647 967
rect 113 933 127 947
rect 153 933 167 947
rect 233 933 247 947
rect 273 933 287 947
rect 373 933 387 947
rect 413 933 427 947
rect 493 933 507 947
rect 533 933 547 947
rect 573 933 587 947
rect 2633 953 2647 967
rect 2772 953 2786 967
rect 2794 953 2808 967
rect 2833 953 2847 967
rect 5193 953 5207 967
rect 1153 933 1167 947
rect 1273 933 1287 947
rect 1313 933 1327 947
rect 1433 933 1447 947
rect 1473 933 1487 947
rect 2313 933 2327 947
rect 2533 933 2547 947
rect 2973 933 2987 947
rect 3013 933 3027 947
rect 3153 933 3167 947
rect 3193 933 3207 947
rect 3433 933 3447 947
rect 3473 933 3487 947
rect 3593 933 3607 947
rect 3633 933 3647 947
rect 3733 933 3747 947
rect 3773 933 3787 947
rect 3893 933 3907 947
rect 3933 933 3947 947
rect 3993 933 4007 947
rect 4153 933 4167 947
rect 4193 933 4207 947
rect 4313 933 4327 947
rect 4373 933 4387 947
rect 4693 933 4707 947
rect 4733 933 4747 947
rect 4793 933 4807 947
rect 4833 933 4847 947
rect 4873 933 4887 947
rect 4993 933 5007 947
rect 5073 933 5087 947
rect 5133 933 5147 947
rect 5173 933 5187 947
rect 5293 933 5307 947
rect 5333 933 5347 947
rect 5453 933 5467 947
rect 5573 933 5587 947
rect 5613 933 5627 947
rect 5653 933 5667 947
rect 5693 933 5707 947
rect 5893 933 5907 947
rect 5933 933 5947 947
rect 693 913 707 927
rect 933 913 947 927
rect 1533 913 1547 927
rect 1593 913 1607 927
rect 1773 913 1787 927
rect 1833 913 1847 927
rect 2013 913 2027 927
rect 2133 913 2147 927
rect 2693 913 2707 927
rect 2773 913 2787 927
rect 3393 913 3407 927
rect 4513 913 4527 927
rect 4573 913 4587 927
rect 6033 893 6047 907
rect 6073 893 6087 907
rect 133 873 147 887
rect 393 873 407 887
rect 553 873 567 887
rect 673 873 687 887
rect 733 873 747 887
rect 1133 873 1147 887
rect 1253 873 1267 887
rect 1293 873 1307 887
rect 1413 873 1427 887
rect 1713 873 1727 887
rect 1953 873 1967 887
rect 2193 873 2207 887
rect 2333 873 2347 887
rect 2373 873 2387 887
rect 2453 873 2467 887
rect 2613 873 2627 887
rect 2993 873 3007 887
rect 3134 873 3148 887
rect 3213 873 3227 887
rect 3492 873 3506 887
rect 3514 873 3528 887
rect 3793 873 3807 887
rect 4013 873 4027 887
rect 4053 873 4067 887
rect 4133 873 4147 887
rect 4213 873 4227 887
rect 4393 873 4407 887
rect 4753 873 4767 887
rect 4813 873 4827 887
rect 5113 873 5127 887
rect 5193 873 5207 887
rect 5393 873 5407 887
rect 5433 873 5447 887
rect 5533 873 5547 887
rect 5673 873 5687 887
rect 5753 873 5767 887
rect 5873 873 5887 887
rect 5933 873 5947 887
rect 6053 873 6067 887
rect 93 853 107 867
rect 313 853 327 867
rect 373 853 387 867
rect 833 853 847 867
rect 893 853 907 867
rect 1013 853 1027 867
rect 1073 853 1087 867
rect 1533 853 1547 867
rect 2713 853 2727 867
rect 2753 853 2767 867
rect 2833 853 2847 867
rect 2873 853 2887 867
rect 3293 853 3307 867
rect 3333 853 3347 867
rect 253 833 267 847
rect 393 833 407 847
rect 553 833 567 847
rect 593 833 607 847
rect 653 833 667 847
rect 1173 833 1187 847
rect 1253 833 1267 847
rect 2413 833 2427 847
rect 2473 834 2487 848
rect 2993 833 3007 847
rect 3393 833 3407 847
rect 3693 833 3707 847
rect 4133 833 4147 847
rect 4853 853 4867 867
rect 4273 833 4287 847
rect 5213 833 5227 847
rect 5433 833 5447 847
rect 5573 833 5587 847
rect 5753 833 5767 847
rect 5953 833 5967 847
rect 133 813 147 827
rect 173 813 187 827
rect 233 813 247 827
rect 453 813 467 827
rect 613 813 627 827
rect 1013 813 1027 827
rect 1193 813 1207 827
rect 2473 812 2487 826
rect 2653 813 2667 827
rect 2693 813 2707 827
rect 2833 813 2847 827
rect 2873 813 2887 827
rect 3013 813 3027 827
rect 3313 813 3327 827
rect 3353 813 3367 827
rect 3493 813 3507 827
rect 93 793 107 807
rect 313 793 327 807
rect 893 793 907 807
rect 933 793 947 807
rect 1073 793 1087 807
rect 1133 793 1147 807
rect 1413 793 1427 807
rect 1953 793 1967 807
rect 2013 793 2027 807
rect 2613 793 2627 807
rect 2973 793 2987 807
rect 3913 793 3927 807
rect 5333 813 5347 827
rect 5473 813 5487 827
rect 4593 793 4607 807
rect 4633 793 4647 807
rect 5653 793 5667 807
rect 5893 793 5907 807
rect 293 773 307 787
rect 493 773 507 787
rect 553 773 567 787
rect 693 773 707 787
rect 773 773 787 787
rect 973 773 987 787
rect 1153 773 1167 787
rect 1193 773 1207 787
rect 1293 773 1307 787
rect 1473 773 1487 787
rect 1533 773 1547 787
rect 1633 773 1647 787
rect 1833 773 1847 787
rect 1913 773 1927 787
rect 3253 773 3267 787
rect 193 753 207 767
rect 253 753 267 767
rect 413 753 427 767
rect 632 753 646 767
rect 1393 753 1407 767
rect 1453 753 1467 767
rect 1713 753 1727 767
rect 1973 753 1987 767
rect 2013 753 2027 767
rect 2253 753 2267 767
rect 2573 753 2587 767
rect 2653 753 2667 767
rect 2733 753 2747 767
rect 2793 753 2807 767
rect 3093 753 3107 767
rect 3193 753 3207 767
rect 3453 773 3467 787
rect 3773 773 3787 787
rect 4373 773 4387 787
rect 4813 773 4827 787
rect 5593 773 5607 787
rect 5693 773 5707 787
rect 3693 753 3707 767
rect 3753 753 3767 767
rect 4054 753 4068 767
rect 4113 753 4127 767
rect 4353 753 4367 767
rect 4473 753 4487 767
rect 4593 753 4607 767
rect 4693 753 4707 767
rect 5753 753 5767 767
rect 5793 753 5807 767
rect 413 713 427 727
rect 453 713 467 727
rect 653 733 667 747
rect 1513 733 1527 747
rect 1633 733 1647 747
rect 973 713 987 727
rect 1013 713 1027 727
rect 1253 713 1267 727
rect 1393 713 1407 727
rect 1533 713 1547 727
rect 1913 733 1927 747
rect 2053 733 2067 747
rect 2233 733 2247 747
rect 2333 733 2347 747
rect 2373 733 2387 747
rect 2633 733 2647 747
rect 2673 733 2687 747
rect 3013 733 3027 747
rect 3233 733 3247 747
rect 3333 733 3347 747
rect 3673 733 3687 747
rect 4173 733 4187 747
rect 4293 733 4307 747
rect 4373 733 4387 747
rect 4853 733 4867 747
rect 4913 733 4927 747
rect 4993 733 5007 747
rect 1973 713 1987 727
rect 2013 713 2027 727
rect 2733 713 2747 727
rect 2773 713 2787 727
rect 3293 713 3307 727
rect 4073 713 4087 727
rect 4113 713 4127 727
rect 4553 713 4567 727
rect 4593 713 4607 727
rect 5693 713 5707 727
rect 5733 713 5747 727
rect 5973 713 5987 727
rect 6013 713 6027 727
rect 113 693 127 707
rect 253 693 267 707
rect 373 693 387 707
rect 613 693 627 707
rect 733 693 747 707
rect 893 693 907 707
rect 1073 693 1087 707
rect 1633 693 1647 707
rect 1713 693 1727 707
rect 2173 693 2187 707
rect 2333 693 2347 707
rect 2473 693 2487 707
rect 2573 693 2587 707
rect 2633 693 2647 707
rect 2693 693 2707 707
rect 2853 693 2867 707
rect 3013 693 3027 707
rect 3133 693 3147 707
rect 3192 693 3206 707
rect 3214 693 3228 707
rect 3573 693 3587 707
rect 3633 693 3647 707
rect 3673 693 3687 707
rect 3773 693 3787 707
rect 3873 693 3887 707
rect 3913 693 3927 707
rect 3973 693 3987 707
rect 4233 693 4247 707
rect 4333 693 4347 707
rect 4373 693 4387 707
rect 4473 693 4487 707
rect 4693 693 4707 707
rect 4773 693 4787 707
rect 4913 693 4927 707
rect 4993 693 5007 707
rect 5093 693 5107 707
rect 5313 693 5327 707
rect 5473 693 5487 707
rect 5573 693 5587 707
rect 5773 693 5787 707
rect 5893 693 5907 707
rect 73 653 87 667
rect 193 653 207 667
rect 493 653 507 667
rect 933 653 947 667
rect 1193 653 1207 667
rect 1253 653 1267 667
rect 1953 653 1967 667
rect 2033 653 2047 667
rect 2073 653 2087 667
rect 2153 653 2167 667
rect 2193 653 2207 667
rect 2293 653 2307 667
rect 2833 653 2847 667
rect 2973 653 2987 667
rect 3113 653 3127 667
rect 3393 653 3407 667
rect 3453 653 3467 667
rect 3793 653 3807 667
rect 3853 653 3867 667
rect 4173 653 4187 667
rect 4293 653 4307 667
rect 4353 653 4367 667
rect 4633 653 4647 667
rect 4813 653 4827 667
rect 5013 653 5027 667
rect 5213 653 5227 667
rect 5273 653 5287 667
rect 5953 653 5967 667
rect 233 633 247 647
rect 273 633 287 647
rect 553 633 567 647
rect 593 633 607 647
rect 793 633 807 647
rect 833 633 847 647
rect 873 633 887 647
rect 1513 633 1527 647
rect 1653 633 1667 647
rect 1693 633 1707 647
rect 1833 633 1847 647
rect 1993 633 2007 647
rect 2613 633 2627 647
rect 3153 633 3167 647
rect 3193 633 3207 647
rect 3313 633 3327 647
rect 3693 633 3707 647
rect 3733 633 3747 647
rect 4153 633 4167 647
rect 4393 633 4407 647
rect 4433 633 4447 647
rect 4673 633 4687 647
rect 4853 633 4867 647
rect 4893 633 4907 647
rect 5373 633 5387 647
rect 5413 633 5427 647
rect 5553 633 5567 647
rect 5593 633 5607 647
rect 5713 633 5727 647
rect 5833 633 5847 647
rect 5873 633 5887 647
rect 5933 633 5947 647
rect 73 613 87 627
rect 173 613 187 627
rect 593 593 607 607
rect 1793 613 1807 627
rect 1953 613 1967 627
rect 2233 613 2247 627
rect 3353 613 3367 627
rect 3453 613 3467 627
rect 3513 613 3527 627
rect 3633 613 3647 627
rect 3673 613 3687 627
rect 5913 613 5927 627
rect 5973 613 5987 627
rect 953 593 967 607
rect 1353 593 1367 607
rect 1653 593 1667 607
rect 1833 593 1847 607
rect 2073 593 2087 607
rect 2533 593 2547 607
rect 2574 593 2588 607
rect 2613 593 2627 607
rect 2853 593 2867 607
rect 3253 593 3267 607
rect 4393 593 4407 607
rect 4853 593 4867 607
rect 4893 593 4907 607
rect 4953 593 4967 607
rect 5013 593 5027 607
rect 373 573 387 587
rect 673 573 687 587
rect 873 573 887 587
rect 2893 573 2907 587
rect 2932 573 2946 587
rect 2954 573 2968 587
rect 3072 573 3086 587
rect 3153 573 3167 587
rect 4113 573 4127 587
rect 4233 573 4247 587
rect 4354 573 4368 587
rect 4553 573 4567 587
rect 4673 573 4687 587
rect 413 553 427 567
rect 573 553 587 567
rect 633 553 647 567
rect 733 553 747 567
rect 1013 553 1027 567
rect 2532 553 2546 567
rect 2573 553 2587 567
rect 3294 553 3308 567
rect 3333 553 3347 567
rect 3613 553 3627 567
rect 3713 553 3727 567
rect 4433 553 4447 567
rect 4533 553 4547 567
rect 4773 553 4787 567
rect 5013 553 5027 567
rect 5833 553 5847 567
rect 5893 553 5907 567
rect 113 533 127 547
rect 213 533 227 547
rect 1033 533 1047 547
rect 1253 533 1267 547
rect 1493 533 1507 547
rect 1573 533 1587 547
rect 1873 533 1887 547
rect 2033 533 2047 547
rect 2153 533 2167 547
rect 2293 533 2307 547
rect 2473 533 2487 547
rect 4753 533 4767 547
rect 4793 533 4807 547
rect 4833 533 4847 547
rect 5273 533 5287 547
rect 5633 533 5647 547
rect 413 513 427 527
rect 1993 513 2007 527
rect 273 493 287 507
rect 693 493 707 507
rect 853 493 867 507
rect 932 493 946 507
rect 954 493 968 507
rect 1073 493 1087 507
rect 1473 493 1487 507
rect 1553 493 1567 507
rect 1793 493 1807 507
rect 2053 493 2067 507
rect 2193 493 2207 507
rect 3193 513 3207 527
rect 3753 513 3767 527
rect 4013 513 4027 527
rect 4513 513 4527 527
rect 4573 513 4587 527
rect 93 473 107 487
rect 333 473 347 487
rect 1233 473 1247 487
rect 3673 473 3687 487
rect 3853 493 3867 507
rect 3953 493 3967 507
rect 4153 493 4167 507
rect 4253 493 4267 507
rect 5093 493 5107 507
rect 3893 473 3907 487
rect 4013 473 4027 487
rect 4433 473 4447 487
rect 5233 473 5247 487
rect 5313 473 5327 487
rect 5693 473 5707 487
rect 5773 473 5787 487
rect 213 453 227 467
rect 433 453 447 467
rect 493 453 507 467
rect 693 453 707 467
rect 993 453 1007 467
rect 1093 453 1107 467
rect 1153 453 1167 467
rect 1393 453 1407 467
rect 2573 453 2587 467
rect 2613 453 2627 467
rect 2773 453 2787 467
rect 3153 453 3167 467
rect 4033 453 4047 467
rect 4373 453 4387 467
rect 4753 453 4767 467
rect 5013 453 5027 467
rect 5293 453 5307 467
rect 5393 453 5407 467
rect 5473 453 5487 467
rect 5533 453 5547 467
rect 5613 453 5627 467
rect 5753 453 5767 467
rect 5893 453 5907 467
rect 5933 453 5947 467
rect 333 433 347 447
rect 373 433 387 447
rect 553 433 567 447
rect 2153 433 2167 447
rect 2293 433 2307 447
rect 4433 433 4447 447
rect 4473 433 4487 447
rect 5593 433 5607 447
rect 233 413 247 427
rect 273 413 287 427
rect 433 413 447 427
rect 953 413 967 427
rect 993 413 1007 427
rect 1073 413 1087 427
rect 1233 413 1247 427
rect 1273 413 1287 427
rect 1393 413 1407 427
rect 1433 413 1447 427
rect 1813 413 1827 427
rect 2193 413 2207 427
rect 2613 413 2627 427
rect 2653 413 2667 427
rect 2773 413 2787 427
rect 3233 413 3247 427
rect 3473 413 3487 427
rect 3713 413 3727 427
rect 4073 413 4087 427
rect 4113 413 4127 427
rect 4373 413 4387 427
rect 4413 413 4427 427
rect 4773 413 4787 427
rect 5173 413 5187 427
rect 5213 413 5227 427
rect 5333 413 5347 427
rect 5393 413 5407 427
rect 5713 413 5727 427
rect 5753 413 5767 427
rect 5893 413 5907 427
rect 5933 413 5947 427
rect 5973 413 5987 427
rect 193 393 207 407
rect 373 393 387 407
rect 633 393 647 407
rect 733 393 747 407
rect 1193 393 1207 407
rect 1493 393 1507 407
rect 1553 393 1567 407
rect 1873 393 1887 407
rect 1933 393 1947 407
rect 2153 393 2167 407
rect 2233 393 2247 407
rect 2373 393 2387 407
rect 2573 393 2587 407
rect 2813 393 2827 407
rect 2873 393 2887 407
rect 2893 393 2907 407
rect 2953 393 2967 407
rect 3093 393 3107 407
rect 3153 393 3167 407
rect 3193 393 3207 407
rect 3753 393 3767 407
rect 3773 393 3787 407
rect 3833 393 3847 407
rect 4153 393 4167 407
rect 4473 393 4487 407
rect 4533 393 4547 407
rect 4813 393 4827 407
rect 5133 393 5147 407
rect 5533 393 5547 407
rect 5593 393 5607 407
rect 213 353 227 367
rect 333 353 347 367
rect 413 353 427 367
rect 573 353 587 367
rect 693 353 707 367
rect 753 353 767 367
rect 853 353 867 367
rect 1093 353 1107 367
rect 1293 353 1307 367
rect 1373 353 1387 367
rect 1473 353 1487 367
rect 1673 353 1687 367
rect 1713 353 1727 367
rect 2053 353 2067 367
rect 2133 353 2147 367
rect 2333 353 2347 367
rect 2473 353 2487 367
rect 2633 353 2647 367
rect 2713 353 2727 367
rect 2753 353 2767 367
rect 2793 353 2807 367
rect 3093 353 3107 367
rect 3373 353 3387 367
rect 3493 353 3507 367
rect 3693 353 3707 367
rect 3953 353 3967 367
rect 4093 353 4107 367
rect 4133 353 4147 367
rect 4393 353 4407 367
rect 4433 353 4447 367
rect 4713 353 4727 367
rect 4753 353 4767 367
rect 5013 353 5027 367
rect 5153 353 5167 367
rect 5233 353 5247 367
rect 5293 353 5307 367
rect 5413 353 5427 367
rect 5693 353 5707 367
rect 5913 353 5927 367
rect 5993 353 6007 367
rect 93 333 107 347
rect 133 333 147 347
rect 1453 333 1467 347
rect 1493 333 1507 347
rect 1553 333 1567 347
rect 1613 333 1627 347
rect 2173 333 2187 347
rect 2213 333 2227 347
rect 2673 333 2687 347
rect 3173 333 3187 347
rect 3213 333 3227 347
rect 3613 333 3627 347
rect 4213 333 4227 347
rect 4253 333 4267 347
rect 4533 333 4547 347
rect 4593 333 4607 347
rect 4873 333 4887 347
rect 4913 333 4927 347
rect 1693 313 1707 327
rect 1853 313 1867 327
rect 2333 313 2347 327
rect 2473 313 2487 327
rect 2633 313 2647 327
rect 2693 313 2707 327
rect 2753 313 2767 327
rect 2793 313 2807 327
rect 2873 313 2887 327
rect 3253 313 3267 327
rect 613 293 627 307
rect 673 293 687 307
rect 493 273 507 287
rect 1033 293 1047 307
rect 1553 293 1567 307
rect 1613 293 1627 307
rect 1933 293 1947 307
rect 1993 293 2007 307
rect 2173 293 2187 307
rect 2233 293 2247 307
rect 2293 293 2307 307
rect 2853 293 2867 307
rect 3133 293 3147 307
rect 3473 293 3487 307
rect 3573 313 3587 327
rect 4673 313 4687 327
rect 4813 313 4827 327
rect 5133 313 5147 327
rect 5193 313 5207 327
rect 5233 313 5247 327
rect 5313 313 5327 327
rect 5873 333 5887 347
rect 5793 313 5807 327
rect 5993 313 6007 327
rect 3753 293 3767 307
rect 4913 293 4927 307
rect 5393 293 5407 307
rect 1013 273 1027 287
rect 1093 273 1107 287
rect 1213 273 1227 287
rect 2213 273 2227 287
rect 2533 273 2547 287
rect 2713 273 2727 287
rect 2753 273 2767 287
rect 3113 273 3127 287
rect 3333 273 3347 287
rect 3673 273 3687 287
rect 4072 273 4086 287
rect 4094 273 4108 287
rect 4633 273 4647 287
rect 5873 273 5887 287
rect 5953 273 5967 287
rect 293 253 307 267
rect 233 233 247 247
rect 673 233 687 247
rect 793 233 807 247
rect 1373 253 1387 267
rect 1453 253 1467 267
rect 1813 253 1827 267
rect 1893 253 1907 267
rect 2373 253 2387 267
rect 2513 253 2527 267
rect 2633 253 2647 267
rect 2673 253 2687 267
rect 3053 253 3067 267
rect 3093 253 3107 267
rect 3613 253 3627 267
rect 3693 253 3707 267
rect 3833 253 3847 267
rect 3933 253 3947 267
rect 4213 253 4227 267
rect 4873 253 4887 267
rect 4913 253 4927 267
rect 5073 253 5087 267
rect 5153 253 5167 267
rect 5313 253 5327 267
rect 5913 253 5927 267
rect 1533 233 1547 247
rect 1773 233 1787 247
rect 2213 233 2227 247
rect 2253 233 2267 247
rect 2453 233 2467 247
rect 2913 233 2927 247
rect 3733 233 3747 247
rect 4293 233 4307 247
rect 5134 233 5148 247
rect 5173 233 5187 247
rect 5553 233 5567 247
rect 5613 233 5627 247
rect 293 213 307 227
rect 233 193 247 207
rect 913 213 927 227
rect 2593 213 2607 227
rect 3573 213 3587 227
rect 3773 213 3787 227
rect 4053 213 4067 227
rect 4213 213 4227 227
rect 4253 213 4267 227
rect 2013 193 2027 207
rect 2053 193 2067 207
rect 2093 193 2107 207
rect 2213 193 2227 207
rect 2253 193 2267 207
rect 2673 193 2687 207
rect 2733 193 2747 207
rect 3053 193 3067 207
rect 3093 193 3107 207
rect 3213 193 3227 207
rect 3253 193 3267 207
rect 4293 193 4307 207
rect 4793 213 4807 227
rect 4873 213 4887 227
rect 5153 213 5167 227
rect 5233 213 5247 227
rect 5313 193 5327 207
rect 5373 193 5387 207
rect 5553 193 5567 207
rect 5613 193 5627 207
rect 5913 193 5927 207
rect 5953 193 5967 207
rect 193 173 207 187
rect 313 173 327 187
rect 673 173 687 187
rect 793 173 807 187
rect 913 173 927 187
rect 1013 173 1027 187
rect 1213 173 1227 187
rect 1253 173 1267 187
rect 1453 173 1467 187
rect 1513 173 1527 187
rect 1753 173 1767 187
rect 2473 173 2487 187
rect 2513 173 2527 187
rect 2573 173 2587 187
rect 2613 173 2627 187
rect 2913 173 2927 187
rect 3393 173 3407 187
rect 3433 173 3447 187
rect 3693 173 3707 187
rect 3733 173 3747 187
rect 3773 173 3787 187
rect 3813 173 3827 187
rect 3933 173 3947 187
rect 4013 173 4027 187
rect 4173 173 4187 187
rect 4213 173 4227 187
rect 4393 173 4407 187
rect 4633 173 4647 187
rect 4953 173 4967 187
rect 5073 173 5087 187
rect 5133 173 5147 187
rect 5253 173 5267 187
rect 5453 173 5467 187
rect 5493 173 5507 187
rect 5693 173 5707 187
rect 4993 153 5007 167
rect 433 133 447 147
rect 493 133 507 147
rect 753 133 767 147
rect 893 133 907 147
rect 1033 133 1047 147
rect 1093 133 1107 147
rect 1573 133 1587 147
rect 1633 133 1647 147
rect 1993 133 2007 147
rect 2073 133 2087 147
rect 2193 133 2207 147
rect 2273 133 2287 147
rect 2733 133 2747 147
rect 2793 133 2807 147
rect 3033 133 3047 147
rect 3113 133 3127 147
rect 3153 133 3167 147
rect 3213 133 3227 147
rect 4453 133 4467 147
rect 4593 133 4607 147
rect 4733 133 4747 147
rect 5373 133 5387 147
rect 5433 133 5447 147
rect 5613 133 5627 147
rect 5673 133 5687 147
rect 5893 133 5907 147
rect 5973 133 5987 147
rect 173 113 187 127
rect 213 113 227 127
rect 253 113 267 127
rect 613 113 627 127
rect 653 113 667 127
rect 713 113 727 127
rect 933 113 947 127
rect 973 113 987 127
rect 1233 113 1247 127
rect 1353 113 1367 127
rect 1473 113 1487 127
rect 1513 113 1527 127
rect 1773 113 1787 127
rect 1893 113 1907 127
rect 2033 113 2047 127
rect 2233 113 2247 127
rect 2373 113 2387 127
rect 2453 113 2467 127
rect 2513 113 2527 127
rect 2553 113 2567 127
rect 3073 113 3087 127
rect 3453 113 3467 127
rect 3573 113 3587 127
rect 3613 113 3627 127
rect 3713 113 3727 127
rect 3753 113 3767 127
rect 3873 113 3887 127
rect 3913 113 3927 127
rect 4033 113 4047 127
rect 4153 113 4167 127
rect 4193 113 4207 127
rect 1633 93 1647 107
rect 1693 93 1707 107
rect 893 73 907 87
rect 933 73 947 87
rect 1293 73 1307 87
rect 1473 73 1487 87
rect 1993 93 2007 107
rect 2273 93 2287 107
rect 3773 93 3787 107
rect 3833 93 3847 107
rect 4873 113 4887 127
rect 4913 113 4927 127
rect 5013 113 5027 127
rect 5053 113 5067 127
rect 5153 113 5167 127
rect 5193 113 5207 127
rect 5853 113 5867 127
rect 4773 93 4787 107
rect 5673 93 5687 107
rect 5753 93 5767 107
rect 5833 93 5847 107
rect 5973 93 5987 107
rect 6033 93 6047 107
rect 2413 73 2427 87
rect 2553 73 2567 87
rect 2813 73 2827 87
rect 3033 73 3047 87
rect 3353 73 3367 87
rect 4153 73 4167 87
rect 4193 73 4207 87
rect 4953 73 4967 87
rect 5053 73 5067 87
rect 5233 73 5247 87
rect 2073 53 2087 67
rect 2173 53 2187 67
rect 3413 53 3427 67
rect 3713 53 3727 67
rect 3913 53 3927 67
rect 5153 53 5167 67
rect 253 33 267 47
rect 333 33 347 47
rect 973 33 987 47
rect 1253 33 1267 47
rect 1513 33 1527 47
rect 2233 33 2247 47
rect 3293 33 3307 47
rect 3333 33 3347 47
rect 3373 33 3387 47
rect 3473 33 3487 47
rect 3573 33 3587 47
rect 5373 33 5387 47
rect 433 13 447 27
rect 2033 13 2047 27
rect 3413 13 3427 27
rect 3453 13 3467 27
rect 3493 13 3507 27
<< metal3 >>
rect 1316 6007 1324 6044
rect 136 5907 144 5973
rect 96 5767 104 5893
rect 176 5847 184 5893
rect 167 5836 184 5847
rect 216 5847 224 5973
rect 267 5896 334 5904
rect 436 5847 444 5953
rect 456 5907 464 5933
rect 616 5907 624 5933
rect 776 5916 824 5924
rect 776 5904 784 5916
rect 716 5900 784 5904
rect 713 5896 784 5900
rect 713 5887 727 5896
rect 556 5860 684 5864
rect 553 5856 687 5860
rect 553 5847 567 5856
rect 673 5847 687 5856
rect 216 5836 233 5847
rect 167 5833 180 5836
rect 220 5833 233 5836
rect 487 5836 513 5844
rect 116 5747 124 5833
rect 236 5667 244 5753
rect 276 5747 284 5833
rect 596 5807 604 5833
rect 636 5807 644 5833
rect 736 5807 744 5833
rect 776 5787 784 5833
rect 796 5767 804 5893
rect 816 5847 824 5916
rect 836 5907 844 5973
rect 896 5887 904 5973
rect 887 5876 904 5887
rect 887 5873 900 5876
rect 856 5856 944 5864
rect 856 5827 864 5856
rect 896 5807 904 5833
rect 936 5807 944 5856
rect 956 5767 964 5893
rect 976 5787 984 5833
rect 1036 5807 1044 5893
rect 116 5627 124 5653
rect 236 5627 244 5653
rect 296 5627 304 5753
rect 436 5627 444 5653
rect 167 5624 180 5627
rect 167 5613 184 5624
rect 287 5613 304 5627
rect 16 4187 24 4913
rect 36 4147 44 5473
rect 96 5447 104 5533
rect 96 4947 104 5373
rect 116 5364 124 5613
rect 136 5427 144 5553
rect 176 5527 184 5613
rect 256 5527 264 5553
rect 136 5387 144 5413
rect 116 5356 144 5364
rect 136 5327 144 5356
rect 136 5316 153 5327
rect 140 5313 153 5316
rect 116 5287 124 5313
rect 176 5284 184 5513
rect 296 5404 304 5613
rect 473 5604 487 5613
rect 473 5600 504 5604
rect 476 5596 504 5600
rect 467 5564 480 5567
rect 467 5560 484 5564
rect 467 5553 487 5560
rect 316 5487 324 5553
rect 473 5547 487 5553
rect 276 5396 304 5404
rect 167 5276 184 5284
rect 116 5047 124 5173
rect 156 5107 164 5273
rect 196 5107 204 5233
rect 236 5107 244 5373
rect 276 5344 284 5396
rect 316 5387 324 5433
rect 416 5427 424 5533
rect 496 5507 504 5596
rect 516 5547 524 5753
rect 556 5667 564 5753
rect 556 5627 564 5653
rect 607 5616 633 5624
rect 696 5567 704 5733
rect 756 5627 764 5653
rect 536 5556 573 5564
rect 536 5544 544 5556
rect 527 5536 544 5544
rect 276 5340 304 5344
rect 276 5336 307 5340
rect 293 5327 307 5336
rect 256 5187 264 5313
rect 376 5287 384 5373
rect 416 5327 424 5413
rect 476 5387 484 5413
rect 447 5384 460 5387
rect 447 5373 464 5384
rect 456 5364 464 5373
rect 456 5356 504 5364
rect 456 5287 464 5313
rect 496 5264 504 5356
rect 476 5256 504 5264
rect 196 4984 204 5093
rect 216 5007 224 5033
rect 176 4980 204 4984
rect 173 4976 204 4980
rect 173 4967 187 4976
rect 56 4427 64 4893
rect 116 4867 124 4953
rect 196 4867 204 4933
rect 256 4927 264 5033
rect 296 5007 304 5033
rect 376 4967 384 5093
rect 413 5084 427 5093
rect 396 5080 427 5084
rect 396 5076 424 5080
rect 396 5007 404 5076
rect 447 5044 460 5047
rect 447 5033 464 5044
rect 276 4807 284 4893
rect 267 4796 284 4807
rect 267 4793 280 4796
rect 216 4767 224 4793
rect 116 4527 124 4633
rect 16 4047 24 4113
rect 36 3887 44 4133
rect 16 3667 24 3773
rect 16 3547 24 3613
rect 36 3147 44 3833
rect 56 3347 64 4373
rect 76 4284 84 4393
rect 96 4367 104 4413
rect 136 4347 144 4373
rect 196 4327 204 4613
rect 236 4587 244 4733
rect 276 4624 284 4753
rect 316 4747 324 4893
rect 376 4867 384 4893
rect 416 4887 424 4913
rect 407 4796 433 4804
rect 356 4767 364 4793
rect 456 4764 464 5033
rect 476 4947 484 5256
rect 556 5187 564 5413
rect 616 5387 624 5513
rect 656 5447 664 5553
rect 776 5527 784 5553
rect 647 5316 673 5324
rect 596 5287 604 5313
rect 540 5104 553 5107
rect 536 5093 553 5104
rect 496 4887 504 5033
rect 536 4927 544 5093
rect 576 5047 584 5153
rect 616 5107 624 5233
rect 676 5147 684 5213
rect 716 5207 724 5373
rect 756 5327 764 5433
rect 776 5387 784 5513
rect 796 5448 804 5613
rect 916 5567 924 5693
rect 1016 5627 1024 5693
rect 996 5507 1004 5553
rect 796 5327 804 5412
rect 796 5287 804 5313
rect 856 5227 864 5473
rect 996 5387 1004 5493
rect 1056 5427 1064 5613
rect 1056 5387 1064 5413
rect 916 5227 924 5373
rect 1040 5324 1053 5327
rect 1036 5313 1053 5324
rect 1016 5287 1024 5313
rect 716 5107 724 5133
rect 607 5096 624 5107
rect 607 5093 620 5096
rect 676 5044 684 5093
rect 676 5036 733 5044
rect 556 4867 564 4953
rect 447 4756 464 4764
rect 267 4616 284 4624
rect 256 4587 264 4613
rect 256 4576 273 4587
rect 260 4573 273 4576
rect 376 4524 384 4713
rect 396 4587 404 4653
rect 436 4647 444 4753
rect 436 4587 444 4633
rect 376 4516 413 4524
rect 216 4407 224 4493
rect 256 4487 264 4513
rect 256 4347 264 4393
rect 296 4387 304 4513
rect 476 4487 484 4853
rect 576 4664 584 4973
rect 616 4967 624 5033
rect 756 5007 764 5093
rect 796 5087 804 5193
rect 836 5107 844 5133
rect 827 5036 853 5044
rect 876 5007 884 5093
rect 976 5087 984 5253
rect 1036 5107 1044 5313
rect 1096 5167 1104 5993
rect 1136 5847 1144 5973
rect 1156 5767 1164 5893
rect 1236 5847 1244 5933
rect 1296 5907 1304 5973
rect 1247 5836 1273 5844
rect 1316 5787 1324 5833
rect 1216 5627 1224 5653
rect 1116 5107 1124 5213
rect 1136 5207 1144 5233
rect 1156 5147 1164 5553
rect 1176 5507 1184 5613
rect 1236 5567 1244 5693
rect 1316 5687 1324 5773
rect 1256 5607 1264 5653
rect 1356 5647 1364 5893
rect 1456 5847 1464 5993
rect 1616 5907 1624 5933
rect 1676 5907 1684 5953
rect 1196 5327 1204 5413
rect 1216 5387 1224 5473
rect 1296 5467 1304 5633
rect 1316 5387 1324 5533
rect 1356 5507 1364 5533
rect 1376 5407 1384 5473
rect 1416 5447 1424 5773
rect 1456 5747 1464 5833
rect 1496 5727 1504 5833
rect 1536 5807 1544 5893
rect 1576 5767 1584 5893
rect 1676 5864 1684 5893
rect 1636 5860 1684 5864
rect 1633 5856 1684 5860
rect 1633 5847 1647 5856
rect 1747 5844 1760 5847
rect 1747 5833 1764 5844
rect 1596 5807 1604 5833
rect 1496 5547 1504 5673
rect 1456 5507 1464 5533
rect 1476 5424 1484 5473
rect 1516 5427 1524 5653
rect 1536 5507 1544 5553
rect 1596 5487 1604 5613
rect 1636 5507 1644 5613
rect 1456 5416 1484 5424
rect 1456 5387 1464 5416
rect 1676 5404 1684 5793
rect 1756 5767 1764 5833
rect 1776 5787 1784 5833
rect 1656 5400 1684 5404
rect 1653 5396 1684 5400
rect 1653 5387 1667 5396
rect 1456 5373 1473 5387
rect 1196 5227 1204 5313
rect 1196 5107 1204 5133
rect 656 4967 664 4993
rect 596 4724 604 4933
rect 656 4807 664 4913
rect 716 4867 724 4973
rect 707 4804 720 4807
rect 707 4800 724 4804
rect 707 4793 727 4800
rect 713 4787 727 4793
rect 596 4716 624 4724
rect 576 4660 604 4664
rect 576 4656 607 4660
rect 593 4647 607 4656
rect 576 4527 584 4613
rect 567 4516 584 4527
rect 567 4513 580 4516
rect 216 4296 284 4304
rect 76 4276 113 4284
rect 216 4284 224 4296
rect 276 4287 284 4296
rect 167 4276 224 4284
rect 287 4276 313 4284
rect 236 4247 244 4273
rect 76 3907 84 4173
rect 116 4067 124 4193
rect 136 4067 144 4173
rect 107 4056 124 4067
rect 107 4053 120 4056
rect 116 3967 124 3993
rect 96 3767 104 3853
rect 116 3727 124 3813
rect 136 3767 144 3873
rect 176 3607 184 4153
rect 216 4107 224 4193
rect 336 4167 344 4333
rect 256 4067 264 4133
rect 296 4067 304 4133
rect 336 4067 344 4113
rect 236 3827 244 3973
rect 276 3944 284 3993
rect 276 3940 304 3944
rect 276 3936 307 3940
rect 293 3927 307 3936
rect 276 3827 284 3893
rect 200 3764 213 3767
rect 196 3753 213 3764
rect 196 3567 204 3753
rect 256 3727 264 3753
rect 216 3647 224 3713
rect 107 3536 133 3544
rect 216 3487 224 3633
rect 316 3587 324 3953
rect 376 3947 384 4413
rect 436 4347 444 4393
rect 576 4367 584 4413
rect 533 4344 547 4353
rect 516 4340 547 4344
rect 516 4336 544 4340
rect 393 4044 407 4053
rect 393 4040 424 4044
rect 396 4036 424 4040
rect 236 3547 244 3573
rect 276 3547 284 3573
rect 336 3504 344 3933
rect 416 3927 424 4036
rect 356 3707 364 3913
rect 436 3867 444 4053
rect 476 4047 484 4293
rect 516 4287 524 4336
rect 496 4056 533 4064
rect 496 4007 504 4056
rect 396 3767 404 3853
rect 456 3784 464 3813
rect 416 3776 464 3784
rect 416 3767 424 3776
rect 407 3756 424 3767
rect 407 3753 420 3756
rect 436 3727 444 3753
rect 476 3687 484 3933
rect 556 3887 564 4253
rect 596 4067 604 4453
rect 616 4267 624 4716
rect 636 4587 644 4633
rect 676 4587 684 4693
rect 716 4587 724 4713
rect 756 4667 764 4893
rect 796 4867 804 4973
rect 836 4824 844 4933
rect 876 4904 884 4993
rect 896 4967 904 5013
rect 867 4896 884 4904
rect 816 4820 844 4824
rect 813 4816 844 4820
rect 813 4807 827 4816
rect 856 4807 864 4893
rect 636 4524 644 4573
rect 796 4527 804 4613
rect 816 4587 824 4733
rect 936 4707 944 5033
rect 856 4587 864 4653
rect 916 4564 924 4673
rect 956 4667 964 4853
rect 1016 4807 1024 5013
rect 1036 5007 1044 5093
rect 1073 5084 1087 5093
rect 1073 5080 1104 5084
rect 1076 5076 1107 5080
rect 1093 5067 1107 5076
rect 1216 5047 1224 5233
rect 1246 5144 1260 5147
rect 1246 5133 1264 5144
rect 1256 5047 1264 5133
rect 1056 4987 1064 5033
rect 976 4764 984 4793
rect 976 4756 1004 4764
rect 996 4627 1004 4756
rect 996 4587 1004 4613
rect 1016 4567 1024 4693
rect 1056 4687 1064 4893
rect 916 4556 953 4564
rect 636 4516 693 4524
rect 616 4127 624 4213
rect 587 4056 604 4067
rect 587 4053 600 4056
rect 636 4007 644 4373
rect 656 4347 664 4413
rect 716 4347 724 4473
rect 756 4287 764 4473
rect 916 4447 924 4556
rect 1016 4556 1033 4567
rect 1020 4553 1033 4556
rect 996 4516 1053 4524
rect 996 4507 1004 4516
rect 987 4496 1004 4507
rect 987 4493 1000 4496
rect 1016 4467 1024 4493
rect 876 4367 884 4393
rect 916 4387 924 4433
rect 1076 4427 1084 5013
rect 1096 4584 1104 4973
rect 1116 4947 1124 5033
rect 1176 4887 1184 4913
rect 1196 4907 1204 4973
rect 1276 4927 1284 5353
rect 1456 5344 1464 5373
rect 1436 5336 1464 5344
rect 1316 5287 1324 5313
rect 1356 5247 1364 5313
rect 1396 5267 1404 5293
rect 1436 5287 1444 5336
rect 1456 5284 1464 5313
rect 1516 5287 1524 5333
rect 1456 5276 1484 5284
rect 1336 5207 1344 5233
rect 1296 5147 1304 5193
rect 1396 5167 1404 5213
rect 1376 5107 1384 5133
rect 1367 5096 1384 5107
rect 1367 5093 1380 5096
rect 1316 4967 1324 5093
rect 1416 5047 1424 5193
rect 1316 4887 1324 4913
rect 1273 4864 1287 4873
rect 1147 4856 1204 4864
rect 1273 4860 1304 4864
rect 1276 4856 1304 4860
rect 1116 4727 1124 4793
rect 1156 4747 1164 4793
rect 1196 4764 1204 4856
rect 1176 4756 1204 4764
rect 1116 4687 1124 4713
rect 1176 4647 1184 4756
rect 1156 4587 1164 4613
rect 1196 4587 1204 4633
rect 1096 4576 1124 4584
rect 1096 4347 1104 4553
rect 1116 4467 1124 4576
rect 1136 4407 1144 4513
rect 1236 4487 1244 4733
rect 1256 4687 1264 4773
rect 1276 4527 1284 4633
rect 1296 4587 1304 4856
rect 1336 4627 1344 4913
rect 1376 4664 1384 4973
rect 1436 4927 1444 5273
rect 1456 5167 1464 5253
rect 1476 5107 1484 5276
rect 1576 5227 1584 5253
rect 1656 5247 1664 5273
rect 1516 5107 1524 5213
rect 1476 5007 1484 5093
rect 1556 5064 1564 5193
rect 1536 5060 1564 5064
rect 1533 5056 1564 5060
rect 1533 5047 1547 5056
rect 1396 4747 1404 4893
rect 1427 4856 1453 4864
rect 1356 4656 1384 4664
rect 1356 4587 1364 4656
rect 1307 4584 1320 4587
rect 1307 4573 1324 4584
rect 1347 4576 1364 4587
rect 1347 4573 1360 4576
rect 1316 4564 1324 4573
rect 1316 4556 1344 4564
rect 807 4336 833 4344
rect 1096 4336 1113 4347
rect 1100 4333 1113 4336
rect 747 4273 764 4287
rect 696 4167 704 4273
rect 756 4247 764 4273
rect 816 4167 824 4273
rect 856 4247 864 4273
rect 496 3727 504 3873
rect 596 3867 604 3993
rect 676 3907 684 4133
rect 813 4064 827 4073
rect 796 4060 827 4064
rect 796 4056 824 4060
rect 796 4044 804 4056
rect 856 4047 864 4113
rect 896 4107 904 4213
rect 936 4127 944 4293
rect 996 4107 1004 4293
rect 1056 4280 1133 4285
rect 1053 4277 1133 4280
rect 1053 4267 1067 4277
rect 1016 4087 1024 4253
rect 1136 4204 1144 4252
rect 1036 4200 1144 4204
rect 1033 4196 1144 4200
rect 1033 4187 1047 4196
rect 767 4036 804 4044
rect 816 3907 824 4033
rect 936 3967 944 4053
rect 636 3844 644 3893
rect 616 3836 644 3844
rect 616 3804 624 3836
rect 596 3796 624 3804
rect 596 3767 604 3796
rect 587 3756 604 3767
rect 587 3753 600 3756
rect 536 3707 544 3753
rect 336 3496 364 3504
rect 116 3447 124 3473
rect 276 3367 284 3413
rect 336 3407 344 3473
rect 356 3347 364 3496
rect 416 3487 424 3593
rect 476 3547 484 3573
rect 516 3547 524 3633
rect 407 3476 424 3487
rect 407 3473 420 3476
rect 467 3476 493 3484
rect 536 3387 544 3473
rect 136 3307 144 3333
rect 256 3307 264 3333
rect 396 3307 404 3333
rect 76 2967 84 3293
rect 116 3187 124 3233
rect 156 3147 164 3233
rect 236 3147 244 3233
rect 276 3187 284 3233
rect 296 3207 304 3293
rect 116 3027 124 3053
rect 76 2956 93 2967
rect 80 2953 93 2956
rect 56 2747 64 2853
rect 47 2736 64 2747
rect 47 2733 60 2736
rect 93 2704 107 2713
rect 47 2700 107 2704
rect 47 2696 104 2700
rect 36 2267 44 2433
rect 76 1884 84 2253
rect 116 2207 124 2913
rect 136 2487 144 2953
rect 156 2907 164 3013
rect 176 2927 184 2953
rect 216 2787 224 3053
rect 296 3027 304 3193
rect 256 2927 264 3013
rect 276 2587 284 2853
rect 316 2724 324 2953
rect 356 2804 364 3153
rect 396 3027 404 3293
rect 416 3187 424 3213
rect 576 3104 584 3673
rect 656 3547 664 3813
rect 716 3707 724 3813
rect 756 3767 764 3893
rect 756 3727 764 3753
rect 796 3707 804 3813
rect 876 3707 884 3813
rect 896 3727 904 3753
rect 696 3567 704 3593
rect 696 3327 704 3353
rect 736 3347 744 3373
rect 636 3187 644 3293
rect 756 3267 764 3673
rect 816 3607 824 3673
rect 856 3527 864 3673
rect 936 3667 944 3893
rect 956 3767 964 3873
rect 976 3827 984 3953
rect 996 3887 1004 3993
rect 1036 3907 1044 4033
rect 976 3687 984 3753
rect 896 3527 904 3653
rect 1016 3647 1024 3733
rect 1056 3684 1064 3853
rect 1076 3707 1084 4173
rect 1156 4147 1164 4473
rect 1176 4227 1184 4433
rect 1096 3907 1104 4033
rect 1156 3827 1164 3853
rect 1136 3727 1144 3753
rect 1056 3676 1084 3684
rect 1076 3667 1084 3676
rect 940 3524 953 3527
rect 936 3513 953 3524
rect 936 3504 944 3513
rect 916 3496 944 3504
rect 676 3227 684 3253
rect 676 3147 684 3213
rect 716 3167 724 3233
rect 776 3207 784 3253
rect 556 3096 584 3104
rect 556 3027 564 3096
rect 796 3067 804 3473
rect 916 3467 924 3496
rect 1076 3487 1084 3653
rect 907 3456 924 3467
rect 907 3453 920 3456
rect 856 3387 864 3453
rect 887 3436 953 3444
rect 1027 3436 1093 3444
rect 1116 3427 1124 3633
rect 1136 3567 1144 3713
rect 1176 3487 1184 3873
rect 1196 3707 1204 4413
rect 1256 4407 1264 4453
rect 1216 4367 1224 4393
rect 1267 4364 1280 4367
rect 1267 4353 1284 4364
rect 1276 4327 1284 4353
rect 1236 4147 1244 4233
rect 1256 4167 1264 4293
rect 1236 4024 1244 4093
rect 1216 4020 1244 4024
rect 1213 4016 1244 4020
rect 1213 4007 1227 4016
rect 1256 3827 1264 4153
rect 1247 3816 1264 3827
rect 1247 3813 1260 3816
rect 1296 3727 1304 4473
rect 1336 4347 1344 4556
rect 1356 4487 1364 4513
rect 1376 4427 1384 4633
rect 1396 4387 1404 4433
rect 1396 4287 1404 4373
rect 1316 4227 1324 4253
rect 1356 4247 1364 4273
rect 1356 4147 1364 4233
rect 1376 4067 1384 4113
rect 1416 4107 1424 4693
rect 1436 4667 1444 4856
rect 1496 4627 1504 4953
rect 1576 4807 1584 5133
rect 1656 5107 1664 5233
rect 1636 4967 1644 5033
rect 1656 5007 1664 5093
rect 1676 4824 1684 4933
rect 1696 4867 1704 5173
rect 1716 5147 1724 5733
rect 1736 5607 1744 5713
rect 1736 5447 1744 5593
rect 1756 5547 1764 5693
rect 1796 5647 1804 5753
rect 1836 5707 1844 5853
rect 1796 5507 1804 5533
rect 1816 5487 1824 5593
rect 1736 5064 1744 5373
rect 1756 5327 1764 5453
rect 1876 5447 1884 5933
rect 1936 5907 1944 5953
rect 2016 5907 2024 5953
rect 2196 5907 2204 5933
rect 2236 5864 2244 5913
rect 2216 5860 2244 5864
rect 2213 5856 2244 5860
rect 2116 5787 2124 5853
rect 2213 5847 2227 5856
rect 2176 5787 2184 5833
rect 1996 5607 2004 5713
rect 1956 5507 1964 5553
rect 1996 5487 2004 5593
rect 2036 5487 2044 5653
rect 2076 5607 2084 5713
rect 2076 5596 2093 5607
rect 2080 5593 2093 5596
rect 2116 5547 2124 5773
rect 2136 5627 2144 5733
rect 2216 5644 2224 5833
rect 2256 5687 2264 5933
rect 2296 5927 2304 5973
rect 2296 5867 2304 5913
rect 2196 5636 2224 5644
rect 2196 5607 2204 5636
rect 2187 5596 2204 5607
rect 2187 5593 2200 5596
rect 2167 5544 2180 5547
rect 2167 5540 2184 5544
rect 2167 5533 2187 5540
rect 2156 5507 2164 5533
rect 2173 5527 2187 5533
rect 2216 5527 2224 5593
rect 2316 5567 2324 5793
rect 2336 5787 2344 5893
rect 2476 5876 2533 5884
rect 2433 5844 2447 5853
rect 2476 5847 2484 5876
rect 2433 5840 2473 5844
rect 2436 5836 2473 5840
rect 2436 5767 2444 5836
rect 2556 5844 2564 5933
rect 2616 5907 2624 5933
rect 2656 5907 2664 5973
rect 2756 5947 2764 5973
rect 2536 5836 2564 5844
rect 2576 5847 2584 5873
rect 2576 5836 2593 5847
rect 2516 5767 2524 5833
rect 2416 5564 2424 5653
rect 2436 5627 2444 5693
rect 2487 5624 2500 5627
rect 2487 5613 2504 5624
rect 2416 5556 2453 5564
rect 1780 5384 1793 5387
rect 1776 5373 1793 5384
rect 1776 5167 1784 5373
rect 1916 5327 1924 5433
rect 1976 5387 1984 5433
rect 1816 5287 1824 5313
rect 1796 5107 1804 5233
rect 1856 5147 1864 5233
rect 1876 5187 1884 5273
rect 1916 5247 1924 5313
rect 1956 5287 1964 5313
rect 1996 5264 2004 5473
rect 2076 5327 2084 5453
rect 2136 5387 2144 5433
rect 2107 5384 2120 5387
rect 2107 5373 2124 5384
rect 2116 5364 2124 5373
rect 2116 5356 2144 5364
rect 2116 5287 2124 5313
rect 1996 5256 2024 5264
rect 1876 5107 1884 5173
rect 1787 5096 1804 5107
rect 1787 5093 1800 5096
rect 1736 5056 1784 5064
rect 1776 5047 1784 5056
rect 1740 5044 1753 5047
rect 1736 5033 1753 5044
rect 1776 5036 1793 5047
rect 1780 5033 1793 5036
rect 1716 4927 1724 4993
rect 1736 4907 1744 5033
rect 1756 4867 1764 4893
rect 1676 4816 1724 4824
rect 1716 4807 1724 4816
rect 1716 4796 1733 4807
rect 1720 4793 1733 4796
rect 1536 4767 1544 4793
rect 1436 4487 1444 4513
rect 1456 4467 1464 4573
rect 1496 4447 1504 4573
rect 1336 3967 1344 4053
rect 1356 3907 1364 3973
rect 1396 3947 1404 3993
rect 1456 3964 1464 4413
rect 1536 4407 1544 4753
rect 1656 4704 1664 4773
rect 1696 4707 1704 4793
rect 1756 4764 1764 4853
rect 1736 4760 1764 4764
rect 1733 4756 1764 4760
rect 1733 4747 1747 4756
rect 1776 4727 1784 4973
rect 1816 4927 1824 5093
rect 1916 5047 1924 5153
rect 1876 4907 1884 4933
rect 1820 4804 1833 4807
rect 1816 4793 1833 4804
rect 1816 4767 1824 4793
rect 1656 4696 1684 4704
rect 1576 4527 1584 4693
rect 1596 4647 1604 4673
rect 1636 4587 1644 4673
rect 1676 4647 1684 4696
rect 1647 4584 1660 4587
rect 1647 4573 1664 4584
rect 1576 4427 1584 4473
rect 1616 4427 1624 4513
rect 1656 4447 1664 4573
rect 1676 4547 1684 4633
rect 1747 4544 1760 4547
rect 1747 4533 1764 4544
rect 1716 4407 1724 4453
rect 1436 3956 1464 3964
rect 1436 3827 1444 3956
rect 1476 3947 1484 4053
rect 1476 3887 1484 3933
rect 1496 3867 1504 4393
rect 1533 4324 1547 4333
rect 1533 4320 1564 4324
rect 1536 4316 1567 4320
rect 1553 4307 1567 4316
rect 1516 4247 1524 4273
rect 1516 4167 1524 4233
rect 1576 4147 1584 4333
rect 1536 3907 1544 4113
rect 1596 3844 1604 4373
rect 1636 4287 1644 4373
rect 1656 4287 1664 4393
rect 1707 4344 1720 4347
rect 1707 4333 1724 4344
rect 1656 4276 1673 4287
rect 1660 4273 1673 4276
rect 1716 4247 1724 4333
rect 1756 4307 1764 4533
rect 1776 4527 1784 4633
rect 1776 4268 1784 4293
rect 1616 4107 1624 4193
rect 1616 4067 1624 4093
rect 1656 3967 1664 4053
rect 1656 3887 1664 3953
rect 1696 3847 1704 4153
rect 1776 4147 1784 4232
rect 1796 4187 1804 4653
rect 1816 4487 1824 4573
rect 1836 4407 1844 4753
rect 1876 4707 1884 4793
rect 1936 4747 1944 4933
rect 1956 4707 1964 5133
rect 1996 5047 2004 5233
rect 2016 4987 2024 5256
rect 2056 5107 2064 5213
rect 2136 5187 2144 5356
rect 2176 5287 2184 5373
rect 2076 5047 2084 5153
rect 2096 5107 2104 5173
rect 2196 5107 2204 5493
rect 2276 5387 2284 5453
rect 2356 5448 2364 5553
rect 2496 5527 2504 5613
rect 2476 5427 2484 5453
rect 2256 5287 2264 5313
rect 2276 5107 2284 5233
rect 2296 5227 2304 5313
rect 2356 5167 2364 5412
rect 2396 5387 2404 5413
rect 2453 5387 2467 5393
rect 2447 5380 2467 5387
rect 2447 5376 2464 5380
rect 2447 5373 2460 5376
rect 2476 5327 2484 5413
rect 2496 5327 2504 5393
rect 2400 5324 2413 5327
rect 2396 5313 2413 5324
rect 2467 5316 2484 5327
rect 2467 5313 2480 5316
rect 2396 5267 2404 5313
rect 2396 5227 2404 5253
rect 2496 5247 2504 5313
rect 2536 5267 2544 5836
rect 2580 5833 2593 5836
rect 2556 5667 2564 5813
rect 2636 5747 2644 5833
rect 2556 5624 2564 5653
rect 2556 5616 2593 5624
rect 2633 5604 2647 5613
rect 2633 5600 2664 5604
rect 2636 5596 2664 5600
rect 2576 5507 2584 5553
rect 2616 5527 2624 5553
rect 2656 5507 2664 5596
rect 2636 5496 2653 5504
rect 2573 5364 2587 5373
rect 2636 5364 2644 5496
rect 2573 5360 2644 5364
rect 2576 5356 2644 5360
rect 2676 5327 2684 5853
rect 2796 5827 2804 5913
rect 2716 5687 2724 5813
rect 2716 5627 2724 5673
rect 2756 5627 2764 5733
rect 2796 5567 2804 5773
rect 2816 5727 2824 5773
rect 2836 5747 2844 5933
rect 2896 5907 2904 5973
rect 2936 5864 2944 5973
rect 2916 5860 2944 5864
rect 2913 5856 2944 5860
rect 2913 5847 2927 5856
rect 2876 5727 2884 5833
rect 2856 5716 2873 5724
rect 2756 5427 2764 5493
rect 2567 5316 2593 5324
rect 2676 5316 2693 5327
rect 2680 5313 2693 5316
rect 2736 5284 2744 5313
rect 2776 5307 2784 5533
rect 2776 5296 2793 5307
rect 2780 5293 2793 5296
rect 2836 5287 2844 5693
rect 2856 5547 2864 5716
rect 2876 5627 2884 5673
rect 2916 5567 2924 5753
rect 2956 5747 2964 5813
rect 3016 5807 3024 5893
rect 3076 5867 3084 5973
rect 3176 5867 3184 5933
rect 3216 5924 3224 5973
rect 3196 5920 3224 5924
rect 3193 5916 3224 5920
rect 3193 5907 3207 5916
rect 3036 5787 3044 5813
rect 2996 5747 3004 5773
rect 2916 5556 2933 5567
rect 2920 5553 2933 5556
rect 2896 5467 2904 5553
rect 2976 5487 2984 5673
rect 2996 5467 3004 5633
rect 3036 5607 3044 5773
rect 3027 5596 3044 5607
rect 3027 5593 3040 5596
rect 3076 5547 3084 5853
rect 3236 5827 3244 5853
rect 3096 5727 3104 5813
rect 3096 5607 3104 5713
rect 3136 5627 3144 5693
rect 3156 5560 3193 5564
rect 3153 5556 3193 5560
rect 3153 5547 3167 5556
rect 3036 5507 3044 5533
rect 2716 5280 2744 5284
rect 2713 5276 2744 5280
rect 2713 5267 2727 5276
rect 2856 5267 2864 5373
rect 2876 5287 2884 5313
rect 2916 5287 2924 5453
rect 3033 5444 3047 5453
rect 3016 5440 3047 5444
rect 3016 5436 3044 5440
rect 3016 5407 3024 5436
rect 2967 5316 2993 5324
rect 2726 5260 2727 5267
rect 2436 5167 2444 5213
rect 2556 5207 2564 5233
rect 2416 5107 2424 5133
rect 2456 5107 2464 5153
rect 2576 5107 2584 5153
rect 2636 5107 2644 5133
rect 2220 5104 2233 5107
rect 2216 5093 2233 5104
rect 2627 5093 2644 5107
rect 1996 4807 2004 4893
rect 2056 4867 2064 4953
rect 2116 4907 2124 5033
rect 2067 4856 2104 4864
rect 2036 4747 2044 4793
rect 1856 4587 1864 4633
rect 1907 4584 1920 4587
rect 1907 4573 1924 4584
rect 1827 4336 1853 4344
rect 1876 4324 1884 4513
rect 1916 4504 1924 4573
rect 1896 4496 1924 4504
rect 1896 4427 1904 4496
rect 1916 4407 1924 4433
rect 1976 4367 1984 4653
rect 2016 4587 2024 4713
rect 2036 4707 2044 4733
rect 2056 4587 2064 4653
rect 2076 4647 2084 4673
rect 2096 4607 2104 4856
rect 2136 4807 2144 4973
rect 2196 4847 2204 5033
rect 2216 4907 2224 5093
rect 2547 5076 2604 5084
rect 2496 5044 2504 5073
rect 2596 5047 2604 5076
rect 2636 5068 2644 5093
rect 2447 5036 2504 5044
rect 2607 5036 2633 5044
rect 2627 5024 2640 5027
rect 2627 5013 2644 5024
rect 2176 4767 2184 4793
rect 2020 4524 2033 4527
rect 2016 4513 2033 4524
rect 2087 4516 2124 4524
rect 2016 4487 2024 4513
rect 2016 4347 2024 4413
rect 1856 4316 1884 4324
rect 1856 4247 1864 4316
rect 1913 4284 1927 4293
rect 1913 4280 1953 4284
rect 1916 4276 1953 4280
rect 1980 4284 1993 4287
rect 1976 4273 1993 4284
rect 1916 4187 1924 4253
rect 1976 4227 1984 4273
rect 1716 4007 1724 4093
rect 1756 3927 1764 4053
rect 1796 3967 1804 4053
rect 1816 3907 1824 4113
rect 1876 4007 1884 4133
rect 1896 3947 1904 4033
rect 1936 4007 1944 4193
rect 1976 4047 1984 4213
rect 2036 4107 2044 4413
rect 1576 3840 1604 3844
rect 1573 3836 1604 3840
rect 1573 3827 1587 3836
rect 1427 3816 1444 3827
rect 1427 3813 1440 3816
rect 1367 3756 1393 3764
rect 1447 3756 1473 3764
rect 1247 3544 1260 3547
rect 1247 3533 1264 3544
rect 1256 3487 1264 3533
rect 836 3307 844 3353
rect 856 3247 864 3333
rect 1176 3267 1184 3413
rect 1216 3387 1224 3453
rect 1276 3267 1284 3693
rect 1336 3387 1344 3573
rect 1396 3547 1404 3573
rect 1436 3347 1444 3693
rect 1456 3427 1464 3593
rect 1496 3547 1504 3813
rect 1716 3767 1724 3873
rect 1876 3827 1884 3853
rect 1556 3584 1564 3753
rect 1596 3707 1604 3753
rect 1596 3667 1604 3693
rect 1676 3687 1684 3753
rect 1756 3587 1764 3813
rect 1907 3756 1933 3764
rect 1856 3727 1864 3753
rect 1547 3576 1564 3584
rect 1607 3584 1620 3587
rect 1607 3573 1624 3584
rect 1536 3547 1544 3573
rect 816 3207 824 3233
rect 956 3187 964 3233
rect 1076 3107 1084 3253
rect 1236 3127 1244 3193
rect 1276 3147 1284 3253
rect 396 3016 413 3027
rect 400 3013 413 3016
rect 680 3024 693 3027
rect 676 3013 693 3024
rect 936 3016 993 3024
rect 456 2907 464 3013
rect 336 2800 364 2804
rect 333 2796 364 2800
rect 333 2787 347 2796
rect 376 2787 384 2813
rect 416 2787 424 2853
rect 536 2747 544 2913
rect 596 2907 604 3013
rect 676 2967 684 3013
rect 716 2927 724 2953
rect 736 2907 744 3013
rect 756 2927 764 2953
rect 767 2916 784 2924
rect 316 2716 353 2724
rect 276 2487 284 2573
rect 336 2507 344 2673
rect 396 2647 404 2713
rect 456 2587 464 2733
rect 576 2507 584 2853
rect 596 2647 604 2893
rect 776 2827 784 2916
rect 647 2776 673 2784
rect 736 2727 744 2813
rect 813 2784 827 2793
rect 787 2780 827 2784
rect 787 2776 824 2780
rect 736 2716 753 2727
rect 740 2713 753 2716
rect 876 2547 884 2993
rect 936 2947 944 3016
rect 960 2964 973 2967
rect 956 2953 973 2964
rect 956 2867 964 2953
rect 916 2827 924 2853
rect 956 2787 964 2853
rect 716 2507 724 2533
rect 216 2367 224 2473
rect 276 2367 284 2473
rect 456 2367 464 2433
rect 96 1907 104 2193
rect 76 1876 104 1884
rect 96 1787 104 1876
rect 96 1467 104 1493
rect 116 1484 124 1953
rect 156 1807 164 1893
rect 176 1744 184 2353
rect 576 2327 584 2493
rect 596 2367 604 2433
rect 596 2307 604 2353
rect 367 2264 380 2267
rect 367 2253 384 2264
rect 196 1927 204 2033
rect 216 1984 224 2173
rect 236 2067 244 2253
rect 376 2227 384 2253
rect 296 1987 304 2013
rect 216 1976 253 1984
rect 356 1984 364 2193
rect 516 2087 524 2213
rect 436 1987 444 2053
rect 356 1976 393 1984
rect 273 1907 287 1913
rect 273 1900 293 1907
rect 276 1896 293 1900
rect 280 1893 293 1896
rect 213 1744 227 1753
rect 176 1736 204 1744
rect 213 1740 253 1744
rect 216 1736 253 1740
rect 116 1480 144 1484
rect 116 1476 147 1480
rect 133 1467 147 1476
rect 136 1307 144 1453
rect 107 1296 124 1304
rect 96 1247 104 1293
rect 96 1047 104 1173
rect 116 1147 124 1296
rect 156 1287 164 1693
rect 196 1587 204 1736
rect 267 1736 293 1744
rect 236 1647 244 1673
rect 220 1464 233 1467
rect 216 1453 233 1464
rect 216 1407 224 1453
rect 256 1404 264 1493
rect 276 1467 284 1513
rect 256 1396 284 1404
rect 156 1247 164 1273
rect 147 1236 164 1247
rect 147 1233 160 1236
rect 196 1227 204 1273
rect 196 1216 213 1227
rect 200 1213 213 1216
rect 220 1164 233 1167
rect 216 1160 233 1164
rect 213 1153 233 1160
rect 213 1147 227 1153
rect 156 1027 164 1133
rect 256 1047 264 1373
rect 276 1027 284 1396
rect 296 1367 304 1393
rect 316 1267 324 1913
rect 356 1907 364 1976
rect 576 1927 584 2213
rect 676 1987 684 2073
rect 696 2067 704 2413
rect 736 2407 744 2433
rect 756 2387 764 2493
rect 796 2407 804 2473
rect 876 2444 884 2533
rect 856 2440 884 2444
rect 853 2436 884 2440
rect 853 2427 867 2436
rect 896 2427 904 2713
rect 1016 2647 1024 3073
rect 1156 3027 1164 3073
rect 1087 3016 1113 3024
rect 1096 2927 1104 2953
rect 1136 2867 1144 2953
rect 1236 2907 1244 3113
rect 1296 3027 1304 3093
rect 1376 3087 1384 3333
rect 1400 3304 1413 3307
rect 1396 3293 1413 3304
rect 1396 3167 1404 3293
rect 1456 3267 1464 3413
rect 1516 3267 1524 3473
rect 1556 3107 1564 3473
rect 1596 3407 1604 3473
rect 1616 3087 1624 3573
rect 1696 3547 1704 3573
rect 1640 3544 1653 3547
rect 1636 3533 1653 3544
rect 1636 3487 1644 3533
rect 1727 3476 1753 3484
rect 1676 3387 1684 3453
rect 1796 3427 1804 3593
rect 1836 3547 1844 3573
rect 1856 3487 1864 3573
rect 1876 3547 1884 3653
rect 1976 3547 1984 3813
rect 2016 3767 2024 3993
rect 2036 3867 2044 3953
rect 2056 3867 2064 4473
rect 2116 4467 2124 4516
rect 2076 4127 2084 4433
rect 2136 4304 2144 4713
rect 2156 4347 2164 4593
rect 2196 4587 2204 4653
rect 2236 4604 2244 4933
rect 2296 4927 2304 5013
rect 2316 4927 2324 4973
rect 2296 4867 2304 4913
rect 2376 4844 2384 4993
rect 2396 4947 2404 5013
rect 2636 4967 2644 5013
rect 2356 4836 2384 4844
rect 2300 4804 2313 4807
rect 2296 4793 2313 4804
rect 2216 4596 2244 4604
rect 2176 4387 2184 4493
rect 2216 4464 2224 4596
rect 2236 4467 2244 4573
rect 2256 4547 2264 4713
rect 2276 4647 2284 4793
rect 2276 4587 2284 4633
rect 2296 4607 2304 4793
rect 2356 4787 2364 4836
rect 2376 4820 2413 4824
rect 2373 4816 2413 4820
rect 2373 4807 2387 4816
rect 2456 4787 2464 4853
rect 2496 4827 2504 4853
rect 2487 4816 2504 4827
rect 2487 4813 2500 4816
rect 2316 4667 2324 4753
rect 2336 4604 2344 4733
rect 2376 4627 2384 4713
rect 2416 4688 2424 4773
rect 2336 4596 2364 4604
rect 2196 4456 2224 4464
rect 2167 4344 2180 4347
rect 2167 4333 2184 4344
rect 2176 4307 2184 4333
rect 2116 4296 2144 4304
rect 2096 4247 2104 4273
rect 2116 4144 2124 4296
rect 2133 4267 2147 4273
rect 2133 4260 2153 4267
rect 2136 4256 2153 4260
rect 2140 4253 2153 4256
rect 2156 4187 2164 4213
rect 2116 4136 2144 4144
rect 2096 4067 2104 4113
rect 2136 4107 2144 4136
rect 2196 4107 2204 4456
rect 2216 4347 2224 4433
rect 2216 4336 2233 4347
rect 2220 4333 2233 4336
rect 2276 4287 2284 4473
rect 2296 4287 2304 4453
rect 2267 4276 2284 4287
rect 2267 4273 2280 4276
rect 2316 4187 2324 4533
rect 2336 4407 2344 4573
rect 2356 4487 2364 4596
rect 2396 4527 2404 4673
rect 2416 4587 2424 4652
rect 2476 4587 2484 4653
rect 2496 4647 2504 4773
rect 2516 4667 2524 4953
rect 2576 4887 2584 4933
rect 2656 4927 2664 5213
rect 2676 4987 2684 5153
rect 2536 4647 2544 4833
rect 2576 4807 2584 4873
rect 2607 4864 2620 4867
rect 2607 4853 2624 4864
rect 2647 4856 2684 4864
rect 2616 4844 2624 4853
rect 2616 4836 2664 4844
rect 2656 4807 2664 4836
rect 2616 4767 2624 4793
rect 2676 4784 2684 4856
rect 2656 4776 2684 4784
rect 2516 4487 2524 4573
rect 2596 4524 2604 4673
rect 2616 4607 2624 4713
rect 2656 4707 2664 4776
rect 2696 4707 2704 5233
rect 2716 4987 2724 5173
rect 2736 5147 2744 5253
rect 2776 5207 2784 5253
rect 2736 5107 2744 5133
rect 2796 5107 2804 5193
rect 2787 5096 2804 5107
rect 2787 5093 2800 5096
rect 2767 5044 2780 5047
rect 2836 5044 2844 5233
rect 2856 5107 2864 5253
rect 2936 5187 2944 5253
rect 2956 5187 2964 5213
rect 2896 5107 2904 5173
rect 2976 5127 2984 5273
rect 2996 5247 3004 5313
rect 3036 5287 3044 5313
rect 3056 5227 3064 5373
rect 2996 5047 3004 5193
rect 3013 5107 3027 5113
rect 3076 5107 3084 5133
rect 3013 5100 3033 5107
rect 3016 5096 3033 5100
rect 3020 5093 3033 5096
rect 3096 5047 3104 5433
rect 3116 5067 3124 5293
rect 3136 5267 3144 5493
rect 3216 5487 3224 5613
rect 3156 5447 3164 5473
rect 3176 5327 3184 5413
rect 3196 5387 3204 5453
rect 3216 5327 3224 5393
rect 3256 5287 3264 5893
rect 3276 5748 3284 5813
rect 3316 5784 3324 5973
rect 3496 5927 3504 5973
rect 3676 5947 3684 5993
rect 3540 5924 3553 5927
rect 3536 5920 3553 5924
rect 3533 5913 3553 5920
rect 3627 5920 3704 5924
rect 3627 5916 3707 5920
rect 3533 5907 3547 5913
rect 3693 5907 3707 5916
rect 3387 5896 3413 5904
rect 3467 5896 3533 5904
rect 3376 5856 3464 5864
rect 3376 5847 3384 5856
rect 3367 5836 3384 5847
rect 3367 5833 3380 5836
rect 3396 5787 3404 5833
rect 3296 5776 3324 5784
rect 3276 5624 3284 5712
rect 3296 5707 3304 5776
rect 3316 5727 3324 5753
rect 3336 5627 3344 5693
rect 3436 5687 3444 5813
rect 3276 5616 3313 5624
rect 3136 5104 3144 5253
rect 3276 5247 3284 5616
rect 3336 5616 3353 5627
rect 3340 5613 3353 5616
rect 3336 5527 3344 5553
rect 3376 5524 3384 5553
rect 3356 5516 3384 5524
rect 3296 5428 3304 5473
rect 3336 5407 3344 5453
rect 3296 5347 3304 5392
rect 3356 5344 3364 5516
rect 3376 5407 3384 5493
rect 3396 5347 3404 5673
rect 3456 5447 3464 5856
rect 3576 5847 3584 5893
rect 3716 5847 3724 5973
rect 3567 5836 3584 5847
rect 3567 5833 3580 5836
rect 3516 5787 3524 5833
rect 3496 5527 3504 5613
rect 3496 5467 3504 5513
rect 3536 5487 3544 5613
rect 3556 5527 3564 5833
rect 3556 5513 3574 5527
rect 3516 5476 3533 5484
rect 3413 5424 3427 5433
rect 3413 5420 3444 5424
rect 3416 5416 3444 5420
rect 3336 5336 3364 5344
rect 3316 5308 3324 5333
rect 3196 5124 3204 5233
rect 3236 5147 3244 5233
rect 3316 5147 3324 5272
rect 3336 5227 3344 5336
rect 3356 5227 3364 5313
rect 3376 5147 3384 5233
rect 3196 5120 3224 5124
rect 3196 5116 3227 5120
rect 3213 5107 3227 5116
rect 3356 5107 3364 5133
rect 3436 5127 3444 5416
rect 3516 5344 3524 5476
rect 3556 5447 3564 5513
rect 3596 5467 3604 5753
rect 3636 5667 3644 5733
rect 3676 5708 3684 5813
rect 3756 5707 3764 5973
rect 3836 5907 3844 5973
rect 4056 5907 4064 6044
rect 4096 5967 4104 6044
rect 3887 5896 3904 5904
rect 3876 5844 3884 5893
rect 3827 5836 3884 5844
rect 3676 5627 3684 5672
rect 3556 5387 3564 5433
rect 3496 5340 3524 5344
rect 3493 5336 3524 5340
rect 3493 5327 3507 5336
rect 3547 5324 3560 5327
rect 3547 5320 3564 5324
rect 3547 5313 3567 5320
rect 3553 5307 3567 5313
rect 3576 5247 3584 5333
rect 3616 5267 3624 5553
rect 3656 5527 3664 5553
rect 3696 5487 3704 5553
rect 3676 5407 3684 5433
rect 3716 5407 3724 5693
rect 3736 5504 3744 5673
rect 3776 5627 3784 5653
rect 3796 5567 3804 5713
rect 3736 5500 3764 5504
rect 3736 5496 3767 5500
rect 3753 5487 3767 5496
rect 3736 5347 3744 5453
rect 3816 5447 3824 5673
rect 3876 5667 3884 5713
rect 3856 5507 3864 5653
rect 3876 5627 3884 5653
rect 3896 5644 3904 5896
rect 3956 5767 3964 5833
rect 3956 5687 3964 5753
rect 3996 5727 4004 5833
rect 4076 5808 4084 5893
rect 3896 5640 3944 5644
rect 3896 5636 3947 5640
rect 3933 5627 3947 5636
rect 3876 5616 3893 5627
rect 3880 5613 3893 5616
rect 3876 5527 3884 5553
rect 3856 5468 3864 5493
rect 3653 5324 3667 5333
rect 3653 5320 3684 5324
rect 3656 5316 3684 5320
rect 3676 5287 3684 5316
rect 3776 5267 3784 5413
rect 3856 5387 3864 5432
rect 3916 5427 3924 5533
rect 4016 5427 4024 5613
rect 4076 5567 4084 5772
rect 4096 5767 4104 5853
rect 4136 5807 4144 5993
rect 4296 5927 4304 5973
rect 4196 5916 4253 5924
rect 4196 5867 4204 5916
rect 4396 5867 4404 5973
rect 4587 5904 4600 5907
rect 4587 5893 4604 5904
rect 4300 5864 4313 5867
rect 4296 5853 4313 5864
rect 4236 5827 4244 5853
rect 4136 5624 4144 5673
rect 4107 5620 4144 5624
rect 4107 5616 4147 5620
rect 4133 5607 4147 5616
rect 3956 5324 3964 5333
rect 4056 5327 4064 5453
rect 3956 5316 3993 5324
rect 3816 5268 3824 5313
rect 3536 5107 3544 5233
rect 3136 5096 3173 5104
rect 2767 5040 2784 5044
rect 2767 5033 2787 5040
rect 2836 5036 2873 5044
rect 2773 5027 2787 5033
rect 2676 4587 2684 4673
rect 2716 4627 2724 4913
rect 2756 4887 2764 4973
rect 2796 4824 2804 4973
rect 2856 4927 2864 5036
rect 2996 5036 3013 5047
rect 3000 5033 3013 5036
rect 2896 4947 2904 4973
rect 2876 4867 2884 4933
rect 2756 4816 2804 4824
rect 2756 4724 2764 4816
rect 2776 4767 2784 4793
rect 2816 4767 2824 4793
rect 2916 4767 2924 4953
rect 2936 4727 2944 5033
rect 2956 4907 2964 4953
rect 3016 4807 3024 4973
rect 3036 4867 3044 4893
rect 2756 4716 2784 4724
rect 2736 4647 2744 4693
rect 2596 4516 2644 4524
rect 2536 4464 2544 4493
rect 2496 4456 2544 4464
rect 2576 4464 2584 4493
rect 2576 4460 2604 4464
rect 2576 4456 2607 4460
rect 2336 4227 2344 4393
rect 2356 4187 2364 4373
rect 2436 4347 2444 4433
rect 2476 4347 2484 4453
rect 2496 4407 2504 4456
rect 2593 4447 2607 4456
rect 2593 4440 2594 4447
rect 2376 4227 2384 4333
rect 2576 4307 2584 4433
rect 2236 4127 2244 4173
rect 2416 4167 2424 4273
rect 2456 4187 2464 4273
rect 2436 4127 2444 4153
rect 2236 4067 2244 4113
rect 2276 4067 2284 4093
rect 2147 4056 2184 4064
rect 2116 3927 2124 3993
rect 2176 3888 2184 4056
rect 2296 4007 2304 4113
rect 2396 4067 2404 4113
rect 2347 3996 2373 4004
rect 2036 3827 2044 3853
rect 2056 3727 2064 3753
rect 2116 3607 2124 3853
rect 2176 3827 2184 3852
rect 2116 3547 2124 3593
rect 1976 3536 1993 3547
rect 1980 3533 1993 3536
rect 2047 3544 2060 3547
rect 2047 3533 2064 3544
rect 1956 3476 2013 3484
rect 1956 3447 1964 3476
rect 2056 3427 2064 3533
rect 2136 3487 2144 3573
rect 2156 3547 2164 3653
rect 2196 3607 2204 3693
rect 2236 3687 2244 3813
rect 2256 3667 2264 3973
rect 2436 3947 2444 4053
rect 2276 3767 2284 3933
rect 2316 3827 2324 3873
rect 2336 3867 2344 3913
rect 2336 3767 2344 3853
rect 2276 3756 2293 3767
rect 2280 3753 2293 3756
rect 2376 3727 2384 3873
rect 2436 3767 2444 3933
rect 2456 3887 2464 4173
rect 2496 4167 2504 4213
rect 2476 3867 2484 3993
rect 2496 3927 2504 4093
rect 2516 3947 2524 4293
rect 2616 4207 2624 4493
rect 2576 4067 2584 4133
rect 2616 4067 2624 4093
rect 2596 3907 2604 3993
rect 2636 3867 2644 4516
rect 2696 4347 2704 4453
rect 2716 4407 2724 4433
rect 2736 4387 2744 4573
rect 2756 4247 2764 4693
rect 2776 4347 2784 4716
rect 2836 4567 2844 4713
rect 3036 4667 3044 4733
rect 3076 4707 3084 5033
rect 3116 4907 3124 5013
rect 3156 4927 3164 5033
rect 3196 5007 3204 5033
rect 3120 4864 3133 4867
rect 3116 4853 3133 4864
rect 3116 4767 3124 4853
rect 2827 4516 2853 4524
rect 2816 4347 2824 4373
rect 2836 4287 2844 4473
rect 2856 4387 2864 4492
rect 2876 4407 2884 4633
rect 2936 4607 2944 4653
rect 3076 4587 3084 4633
rect 3033 4564 3047 4573
rect 3016 4560 3047 4564
rect 3016 4556 3044 4560
rect 3016 4528 3024 4556
rect 2956 4467 2964 4493
rect 2676 4127 2684 4193
rect 2736 4107 2744 4213
rect 2776 4147 2784 4193
rect 2796 4167 2804 4273
rect 2716 3907 2724 4053
rect 2736 4007 2744 4093
rect 2776 4067 2784 4133
rect 2800 4044 2813 4047
rect 2796 4033 2813 4044
rect 2736 3996 2753 4007
rect 2740 3993 2753 3996
rect 2796 3947 2804 4033
rect 2476 3827 2484 3853
rect 2756 3767 2764 3873
rect 2436 3756 2453 3767
rect 2440 3753 2453 3756
rect 2496 3727 2504 3753
rect 2276 3487 2284 3713
rect 2296 3547 2304 3673
rect 2336 3587 2344 3673
rect 2336 3547 2344 3573
rect 2176 3427 2184 3453
rect 1707 3296 1733 3304
rect 1756 3207 1764 3233
rect 1876 3207 1884 3233
rect 1653 3124 1667 3133
rect 1653 3120 1684 3124
rect 1656 3116 1684 3120
rect 1436 3027 1444 3073
rect 1076 2747 1084 2853
rect 936 2407 944 2473
rect 976 2387 984 2493
rect 1076 2487 1084 2613
rect 1136 2587 1144 2733
rect 1196 2587 1204 2773
rect 1276 2547 1284 2933
rect 1316 2908 1324 2953
rect 1336 2927 1344 3013
rect 1473 3004 1487 3013
rect 1473 3000 1513 3004
rect 1476 2996 1513 3000
rect 1440 2964 1453 2967
rect 1436 2953 1453 2964
rect 1316 2747 1324 2872
rect 1436 2867 1444 2953
rect 1476 2927 1484 2996
rect 1507 2964 1520 2967
rect 1507 2953 1524 2964
rect 1516 2904 1524 2953
rect 1516 2896 1544 2904
rect 1496 2747 1504 2853
rect 1376 2707 1384 2733
rect 1436 2707 1444 2733
rect 1316 2507 1324 2613
rect 1436 2607 1444 2693
rect 1536 2527 1544 2896
rect 1556 2887 1564 2913
rect 1493 2507 1507 2513
rect 1120 2504 1133 2507
rect 1116 2493 1133 2504
rect 1247 2496 1273 2504
rect 1487 2500 1507 2507
rect 1487 2496 1504 2500
rect 1487 2493 1500 2496
rect 996 2407 1004 2433
rect 1116 2407 1124 2493
rect 1176 2367 1184 2493
rect 767 2296 784 2304
rect 756 2267 764 2293
rect 776 2267 784 2296
rect 916 2276 973 2284
rect 776 2256 793 2267
rect 780 2253 793 2256
rect 916 2227 924 2276
rect 1073 2264 1087 2273
rect 1073 2260 1113 2264
rect 1076 2256 1113 2260
rect 736 2167 744 2193
rect 736 2127 744 2153
rect 976 2107 984 2213
rect 1096 2087 1104 2193
rect 1136 2127 1144 2193
rect 1156 2067 1164 2253
rect 1207 2224 1220 2227
rect 1207 2213 1224 2224
rect 696 1987 704 2053
rect 856 1987 864 2033
rect 696 1976 713 1987
rect 700 1973 713 1976
rect 800 1984 813 1987
rect 796 1973 813 1984
rect 796 1927 804 1973
rect 467 1916 493 1924
rect 627 1916 653 1924
rect 376 1527 384 1833
rect 416 1756 473 1764
rect 416 1707 424 1756
rect 476 1587 484 1693
rect 536 1647 544 1813
rect 576 1747 584 1793
rect 616 1747 624 1773
rect 596 1647 604 1673
rect 636 1587 644 1673
rect 336 1367 344 1473
rect 376 1387 384 1513
rect 436 1487 444 1553
rect 436 1387 444 1473
rect 376 1376 393 1387
rect 380 1373 393 1376
rect 476 1364 484 1573
rect 516 1387 524 1413
rect 576 1387 584 1533
rect 516 1376 533 1387
rect 520 1373 533 1376
rect 456 1356 484 1364
rect 116 947 124 1013
rect 156 947 164 973
rect 96 807 104 853
rect 136 827 144 873
rect 76 627 84 653
rect 116 547 124 693
rect 176 627 184 813
rect 196 667 204 753
rect 216 547 224 1013
rect 236 947 244 993
rect 316 987 324 1253
rect 356 1227 364 1253
rect 356 1216 373 1227
rect 360 1213 373 1216
rect 336 1127 344 1213
rect 456 1107 464 1356
rect 616 1307 624 1393
rect 656 1327 664 1793
rect 756 1787 764 1873
rect 916 1827 924 1913
rect 956 1887 964 1913
rect 976 1847 984 1973
rect 1020 1924 1033 1927
rect 1016 1913 1033 1924
rect 1016 1887 1024 1913
rect 1156 1827 1164 1953
rect 873 1744 887 1753
rect 873 1740 913 1744
rect 876 1736 913 1740
rect 927 1736 953 1744
rect 676 1547 684 1693
rect 736 1467 744 1533
rect 816 1464 824 1593
rect 896 1567 904 1673
rect 796 1460 824 1464
rect 793 1456 824 1460
rect 793 1447 807 1456
rect 616 1247 624 1293
rect 676 1247 684 1273
rect 756 1227 764 1293
rect 756 1216 773 1227
rect 760 1213 773 1216
rect 496 1027 504 1153
rect 536 1127 544 1153
rect 616 1067 624 1093
rect 276 947 284 973
rect 236 827 244 933
rect 256 767 264 833
rect 256 707 264 753
rect 276 664 284 933
rect 316 867 324 973
rect 376 947 384 973
rect 536 947 544 1033
rect 636 1027 644 1173
rect 836 1164 844 1473
rect 893 1467 907 1473
rect 893 1460 913 1467
rect 896 1456 913 1460
rect 900 1453 913 1456
rect 936 1407 944 1533
rect 967 1464 980 1467
rect 967 1453 984 1464
rect 976 1407 984 1453
rect 896 1367 904 1393
rect 896 1327 904 1353
rect 916 1167 924 1293
rect 936 1227 944 1273
rect 947 1216 973 1224
rect 807 1156 844 1164
rect 400 944 413 947
rect 396 933 413 944
rect 587 944 600 947
rect 587 933 604 944
rect 396 924 404 933
rect 376 916 404 924
rect 376 867 384 916
rect 396 847 404 873
rect 327 804 340 807
rect 327 793 344 804
rect 256 656 284 664
rect 256 647 264 656
rect 296 647 304 773
rect 247 636 264 647
rect 247 633 260 636
rect 287 636 304 647
rect 287 633 300 636
rect 127 536 144 544
rect 96 347 104 473
rect 136 347 144 536
rect 216 427 224 453
rect 276 427 284 493
rect 336 487 344 793
rect 416 727 424 753
rect 456 727 464 813
rect 496 787 504 933
rect 556 847 564 873
rect 596 847 604 933
rect 556 787 564 833
rect 376 587 384 693
rect 416 567 424 713
rect 616 707 624 813
rect 636 767 644 953
rect 696 927 704 973
rect 687 876 733 884
rect 656 747 664 833
rect 776 787 784 1033
rect 836 867 844 1156
rect 896 867 904 1153
rect 936 807 944 913
rect 996 884 1004 1813
rect 1156 1724 1164 1773
rect 1136 1720 1164 1724
rect 1133 1716 1164 1720
rect 1133 1707 1147 1716
rect 1073 1664 1087 1673
rect 1073 1660 1133 1664
rect 1076 1656 1133 1660
rect 1196 1627 1204 2113
rect 1216 2107 1224 2213
rect 1236 2127 1244 2433
rect 1216 2007 1224 2093
rect 1296 2027 1304 2373
rect 1316 2227 1324 2333
rect 1336 2104 1344 2433
rect 1376 2367 1384 2433
rect 1436 2347 1444 2493
rect 1496 2407 1504 2433
rect 1396 2307 1404 2333
rect 1387 2256 1413 2264
rect 1316 2096 1344 2104
rect 1316 2047 1324 2096
rect 1216 1967 1224 1993
rect 1236 1847 1244 1913
rect 1256 1747 1264 1973
rect 1316 1824 1324 1993
rect 1336 1987 1344 2053
rect 1376 1987 1384 2013
rect 1356 1847 1364 1893
rect 1316 1816 1333 1824
rect 1336 1787 1344 1813
rect 1247 1736 1264 1747
rect 1247 1733 1260 1736
rect 1287 1744 1300 1747
rect 1287 1733 1304 1744
rect 1056 1367 1064 1453
rect 1056 1164 1064 1353
rect 1096 1327 1104 1453
rect 1156 1327 1164 1393
rect 1176 1224 1184 1253
rect 1136 1216 1184 1224
rect 1136 1184 1144 1216
rect 1107 1176 1144 1184
rect 1056 1156 1084 1164
rect 1076 1047 1084 1156
rect 1156 1067 1164 1173
rect 1176 947 1184 973
rect 1167 933 1184 947
rect 976 876 1004 884
rect 336 447 344 473
rect 216 416 233 427
rect 220 413 233 416
rect 196 367 204 393
rect 196 356 213 367
rect 200 353 213 356
rect 236 207 244 233
rect 180 184 193 187
rect 176 173 193 184
rect 176 127 184 173
rect 276 144 284 413
rect 376 407 384 433
rect 416 367 424 513
rect 496 467 504 653
rect 436 427 444 453
rect 556 447 564 633
rect 596 607 604 633
rect 576 367 584 553
rect 636 407 644 553
rect 296 227 304 253
rect 296 187 304 213
rect 296 176 313 187
rect 300 173 313 176
rect 236 136 284 144
rect 236 127 244 136
rect 227 116 244 127
rect 227 113 240 116
rect 256 47 264 113
rect 336 47 344 353
rect 676 324 684 573
rect 696 507 704 773
rect 896 707 904 793
rect 936 724 944 793
rect 976 787 984 876
rect 1016 827 1024 853
rect 1076 807 1084 853
rect 1136 807 1144 873
rect 1176 847 1184 933
rect 1196 827 1204 1613
rect 1256 1567 1264 1673
rect 1296 1647 1304 1733
rect 1316 1627 1324 1733
rect 1336 1607 1344 1773
rect 1276 1447 1284 1533
rect 1336 1447 1344 1593
rect 1256 1227 1264 1293
rect 1316 1167 1324 1273
rect 1276 1127 1284 1153
rect 1276 1047 1284 1113
rect 1236 887 1244 1033
rect 1256 947 1264 973
rect 1316 947 1324 1033
rect 1256 936 1273 947
rect 1260 933 1273 936
rect 1236 876 1253 887
rect 1240 873 1253 876
rect 936 716 973 724
rect 736 567 744 693
rect 807 636 833 644
rect 876 587 884 633
rect 936 507 944 653
rect 956 507 964 593
rect 1016 567 1024 713
rect 1076 707 1084 793
rect 696 367 704 453
rect 747 404 760 407
rect 747 393 764 404
rect 756 367 764 393
rect 856 367 864 493
rect 956 427 964 493
rect 996 427 1004 453
rect 656 316 684 324
rect 496 147 504 273
rect 436 27 444 133
rect 616 127 624 293
rect 656 127 664 316
rect 1036 307 1044 533
rect 1076 427 1084 493
rect 1156 467 1164 773
rect 1196 667 1204 773
rect 1256 727 1264 833
rect 1296 787 1304 873
rect 1256 547 1264 653
rect 1356 607 1364 1333
rect 1376 1327 1384 1453
rect 1396 1347 1404 1853
rect 1416 1544 1424 2093
rect 1456 1687 1464 2313
rect 1476 2267 1484 2353
rect 1496 2207 1504 2393
rect 1476 2067 1484 2153
rect 1536 2107 1544 2373
rect 1596 2327 1604 2893
rect 1636 2887 1644 2953
rect 1676 2867 1684 3116
rect 1816 3107 1824 3193
rect 1916 3167 1924 3193
rect 1876 3107 1884 3153
rect 1736 3027 1744 3073
rect 1816 3047 1824 3093
rect 1760 3024 1773 3027
rect 1756 3013 1773 3024
rect 1716 2907 1724 2953
rect 1756 2907 1764 3013
rect 1816 2967 1824 2993
rect 1807 2956 1824 2967
rect 1807 2953 1820 2956
rect 1876 2947 1884 3093
rect 1936 2947 1944 3133
rect 1876 2936 1893 2947
rect 1880 2933 1893 2936
rect 1976 2924 1984 3013
rect 1996 3004 2004 3393
rect 2116 3267 2124 3393
rect 2256 3307 2264 3433
rect 2376 3407 2384 3613
rect 2396 3516 2433 3524
rect 2396 3427 2404 3516
rect 2456 3467 2464 3673
rect 2596 3607 2604 3753
rect 2496 3387 2504 3453
rect 2516 3407 2524 3513
rect 2056 3184 2064 3233
rect 2056 3176 2124 3184
rect 2076 3027 2084 3153
rect 2027 3016 2053 3024
rect 2076 3013 2093 3027
rect 2076 3004 2084 3013
rect 1996 2996 2024 3004
rect 1956 2916 1984 2924
rect 1736 2787 1744 2833
rect 1627 2776 1653 2784
rect 1727 2776 1744 2787
rect 1727 2773 1740 2776
rect 1636 2367 1644 2653
rect 1736 2627 1744 2713
rect 1656 2527 1664 2613
rect 1836 2607 1844 2853
rect 1956 2807 1964 2916
rect 2016 2847 2024 2996
rect 2036 2996 2084 3004
rect 2036 2827 2044 2996
rect 2076 2827 2084 2933
rect 2116 2927 2124 3176
rect 2156 3147 2164 3253
rect 2256 3187 2264 3293
rect 2296 3267 2304 3373
rect 2296 3207 2304 3253
rect 2336 3107 2344 3333
rect 2396 3307 2404 3333
rect 2556 3327 2564 3553
rect 2596 3327 2604 3353
rect 2376 3187 2384 3233
rect 2416 3207 2424 3233
rect 2136 2967 2144 3073
rect 2396 3027 2404 3073
rect 2167 3016 2193 3024
rect 2247 3016 2304 3024
rect 2176 2904 2184 2953
rect 2216 2927 2224 2953
rect 2256 2907 2264 2953
rect 2156 2896 2184 2904
rect 2156 2827 2164 2896
rect 2236 2787 2244 2873
rect 2296 2787 2304 3016
rect 2367 3024 2380 3027
rect 2367 3013 2384 3024
rect 2376 2827 2384 3013
rect 2416 2967 2424 3113
rect 2436 3027 2444 3073
rect 2476 2967 2484 3133
rect 2516 3087 2524 3293
rect 2616 3087 2624 3253
rect 2636 3164 2644 3753
rect 2716 3647 2724 3753
rect 2756 3727 2764 3753
rect 2796 3687 2804 3933
rect 2856 3867 2864 4273
rect 2896 3827 2904 4033
rect 2916 3907 2924 4253
rect 2936 3827 2944 4193
rect 2956 4187 2964 4413
rect 2976 4227 2984 4413
rect 3016 4407 3024 4492
rect 3056 4447 3064 4513
rect 2996 4347 3004 4393
rect 3096 4367 3104 4493
rect 2996 4227 3004 4333
rect 3036 4307 3044 4353
rect 3096 4304 3104 4353
rect 3116 4347 3124 4753
rect 3156 4748 3164 4793
rect 3136 4407 3144 4513
rect 3156 4427 3164 4712
rect 3176 4327 3184 4853
rect 3196 4727 3204 4793
rect 3216 4707 3224 4973
rect 3236 4907 3244 4993
rect 3216 4527 3224 4613
rect 3236 4467 3244 4573
rect 3256 4487 3264 4853
rect 3276 4747 3284 5033
rect 3300 5024 3313 5027
rect 3296 5013 3313 5024
rect 3296 4907 3304 5013
rect 3413 5004 3427 5013
rect 3356 5000 3427 5004
rect 3353 4996 3424 5000
rect 3353 4987 3367 4996
rect 3366 4980 3367 4987
rect 3376 4947 3384 4973
rect 3307 4804 3320 4807
rect 3307 4793 3324 4804
rect 3316 4767 3324 4793
rect 3336 4747 3344 4793
rect 3196 4387 3204 4433
rect 3096 4300 3164 4304
rect 3096 4296 3167 4300
rect 3153 4287 3167 4296
rect 3016 4124 3024 4233
rect 2996 4116 3024 4124
rect 2996 4044 3004 4116
rect 3036 4107 3044 4253
rect 3116 4227 3124 4273
rect 2976 4036 3004 4044
rect 2976 4007 2984 4036
rect 2976 3996 2993 4007
rect 2980 3993 2993 3996
rect 2856 3767 2864 3813
rect 3056 3784 3064 4213
rect 3196 4107 3204 4273
rect 3096 4067 3104 4093
rect 3136 4067 3144 4093
rect 3116 3967 3124 3993
rect 3036 3780 3064 3784
rect 3033 3776 3064 3780
rect 3033 3767 3047 3776
rect 3076 3767 3084 3853
rect 2856 3756 2873 3767
rect 2860 3753 2873 3756
rect 2916 3727 2924 3753
rect 2756 3627 2764 3673
rect 2656 3527 2664 3593
rect 2796 3547 2804 3633
rect 2836 3547 2844 3573
rect 2827 3484 2840 3487
rect 2827 3473 2844 3484
rect 2636 3156 2664 3164
rect 2593 3004 2607 3013
rect 2633 3004 2647 3013
rect 2593 3000 2647 3004
rect 2596 2996 2644 3000
rect 2476 2956 2493 2967
rect 2480 2953 2493 2956
rect 2416 2907 2424 2953
rect 2616 2907 2624 2953
rect 2656 2847 2664 3156
rect 2676 3067 2684 3473
rect 2736 3307 2744 3473
rect 2716 3207 2724 3233
rect 2756 3187 2764 3233
rect 2796 3207 2804 3413
rect 2836 3347 2844 3473
rect 2836 3207 2844 3233
rect 2696 3147 2704 3173
rect 2856 3167 2864 3713
rect 3096 3687 3104 3713
rect 2956 3607 2964 3633
rect 2996 3547 3004 3573
rect 3076 3544 3084 3653
rect 3096 3607 3104 3633
rect 3116 3587 3124 3813
rect 3136 3648 3144 3813
rect 3176 3767 3184 3993
rect 3216 3924 3224 4313
rect 3236 4127 3244 4213
rect 3276 4207 3284 4453
rect 3296 4407 3304 4693
rect 3316 4487 3324 4653
rect 3356 4587 3364 4693
rect 3376 4687 3384 4733
rect 3416 4627 3424 4933
rect 3436 4707 3444 4953
rect 3456 4807 3464 4913
rect 3516 4907 3524 5033
rect 3496 4768 3504 4793
rect 3476 4667 3484 4713
rect 3496 4667 3504 4732
rect 3536 4687 3544 4813
rect 3556 4667 3564 5133
rect 3656 5107 3664 5153
rect 3676 5147 3684 5233
rect 3716 5107 3724 5233
rect 3707 5096 3724 5107
rect 3707 5093 3720 5096
rect 3396 4616 3413 4624
rect 3336 4447 3344 4513
rect 3316 4347 3324 4413
rect 3396 4387 3404 4616
rect 3476 4587 3484 4613
rect 3536 4547 3544 4613
rect 3576 4524 3584 5093
rect 3596 4707 3604 5033
rect 3636 5007 3644 5093
rect 3687 5044 3700 5047
rect 3687 5040 3704 5044
rect 3687 5033 3707 5040
rect 3693 5027 3707 5033
rect 3656 4867 3664 4973
rect 3596 4693 3613 4707
rect 3596 4587 3604 4693
rect 3636 4587 3644 4713
rect 3676 4627 3684 4753
rect 3696 4667 3704 4813
rect 3736 4747 3744 5133
rect 3816 5107 3824 5232
rect 3787 5104 3800 5107
rect 3787 5093 3804 5104
rect 3796 5084 3804 5093
rect 3796 5076 3884 5084
rect 3876 5047 3884 5076
rect 3796 5007 3804 5033
rect 3856 4987 3864 5033
rect 3896 5007 3904 5133
rect 3733 4644 3747 4653
rect 3716 4640 3747 4644
rect 3716 4636 3744 4640
rect 3716 4587 3724 4636
rect 3756 4627 3764 4953
rect 3796 4867 3804 4953
rect 3916 4904 3924 4993
rect 3936 4947 3944 5213
rect 3956 5107 3964 5316
rect 4047 5316 4064 5327
rect 4047 5313 4060 5316
rect 4076 5227 4084 5413
rect 4116 5227 4124 5373
rect 4156 5327 4164 5433
rect 4176 5427 4184 5773
rect 4196 5407 4204 5793
rect 4236 5788 4244 5813
rect 4276 5787 4284 5833
rect 4296 5807 4304 5853
rect 4216 5544 4224 5653
rect 4236 5567 4244 5752
rect 4296 5727 4304 5793
rect 4296 5607 4304 5713
rect 4216 5536 4244 5544
rect 4216 5384 4224 5513
rect 4187 5376 4224 5384
rect 4236 5348 4244 5536
rect 4207 5316 4233 5324
rect 4256 5287 4264 5593
rect 4376 5567 4384 5653
rect 4396 5627 4404 5853
rect 4476 5727 4484 5813
rect 3996 5107 4004 5213
rect 3896 4896 3924 4904
rect 3896 4827 3904 4896
rect 3796 4816 3833 4824
rect 3796 4767 3804 4816
rect 3976 4807 3984 4973
rect 4016 4907 4024 5013
rect 4056 4907 4064 5133
rect 4076 4867 4084 5153
rect 4096 5047 4104 5133
rect 4116 5007 4124 5093
rect 4156 5007 4164 5093
rect 4196 5004 4204 5213
rect 4276 5168 4284 5373
rect 4316 5327 4324 5413
rect 4336 5387 4344 5513
rect 4376 5327 4384 5433
rect 4367 5316 4384 5327
rect 4367 5313 4380 5316
rect 4276 5107 4284 5132
rect 4240 5104 4253 5107
rect 4236 5093 4253 5104
rect 4276 5096 4293 5107
rect 4280 5093 4293 5096
rect 4236 5047 4244 5093
rect 4300 5044 4313 5047
rect 4296 5033 4313 5044
rect 4196 4996 4224 5004
rect 4007 4856 4033 4864
rect 4136 4807 4144 4933
rect 4067 4796 4093 4804
rect 3936 4747 3944 4793
rect 3796 4584 3804 4693
rect 3856 4604 3864 4733
rect 3916 4647 3924 4673
rect 3856 4596 3904 4604
rect 3896 4587 3904 4596
rect 3767 4576 3804 4584
rect 3847 4576 3873 4584
rect 3896 4576 3913 4587
rect 3900 4573 3913 4576
rect 3556 4516 3584 4524
rect 3456 4467 3464 4513
rect 3556 4487 3564 4516
rect 3416 4347 3424 4433
rect 3456 4347 3464 4393
rect 3307 4336 3324 4347
rect 3307 4333 3320 4336
rect 3396 4247 3404 4273
rect 3356 4187 3364 4233
rect 3376 4147 3384 4173
rect 3436 4167 3444 4273
rect 3456 4167 3464 4333
rect 3496 4187 3504 4293
rect 3516 4207 3524 4473
rect 3547 4444 3560 4447
rect 3547 4433 3564 4444
rect 3556 4307 3564 4433
rect 3576 4187 3584 4493
rect 3616 4467 3624 4513
rect 3316 4067 3324 4133
rect 3260 4064 3273 4067
rect 3256 4053 3273 4064
rect 3256 3927 3264 4053
rect 3336 4007 3344 4113
rect 3376 4047 3384 4133
rect 3296 3967 3304 3993
rect 3436 3984 3444 4033
rect 3396 3976 3444 3984
rect 3396 3964 3404 3976
rect 3367 3956 3404 3964
rect 3216 3916 3244 3924
rect 3216 3767 3224 3893
rect 3236 3867 3244 3916
rect 3316 3827 3324 3873
rect 3247 3816 3273 3824
rect 3376 3767 3384 3853
rect 3436 3827 3444 3873
rect 3320 3764 3333 3767
rect 3316 3760 3333 3764
rect 3313 3753 3333 3760
rect 3313 3747 3327 3753
rect 3076 3536 3113 3544
rect 2876 3407 2884 3473
rect 2956 3447 2964 3533
rect 3136 3487 3144 3612
rect 3156 3547 3164 3593
rect 2976 3407 2984 3473
rect 2876 3367 2884 3393
rect 3036 3307 3044 3413
rect 3136 3307 3144 3373
rect 3196 3367 3204 3633
rect 3236 3547 3244 3613
rect 3276 3487 3284 3593
rect 3316 3547 3324 3633
rect 3276 3476 3293 3487
rect 3280 3473 3293 3476
rect 3256 3347 3264 3453
rect 2876 3207 2884 3233
rect 2696 3027 2704 3133
rect 2687 3016 2704 3027
rect 2687 3013 2700 3016
rect 2076 2776 2113 2784
rect 2076 2747 2084 2776
rect 1656 2427 1664 2513
rect 1836 2487 1844 2533
rect 1876 2507 1884 2533
rect 1936 2507 1944 2733
rect 1927 2496 1944 2507
rect 1996 2507 2004 2693
rect 1996 2496 2013 2507
rect 1927 2493 1940 2496
rect 2000 2493 2013 2496
rect 2096 2504 2104 2713
rect 2236 2667 2244 2773
rect 2353 2724 2367 2733
rect 2376 2724 2384 2813
rect 2353 2720 2393 2724
rect 2356 2716 2393 2720
rect 2156 2507 2164 2633
rect 2067 2496 2104 2504
rect 2180 2504 2193 2507
rect 2176 2493 2193 2504
rect 2113 2484 2127 2493
rect 2176 2484 2184 2493
rect 2113 2480 2184 2484
rect 2116 2476 2184 2480
rect 1716 2427 1724 2473
rect 1736 2456 1793 2464
rect 1736 2427 1744 2456
rect 1853 2444 1867 2453
rect 1853 2440 1993 2444
rect 1856 2436 1993 2440
rect 1716 2416 1733 2427
rect 1720 2413 1733 2416
rect 1776 2387 1784 2413
rect 1816 2347 1824 2393
rect 1976 2307 1984 2353
rect 1636 2267 1644 2293
rect 1756 2267 1764 2293
rect 1580 2264 1593 2267
rect 1576 2253 1593 2264
rect 1576 2167 1584 2253
rect 1813 2244 1827 2253
rect 1796 2240 1827 2244
rect 1796 2236 1824 2240
rect 1600 2204 1613 2207
rect 1596 2200 1613 2204
rect 1593 2193 1613 2200
rect 1667 2196 1693 2204
rect 1796 2204 1804 2236
rect 1767 2196 1804 2204
rect 1593 2187 1607 2193
rect 1816 2167 1824 2213
rect 1896 2167 1904 2193
rect 1936 2167 1944 2193
rect 1476 1987 1484 2053
rect 1527 1984 1540 1987
rect 1527 1973 1544 1984
rect 1536 1907 1544 1973
rect 1556 1927 1564 2073
rect 1416 1536 1444 1544
rect 1436 1287 1444 1536
rect 1376 1067 1384 1173
rect 1436 947 1444 1093
rect 1416 807 1424 873
rect 1456 767 1464 1673
rect 1476 1587 1484 1733
rect 1536 1687 1544 1773
rect 1576 1687 1584 2153
rect 1976 2144 1984 2293
rect 2116 2267 2124 2293
rect 2107 2256 2124 2267
rect 2107 2253 2120 2256
rect 1956 2136 1984 2144
rect 1616 1867 1624 2073
rect 1696 1996 1773 2004
rect 1696 1967 1704 1996
rect 1847 1996 1893 2004
rect 1636 1920 1713 1924
rect 1633 1916 1713 1920
rect 1633 1907 1647 1916
rect 1676 1867 1684 1893
rect 1676 1807 1684 1853
rect 1627 1676 1653 1684
rect 1696 1647 1704 1673
rect 1736 1627 1744 1793
rect 1496 1307 1504 1453
rect 1556 1407 1564 1533
rect 1656 1467 1664 1493
rect 1516 1347 1524 1393
rect 1616 1367 1624 1453
rect 1676 1407 1684 1533
rect 1736 1407 1744 1613
rect 1756 1487 1764 1593
rect 1776 1527 1784 1833
rect 1836 1807 1844 1953
rect 1893 1944 1907 1953
rect 1893 1940 1924 1944
rect 1896 1936 1924 1940
rect 1896 1824 1904 1893
rect 1916 1867 1924 1936
rect 1916 1827 1924 1853
rect 1956 1847 1964 2136
rect 2076 2127 2084 2213
rect 2116 2087 2124 2213
rect 1993 1984 2007 1993
rect 1993 1980 2033 1984
rect 1996 1976 2033 1980
rect 2116 1984 2124 2073
rect 2087 1976 2124 1984
rect 2067 1924 2080 1927
rect 2067 1913 2084 1924
rect 1876 1816 1904 1824
rect 1876 1787 1884 1816
rect 1893 1784 1907 1793
rect 1976 1784 1984 1913
rect 1893 1780 1984 1784
rect 1896 1776 1984 1780
rect 1836 1736 1873 1744
rect 1816 1567 1824 1733
rect 1836 1627 1844 1736
rect 1900 1744 1913 1747
rect 1896 1733 1913 1744
rect 1856 1607 1864 1673
rect 1896 1647 1904 1733
rect 2036 1607 2044 1693
rect 1736 1393 1753 1407
rect 1736 1347 1744 1393
rect 1476 787 1484 933
rect 1516 927 1524 1053
rect 1596 1047 1604 1213
rect 1636 1187 1644 1313
rect 1776 1307 1784 1453
rect 1816 1267 1824 1453
rect 1696 1167 1704 1253
rect 1876 1227 1884 1513
rect 1896 1407 1904 1473
rect 1916 1347 1924 1573
rect 1956 1484 1964 1593
rect 2056 1587 2064 1813
rect 2076 1684 2084 1913
rect 2096 1907 2104 1976
rect 2116 1867 2124 1953
rect 2116 1744 2124 1853
rect 2136 1827 2144 2113
rect 2176 1824 2184 2413
rect 2216 2404 2224 2633
rect 2196 2396 2224 2404
rect 2196 2307 2204 2396
rect 2236 2367 2244 2653
rect 2276 2327 2284 2593
rect 2356 2507 2364 2533
rect 2316 2407 2324 2493
rect 2436 2427 2444 2713
rect 2476 2687 2484 2773
rect 2516 2727 2524 2813
rect 2556 2627 2564 2713
rect 2656 2607 2664 2833
rect 2676 2807 2684 2953
rect 2716 2807 2724 2833
rect 2656 2507 2664 2593
rect 2576 2500 2613 2504
rect 2573 2496 2613 2500
rect 2573 2487 2587 2496
rect 2696 2447 2704 2613
rect 2416 2416 2433 2424
rect 2276 2167 2284 2273
rect 2276 2067 2284 2153
rect 2316 1967 2324 2313
rect 2336 2047 2344 2413
rect 2376 2287 2384 2353
rect 2416 2267 2424 2416
rect 2496 2367 2504 2413
rect 2536 2227 2544 2433
rect 2596 2227 2604 2333
rect 2376 2027 2384 2213
rect 2636 2087 2644 2433
rect 2696 2287 2704 2433
rect 2636 2064 2644 2073
rect 2636 2056 2664 2064
rect 2456 1987 2464 2013
rect 2400 1984 2413 1987
rect 2396 1973 2413 1984
rect 2176 1816 2204 1824
rect 2096 1736 2124 1744
rect 2096 1707 2104 1736
rect 2076 1676 2104 1684
rect 2096 1547 2104 1676
rect 2136 1607 2144 1733
rect 2176 1527 2184 1593
rect 1993 1504 2007 1513
rect 1936 1476 1964 1484
rect 1976 1500 2007 1504
rect 1976 1496 2004 1500
rect 1936 1387 1944 1476
rect 1976 1447 1984 1496
rect 2033 1464 2047 1473
rect 2116 1467 2124 1493
rect 2033 1460 2073 1464
rect 2036 1456 2073 1460
rect 1967 1436 1984 1447
rect 1967 1433 1980 1436
rect 2176 1407 2184 1513
rect 1960 1384 1973 1387
rect 1956 1373 1973 1384
rect 1956 1347 1964 1373
rect 1896 1227 1904 1253
rect 1896 1216 1913 1227
rect 1900 1213 1913 1216
rect 1736 1127 1744 1153
rect 1776 1127 1784 1173
rect 1776 927 1784 1033
rect 1836 927 1844 1053
rect 1956 1027 1964 1333
rect 2056 1187 2064 1393
rect 2136 1367 2144 1393
rect 2176 1287 2184 1393
rect 2047 1176 2064 1187
rect 2047 1173 2060 1176
rect 2093 1164 2107 1173
rect 2093 1160 2124 1164
rect 2096 1156 2124 1160
rect 2116 1127 2124 1156
rect 1516 913 1533 927
rect 1556 916 1593 924
rect 1516 764 1524 913
rect 1556 904 1564 916
rect 1536 896 1564 904
rect 1536 867 1544 896
rect 1496 756 1524 764
rect 1396 727 1404 753
rect 1496 547 1504 756
rect 1516 647 1524 733
rect 1536 727 1544 773
rect 1636 747 1644 773
rect 1716 767 1724 873
rect 1916 787 1924 1013
rect 2016 927 2024 1033
rect 1956 807 1964 873
rect 1636 707 1644 733
rect 1716 647 1724 693
rect 1836 647 1844 773
rect 2016 767 2024 793
rect 1707 636 1724 647
rect 1707 633 1720 636
rect 1656 607 1664 633
rect 1096 367 1104 453
rect 1236 427 1244 473
rect 1396 427 1404 453
rect 1447 424 1460 427
rect 1447 413 1464 424
rect 1273 404 1287 413
rect 1207 400 1287 404
rect 1207 396 1284 400
rect 676 247 684 293
rect 676 187 684 233
rect 796 187 804 233
rect 916 187 924 213
rect 1016 187 1024 273
rect 1036 147 1044 293
rect 1096 147 1104 273
rect 1216 187 1224 273
rect 1213 164 1227 173
rect 1213 160 1244 164
rect 1216 156 1244 160
rect 716 140 753 144
rect 713 136 753 140
rect 713 127 727 136
rect 896 87 904 133
rect 1236 127 1244 156
rect 936 87 944 113
rect 976 47 984 113
rect 1256 47 1264 173
rect 1296 87 1304 353
rect 1376 267 1384 353
rect 1456 347 1464 413
rect 1476 367 1484 493
rect 1496 407 1504 533
rect 1556 407 1564 493
rect 1507 336 1553 344
rect 1516 296 1553 304
rect 1376 127 1384 253
rect 1456 187 1464 253
rect 1516 187 1524 296
rect 1367 116 1384 127
rect 1367 113 1380 116
rect 1476 87 1484 113
rect 1516 47 1524 113
rect 1536 104 1544 233
rect 1576 147 1584 533
rect 1796 507 1804 613
rect 1836 607 1844 633
rect 1656 380 1724 384
rect 1656 376 1727 380
rect 1656 344 1664 376
rect 1713 367 1727 376
rect 1687 364 1700 367
rect 1687 353 1704 364
rect 1627 336 1664 344
rect 1696 327 1704 353
rect 1616 147 1624 293
rect 1816 267 1824 413
rect 1876 407 1884 533
rect 1916 407 1924 733
rect 1976 727 1984 753
rect 2016 727 2024 753
rect 2036 667 2044 1013
rect 2076 824 2084 1073
rect 2116 1047 2124 1113
rect 2136 1068 2144 1253
rect 2196 1244 2204 1816
rect 2276 1747 2284 1833
rect 2267 1676 2304 1684
rect 2216 1567 2224 1673
rect 2256 1507 2264 1613
rect 2216 1287 2224 1353
rect 2276 1327 2284 1653
rect 2296 1627 2304 1676
rect 2316 1667 2324 1953
rect 2396 1907 2404 1973
rect 2356 1747 2364 1893
rect 2373 1864 2387 1873
rect 2373 1860 2404 1864
rect 2376 1856 2404 1860
rect 2316 1467 2324 1493
rect 2196 1236 2224 1244
rect 2196 1067 2204 1213
rect 2216 1167 2224 1236
rect 2296 1164 2304 1213
rect 2336 1164 2344 1373
rect 2356 1267 2364 1493
rect 2376 1307 2384 1653
rect 2396 1647 2404 1856
rect 2436 1847 2444 1913
rect 2476 1827 2484 1893
rect 2396 1407 2404 1453
rect 2416 1407 2424 1533
rect 2496 1304 2504 2033
rect 2520 1964 2533 1967
rect 2516 1953 2533 1964
rect 2516 1867 2524 1953
rect 2596 1884 2604 1953
rect 2576 1876 2604 1884
rect 2576 1827 2584 1876
rect 2556 1767 2564 1793
rect 2596 1747 2604 1773
rect 2516 1687 2524 1733
rect 2516 1676 2533 1687
rect 2520 1673 2533 1676
rect 2576 1627 2584 1673
rect 2616 1647 2624 1833
rect 2656 1784 2664 2056
rect 2716 1927 2724 2053
rect 2647 1776 2664 1784
rect 2636 1687 2644 1773
rect 2596 1447 2604 1473
rect 2547 1436 2584 1444
rect 2576 1424 2584 1436
rect 2576 1420 2624 1424
rect 2576 1416 2627 1420
rect 2613 1407 2627 1416
rect 2596 1304 2604 1373
rect 2636 1307 2644 1593
rect 2676 1387 2684 1733
rect 2736 1627 2744 3153
rect 2756 2647 2764 3053
rect 2796 3027 2804 3073
rect 2816 2967 2824 3133
rect 2916 3027 2924 3093
rect 2936 3067 2944 3293
rect 3096 3256 3184 3264
rect 3096 3224 3104 3256
rect 3076 3216 3104 3224
rect 3076 3204 3084 3216
rect 3116 3207 3124 3233
rect 3047 3196 3084 3204
rect 3156 3187 3164 3233
rect 3176 3187 3184 3256
rect 2956 3027 2964 3113
rect 2847 3024 2860 3027
rect 2847 3013 2864 3024
rect 2776 2787 2784 2933
rect 2856 2927 2864 3013
rect 3056 2967 3064 3073
rect 3096 3027 3104 3133
rect 3136 3067 3144 3093
rect 3136 3027 3144 3053
rect 3216 3027 3224 3093
rect 3236 3027 3244 3293
rect 3316 3247 3324 3433
rect 3356 3407 3364 3673
rect 3456 3647 3464 3753
rect 3476 3727 3484 4133
rect 3536 3887 3544 4173
rect 3636 4147 3644 4473
rect 3676 4467 3684 4573
rect 3867 4516 3893 4524
rect 3736 4467 3744 4513
rect 3696 4407 3704 4433
rect 3776 4367 3784 4493
rect 3676 4187 3684 4333
rect 3556 4007 3564 4133
rect 3736 4107 3744 4353
rect 3796 4307 3804 4473
rect 3816 4347 3824 4433
rect 3787 4296 3804 4307
rect 3787 4293 3800 4296
rect 3756 4127 3764 4233
rect 3816 4227 3824 4333
rect 3796 4167 3804 4193
rect 3856 4187 3864 4393
rect 3936 4387 3944 4493
rect 3956 4407 3964 4713
rect 3976 4467 3984 4713
rect 4016 4487 4024 4633
rect 4036 4587 4044 4613
rect 4056 4544 4064 4753
rect 4076 4627 4084 4733
rect 4096 4627 4104 4753
rect 4136 4727 4144 4793
rect 4156 4667 4164 4713
rect 4176 4647 4184 4733
rect 4216 4727 4224 4996
rect 4276 4987 4284 5033
rect 4296 5007 4304 5033
rect 4196 4587 4204 4693
rect 4036 4536 4064 4544
rect 4036 4467 4044 4536
rect 4056 4487 4064 4513
rect 3913 4284 3927 4293
rect 3996 4287 4004 4373
rect 3913 4280 3953 4284
rect 3916 4276 3953 4280
rect 3956 4127 3964 4273
rect 3756 4067 3764 4113
rect 3856 4067 3864 4113
rect 4036 4067 4044 4393
rect 4096 4387 4104 4473
rect 4116 4427 4124 4573
rect 4156 4467 4164 4573
rect 4176 4407 4184 4493
rect 4236 4487 4244 4913
rect 4296 4807 4304 4993
rect 4316 4927 4324 4993
rect 4336 4967 4344 5253
rect 4356 4967 4364 5093
rect 4396 5064 4404 5493
rect 4416 5467 4424 5653
rect 4536 5627 4544 5773
rect 4576 5707 4584 5833
rect 4596 5787 4604 5893
rect 4616 5764 4624 5993
rect 4796 5976 4864 5984
rect 4796 5947 4804 5976
rect 4856 5964 4864 5976
rect 4856 5956 4884 5964
rect 4656 5907 4664 5933
rect 4836 5907 4844 5953
rect 4776 5896 4833 5904
rect 4776 5867 4784 5896
rect 4876 5867 4884 5956
rect 4916 5864 4924 5973
rect 4956 5947 4964 5973
rect 5176 5964 5184 5993
rect 5176 5956 5204 5964
rect 4953 5927 4967 5933
rect 4953 5920 4973 5927
rect 4956 5916 4973 5920
rect 4960 5913 4973 5916
rect 5013 5904 5027 5913
rect 4976 5900 5027 5904
rect 5133 5904 5147 5913
rect 5133 5900 5173 5904
rect 4976 5896 5024 5900
rect 5136 5896 5173 5900
rect 4916 5856 4953 5864
rect 4596 5756 4624 5764
rect 4596 5667 4604 5756
rect 4480 5624 4493 5627
rect 4476 5613 4493 5624
rect 4416 5127 4424 5213
rect 4456 5147 4464 5513
rect 4476 5447 4484 5613
rect 4567 5556 4593 5564
rect 4516 5467 4524 5533
rect 4556 5407 4564 5553
rect 4616 5427 4624 5733
rect 4656 5727 4664 5773
rect 4656 5627 4664 5653
rect 4696 5627 4704 5753
rect 4656 5487 4664 5613
rect 4716 5507 4724 5573
rect 4513 5384 4527 5393
rect 4487 5380 4527 5384
rect 4487 5376 4524 5380
rect 4607 5376 4633 5384
rect 4476 5248 4484 5373
rect 4556 5267 4564 5333
rect 4636 5307 4644 5373
rect 4656 5347 4664 5413
rect 4676 5327 4684 5493
rect 4696 5407 4704 5473
rect 4736 5447 4744 5813
rect 4756 5507 4764 5773
rect 4796 5707 4804 5853
rect 4776 5607 4784 5673
rect 4816 5647 4824 5693
rect 4807 5636 4824 5647
rect 4807 5633 4820 5636
rect 4836 5547 4844 5733
rect 4876 5727 4884 5853
rect 4856 5607 4864 5713
rect 4787 5524 4800 5527
rect 4787 5513 4804 5524
rect 4796 5447 4804 5513
rect 4916 5508 4924 5793
rect 4696 5376 4773 5384
rect 4376 5056 4404 5064
rect 4336 4887 4344 4953
rect 4376 4927 4384 5056
rect 4416 5044 4424 5113
rect 4476 5087 4484 5212
rect 4396 5040 4424 5044
rect 4393 5036 4424 5040
rect 4393 5027 4407 5036
rect 4436 4987 4444 5013
rect 4516 4984 4524 5173
rect 4596 5107 4604 5133
rect 4553 5084 4567 5093
rect 4636 5084 4644 5253
rect 4696 5227 4704 5376
rect 4727 5316 4753 5324
rect 4716 5244 4724 5292
rect 4716 5240 4744 5244
rect 4716 5236 4747 5240
rect 4733 5227 4747 5236
rect 4696 5147 4704 5213
rect 4553 5080 4584 5084
rect 4556 5076 4584 5080
rect 4536 5008 4544 5033
rect 4576 4987 4584 5076
rect 4616 5076 4644 5084
rect 4616 5064 4624 5076
rect 4596 5056 4624 5064
rect 4596 5007 4604 5056
rect 4627 5036 4653 5044
rect 4496 4976 4524 4984
rect 4496 4907 4504 4976
rect 4356 4807 4364 4853
rect 4256 4747 4264 4793
rect 4296 4727 4304 4793
rect 4296 4667 4304 4713
rect 4336 4667 4344 4733
rect 4356 4587 4364 4613
rect 4327 4584 4340 4587
rect 4327 4573 4344 4584
rect 4336 4564 4344 4573
rect 4336 4556 4364 4564
rect 4296 4487 4304 4513
rect 4156 4347 4164 4373
rect 4076 4187 4084 4333
rect 4116 4107 4124 4333
rect 4176 4287 4184 4393
rect 4136 4247 4144 4273
rect 4216 4247 4224 4453
rect 4296 4407 4304 4473
rect 4256 4347 4264 4393
rect 4156 4067 4164 4093
rect 3747 4056 3764 4067
rect 3747 4053 3760 4056
rect 3907 4064 3920 4067
rect 3907 4053 3924 4064
rect 3596 3907 3604 3993
rect 3696 3967 3704 4053
rect 3727 4004 3740 4007
rect 3727 3993 3744 4004
rect 3736 3947 3744 3993
rect 3536 3827 3544 3873
rect 3516 3727 3524 3753
rect 3556 3667 3564 3753
rect 3396 3547 3404 3593
rect 3456 3547 3464 3633
rect 3596 3627 3604 3813
rect 3636 3707 3644 3893
rect 3716 3887 3724 3913
rect 3696 3827 3704 3853
rect 3716 3767 3724 3873
rect 3836 3867 3844 3973
rect 3876 3947 3884 3993
rect 3916 3967 3924 4053
rect 3676 3667 3684 3753
rect 3776 3687 3784 3753
rect 3447 3536 3464 3547
rect 3447 3533 3460 3536
rect 3416 3447 3424 3473
rect 3356 3307 3364 3393
rect 3556 3387 3564 3473
rect 3376 3307 3384 3373
rect 3576 3367 3584 3533
rect 3496 3307 3504 3333
rect 3596 3307 3604 3573
rect 3633 3547 3647 3553
rect 3627 3540 3647 3547
rect 3627 3536 3644 3540
rect 3627 3533 3640 3536
rect 3647 3476 3673 3484
rect 3696 3407 3704 3553
rect 3736 3547 3744 3613
rect 3736 3536 3753 3547
rect 3740 3533 3753 3536
rect 3776 3487 3784 3573
rect 3796 3547 3804 3693
rect 3836 3687 3844 3813
rect 3856 3667 3864 3733
rect 3856 3547 3864 3613
rect 3876 3607 3884 3853
rect 3936 3827 3944 3933
rect 3996 3927 4004 4053
rect 4016 3907 4024 3973
rect 4056 3967 4064 3993
rect 3916 3727 3924 3753
rect 3856 3536 3873 3547
rect 3860 3533 3873 3536
rect 3896 3487 3904 3573
rect 3936 3547 3944 3693
rect 3956 3687 3964 3753
rect 3996 3727 4004 3773
rect 4056 3667 4064 3873
rect 4076 3827 4084 3913
rect 4156 3887 4164 4053
rect 4193 4044 4207 4053
rect 4193 4040 4224 4044
rect 4196 4036 4224 4040
rect 4216 4007 4224 4036
rect 4216 3867 4224 3993
rect 4256 3887 4264 4233
rect 4296 3947 4304 4273
rect 4316 4207 4324 4473
rect 4336 4067 4344 4493
rect 4356 4447 4364 4556
rect 4376 4467 4384 4873
rect 4416 4867 4424 4893
rect 4467 4864 4480 4867
rect 4467 4853 4484 4864
rect 4396 4796 4433 4804
rect 4396 4668 4404 4796
rect 4416 4627 4424 4753
rect 4476 4747 4484 4853
rect 4496 4644 4504 4713
rect 4516 4707 4524 4933
rect 4476 4636 4504 4644
rect 4396 4528 4404 4613
rect 4476 4604 4484 4636
rect 4536 4607 4544 4972
rect 4676 4927 4684 5113
rect 4716 4907 4724 5193
rect 4756 5047 4764 5233
rect 4796 5107 4804 5313
rect 4836 5207 4844 5493
rect 4916 5327 4924 5472
rect 4860 5324 4873 5327
rect 4856 5313 4873 5324
rect 4856 5227 4864 5313
rect 4836 5107 4844 5133
rect 4876 5107 4884 5153
rect 4796 5064 4804 5093
rect 4796 5056 4844 5064
rect 4836 5047 4844 5056
rect 4836 5036 4853 5047
rect 4840 5033 4853 5036
rect 4896 5024 4904 5233
rect 4916 5227 4924 5273
rect 4936 5168 4944 5673
rect 4956 5627 4964 5853
rect 4976 5787 4984 5896
rect 5196 5867 5204 5956
rect 5216 5907 5224 5973
rect 5256 5967 5264 5993
rect 5256 5927 5264 5953
rect 5120 5864 5133 5867
rect 5116 5853 5133 5864
rect 4976 5687 4984 5773
rect 5036 5767 5044 5853
rect 5116 5807 5124 5853
rect 4996 5627 5004 5673
rect 4960 5564 4973 5567
rect 4956 5560 4973 5564
rect 4953 5553 4973 5560
rect 4953 5547 4967 5553
rect 5036 5507 5044 5753
rect 5156 5704 5164 5773
rect 5136 5696 5164 5704
rect 5096 5527 5104 5693
rect 5116 5507 5124 5593
rect 5136 5567 5144 5696
rect 5176 5627 5184 5673
rect 5136 5556 5153 5567
rect 5140 5553 5153 5556
rect 5236 5527 5244 5853
rect 5296 5808 5304 5973
rect 5336 5967 5344 6044
rect 5356 6036 5384 6044
rect 5416 6036 5444 6044
rect 5356 5987 5364 6036
rect 5416 5964 5424 6036
rect 5476 5967 5484 6044
rect 5416 5956 5444 5964
rect 5376 5927 5384 5953
rect 5396 5904 5404 5933
rect 5356 5896 5404 5904
rect 5356 5867 5364 5896
rect 5276 5687 5284 5753
rect 5296 5667 5304 5772
rect 5316 5724 5324 5853
rect 5396 5827 5404 5853
rect 5436 5827 5444 5956
rect 5516 5847 5524 5993
rect 5416 5747 5424 5793
rect 5476 5787 5484 5833
rect 5316 5716 5333 5724
rect 5296 5627 5304 5653
rect 5336 5627 5344 5713
rect 5256 5564 5264 5593
rect 5256 5556 5304 5564
rect 4876 5016 4904 5024
rect 4796 4948 4804 4973
rect 4556 4807 4564 4893
rect 4660 4864 4673 4867
rect 4656 4853 4673 4864
rect 4556 4687 4564 4753
rect 4596 4747 4604 4793
rect 4636 4747 4644 4853
rect 4656 4807 4664 4853
rect 4713 4844 4727 4853
rect 4713 4840 4764 4844
rect 4716 4836 4764 4840
rect 4696 4767 4704 4793
rect 4736 4747 4744 4793
rect 4756 4787 4764 4836
rect 4756 4776 4773 4787
rect 4760 4773 4773 4776
rect 4796 4724 4804 4912
rect 4776 4716 4804 4724
rect 4476 4596 4504 4604
rect 4496 4587 4504 4596
rect 4356 4247 4364 4433
rect 4376 4347 4384 4393
rect 4396 4304 4404 4492
rect 4456 4467 4464 4573
rect 4496 4447 4504 4573
rect 4496 4407 4504 4433
rect 4536 4307 4544 4453
rect 4576 4428 4584 4693
rect 4716 4687 4724 4713
rect 4776 4647 4784 4716
rect 4816 4647 4824 4933
rect 4856 4927 4864 4993
rect 4876 4947 4884 5016
rect 4836 4887 4844 4913
rect 4876 4768 4884 4873
rect 4836 4667 4844 4753
rect 4616 4507 4624 4593
rect 4733 4587 4747 4593
rect 4733 4580 4753 4587
rect 4736 4576 4753 4580
rect 4740 4573 4753 4576
rect 4807 4576 4844 4584
rect 4576 4347 4584 4392
rect 4376 4296 4404 4304
rect 4376 4107 4384 4296
rect 4396 4247 4404 4273
rect 4436 4247 4444 4273
rect 4616 4267 4624 4493
rect 4656 4467 4664 4493
rect 4696 4487 4704 4553
rect 4736 4467 4744 4513
rect 4436 4067 4444 4113
rect 4336 4056 4353 4067
rect 4340 4053 4353 4056
rect 4316 3967 4324 4053
rect 4136 3827 4144 3853
rect 4127 3816 4144 3827
rect 4127 3813 4140 3816
rect 4156 3787 4164 3833
rect 4176 3607 4184 3813
rect 4276 3767 4284 3853
rect 4236 3727 4244 3753
rect 4316 3727 4324 3953
rect 4336 3947 4344 3993
rect 4356 3687 4364 3853
rect 4416 3827 4424 3933
rect 4456 3904 4464 4173
rect 4496 4067 4504 4233
rect 4576 4107 4584 4213
rect 4656 4187 4664 4453
rect 4696 4367 4704 4393
rect 4736 4367 4744 4413
rect 4676 4207 4684 4233
rect 4696 4187 4704 4353
rect 4653 4067 4667 4073
rect 4487 4056 4504 4067
rect 4487 4053 4500 4056
rect 4647 4060 4667 4067
rect 4647 4056 4664 4060
rect 4647 4053 4660 4056
rect 4436 3896 4464 3904
rect 4436 3767 4444 3896
rect 4456 3827 4464 3873
rect 3927 3536 3944 3547
rect 3927 3533 3940 3536
rect 4056 3504 4064 3593
rect 4236 3547 4244 3673
rect 4356 3547 4364 3673
rect 4396 3667 4404 3753
rect 4456 3744 4464 3813
rect 4436 3736 4464 3744
rect 4167 3536 4193 3544
rect 4207 3536 4224 3544
rect 4036 3500 4064 3504
rect 4033 3496 4064 3500
rect 4216 3504 4224 3536
rect 4380 3544 4393 3547
rect 4376 3533 4393 3544
rect 4376 3524 4384 3533
rect 4327 3516 4384 3524
rect 4216 3496 4253 3504
rect 4033 3487 4047 3496
rect 4227 3484 4240 3487
rect 4227 3473 4244 3484
rect 4387 3484 4400 3487
rect 4387 3480 4404 3484
rect 4387 3473 4407 3480
rect 3996 3447 4004 3473
rect 3347 3296 3364 3307
rect 3347 3293 3360 3296
rect 3436 3260 3524 3264
rect 3433 3256 3524 3260
rect 3433 3247 3447 3256
rect 3516 3247 3524 3256
rect 3367 3236 3393 3244
rect 3527 3236 3553 3244
rect 3476 3207 3484 3233
rect 3636 3207 3644 3373
rect 3956 3347 3964 3433
rect 3700 3304 3713 3307
rect 3696 3293 3713 3304
rect 3696 3247 3704 3293
rect 3776 3247 3784 3333
rect 3996 3324 4004 3433
rect 4076 3407 4084 3473
rect 4236 3467 4244 3473
rect 4236 3456 4253 3467
rect 4240 3453 4253 3456
rect 4316 3367 4324 3473
rect 4393 3467 4407 3473
rect 4436 3427 4444 3736
rect 4496 3707 4504 3993
rect 4596 3927 4604 4053
rect 4716 4007 4724 4113
rect 4736 4067 4744 4293
rect 4776 4127 4784 4433
rect 4796 4344 4804 4453
rect 4836 4427 4844 4576
rect 4856 4447 4864 4713
rect 4876 4627 4884 4732
rect 4876 4407 4884 4553
rect 4896 4408 4904 4993
rect 4916 4708 4924 4953
rect 4936 4804 4944 5132
rect 4956 5107 4964 5473
rect 4956 4867 4964 4933
rect 4976 4907 4984 5493
rect 4996 5387 5004 5413
rect 5036 5264 5044 5373
rect 5056 5327 5064 5413
rect 5087 5376 5113 5384
rect 5096 5267 5104 5313
rect 5016 5256 5044 5264
rect 5016 5147 5024 5256
rect 5036 5187 5044 5213
rect 5116 5107 5124 5133
rect 4996 4927 5004 5033
rect 5036 4987 5044 5093
rect 5056 4967 5064 5033
rect 5136 4987 5144 5193
rect 5156 5107 5164 5253
rect 5176 5147 5184 5373
rect 5196 5327 5204 5453
rect 5236 5327 5244 5453
rect 5276 5307 5284 5533
rect 5296 5347 5304 5556
rect 5336 5467 5344 5553
rect 5376 5467 5384 5693
rect 5456 5627 5464 5693
rect 5416 5524 5424 5613
rect 5436 5527 5444 5553
rect 5396 5516 5424 5524
rect 5316 5344 5324 5433
rect 5356 5387 5364 5433
rect 5316 5336 5344 5344
rect 5336 5324 5344 5336
rect 5396 5327 5404 5516
rect 5436 5487 5444 5513
rect 5496 5507 5504 5593
rect 5456 5404 5464 5493
rect 5516 5447 5524 5793
rect 5556 5707 5564 5933
rect 5776 5907 5784 5933
rect 5587 5896 5613 5904
rect 5636 5807 5644 5833
rect 5533 5544 5547 5553
rect 5576 5547 5584 5673
rect 5736 5667 5744 5893
rect 5913 5884 5927 5893
rect 5913 5880 5944 5884
rect 5916 5876 5944 5880
rect 5896 5807 5904 5833
rect 5776 5627 5784 5673
rect 5720 5624 5733 5627
rect 5716 5613 5733 5624
rect 5533 5540 5573 5544
rect 5536 5536 5573 5540
rect 5616 5507 5624 5533
rect 5436 5400 5464 5404
rect 5433 5396 5464 5400
rect 5433 5387 5447 5396
rect 5336 5316 5364 5324
rect 5196 5187 5204 5273
rect 4956 4856 4973 4867
rect 4960 4853 4973 4856
rect 5056 4807 5064 4833
rect 4936 4796 4964 4804
rect 4936 4707 4944 4773
rect 4956 4727 4964 4796
rect 5047 4796 5064 4807
rect 5047 4793 5060 4796
rect 4996 4747 5004 4793
rect 5036 4767 5044 4793
rect 4916 4587 4924 4672
rect 5036 4647 5044 4713
rect 5056 4667 5064 4733
rect 5076 4647 5084 4973
rect 5096 4667 5104 4893
rect 5136 4807 5144 4893
rect 5116 4707 5124 4733
rect 5156 4687 5164 4933
rect 5196 4847 5204 4973
rect 5196 4807 5204 4833
rect 5187 4796 5204 4807
rect 5216 4804 5224 5153
rect 5236 4824 5244 5133
rect 5276 5107 5284 5193
rect 5296 5147 5304 5233
rect 5316 5107 5324 5313
rect 5356 5307 5364 5316
rect 5356 5296 5373 5307
rect 5360 5293 5373 5296
rect 5256 4947 5264 5033
rect 5356 4907 5364 5273
rect 5456 5267 5464 5313
rect 5476 5147 5484 5373
rect 5496 5327 5504 5413
rect 5576 5287 5584 5493
rect 5596 5387 5604 5413
rect 5636 5344 5644 5593
rect 5616 5340 5644 5344
rect 5613 5336 5644 5340
rect 5613 5327 5627 5336
rect 5656 5327 5664 5553
rect 5716 5547 5724 5613
rect 5407 5096 5433 5104
rect 5513 5104 5527 5113
rect 5487 5100 5527 5104
rect 5487 5096 5524 5100
rect 5236 4816 5264 4824
rect 5256 4807 5264 4816
rect 5216 4796 5244 4804
rect 5256 4796 5273 4807
rect 5187 4793 5200 4796
rect 5236 4707 5244 4796
rect 5260 4793 5273 4796
rect 4956 4587 4964 4633
rect 4796 4336 4833 4344
rect 4896 4287 4904 4372
rect 4976 4347 4984 4533
rect 4996 4364 5004 4613
rect 5056 4587 5064 4613
rect 5236 4587 5244 4613
rect 5080 4584 5093 4587
rect 5076 4573 5093 4584
rect 5076 4544 5084 4573
rect 5193 4564 5207 4573
rect 5256 4564 5264 4713
rect 5193 4560 5264 4564
rect 5196 4556 5264 4560
rect 5056 4536 5084 4544
rect 5276 4544 5284 4693
rect 5296 4627 5304 4853
rect 5327 4804 5340 4807
rect 5327 4793 5344 4804
rect 5276 4540 5304 4544
rect 5276 4536 5307 4540
rect 5036 4467 5044 4513
rect 4996 4356 5024 4364
rect 4976 4333 4993 4347
rect 4840 4284 4853 4287
rect 4836 4280 4853 4284
rect 4833 4273 4853 4280
rect 4833 4267 4847 4273
rect 4836 4167 4844 4253
rect 4956 4227 4964 4333
rect 4976 4307 4984 4333
rect 5016 4287 5024 4356
rect 5056 4287 5064 4536
rect 5293 4527 5307 4536
rect 5076 4427 5084 4493
rect 5116 4467 5124 4513
rect 5216 4487 5224 4513
rect 5096 4347 5104 4373
rect 4736 4056 4753 4067
rect 4740 4053 4753 4056
rect 4716 3993 4733 4007
rect 4656 3967 4664 3993
rect 4716 3967 4724 3993
rect 4576 3916 4593 3924
rect 4536 3627 4544 3813
rect 4576 3767 4584 3916
rect 4776 3884 4784 3973
rect 4796 3907 4804 4053
rect 4836 3927 4844 4153
rect 4896 4067 4904 4173
rect 4936 4067 4944 4193
rect 4756 3880 4784 3884
rect 4753 3876 4784 3880
rect 4616 3827 4624 3873
rect 4753 3867 4767 3876
rect 4916 3867 4924 3973
rect 4766 3860 4767 3867
rect 4607 3816 4624 3827
rect 4607 3813 4620 3816
rect 4716 3816 4753 3824
rect 4616 3707 4624 3753
rect 4516 3547 4524 3593
rect 4556 3547 4564 3573
rect 4656 3547 4664 3813
rect 4716 3707 4724 3816
rect 4776 3767 4784 3853
rect 4736 3727 4744 3753
rect 4816 3707 4824 3833
rect 4853 3827 4867 3833
rect 4853 3820 4873 3827
rect 4856 3816 4873 3820
rect 4860 3813 4873 3816
rect 4916 3767 4924 3853
rect 4907 3756 4924 3767
rect 4907 3753 4920 3756
rect 4856 3727 4864 3753
rect 4696 3547 4704 3573
rect 4476 3504 4484 3533
rect 4476 3496 4564 3504
rect 4556 3484 4564 3496
rect 4736 3487 4744 3593
rect 4836 3547 4844 3613
rect 4936 3567 4944 3813
rect 4956 3667 4964 3933
rect 4976 3588 4984 4253
rect 4996 3847 5004 4233
rect 5036 3967 5044 4053
rect 5056 4007 5064 4273
rect 5076 4107 5084 4193
rect 5116 4127 5124 4453
rect 5156 4388 5164 4453
rect 5176 4367 5184 4453
rect 5160 4366 5184 4367
rect 5167 4356 5184 4366
rect 5167 4353 5180 4356
rect 5156 4287 5164 4313
rect 5156 4276 5173 4287
rect 5160 4273 5173 4276
rect 5136 4147 5144 4233
rect 5216 4187 5224 4273
rect 5236 4267 5244 4333
rect 5076 4067 5084 4093
rect 5056 3847 5064 3913
rect 4996 3836 5013 3847
rect 5000 3833 5013 3836
rect 5116 3767 5124 4073
rect 5156 4007 5164 4113
rect 5256 4067 5264 4473
rect 5316 4427 5324 4713
rect 5336 4707 5344 4793
rect 5356 4587 5364 4893
rect 5396 4864 5404 4933
rect 5416 4907 5424 5033
rect 5436 4927 5444 4973
rect 5396 4856 5433 4864
rect 5476 4807 5484 4973
rect 5467 4796 5484 4807
rect 5467 4793 5480 4796
rect 5376 4667 5384 4753
rect 5396 4587 5404 4633
rect 5247 4056 5264 4067
rect 5247 4053 5260 4056
rect 5156 3996 5173 4007
rect 5160 3993 5173 3996
rect 5136 3967 5144 3993
rect 5196 3967 5204 4053
rect 5276 4027 5284 4413
rect 5316 4287 5324 4373
rect 5336 4287 5344 4513
rect 5336 4276 5353 4287
rect 5340 4273 5353 4276
rect 5296 3987 5304 4273
rect 5396 4268 5404 4453
rect 5396 4107 5404 4232
rect 5416 4147 5424 4673
rect 5436 4127 5444 4693
rect 5456 4387 5464 4793
rect 5496 4784 5504 5033
rect 5676 4987 5684 5493
rect 5696 5127 5704 5473
rect 5776 5467 5784 5513
rect 5696 5047 5704 5113
rect 5716 5107 5724 5433
rect 5776 5407 5784 5453
rect 5816 5407 5824 5653
rect 5840 5624 5853 5627
rect 5836 5613 5853 5624
rect 5836 5588 5844 5613
rect 5836 5447 5844 5552
rect 5896 5527 5904 5613
rect 5936 5447 5944 5876
rect 5956 5467 5964 5553
rect 5916 5387 5924 5413
rect 5516 4867 5524 4893
rect 5516 4856 5533 4867
rect 5520 4853 5533 4856
rect 5476 4776 5504 4784
rect 5476 4707 5484 4776
rect 5496 4587 5504 4673
rect 5476 4467 5484 4513
rect 5496 4447 5504 4573
rect 5516 4527 5524 4753
rect 5536 4587 5544 4793
rect 5576 4747 5584 4853
rect 5636 4747 5644 4793
rect 5656 4724 5664 4953
rect 5736 4907 5744 5373
rect 5976 5347 5984 5793
rect 5996 5627 6004 5653
rect 6033 5604 6047 5613
rect 6016 5600 6047 5604
rect 6016 5596 6044 5600
rect 6016 5527 6024 5596
rect 6076 5547 6084 5853
rect 5996 5427 6004 5453
rect 5796 5287 5804 5313
rect 5896 5227 5904 5313
rect 5936 5287 5944 5313
rect 5753 5084 5767 5093
rect 5753 5080 5804 5084
rect 5756 5076 5804 5080
rect 5636 4716 5664 4724
rect 5516 4487 5524 4513
rect 5456 4167 5464 4333
rect 5496 4287 5504 4373
rect 5496 4273 5513 4287
rect 5476 4247 5484 4273
rect 5496 4227 5504 4273
rect 5333 4067 5347 4073
rect 5516 4067 5524 4153
rect 5556 4084 5564 4453
rect 5616 4447 5624 4693
rect 5636 4564 5644 4716
rect 5676 4587 5684 4893
rect 5756 4727 5764 4813
rect 5733 4587 5747 4593
rect 5727 4580 5747 4587
rect 5727 4576 5744 4580
rect 5727 4573 5740 4576
rect 5636 4556 5664 4564
rect 5656 4464 5664 4556
rect 5676 4487 5684 4573
rect 5756 4527 5764 4653
rect 5747 4516 5764 4527
rect 5747 4513 5760 4516
rect 5656 4456 5684 4464
rect 5576 4287 5584 4393
rect 5596 4347 5604 4433
rect 5596 4336 5613 4347
rect 5600 4333 5613 4336
rect 5576 4276 5593 4287
rect 5580 4273 5593 4276
rect 5536 4076 5564 4084
rect 5333 4060 5353 4067
rect 5336 4056 5353 4060
rect 5340 4053 5353 4056
rect 5393 4044 5407 4053
rect 5433 4044 5447 4053
rect 5393 4040 5447 4044
rect 5396 4036 5444 4040
rect 5253 3964 5267 3973
rect 5336 3967 5344 3993
rect 5236 3960 5267 3964
rect 5236 3956 5264 3960
rect 5196 3867 5204 3953
rect 5236 3947 5244 3956
rect 5227 3936 5244 3947
rect 5227 3933 5240 3936
rect 5156 3827 5164 3853
rect 4556 3476 4633 3484
rect 3996 3320 4024 3324
rect 3996 3316 4027 3320
rect 4013 3307 4027 3316
rect 3887 3296 3913 3304
rect 3976 3247 3984 3293
rect 4056 3247 4064 3353
rect 4176 3247 4184 3333
rect 4356 3327 4364 3353
rect 4256 3296 4273 3304
rect 3976 3236 3993 3247
rect 3980 3233 3993 3236
rect 4047 3236 4064 3247
rect 4047 3233 4060 3236
rect 3736 3207 3744 3233
rect 4176 3147 4184 3233
rect 4216 3207 4224 3233
rect 3396 3027 3404 3053
rect 3496 3027 3504 3073
rect 3676 3027 3684 3073
rect 3816 3027 3824 3073
rect 3856 3027 3864 3053
rect 3236 3016 3253 3027
rect 3240 3013 3253 3016
rect 3327 3016 3353 3024
rect 3727 3024 3740 3027
rect 3727 3013 3744 3024
rect 3487 2956 3513 2964
rect 2936 2927 2944 2953
rect 2856 2867 2864 2913
rect 3196 2847 3204 2953
rect 2776 2776 2793 2787
rect 2780 2773 2793 2776
rect 2773 2724 2787 2733
rect 2773 2720 2813 2724
rect 2776 2716 2813 2720
rect 2856 2687 2864 2713
rect 2756 2367 2764 2593
rect 2896 2587 2904 2773
rect 2956 2647 2964 2773
rect 2996 2507 3004 2693
rect 3036 2607 3044 2733
rect 3076 2547 3084 2813
rect 3236 2787 3244 2833
rect 3156 2667 3164 2773
rect 3256 2727 3264 2853
rect 3316 2727 3324 2953
rect 3436 2727 3444 2813
rect 3476 2787 3484 2913
rect 3536 2847 3544 3013
rect 3736 2967 3744 3013
rect 3807 2956 3864 2964
rect 3656 2907 3664 2953
rect 3856 2927 3864 2956
rect 3467 2776 3484 2787
rect 3467 2773 3480 2776
rect 3627 2776 3653 2784
rect 3307 2716 3324 2727
rect 3307 2713 3320 2716
rect 3476 2687 3484 2713
rect 3156 2627 3164 2653
rect 3036 2507 3044 2533
rect 2756 2327 2764 2353
rect 2756 2287 2764 2313
rect 2816 2267 2824 2473
rect 2836 2307 2844 2353
rect 2876 2347 2884 2473
rect 2976 2384 2984 2433
rect 2976 2376 3004 2384
rect 2896 2267 2904 2293
rect 2813 2204 2827 2213
rect 2916 2207 2924 2313
rect 2956 2227 2964 2333
rect 2813 2200 2873 2204
rect 2816 2196 2873 2200
rect 2956 2067 2964 2213
rect 2956 1967 2964 2053
rect 2996 1987 3004 2376
rect 3016 2227 3024 2413
rect 2880 1964 2893 1967
rect 2876 1953 2893 1964
rect 2776 1847 2784 1913
rect 2876 1807 2884 1953
rect 2776 1567 2784 1633
rect 2816 1607 2824 1733
rect 2836 1627 2844 1673
rect 2736 1467 2744 1493
rect 2776 1467 2784 1553
rect 2756 1327 2764 1393
rect 2476 1296 2504 1304
rect 2576 1296 2604 1304
rect 2380 1164 2393 1167
rect 2267 1156 2304 1164
rect 2316 1156 2344 1164
rect 2316 1064 2324 1156
rect 2376 1153 2393 1164
rect 2316 1056 2344 1064
rect 2136 927 2144 1032
rect 2056 816 2084 824
rect 2056 747 2064 816
rect 2156 667 2164 1053
rect 2216 887 2224 973
rect 2207 876 2224 887
rect 2207 873 2220 876
rect 2256 767 2264 1013
rect 2296 947 2304 993
rect 2316 964 2324 1033
rect 2336 1007 2344 1056
rect 2356 1027 2364 1133
rect 2376 1067 2384 1153
rect 2316 956 2344 964
rect 2296 936 2313 947
rect 2300 933 2313 936
rect 2336 887 2344 956
rect 2396 887 2404 1033
rect 2387 876 2404 887
rect 2436 887 2444 973
rect 2436 876 2453 887
rect 2387 873 2400 876
rect 2440 873 2453 876
rect 2376 747 2384 873
rect 2476 848 2484 1296
rect 2496 1047 2504 1253
rect 2187 704 2200 707
rect 2187 693 2204 704
rect 2196 667 2204 693
rect 1956 627 1964 653
rect 1996 527 2004 633
rect 2036 547 2044 653
rect 2076 607 2084 653
rect 2236 627 2244 733
rect 2336 707 2344 733
rect 1916 396 1933 407
rect 1920 393 1933 396
rect 2056 367 2064 493
rect 2156 447 2164 533
rect 2156 407 2164 433
rect 2196 427 2204 493
rect 2236 407 2244 613
rect 2296 547 2304 653
rect 2133 344 2147 353
rect 2133 340 2173 344
rect 2136 336 2173 340
rect 1853 304 1867 313
rect 1853 300 1933 304
rect 1856 296 1933 300
rect 1696 236 1773 244
rect 1616 136 1633 147
rect 1620 133 1633 136
rect 1696 107 1704 236
rect 1767 184 1780 187
rect 1767 173 1784 184
rect 1776 127 1784 173
rect 1896 127 1904 253
rect 1996 207 2004 293
rect 1996 196 2013 207
rect 2000 193 2013 196
rect 2067 196 2093 204
rect 2176 147 2184 293
rect 2216 287 2224 333
rect 2236 307 2244 393
rect 2296 307 2304 433
rect 2336 327 2344 353
rect 2216 207 2224 233
rect 2256 207 2264 233
rect 2296 147 2304 293
rect 2376 267 2384 393
rect 2176 133 2193 147
rect 2287 136 2304 147
rect 2287 133 2300 136
rect 1996 107 2004 133
rect 1536 96 1633 104
rect 2036 27 2044 113
rect 2076 67 2084 133
rect 2176 67 2184 133
rect 2236 47 2244 113
rect 2276 107 2284 133
rect 2376 127 2384 253
rect 2416 244 2424 833
rect 2476 707 2484 812
rect 2536 607 2544 933
rect 2576 767 2584 1296
rect 2656 1187 2664 1313
rect 2656 1127 2664 1173
rect 2636 887 2644 953
rect 2627 876 2644 887
rect 2627 873 2640 876
rect 2576 607 2584 693
rect 2616 647 2624 793
rect 2656 767 2664 813
rect 2676 747 2684 993
rect 2696 827 2704 913
rect 2716 867 2724 1053
rect 2736 1007 2744 1253
rect 2816 1184 2824 1533
rect 2856 1267 2864 1593
rect 2876 1547 2884 1693
rect 2896 1507 2904 1813
rect 2996 1807 3004 1973
rect 3076 1927 3084 2333
rect 3116 2107 3124 2613
rect 3176 2507 3184 2573
rect 3136 2424 3144 2493
rect 3167 2444 3180 2447
rect 3167 2433 3184 2444
rect 3136 2416 3164 2424
rect 3136 2267 3144 2333
rect 3156 2087 3164 2416
rect 3176 2407 3184 2433
rect 3216 2367 3224 2433
rect 3176 2207 3184 2353
rect 3236 2324 3244 2393
rect 3256 2348 3264 2473
rect 3316 2367 3324 2473
rect 3236 2316 3253 2324
rect 3256 2267 3264 2312
rect 2936 1767 2944 1793
rect 3016 1627 3024 1873
rect 3076 1767 3084 1913
rect 3120 1904 3133 1907
rect 3116 1900 3133 1904
rect 3113 1893 3133 1900
rect 3113 1887 3127 1893
rect 3216 1847 3224 2153
rect 3196 1747 3204 1773
rect 3216 1627 3224 1673
rect 3236 1607 3244 2193
rect 3256 2167 3264 2253
rect 3313 2204 3327 2213
rect 3287 2200 3327 2204
rect 3287 2196 3324 2200
rect 3256 1967 3264 2113
rect 3356 2067 3364 2333
rect 3316 1967 3324 2053
rect 2876 1467 2884 1493
rect 2996 1467 3004 1493
rect 3036 1467 3044 1533
rect 2933 1384 2947 1393
rect 2907 1380 2947 1384
rect 2907 1376 2944 1380
rect 2896 1327 2904 1373
rect 3016 1287 3024 1393
rect 2896 1227 2904 1273
rect 2816 1176 2844 1184
rect 2756 987 2764 1153
rect 2796 1067 2804 1153
rect 2756 867 2764 973
rect 2836 967 2844 1176
rect 2776 927 2784 953
rect 2796 767 2804 953
rect 2876 867 2884 1153
rect 2836 827 2844 853
rect 2876 827 2884 853
rect 2636 707 2644 733
rect 2736 727 2744 753
rect 2773 704 2787 713
rect 2840 704 2853 707
rect 2707 700 2787 704
rect 2707 696 2784 700
rect 2836 693 2853 704
rect 2836 667 2844 693
rect 2476 367 2484 533
rect 2476 327 2484 353
rect 2536 287 2544 553
rect 2576 467 2584 553
rect 2616 467 2624 593
rect 2616 427 2624 453
rect 2776 427 2784 453
rect 2640 424 2653 427
rect 2636 413 2653 424
rect 2636 404 2644 413
rect 2587 396 2644 404
rect 2396 236 2424 244
rect 2396 144 2404 236
rect 2396 136 2424 144
rect 2416 87 2424 136
rect 2456 127 2464 233
rect 2516 187 2524 253
rect 2576 187 2584 393
rect 2767 356 2793 364
rect 2636 327 2644 353
rect 2676 267 2684 333
rect 2716 327 2724 353
rect 2707 316 2724 327
rect 2707 313 2720 316
rect 2756 287 2764 313
rect 2593 204 2607 213
rect 2636 204 2644 253
rect 2593 200 2624 204
rect 2596 196 2627 200
rect 2636 196 2673 204
rect 2613 187 2627 196
rect 2476 124 2484 173
rect 2476 116 2513 124
rect 2556 87 2564 113
rect 2716 -16 2724 273
rect 2736 147 2744 193
rect 2796 147 2804 313
rect 2816 87 2824 393
rect 2856 307 2864 593
rect 2896 407 2904 573
rect 2876 327 2884 393
rect 2916 247 2924 1253
rect 3056 1227 3064 1273
rect 3036 1127 3044 1173
rect 2936 587 2944 1013
rect 2976 947 2984 973
rect 2996 847 3004 873
rect 3016 827 3024 933
rect 2976 667 2984 793
rect 3016 707 3024 733
rect 3076 587 3084 1593
rect 3096 1267 3104 1493
rect 3176 1447 3184 1553
rect 3116 1327 3124 1433
rect 3096 767 3104 1213
rect 3156 1047 3164 1293
rect 3176 1187 3184 1313
rect 3156 947 3164 1033
rect 3176 1027 3184 1173
rect 3216 1087 3224 1573
rect 3256 1127 3264 1573
rect 3276 1287 3284 1833
rect 3356 1747 3364 1833
rect 3376 1807 3384 2353
rect 3396 2127 3404 2673
rect 3456 2444 3464 2513
rect 3447 2440 3484 2444
rect 3447 2436 3487 2440
rect 3473 2427 3487 2436
rect 3516 2367 3524 2773
rect 3756 2744 3764 2913
rect 3736 2740 3764 2744
rect 3733 2736 3764 2740
rect 3733 2727 3747 2736
rect 3776 2727 3784 2853
rect 3936 2844 3944 3053
rect 3956 2967 3964 3093
rect 3987 3024 4000 3027
rect 3987 3013 4004 3024
rect 4027 3016 4053 3024
rect 3996 3004 4004 3013
rect 3996 2996 4044 3004
rect 3936 2836 3964 2844
rect 3856 2776 3913 2784
rect 3596 2647 3604 2713
rect 3636 2687 3644 2713
rect 3653 2504 3667 2513
rect 3736 2507 3744 2673
rect 3796 2647 3804 2773
rect 3856 2647 3864 2776
rect 3936 2764 3944 2793
rect 3916 2756 3944 2764
rect 3916 2744 3924 2756
rect 3896 2740 3924 2744
rect 3893 2736 3924 2740
rect 3893 2727 3907 2736
rect 3956 2727 3964 2836
rect 3996 2807 4004 2933
rect 4036 2907 4044 2996
rect 4156 2967 4164 3073
rect 4116 2927 4124 2953
rect 4236 2907 4244 3113
rect 4036 2787 4044 2853
rect 4196 2787 4204 2873
rect 4256 2827 4264 3296
rect 4313 3304 4327 3313
rect 4396 3307 4404 3353
rect 4287 3300 4327 3304
rect 4287 3296 4324 3300
rect 4476 3264 4484 3473
rect 4536 3447 4544 3473
rect 4560 3304 4573 3307
rect 4456 3260 4484 3264
rect 4453 3256 4484 3260
rect 4556 3293 4573 3304
rect 4686 3293 4687 3300
rect 4276 3128 4284 3253
rect 4453 3247 4467 3256
rect 4276 3027 4284 3092
rect 4296 2907 4304 2953
rect 4316 2887 4324 3013
rect 4356 2907 4364 3133
rect 4376 3027 4384 3193
rect 4496 3167 4504 3233
rect 4556 3207 4564 3293
rect 4673 3284 4687 3293
rect 4673 3280 4704 3284
rect 4676 3276 4704 3280
rect 4596 3187 4604 3233
rect 4636 3207 4644 3233
rect 4636 3167 4644 3193
rect 4696 3107 4704 3276
rect 4756 3247 4764 3453
rect 4796 3427 4804 3533
rect 4836 3367 4844 3413
rect 4813 3307 4827 3313
rect 4807 3300 4827 3307
rect 4807 3296 4824 3300
rect 4807 3293 4820 3296
rect 4836 3247 4844 3353
rect 4876 3327 4884 3533
rect 4940 3524 4953 3527
rect 4936 3513 4953 3524
rect 4936 3447 4944 3513
rect 4976 3467 4984 3552
rect 5036 3527 5044 3673
rect 4996 3387 5004 3513
rect 4936 3327 4944 3373
rect 5056 3347 5064 3613
rect 5076 3387 5084 3753
rect 5096 3427 5104 3733
rect 5156 3647 5164 3813
rect 5196 3627 5204 3813
rect 5236 3707 5244 3913
rect 5256 3887 5264 3933
rect 5353 3827 5367 3833
rect 5347 3820 5367 3827
rect 5347 3816 5364 3820
rect 5347 3813 5360 3816
rect 5296 3776 5344 3784
rect 5156 3547 5164 3593
rect 5196 3547 5204 3573
rect 5176 3407 5184 3473
rect 4867 3316 4884 3327
rect 4867 3313 4880 3316
rect 4756 3236 4773 3247
rect 4760 3233 4773 3236
rect 4827 3236 4844 3247
rect 4827 3233 4840 3236
rect 4776 3207 4784 3233
rect 4436 3027 4444 3073
rect 4376 3013 4393 3027
rect 4376 2887 4384 3013
rect 4416 2907 4424 2953
rect 4516 2847 4524 2953
rect 4576 2907 4584 2993
rect 4256 2787 4264 2813
rect 4396 2787 4404 2813
rect 4556 2787 4564 2873
rect 4247 2776 4264 2787
rect 4247 2773 4260 2776
rect 3947 2716 3964 2727
rect 3947 2713 3960 2716
rect 3653 2500 3693 2504
rect 3656 2496 3693 2500
rect 3820 2504 3833 2507
rect 3816 2493 3833 2504
rect 3860 2504 3873 2507
rect 3856 2493 3873 2504
rect 3816 2447 3824 2493
rect 3856 2484 3864 2493
rect 3836 2476 3864 2484
rect 3576 2347 3584 2413
rect 3416 2287 3424 2313
rect 3456 2264 3464 2273
rect 3456 2256 3493 2264
rect 3396 1987 3404 2113
rect 3456 1987 3464 2256
rect 3816 2227 3824 2393
rect 3836 2367 3844 2476
rect 3896 2447 3904 2673
rect 3976 2647 3984 2713
rect 4156 2667 4164 2773
rect 4227 2716 4253 2724
rect 4296 2567 4304 2713
rect 4336 2547 4344 2773
rect 4233 2504 4247 2513
rect 4356 2507 4364 2553
rect 4396 2507 4404 2533
rect 4496 2527 4504 2713
rect 4576 2567 4584 2893
rect 4596 2647 4604 2953
rect 3993 2484 4007 2493
rect 4216 2500 4247 2504
rect 4216 2496 4244 2500
rect 3993 2480 4024 2484
rect 3996 2476 4024 2480
rect 3856 2407 3864 2433
rect 3976 2347 3984 2433
rect 4016 2367 4024 2476
rect 4216 2484 4224 2496
rect 4187 2476 4224 2484
rect 3916 2267 3924 2333
rect 3976 2287 3984 2333
rect 4056 2327 4064 2433
rect 4056 2287 4064 2313
rect 3616 2187 3624 2213
rect 3673 2204 3687 2213
rect 3673 2200 3704 2204
rect 3676 2196 3704 2200
rect 3487 2176 3553 2184
rect 3396 1976 3413 1987
rect 3400 1973 3413 1976
rect 3313 1724 3327 1733
rect 3313 1720 3393 1724
rect 3316 1716 3393 1720
rect 3307 1676 3333 1684
rect 3376 1647 3384 1673
rect 3296 1547 3304 1633
rect 3336 1404 3344 1473
rect 3376 1447 3384 1553
rect 3416 1527 3424 1733
rect 3436 1647 3444 1893
rect 3496 1867 3504 2093
rect 3696 2067 3704 2196
rect 3736 2107 3744 2213
rect 4216 2207 4224 2313
rect 3456 1747 3464 1853
rect 3476 1807 3484 1833
rect 3516 1787 3524 1913
rect 3456 1736 3473 1747
rect 3460 1733 3473 1736
rect 3576 1707 3584 2053
rect 3696 2007 3704 2053
rect 3696 1967 3704 1993
rect 3596 1827 3604 1953
rect 3636 1707 3644 1813
rect 3767 1744 3780 1747
rect 3767 1733 3784 1744
rect 3536 1667 3544 1693
rect 3456 1464 3464 1613
rect 3456 1456 3484 1464
rect 3307 1400 3344 1404
rect 3307 1396 3347 1400
rect 3333 1387 3347 1396
rect 3420 1384 3433 1387
rect 3416 1373 3433 1384
rect 3416 1287 3424 1373
rect 3396 1167 3404 1193
rect 3476 1167 3484 1456
rect 3396 1156 3413 1167
rect 3400 1153 3413 1156
rect 3467 1156 3484 1167
rect 3467 1153 3480 1156
rect 3196 947 3204 973
rect 3216 924 3224 1073
rect 3296 1047 3304 1153
rect 3376 1087 3384 1153
rect 3476 1067 3484 1093
rect 3196 916 3224 924
rect 3136 707 3144 873
rect 3196 864 3204 916
rect 3227 884 3240 887
rect 3227 873 3244 884
rect 3196 856 3224 864
rect 3196 707 3204 753
rect 3216 724 3224 856
rect 3236 747 3244 873
rect 3256 787 3264 1013
rect 3296 727 3304 853
rect 3216 716 3244 724
rect 3113 644 3127 653
rect 3216 647 3224 693
rect 3113 640 3153 644
rect 3116 636 3153 640
rect 3207 636 3224 647
rect 3207 633 3220 636
rect 2956 407 2964 573
rect 3076 407 3084 573
rect 3156 467 3164 573
rect 3196 407 3204 513
rect 3236 427 3244 716
rect 3316 647 3324 813
rect 3336 747 3344 853
rect 3356 827 3364 1033
rect 3396 927 3404 973
rect 3436 947 3444 993
rect 3476 947 3484 993
rect 3496 924 3504 1533
rect 3536 1507 3544 1653
rect 3776 1647 3784 1733
rect 3836 1627 3844 1893
rect 3856 1747 3864 2073
rect 3956 1907 3964 1953
rect 3896 1767 3904 1813
rect 4036 1807 4044 2193
rect 4236 2107 4244 2473
rect 4436 2447 4444 2473
rect 4427 2436 4444 2447
rect 4427 2433 4440 2436
rect 4256 2287 4264 2353
rect 4336 2324 4344 2433
rect 4496 2427 4504 2513
rect 4576 2427 4584 2493
rect 4496 2416 4513 2427
rect 4500 2413 4513 2416
rect 4567 2416 4584 2427
rect 4567 2413 4580 2416
rect 4636 2387 4644 3073
rect 4696 2967 4704 3093
rect 4856 3087 4864 3253
rect 4896 3227 4904 3313
rect 5096 3307 5104 3333
rect 4976 3227 4984 3293
rect 5136 3247 5144 3333
rect 5216 3247 5224 3413
rect 5127 3236 5144 3247
rect 5127 3233 5140 3236
rect 4896 3187 4904 3213
rect 5076 3207 5084 3233
rect 5216 3147 5224 3233
rect 4896 3027 4904 3053
rect 4976 3027 4984 3053
rect 5016 3027 5024 3073
rect 5193 3027 5207 3033
rect 5187 3020 5207 3027
rect 5187 3016 5204 3020
rect 5187 3013 5200 3016
rect 4656 2807 4664 2833
rect 4696 2807 4704 2833
rect 4736 2807 4744 3013
rect 4776 2847 4784 2953
rect 4856 2867 4864 3013
rect 4876 2907 4884 2953
rect 5016 2907 5024 3013
rect 4776 2787 4784 2833
rect 5116 2807 5124 2953
rect 5136 2887 5144 3013
rect 5216 3007 5224 3133
rect 5236 2964 5244 3633
rect 5296 3584 5304 3776
rect 5336 3767 5344 3776
rect 5336 3756 5353 3767
rect 5340 3753 5353 3756
rect 5316 3687 5324 3753
rect 5396 3684 5404 3993
rect 5496 3967 5504 3993
rect 5456 3827 5464 3873
rect 5476 3767 5484 3893
rect 5376 3676 5404 3684
rect 5376 3627 5384 3676
rect 5436 3647 5444 3753
rect 5476 3687 5484 3753
rect 5396 3587 5404 3633
rect 5296 3576 5313 3584
rect 5316 3487 5324 3573
rect 5356 3547 5364 3573
rect 5396 3547 5404 3573
rect 5436 3547 5444 3573
rect 5416 3447 5424 3473
rect 5256 3247 5264 3373
rect 5376 3307 5384 3413
rect 5416 3407 5424 3433
rect 5316 3267 5324 3293
rect 5316 3256 5333 3267
rect 5320 3253 5333 3256
rect 5256 3107 5264 3233
rect 5336 3007 5344 3253
rect 5416 3207 5424 3393
rect 5496 3367 5504 3913
rect 5516 3447 5524 3933
rect 5536 3587 5544 4076
rect 5576 4067 5584 4153
rect 5596 4147 5604 4233
rect 5567 4056 5584 4067
rect 5567 4053 5580 4056
rect 5616 4044 5624 4173
rect 5636 4067 5644 4193
rect 5656 4167 5664 4273
rect 5676 4167 5684 4456
rect 5656 4127 5664 4153
rect 5696 4144 5704 4493
rect 5716 4187 5724 4433
rect 5736 4344 5744 4473
rect 5756 4407 5764 4473
rect 5776 4407 5784 5033
rect 5796 4867 5804 5076
rect 5847 4804 5860 4807
rect 5847 4793 5864 4804
rect 5796 4767 5804 4793
rect 5856 4687 5864 4793
rect 5816 4527 5824 4653
rect 5876 4647 5884 4973
rect 5916 4907 5924 5113
rect 5936 4947 5944 5233
rect 5956 4927 5964 5273
rect 5976 5088 5984 5173
rect 6036 5147 6044 5333
rect 6076 5127 6084 5493
rect 5976 4944 5984 5052
rect 5996 4987 6004 5013
rect 6036 4987 6044 5013
rect 5976 4940 6004 4944
rect 5976 4936 6007 4940
rect 5993 4927 6007 4936
rect 5933 4867 5947 4873
rect 5933 4860 5953 4867
rect 5936 4856 5953 4860
rect 5940 4853 5953 4856
rect 5916 4667 5924 4853
rect 5996 4824 6004 4853
rect 5956 4816 6004 4824
rect 5936 4767 5944 4793
rect 5956 4664 5964 4816
rect 5976 4687 5984 4793
rect 5936 4656 5964 4664
rect 5896 4587 5904 4613
rect 5847 4584 5860 4587
rect 5847 4573 5864 4584
rect 5887 4584 5904 4587
rect 5887 4576 5924 4584
rect 5887 4573 5900 4576
rect 5856 4564 5864 4573
rect 5856 4560 5904 4564
rect 5856 4556 5907 4560
rect 5893 4547 5907 4556
rect 5856 4467 5864 4493
rect 5833 4347 5847 4353
rect 5736 4336 5784 4344
rect 5776 4304 5784 4336
rect 5827 4340 5847 4347
rect 5827 4336 5844 4340
rect 5827 4333 5840 4336
rect 5776 4296 5824 4304
rect 5816 4287 5824 4296
rect 5816 4276 5833 4287
rect 5820 4273 5833 4276
rect 5796 4247 5804 4273
rect 5876 4247 5884 4393
rect 5916 4387 5924 4576
rect 5936 4524 5944 4656
rect 6016 4547 6024 4813
rect 6036 4627 6044 4933
rect 6056 4787 6064 4813
rect 6056 4687 6064 4713
rect 6076 4667 6084 5073
rect 5936 4516 5973 4524
rect 5936 4347 5944 4516
rect 5916 4247 5924 4273
rect 5696 4136 5724 4144
rect 5696 4067 5704 4113
rect 5636 4056 5653 4067
rect 5640 4053 5653 4056
rect 5616 4036 5644 4044
rect 5576 3607 5584 3993
rect 5636 3927 5644 4036
rect 5636 3707 5644 3813
rect 5596 3487 5604 3573
rect 5556 3347 5564 3473
rect 5556 3307 5564 3333
rect 5396 3107 5404 3133
rect 5436 3027 5444 3113
rect 5456 3027 5464 3093
rect 5476 3087 5484 3293
rect 5496 3107 5504 3253
rect 5536 3187 5544 3233
rect 5576 3207 5584 3233
rect 5516 3027 5524 3113
rect 5456 3016 5473 3027
rect 5460 3013 5473 3016
rect 5407 3004 5420 3007
rect 5407 2993 5424 3004
rect 5207 2956 5244 2964
rect 5256 2967 5264 2993
rect 5256 2956 5273 2967
rect 5260 2953 5273 2956
rect 5416 2964 5424 2993
rect 5416 2956 5453 2964
rect 5313 2944 5327 2953
rect 5296 2940 5327 2944
rect 5296 2936 5324 2940
rect 5060 2804 5073 2807
rect 5056 2793 5073 2804
rect 4656 2507 4664 2653
rect 4696 2507 4704 2673
rect 4736 2547 4744 2733
rect 4780 2724 4793 2727
rect 4776 2720 4793 2724
rect 4773 2713 4793 2720
rect 4847 2724 4860 2727
rect 4847 2713 4864 2724
rect 4773 2707 4787 2713
rect 4856 2687 4864 2713
rect 4816 2507 4824 2533
rect 4836 2447 4844 2653
rect 4856 2507 4864 2633
rect 4896 2627 4904 2673
rect 4976 2667 4984 2773
rect 5056 2727 5064 2793
rect 5156 2747 5164 2853
rect 5216 2807 5224 2833
rect 5136 2548 5144 2733
rect 5256 2687 5264 2793
rect 5296 2667 5304 2936
rect 5556 2927 5564 2953
rect 5316 2804 5324 2873
rect 5336 2824 5344 2893
rect 5336 2816 5364 2824
rect 5316 2800 5344 2804
rect 5316 2796 5347 2800
rect 5333 2787 5347 2796
rect 5356 2727 5364 2816
rect 5396 2727 5404 2913
rect 5547 2804 5560 2807
rect 5547 2793 5564 2804
rect 5493 2784 5507 2793
rect 5493 2780 5524 2784
rect 5496 2776 5524 2780
rect 5296 2547 5304 2653
rect 5067 2516 5133 2524
rect 4996 2487 5004 2513
rect 5200 2484 5213 2487
rect 5196 2473 5213 2484
rect 4676 2407 4684 2433
rect 4327 2316 4344 2324
rect 4316 2287 4324 2313
rect 4436 2267 4444 2373
rect 4576 2307 4584 2333
rect 4056 1847 4064 1913
rect 4076 1824 4084 1973
rect 4116 1827 4124 1973
rect 4176 1967 4184 2093
rect 4196 1956 4233 1964
rect 4196 1944 4204 1956
rect 4156 1940 4204 1944
rect 4153 1936 4204 1940
rect 4153 1927 4167 1936
rect 4056 1816 4084 1824
rect 3936 1687 3944 1733
rect 4056 1687 4064 1816
rect 4276 1807 4284 2213
rect 4516 2207 4524 2293
rect 4573 2287 4587 2293
rect 4573 2280 4593 2287
rect 4576 2276 4593 2280
rect 4580 2273 4593 2276
rect 4620 2284 4633 2287
rect 4616 2273 4633 2284
rect 4616 2264 4624 2273
rect 4567 2256 4624 2264
rect 4416 2167 4424 2193
rect 4156 1767 4164 1793
rect 4196 1767 4204 1793
rect 4316 1707 4324 2073
rect 4376 1927 4384 1973
rect 4456 1964 4464 2193
rect 4576 2144 4584 2213
rect 4576 2136 4604 2144
rect 4456 1956 4484 1964
rect 4367 1913 4384 1927
rect 4376 1847 4384 1913
rect 4436 1827 4444 1913
rect 4476 1807 4484 1956
rect 3927 1676 3944 1687
rect 3927 1673 3940 1676
rect 3836 1587 3844 1613
rect 3876 1607 3884 1673
rect 4056 1607 4064 1673
rect 3513 1464 3527 1473
rect 3596 1467 3604 1493
rect 3513 1460 3553 1464
rect 3516 1456 3553 1460
rect 3596 1347 3604 1453
rect 3596 1307 3604 1333
rect 3656 1327 3664 1513
rect 3736 1467 3744 1553
rect 4096 1467 4104 1553
rect 3680 1464 3693 1467
rect 3676 1453 3693 1464
rect 3676 1407 3684 1453
rect 3696 1436 3793 1444
rect 3696 1307 3704 1436
rect 3716 1367 3724 1393
rect 3756 1347 3764 1393
rect 3856 1384 3864 1433
rect 3816 1376 3864 1384
rect 3816 1364 3824 1376
rect 3787 1356 3824 1364
rect 3736 1336 3753 1344
rect 3516 1087 3524 1213
rect 3696 1187 3704 1293
rect 3636 1067 3644 1173
rect 3476 916 3504 924
rect 3396 667 3404 833
rect 3456 667 3464 773
rect 3300 644 3313 647
rect 3296 633 3313 644
rect 3076 396 3093 407
rect 3080 393 3093 396
rect 3096 267 3104 353
rect 3156 347 3164 393
rect 3256 364 3264 593
rect 3296 567 3304 633
rect 3367 616 3453 624
rect 3216 360 3264 364
rect 3213 356 3264 360
rect 3213 347 3227 356
rect 3156 336 3173 347
rect 3160 333 3173 336
rect 3056 207 3064 253
rect 3116 207 3124 273
rect 3107 196 3124 207
rect 3107 193 3120 196
rect 3136 184 3144 293
rect 3256 207 3264 313
rect 3336 287 3344 553
rect 3476 427 3484 916
rect 3516 887 3524 993
rect 3596 947 3604 973
rect 3636 947 3644 993
rect 3496 827 3504 873
rect 3696 847 3704 1173
rect 3736 947 3744 1336
rect 3976 1327 3984 1393
rect 3836 1227 3844 1273
rect 3776 947 3784 1013
rect 3816 887 3824 1133
rect 3876 1087 3884 1313
rect 3807 876 3824 887
rect 3807 873 3820 876
rect 3696 767 3704 833
rect 3676 707 3684 733
rect 3516 696 3573 704
rect 3516 627 3524 696
rect 3636 627 3644 693
rect 3756 664 3764 753
rect 3776 707 3784 773
rect 3876 707 3884 1073
rect 3896 947 3904 973
rect 3916 807 3924 1213
rect 3956 1127 3964 1153
rect 3976 1107 3984 1213
rect 3936 947 3944 1093
rect 3996 947 4004 1153
rect 4016 1127 4024 1353
rect 4076 1347 4084 1393
rect 4136 1287 4144 1693
rect 4316 1627 4324 1693
rect 4216 1467 4224 1493
rect 4356 1467 4364 1793
rect 4416 1527 4424 1573
rect 4456 1547 4464 1773
rect 4496 1607 4504 1973
rect 4556 1767 4564 1913
rect 4496 1544 4504 1593
rect 4488 1536 4504 1544
rect 4433 1467 4447 1473
rect 4267 1464 4280 1467
rect 4356 1464 4373 1467
rect 4267 1453 4284 1464
rect 4176 1407 4184 1453
rect 4276 1407 4284 1453
rect 4336 1456 4373 1464
rect 4176 1396 4193 1407
rect 4180 1393 4193 1396
rect 4136 1247 4144 1273
rect 4093 1224 4107 1233
rect 4256 1227 4264 1253
rect 4076 1220 4107 1224
rect 4076 1216 4104 1220
rect 4076 1167 4084 1216
rect 4296 1187 4304 1273
rect 4076 1127 4084 1153
rect 4016 1007 4024 1113
rect 4056 887 4064 1013
rect 4136 947 4144 1173
rect 4336 1107 4344 1456
rect 4360 1453 4373 1456
rect 4427 1460 4447 1467
rect 4427 1456 4444 1460
rect 4427 1453 4440 1456
rect 4436 1367 4444 1393
rect 4396 1227 4404 1273
rect 4456 1187 4464 1253
rect 4376 1127 4384 1153
rect 4416 1107 4424 1153
rect 4136 936 4153 947
rect 4140 933 4153 936
rect 4207 944 4220 947
rect 4207 933 4224 944
rect 4216 887 4224 933
rect 4016 724 4024 873
rect 4056 767 4064 873
rect 4136 847 4144 873
rect 4276 847 4284 1033
rect 4316 947 4324 1013
rect 4376 887 4384 933
rect 4376 873 4393 887
rect 4376 787 4384 873
rect 4476 767 4484 1533
rect 4536 1487 4544 1733
rect 4596 1687 4604 2136
rect 4616 2007 4624 2193
rect 4656 2147 4664 2213
rect 4736 2207 4744 2433
rect 4776 2267 4784 2373
rect 4916 2367 4924 2433
rect 4736 2196 4753 2207
rect 4740 2193 4753 2196
rect 4756 2167 4764 2193
rect 4796 2147 4804 2213
rect 4676 1967 4684 1993
rect 4736 1967 4744 2093
rect 4816 1927 4824 2053
rect 4836 1987 4844 2113
rect 4876 2107 4884 2213
rect 4936 2107 4944 2473
rect 5076 2267 5084 2293
rect 5116 2267 5124 2433
rect 5067 2256 5084 2267
rect 5067 2253 5080 2256
rect 4996 2127 5004 2213
rect 5196 2207 5204 2473
rect 5256 2427 5264 2533
rect 5307 2484 5320 2487
rect 5307 2473 5324 2484
rect 5256 2416 5273 2427
rect 5260 2413 5273 2416
rect 5236 2347 5244 2413
rect 5316 2407 5324 2473
rect 5256 2280 5293 2284
rect 5253 2276 5293 2280
rect 5253 2267 5267 2276
rect 5336 2244 5344 2273
rect 5287 2236 5344 2244
rect 5356 2227 5364 2593
rect 5396 2507 5404 2633
rect 5436 2627 5444 2733
rect 5516 2687 5524 2776
rect 5556 2747 5564 2793
rect 5576 2607 5584 3153
rect 5616 2664 5624 3433
rect 5636 3087 5644 3593
rect 5676 3584 5684 3953
rect 5716 3887 5724 4136
rect 5736 3967 5744 4153
rect 5836 4067 5844 4093
rect 5876 4067 5884 4173
rect 5936 4084 5944 4333
rect 5976 4287 5984 4373
rect 5967 4276 5984 4287
rect 5967 4273 5980 4276
rect 5916 4076 5944 4084
rect 5896 4027 5904 4053
rect 5867 3996 5904 4004
rect 5796 3827 5804 3993
rect 5896 3984 5904 3996
rect 5916 3987 5924 4076
rect 5940 4064 5953 4067
rect 5936 4053 5953 4064
rect 5936 4027 5944 4053
rect 5976 4044 5984 4153
rect 5996 4147 6004 4473
rect 6016 4167 6024 4333
rect 6036 4148 6044 4453
rect 5996 4067 6004 4093
rect 5976 4036 6004 4044
rect 5960 4004 5973 4007
rect 5956 4000 5973 4004
rect 5953 3993 5973 4000
rect 5953 3987 5967 3993
rect 5896 3976 5913 3984
rect 5876 3827 5884 3953
rect 5736 3727 5744 3753
rect 5776 3727 5784 3753
rect 5656 3576 5684 3584
rect 5656 3447 5664 3576
rect 5756 3547 5764 3693
rect 5796 3587 5804 3813
rect 5836 3547 5844 3693
rect 5876 3608 5884 3813
rect 5916 3667 5924 3813
rect 5876 3547 5884 3572
rect 5687 3536 5713 3544
rect 5747 3476 5773 3484
rect 5916 3484 5924 3593
rect 5936 3547 5944 3933
rect 5996 3907 6004 4036
rect 5956 3587 5964 3853
rect 5867 3476 5924 3484
rect 5696 3347 5704 3453
rect 5893 3444 5907 3453
rect 5893 3440 5924 3444
rect 5896 3436 5924 3440
rect 5856 3307 5864 3333
rect 5656 3264 5664 3293
rect 5656 3260 5684 3264
rect 5656 3256 5687 3260
rect 5673 3247 5687 3256
rect 5716 3207 5724 3233
rect 5656 3027 5664 3093
rect 5656 3016 5673 3027
rect 5660 3013 5673 3016
rect 5636 2807 5644 2833
rect 5696 2807 5704 3053
rect 5736 3027 5744 3073
rect 5776 3067 5784 3293
rect 5876 3247 5884 3413
rect 5916 3404 5924 3436
rect 5896 3396 5924 3404
rect 5896 3284 5904 3396
rect 5896 3276 5924 3284
rect 5836 3207 5844 3233
rect 5916 3104 5924 3276
rect 5896 3096 5924 3104
rect 5727 3016 5744 3027
rect 5727 3013 5740 3016
rect 5787 3016 5813 3024
rect 5836 2967 5844 3093
rect 5687 2796 5704 2807
rect 5687 2793 5700 2796
rect 5636 2707 5644 2793
rect 5616 2656 5644 2664
rect 5636 2587 5644 2656
rect 5436 2507 5444 2533
rect 5736 2507 5744 2853
rect 5896 2847 5904 3096
rect 5936 3084 5944 3533
rect 5996 3487 6004 3573
rect 5956 3247 5964 3413
rect 5996 3367 6004 3473
rect 6036 3388 6044 4112
rect 5976 3247 5984 3333
rect 5976 3236 5993 3247
rect 5980 3233 5993 3236
rect 5916 3076 5944 3084
rect 5836 2787 5844 2833
rect 5827 2776 5844 2787
rect 5827 2773 5840 2776
rect 5856 2707 5864 2733
rect 5896 2687 5904 2733
rect 5736 2493 5753 2507
rect 5476 2407 5484 2473
rect 5536 2407 5544 2433
rect 5596 2407 5604 2433
rect 5616 2407 5624 2493
rect 5667 2436 5693 2444
rect 5716 2407 5724 2493
rect 5507 2384 5520 2387
rect 5507 2373 5524 2384
rect 5416 2267 5424 2293
rect 5436 2167 5444 2193
rect 4876 1847 4884 1973
rect 4936 1967 4944 2093
rect 4676 1747 4684 1773
rect 4776 1684 4784 1733
rect 4956 1687 4964 1833
rect 4996 1787 5004 1953
rect 5116 1847 5124 1913
rect 5196 1887 5204 2113
rect 5236 1987 5244 2053
rect 5276 1987 5284 2013
rect 5256 1887 5264 1913
rect 5127 1836 5144 1844
rect 4747 1676 4784 1684
rect 4536 1387 4544 1473
rect 4596 1387 4604 1553
rect 4656 1487 4664 1673
rect 4696 1547 4704 1673
rect 4536 1376 4553 1387
rect 4540 1373 4553 1376
rect 4536 1247 4544 1333
rect 4656 1287 4664 1433
rect 4696 1387 4704 1473
rect 4576 1247 4584 1273
rect 4696 1247 4704 1273
rect 4720 1244 4733 1247
rect 4716 1233 4733 1244
rect 4716 1224 4724 1233
rect 4676 1216 4724 1224
rect 4496 1147 4504 1213
rect 4676 1187 4684 1216
rect 4516 927 4524 1033
rect 4576 927 4584 1053
rect 4696 947 4704 993
rect 4736 947 4744 1173
rect 4756 1007 4764 1633
rect 4856 1547 4864 1673
rect 4996 1627 5004 1673
rect 5036 1607 5044 1673
rect 5096 1627 5104 1733
rect 5136 1687 5144 1836
rect 5296 1827 5304 1913
rect 5356 1867 5364 2153
rect 5396 2027 5404 2153
rect 5396 1944 5404 2013
rect 5436 1967 5444 2053
rect 5476 1967 5484 2093
rect 5516 2067 5524 2373
rect 5556 2207 5564 2333
rect 5596 2207 5604 2393
rect 5716 2367 5724 2393
rect 5736 2307 5744 2493
rect 5860 2484 5873 2487
rect 5856 2473 5873 2484
rect 5756 2327 5764 2433
rect 5816 2367 5824 2473
rect 5647 2256 5673 2264
rect 5776 2107 5784 2353
rect 5816 2267 5824 2313
rect 5856 2287 5864 2473
rect 5916 2307 5924 3076
rect 5936 3007 5944 3053
rect 6016 3027 6024 3053
rect 5960 3024 5973 3027
rect 5956 3013 5973 3024
rect 5956 2927 5964 3013
rect 5936 2807 5944 2833
rect 5976 2807 5984 2893
rect 5976 2707 5984 2793
rect 5876 2207 5884 2293
rect 5907 2264 5920 2267
rect 5907 2253 5924 2264
rect 5916 2207 5924 2253
rect 5807 2196 5833 2204
rect 5876 2167 5884 2193
rect 5756 1967 5764 2073
rect 5816 1967 5824 2093
rect 5756 1956 5773 1967
rect 5760 1953 5773 1956
rect 5396 1936 5444 1944
rect 5436 1907 5444 1936
rect 5396 1867 5404 1893
rect 5296 1747 5304 1773
rect 5456 1747 5464 1773
rect 5496 1747 5504 1813
rect 5536 1787 5544 1953
rect 5656 1847 5664 1913
rect 5616 1747 5624 1833
rect 5736 1767 5744 1793
rect 5796 1767 5804 1833
rect 5876 1767 5884 2113
rect 5916 1807 5924 2193
rect 5956 2184 5964 2293
rect 5996 2267 6004 2433
rect 5936 2176 5964 2184
rect 5176 1607 5184 1673
rect 5216 1647 5224 1733
rect 5253 1724 5267 1733
rect 5236 1720 5267 1724
rect 5236 1716 5264 1720
rect 5236 1687 5244 1716
rect 5487 1676 5513 1684
rect 4776 1407 4784 1513
rect 4816 1467 4824 1533
rect 4956 1467 4964 1533
rect 5036 1527 5044 1593
rect 4867 1464 4880 1467
rect 4867 1453 4884 1464
rect 4956 1456 4973 1467
rect 4960 1453 4973 1456
rect 4876 1407 4884 1453
rect 4776 1396 4793 1407
rect 4780 1393 4793 1396
rect 4836 1347 4844 1373
rect 4816 1187 4824 1273
rect 4856 1227 4864 1253
rect 5016 1227 5024 1273
rect 5076 1267 5084 1533
rect 5096 1467 5104 1513
rect 5136 1467 5144 1493
rect 5096 1327 5104 1453
rect 5176 1407 5184 1453
rect 5176 1396 5193 1407
rect 5180 1393 5193 1396
rect 5156 1344 5164 1393
rect 5156 1336 5184 1344
rect 5136 1227 5144 1253
rect 5156 1224 5164 1313
rect 5176 1267 5184 1336
rect 5156 1216 5173 1224
rect 4816 1147 4824 1173
rect 4876 1027 4884 1153
rect 4996 1087 5004 1153
rect 5116 1127 5124 1153
rect 5156 1087 5164 1153
rect 4836 947 4844 1013
rect 4876 947 4884 973
rect 4340 764 4353 767
rect 4336 753 4353 764
rect 4116 727 4124 753
rect 4016 716 4073 724
rect 3927 696 3973 704
rect 4176 667 4184 733
rect 3756 656 3793 664
rect 3680 644 3693 647
rect 3676 640 3693 644
rect 3673 633 3693 640
rect 3747 644 3760 647
rect 3747 633 3764 644
rect 3673 627 3687 633
rect 3116 176 3144 184
rect 2696 -24 2724 -16
rect 2916 -24 2924 173
rect 3116 147 3124 176
rect 3216 164 3224 193
rect 3156 160 3224 164
rect 3153 156 3224 160
rect 3153 147 3167 156
rect 3176 136 3213 144
rect 3036 87 3044 133
rect 3176 124 3184 136
rect 3087 116 3184 124
rect 3296 76 3353 84
rect 3296 47 3304 76
rect 3376 47 3384 353
rect 3407 176 3433 184
rect 3476 127 3484 293
rect 3467 113 3484 127
rect 3336 -24 3344 33
rect 3416 27 3424 53
rect 3476 47 3484 113
rect 3496 27 3504 353
rect 3616 347 3624 553
rect 3576 227 3584 313
rect 3676 287 3684 473
rect 3716 427 3724 553
rect 3756 527 3764 633
rect 3776 407 3784 656
rect 3856 507 3864 653
rect 3896 536 4044 544
rect 3896 487 3904 536
rect 3696 267 3704 353
rect 3756 307 3764 393
rect 3836 267 3844 393
rect 3956 367 3964 493
rect 4016 487 4024 513
rect 3616 127 3624 253
rect 3736 187 3744 233
rect 3776 187 3784 213
rect 3936 187 3944 253
rect 4016 187 4024 473
rect 4036 467 4044 536
rect 4116 427 4124 573
rect 4156 507 4164 633
rect 4236 587 4244 693
rect 4296 667 4304 733
rect 4336 707 4344 753
rect 4376 707 4384 733
rect 4356 587 4364 653
rect 4396 607 4404 633
rect 4436 567 4444 633
rect 4076 287 4084 413
rect 4156 367 4164 393
rect 4147 356 4164 367
rect 4147 353 4160 356
rect 4096 287 4104 353
rect 4256 347 4264 493
rect 4436 487 4444 553
rect 4376 427 4384 453
rect 4476 447 4484 693
rect 4556 587 4564 713
rect 4433 427 4447 433
rect 4427 420 4447 427
rect 4427 416 4444 420
rect 4427 413 4440 416
rect 4516 404 4524 513
rect 4536 407 4544 553
rect 4576 527 4584 913
rect 4796 887 4804 933
rect 4796 876 4813 887
rect 4800 873 4813 876
rect 4596 767 4604 793
rect 4596 727 4604 753
rect 4636 667 4644 793
rect 4696 707 4704 753
rect 4676 587 4684 633
rect 4756 547 4764 873
rect 4776 567 4784 693
rect 4816 667 4824 773
rect 4856 747 4864 853
rect 4916 747 4924 1073
rect 4916 664 4924 693
rect 4836 656 4924 664
rect 4836 547 4844 656
rect 4856 607 4864 633
rect 4896 607 4904 633
rect 4956 607 4964 973
rect 4996 947 5004 993
rect 5176 987 5184 1213
rect 5193 947 5207 953
rect 5120 944 5133 947
rect 5116 933 5133 944
rect 5187 940 5207 947
rect 5187 936 5204 940
rect 5187 933 5200 936
rect 4996 707 5004 733
rect 5076 707 5084 933
rect 5116 887 5124 933
rect 5216 887 5224 1173
rect 5236 1067 5244 1573
rect 5276 1307 5284 1673
rect 5316 1647 5324 1673
rect 5436 1627 5444 1673
rect 5596 1647 5604 1673
rect 5356 1447 5364 1573
rect 5496 1447 5504 1633
rect 5616 1447 5624 1553
rect 5776 1547 5784 1693
rect 5736 1467 5744 1533
rect 5356 1436 5373 1447
rect 5360 1433 5373 1436
rect 5316 1327 5324 1433
rect 5436 1267 5444 1393
rect 5616 1387 5624 1433
rect 5676 1387 5684 1433
rect 5293 1224 5307 1233
rect 5293 1220 5324 1224
rect 5296 1216 5324 1220
rect 5316 1167 5324 1216
rect 5207 876 5224 887
rect 5207 873 5220 876
rect 5076 696 5093 707
rect 5080 693 5093 696
rect 5016 607 5024 653
rect 5016 567 5024 593
rect 4756 467 4764 533
rect 4796 427 4804 533
rect 5096 507 5104 693
rect 5216 667 5224 833
rect 5236 664 5244 1053
rect 5296 947 5304 973
rect 5336 827 5344 933
rect 5236 656 5273 664
rect 5276 547 5284 653
rect 5316 487 5324 693
rect 5356 647 5364 1213
rect 5476 1167 5484 1273
rect 5516 1167 5524 1293
rect 5556 1227 5564 1253
rect 5676 1227 5684 1313
rect 5776 1244 5784 1533
rect 5816 1307 5824 1693
rect 5856 1287 5864 1393
rect 5896 1327 5904 1393
rect 5776 1236 5813 1244
rect 5896 1244 5904 1273
rect 5936 1267 5944 2176
rect 5956 1507 5964 2053
rect 5976 1827 5984 2153
rect 5976 1747 5984 1813
rect 5996 1467 6004 1493
rect 6036 1467 6044 3352
rect 6016 1347 6024 1393
rect 5996 1336 6013 1344
rect 5867 1236 5904 1244
rect 5436 1087 5444 1153
rect 5396 887 5404 1073
rect 5467 944 5480 947
rect 5467 933 5484 944
rect 5407 876 5433 884
rect 5436 647 5444 833
rect 5476 827 5484 933
rect 5536 887 5544 1073
rect 5476 707 5484 813
rect 5556 647 5564 1113
rect 5576 947 5584 1153
rect 5616 947 5624 1213
rect 5576 707 5584 833
rect 5656 807 5664 933
rect 5696 887 5704 933
rect 5687 876 5704 887
rect 5687 873 5700 876
rect 5756 847 5764 873
rect 5596 647 5604 773
rect 5696 727 5704 773
rect 5796 767 5804 1173
rect 5856 887 5864 1233
rect 5996 1227 6004 1336
rect 5987 1216 6004 1227
rect 5987 1213 6000 1216
rect 5936 947 5944 1153
rect 5856 876 5873 887
rect 5860 873 5873 876
rect 5896 807 5904 933
rect 6016 924 6024 1253
rect 5996 916 6024 924
rect 5876 796 5893 804
rect 5756 727 5764 753
rect 5747 716 5764 727
rect 5747 713 5760 716
rect 5356 636 5373 647
rect 5360 633 5373 636
rect 5427 636 5444 647
rect 5427 633 5440 636
rect 4787 413 4804 427
rect 4487 396 4524 404
rect 4447 356 4504 364
rect 4216 267 4224 333
rect 3696 144 3704 173
rect 3696 136 3744 144
rect 3576 47 3584 113
rect 3716 67 3724 113
rect 3736 104 3744 136
rect 3816 124 3824 173
rect 4056 127 4064 213
rect 4216 187 4224 213
rect 4173 164 4187 173
rect 4256 164 4264 213
rect 4296 207 4304 233
rect 4396 187 4404 353
rect 4496 344 4504 356
rect 4727 356 4753 364
rect 4496 336 4533 344
rect 4607 340 4684 344
rect 4607 336 4687 340
rect 4673 327 4687 336
rect 4636 187 4644 273
rect 4796 227 4804 413
rect 4816 327 4824 393
rect 5016 367 5024 453
rect 5236 444 5244 473
rect 5407 456 5473 464
rect 5547 456 5613 464
rect 5216 440 5244 444
rect 5213 436 5244 440
rect 5213 427 5227 436
rect 4876 267 4884 333
rect 4916 307 4924 333
rect 5136 327 5144 393
rect 5156 267 5164 353
rect 4173 160 4264 164
rect 4176 156 4264 160
rect 3767 116 3824 124
rect 3836 120 3873 124
rect 3833 116 3873 120
rect 3833 107 3847 116
rect 4047 116 4064 127
rect 4047 113 4060 116
rect 3736 96 3773 104
rect 3916 67 3924 113
rect 4156 87 4164 113
rect 4196 87 4204 113
rect 3456 -24 3464 13
rect 4456 -24 4464 133
rect 4596 -24 4604 133
rect 4736 -24 4744 133
rect 4876 127 4884 213
rect 4916 127 4924 253
rect 5076 187 5084 253
rect 5176 247 5184 413
rect 5296 367 5304 453
rect 5320 424 5333 427
rect 5316 413 5333 424
rect 5593 424 5607 433
rect 5576 420 5607 424
rect 5576 416 5604 420
rect 5236 327 5244 353
rect 5316 327 5324 413
rect 5396 367 5404 413
rect 5576 404 5584 416
rect 5547 396 5584 404
rect 5636 404 5644 533
rect 5607 396 5644 404
rect 5396 353 5413 367
rect 5136 187 5144 233
rect 4776 -24 4784 93
rect 4956 87 4964 173
rect 4996 127 5004 153
rect 5156 127 5164 213
rect 5196 127 5204 313
rect 5316 267 5324 313
rect 5396 307 5404 353
rect 5553 224 5567 233
rect 5536 220 5567 224
rect 5596 224 5604 393
rect 5696 367 5704 473
rect 5716 427 5724 633
rect 5776 487 5784 693
rect 5756 427 5764 453
rect 5796 327 5804 753
rect 5876 647 5884 796
rect 5907 704 5920 707
rect 5907 693 5924 704
rect 5836 567 5844 633
rect 5916 627 5924 693
rect 5936 647 5944 873
rect 5956 667 5964 833
rect 5996 727 6004 916
rect 5996 713 6013 727
rect 5976 627 5984 713
rect 5896 467 5904 553
rect 5936 427 5944 453
rect 5976 427 5984 613
rect 5876 287 5884 333
rect 5896 264 5904 413
rect 5996 384 6004 713
rect 5976 376 6004 384
rect 5976 364 5984 376
rect 5927 356 5984 364
rect 5996 327 6004 353
rect 5896 256 5913 264
rect 5627 236 5704 244
rect 5536 216 5564 220
rect 5596 216 5624 224
rect 5236 187 5244 213
rect 5387 200 5464 204
rect 5387 196 5467 200
rect 5236 176 5253 187
rect 5240 173 5253 176
rect 4996 116 5013 127
rect 5000 113 5013 116
rect 5056 87 5064 113
rect 5156 67 5164 113
rect 5316 84 5324 193
rect 5453 187 5467 196
rect 5536 184 5544 216
rect 5616 207 5624 216
rect 5507 176 5544 184
rect 5556 144 5564 193
rect 5616 164 5624 193
rect 5696 187 5704 236
rect 5916 207 5924 253
rect 5956 207 5964 273
rect 5616 156 5644 164
rect 5447 136 5564 144
rect 5636 144 5644 156
rect 5636 136 5673 144
rect 5856 140 5893 144
rect 5853 136 5893 140
rect 5247 76 5324 84
rect 5376 47 5384 133
rect 5613 124 5627 133
rect 5853 127 5867 136
rect 5613 120 5664 124
rect 5616 116 5664 120
rect 5656 107 5664 116
rect 5976 107 5984 133
rect 6036 107 6044 893
rect 6056 887 6064 4533
rect 6076 4168 6084 4613
rect 6076 3587 6084 4132
rect 6076 907 6084 3373
rect 5656 96 5673 107
rect 5660 93 5673 96
rect 5767 96 5833 104
use NOR2X1  _760_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727495070
transform 1 0 4870 0 1 270
box -6 -8 86 272
use INVX1  _761_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727493700
transform 1 0 3690 0 1 270
box -6 -8 66 272
use NOR2X1  _762_
timestamp 1727495070
transform 1 0 3170 0 1 270
box -6 -8 86 272
use OAI21X1  _763_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727498925
transform 1 0 4370 0 -1 790
box -6 -8 106 272
use INVX2  _764_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727493898
transform -1 0 2850 0 -1 1830
box -6 -8 66 272
use NOR2X1  _765_
timestamp 1727495070
transform -1 0 1990 0 1 1310
box -6 -8 86 272
use AOI22X1  _766_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487144
transform -1 0 2050 0 -1 790
box -6 -8 126 272
use OAI21X1  _767_
timestamp 1727498925
transform -1 0 4450 0 1 270
box -6 -8 106 272
use INVX1  _768_
timestamp 1727493700
transform 1 0 4010 0 -1 270
box -6 -8 66 272
use INVX1  _769_
timestamp 1727493700
transform 1 0 4750 0 1 270
box -6 -8 66 272
use NAND2X1  _770_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727494699
transform -1 0 4930 0 -1 270
box -6 -8 86 272
use OAI21X1  _771_
timestamp 1727498925
transform -1 0 5090 0 -1 270
box -6 -8 106 272
use AOI22X1  _772_
timestamp 1727487144
transform -1 0 2290 0 -1 270
box -6 -8 126 272
use OAI21X1  _773_
timestamp 1727498925
transform -1 0 4230 0 -1 270
box -6 -8 106 272
use NOR2X1  _774_
timestamp 1727495070
transform 1 0 4210 0 1 270
box -6 -8 86 272
use OAI21X1  _775_
timestamp 1727498925
transform 1 0 3670 0 -1 790
box -6 -8 106 272
use AOI22X1  _776_
timestamp 1727487144
transform 1 0 2150 0 1 270
box -6 -8 126 272
use OAI21X1  _777_
timestamp 1727498925
transform -1 0 4150 0 1 270
box -6 -8 106 272
use INVX1  _778_
timestamp 1727493700
transform 1 0 3430 0 -1 270
box -6 -8 66 272
use NAND2X1  _779_
timestamp 1727494699
transform -1 0 3630 0 -1 270
box -6 -8 86 272
use OAI21X1  _780_
timestamp 1727498925
transform -1 0 3950 0 -1 270
box -6 -8 106 272
use AOI22X1  _781_
timestamp 1727487144
transform 1 0 1990 0 -1 270
box -6 -8 126 272
use OAI21X1  _782_
timestamp 1727498925
transform -1 0 3790 0 -1 270
box -6 -8 106 272
use INVX2  _783_
timestamp 1727493898
transform -1 0 3490 0 1 4430
box -6 -8 66 272
use NAND2X1  _784_
timestamp 1727494699
transform -1 0 2650 0 -1 3910
box -6 -8 86 272
use OAI21X1  _785_
timestamp 1727498925
transform -1 0 4470 0 -1 3910
box -6 -8 106 272
use INVX2  _786_
timestamp 1727493898
transform -1 0 3250 0 1 4430
box -6 -8 66 272
use NAND2X1  _787_
timestamp 1727494699
transform -1 0 4610 0 -1 4950
box -6 -8 86 272
use OAI21X1  _788_
timestamp 1727498925
transform 1 0 4670 0 -1 4950
box -6 -8 106 272
use INVX2  _789_
timestamp 1727493898
transform -1 0 3550 0 1 4950
box -6 -8 66 272
use NAND2X1  _790_
timestamp 1727494699
transform -1 0 4170 0 1 4950
box -6 -8 86 272
use OAI21X1  _791_
timestamp 1727498925
transform -1 0 4330 0 1 4950
box -6 -8 106 272
use INVX2  _792_
timestamp 1727493898
transform -1 0 5470 0 -1 4950
box -6 -8 66 272
use NAND2X1  _793_
timestamp 1727494699
transform -1 0 4310 0 -1 4950
box -6 -8 86 272
use OAI21X1  _794_
timestamp 1727498925
transform -1 0 4470 0 -1 4950
box -6 -8 106 272
use NAND2X1  _795_
timestamp 1727494699
transform 1 0 2710 0 -1 3910
box -6 -8 86 272
use OAI21X1  _796_
timestamp 1727498925
transform -1 0 2950 0 -1 3910
box -6 -8 106 272
use NAND2X1  _797_
timestamp 1727494699
transform 1 0 1670 0 -1 3910
box -6 -8 86 272
use OAI21X1  _798_
timestamp 1727498925
transform -1 0 2490 0 -1 4430
box -6 -8 106 272
use NAND2X1  _799_
timestamp 1727494699
transform 1 0 1750 0 1 3910
box -6 -8 86 272
use OAI21X1  _800_
timestamp 1727498925
transform -1 0 3350 0 1 3910
box -6 -8 106 272
use NAND2X1  _801_
timestamp 1727494699
transform 1 0 1610 0 1 3910
box -6 -8 86 272
use OAI21X1  _802_
timestamp 1727498925
transform -1 0 3470 0 -1 4430
box -6 -8 106 272
use INVX1  _803_
timestamp 1727493700
transform -1 0 1910 0 -1 3390
box -6 -8 66 272
use NAND2X1  _804_
timestamp 1727494699
transform -1 0 2450 0 -1 2870
box -6 -8 86 272
use OAI21X1  _805_
timestamp 1727498925
transform 1 0 2170 0 1 2870
box -6 -8 106 272
use INVX1  _806_
timestamp 1727493700
transform 1 0 1470 0 -1 2350
box -6 -8 66 272
use NAND2X1  _807_
timestamp 1727494699
transform 1 0 1890 0 -1 2350
box -6 -8 86 272
use OAI21X1  _808_
timestamp 1727498925
transform 1 0 1590 0 -1 2350
box -6 -8 106 272
use INVX1  _809_
timestamp 1727493700
transform 1 0 970 0 1 2870
box -6 -8 66 272
use NAND2X1  _810_
timestamp 1727494699
transform 1 0 2510 0 -1 2870
box -6 -8 86 272
use OAI21X1  _811_
timestamp 1727498925
transform 1 0 1090 0 1 2870
box -6 -8 106 272
use INVX1  _812_
timestamp 1727493700
transform -1 0 770 0 -1 2350
box -6 -8 66 272
use NAND2X1  _813_
timestamp 1727494699
transform 1 0 1470 0 1 1830
box -6 -8 86 272
use OAI21X1  _814_
timestamp 1727498925
transform -1 0 1170 0 -1 2350
box -6 -8 106 272
use INVX1  _815_
timestamp 1727493700
transform -1 0 270 0 -1 1830
box -6 -8 66 272
use NAND2X1  _816_
timestamp 1727494699
transform -1 0 1590 0 -1 1830
box -6 -8 86 272
use OAI21X1  _817_
timestamp 1727498925
transform 1 0 570 0 -1 1830
box -6 -8 106 272
use INVX1  _818_
timestamp 1727493700
transform -1 0 930 0 -1 1830
box -6 -8 66 272
use NAND2X1  _819_
timestamp 1727494699
transform 1 0 1650 0 -1 1830
box -6 -8 86 272
use OAI21X1  _820_
timestamp 1727498925
transform 1 0 1230 0 -1 1830
box -6 -8 106 272
use INVX1  _821_
timestamp 1727493700
transform 1 0 1130 0 1 790
box -6 -8 66 272
use NAND2X1  _822_
timestamp 1727494699
transform -1 0 1750 0 -1 1310
box -6 -8 86 272
use OAI21X1  _823_
timestamp 1727498925
transform 1 0 1250 0 1 790
box -6 -8 106 272
use INVX1  _824_
timestamp 1727493700
transform 1 0 770 0 -1 1310
box -6 -8 66 272
use NAND2X1  _825_
timestamp 1727494699
transform 1 0 1050 0 1 1310
box -6 -8 86 272
use OAI21X1  _826_
timestamp 1727498925
transform 1 0 890 0 1 1310
box -6 -8 106 272
use INVX1  _827_
timestamp 1727493700
transform 1 0 3970 0 1 2350
box -6 -8 66 272
use NAND2X1  _828_
timestamp 1727494699
transform -1 0 3750 0 1 2350
box -6 -8 86 272
use OAI21X1  _829_
timestamp 1727498925
transform -1 0 3910 0 1 2350
box -6 -8 106 272
use INVX1  _830_
timestamp 1727493700
transform 1 0 4070 0 1 1310
box -6 -8 66 272
use NAND2X1  _831_
timestamp 1727494699
transform -1 0 3610 0 1 1310
box -6 -8 86 272
use OAI21X1  _832_
timestamp 1727498925
transform -1 0 3770 0 1 1310
box -6 -8 106 272
use INVX1  _833_
timestamp 1727493700
transform 1 0 3190 0 -1 1830
box -6 -8 66 272
use NAND2X1  _834_
timestamp 1727494699
transform 1 0 3410 0 1 1830
box -6 -8 86 272
use OAI21X1  _835_
timestamp 1727498925
transform 1 0 3310 0 -1 1830
box -6 -8 106 272
use INVX1  _836_
timestamp 1727493700
transform 1 0 2450 0 1 790
box -6 -8 66 272
use NAND2X1  _837_
timestamp 1727494699
transform 1 0 2310 0 1 1310
box -6 -8 86 272
use OAI21X1  _838_
timestamp 1727498925
transform -1 0 2390 0 1 790
box -6 -8 106 272
use INVX1  _839_
timestamp 1727493700
transform -1 0 5630 0 -1 1830
box -6 -8 66 272
use NAND2X1  _840_
timestamp 1727494699
transform -1 0 5050 0 -1 1830
box -6 -8 86 272
use OAI21X1  _841_
timestamp 1727498925
transform -1 0 5510 0 -1 1830
box -6 -8 106 272
use INVX1  _842_
timestamp 1727493700
transform 1 0 5410 0 -1 2350
box -6 -8 66 272
use NAND2X1  _843_
timestamp 1727494699
transform 1 0 4830 0 1 1830
box -6 -8 86 272
use OAI21X1  _844_
timestamp 1727498925
transform -1 0 5310 0 1 1830
box -6 -8 106 272
use INVX1  _845_
timestamp 1727493700
transform -1 0 5030 0 -1 1310
box -6 -8 66 272
use NAND2X1  _846_
timestamp 1727494699
transform 1 0 5090 0 1 1310
box -6 -8 86 272
use OAI21X1  _847_
timestamp 1727498925
transform -1 0 5190 0 -1 1310
box -6 -8 106 272
use INVX1  _848_
timestamp 1727493700
transform 1 0 5550 0 -1 1310
box -6 -8 66 272
use NAND2X1  _849_
timestamp 1727494699
transform -1 0 5190 0 -1 1830
box -6 -8 86 272
use OAI21X1  _850_
timestamp 1727498925
transform 1 0 5250 0 -1 1830
box -6 -8 106 272
use INVX1  _851_
timestamp 1727493700
transform 1 0 1730 0 -1 3390
box -6 -8 66 272
use NAND3X1  _852_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727494898
transform -1 0 1610 0 -1 3910
box -6 -8 106 272
use OAI21X1  _853_
timestamp 1727498925
transform -1 0 1570 0 1 3390
box -6 -8 106 272
use INVX1  _854_
timestamp 1727493700
transform 1 0 1710 0 -1 2870
box -6 -8 66 272
use NAND2X1  _855_
timestamp 1727494699
transform -1 0 1210 0 1 4430
box -6 -8 86 272
use NAND2X1  _856_
timestamp 1727494699
transform 1 0 1350 0 -1 4430
box -6 -8 86 272
use NOR2X1  _857_
timestamp 1727495070
transform 1 0 1210 0 -1 4430
box -6 -8 86 272
use INVX1  _858_
timestamp 1727493700
transform 1 0 1230 0 -1 3910
box -6 -8 66 272
use INVX1  _859_
timestamp 1727493700
transform -1 0 1170 0 -1 3910
box -6 -8 66 272
use INVX2  _860_
timestamp 1727493898
transform -1 0 4410 0 1 5470
box -6 -8 66 272
use OAI21X1  _861_
timestamp 1727498925
transform -1 0 1370 0 1 4430
box -6 -8 106 272
use NAND3X1  _862_
timestamp 1727494898
transform -1 0 1450 0 -1 3910
box -6 -8 106 272
use OAI21X1  _863_
timestamp 1727498925
transform -1 0 1510 0 1 2870
box -6 -8 106 272
use INVX1  _864_
timestamp 1727493700
transform -1 0 790 0 -1 2870
box -6 -8 66 272
use NAND2X1  _865_
timestamp 1727494699
transform 1 0 1530 0 -1 4950
box -6 -8 86 272
use NAND2X1  _866_
timestamp 1727494699
transform -1 0 1370 0 -1 5470
box -6 -8 86 272
use NOR2X1  _867_
timestamp 1727495070
transform 1 0 1270 0 -1 4950
box -6 -8 86 272
use AOI22X1  _868_
timestamp 1727487144
transform 1 0 950 0 1 4430
box -6 -8 126 272
use OAI21X1  _869_
timestamp 1727498925
transform 1 0 790 0 1 4430
box -6 -8 106 272
use INVX1  _870_
timestamp 1727493700
transform 1 0 1410 0 -1 4950
box -6 -8 66 272
use AND2X2  _871_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487319
transform -1 0 1530 0 -1 5470
box -6 -8 106 273
use NAND3X1  _872_
timestamp 1727494898
transform -1 0 1090 0 1 4950
box -6 -8 106 272
use INVX1  _873_
timestamp 1727493700
transform -1 0 570 0 1 4430
box -6 -8 66 272
use NAND3X1  _874_
timestamp 1727494898
transform -1 0 730 0 1 4430
box -6 -8 106 272
use NAND3X1  _875_
timestamp 1727494898
transform 1 0 810 0 -1 4430
box -6 -8 106 272
use INVX1  _876_
timestamp 1727493700
transform -1 0 450 0 -1 4430
box -6 -8 66 272
use AOI21X1  _877_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487319
transform -1 0 750 0 -1 4430
box -6 -8 106 272
use NOR2X1  _878_
timestamp 1727495070
transform -1 0 590 0 -1 4430
box -6 -8 86 272
use NAND2X1  _879_
timestamp 1727494699
transform -1 0 610 0 1 2870
box -6 -8 86 272
use OAI21X1  _880_
timestamp 1727498925
transform -1 0 770 0 1 2870
box -6 -8 106 272
use INVX1  _881_
timestamp 1727493700
transform -1 0 610 0 1 2350
box -6 -8 66 272
use NAND2X1  _882_
timestamp 1727494699
transform 1 0 1830 0 -1 4950
box -6 -8 86 272
use AOI21X1  _883_
timestamp 1727487319
transform 1 0 1110 0 -1 4950
box -6 -8 106 272
use NAND2X1  _884_
timestamp 1727494699
transform 1 0 1310 0 1 4950
box -6 -8 86 272
use NAND2X1  _885_
timestamp 1727494699
transform 1 0 1590 0 1 5470
box -6 -8 86 272
use NOR2X1  _886_
timestamp 1727495070
transform 1 0 1310 0 1 5470
box -6 -8 86 272
use AOI22X1  _887_
timestamp 1727487144
transform 1 0 1730 0 1 5470
box -6 -8 126 272
use OAI21X1  _888_
timestamp 1727498925
transform -1 0 1250 0 1 5470
box -6 -8 106 272
use INVX1  _889_
timestamp 1727493700
transform -1 0 930 0 -1 5470
box -6 -8 66 272
use AND2X2  _890_
timestamp 1727487319
transform -1 0 2010 0 1 5470
box -6 -8 106 273
use NAND2X1  _891_
timestamp 1727494699
transform -1 0 1070 0 -1 5470
box -6 -8 86 272
use INVX1  _892_
timestamp 1727493700
transform -1 0 930 0 1 5470
box -6 -8 66 272
use NAND3X1  _893_
timestamp 1727494898
transform -1 0 650 0 -1 5470
box -6 -8 106 272
use NAND3X1  _894_
timestamp 1727494898
transform -1 0 610 0 1 4950
box -6 -8 106 272
use OAI21X1  _895_
timestamp 1727498925
transform 1 0 950 0 -1 4950
box -6 -8 106 272
use AOI21X1  _896_
timestamp 1727487319
transform -1 0 810 0 -1 5470
box -6 -8 106 272
use INVX2  _897_
timestamp 1727493898
transform -1 0 1670 0 1 4950
box -6 -8 66 272
use OAI21X1  _898_
timestamp 1727498925
transform -1 0 1230 0 -1 5470
box -6 -8 106 272
use INVX2  _899_
timestamp 1727493898
transform 1 0 3010 0 -1 4950
box -6 -8 66 272
use INVX1  _900_
timestamp 1727493700
transform 1 0 3190 0 1 5470
box -6 -8 66 272
use OAI21X1  _901_
timestamp 1727498925
transform -1 0 1550 0 1 4950
box -6 -8 106 272
use AOI21X1  _902_
timestamp 1727487319
transform -1 0 1250 0 1 4950
box -6 -8 106 272
use OAI21X1  _903_
timestamp 1727498925
transform 1 0 790 0 -1 4950
box -6 -8 106 272
use NAND3X1  _904_
timestamp 1727494898
transform -1 0 450 0 1 4430
box -6 -8 106 272
use INVX1  _905_
timestamp 1727493700
transform -1 0 130 0 1 4430
box -6 -8 66 272
use NAND3X1  _906_
timestamp 1727494898
transform -1 0 770 0 1 4950
box -6 -8 106 272
use OAI21X1  _907_
timestamp 1727498925
transform -1 0 730 0 -1 4950
box -6 -8 106 272
use NAND3X1  _908_
timestamp 1727494898
transform -1 0 290 0 1 4430
box -6 -8 106 272
use AOI21X1  _909_
timestamp 1727487319
transform 1 0 230 0 -1 4430
box -6 -8 106 272
use NAND3X1  _910_
timestamp 1727494898
transform -1 0 170 0 -1 4430
box -6 -8 106 272
use NAND2X1  _911_
timestamp 1727494699
transform -1 0 470 0 1 2870
box -6 -8 86 272
use OAI22X1  _912_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727495774
transform -1 0 430 0 -1 2870
box -6 -8 126 272
use INVX1  _913_
timestamp 1727493700
transform 1 0 70 0 -1 2350
box -6 -8 66 272
use INVX1  _914_
timestamp 1727493700
transform 1 0 390 0 -1 3390
box -6 -8 66 272
use AOI21X1  _915_
timestamp 1727487319
transform 1 0 830 0 1 4950
box -6 -8 106 272
use OAI21X1  _916_
timestamp 1727498925
transform -1 0 450 0 1 4950
box -6 -8 106 272
use OAI21X1  _917_
timestamp 1727498925
transform 1 0 990 0 1 5470
box -6 -8 106 272
use AND2X2  _918_
timestamp 1727487319
transform 1 0 2290 0 -1 5990
box -6 -8 106 273
use NAND2X1  _919_
timestamp 1727494699
transform 1 0 1730 0 -1 5990
box -6 -8 86 272
use AOI22X1  _920_
timestamp 1727487144
transform -1 0 2190 0 1 5470
box -6 -8 126 272
use INVX1  _921_
timestamp 1727493700
transform 1 0 1150 0 -1 5990
box -6 -8 66 272
use NAND2X1  _922_
timestamp 1727494699
transform -1 0 1510 0 -1 5990
box -6 -8 86 272
use INVX1  _923_
timestamp 1727493700
transform 1 0 1030 0 -1 5990
box -6 -8 66 272
use NAND3X1  _924_
timestamp 1727494898
transform -1 0 650 0 -1 5990
box -6 -8 106 272
use NAND2X1  _925_
timestamp 1727494699
transform -1 0 2230 0 -1 5990
box -6 -8 86 272
use NOR2X1  _926_
timestamp 1727495070
transform 1 0 1450 0 1 5470
box -6 -8 86 272
use OAI21X1  _927_
timestamp 1727498925
transform -1 0 810 0 -1 5990
box -6 -8 106 272
use AOI21X1  _928_
timestamp 1727487319
transform 1 0 550 0 1 5470
box -6 -8 106 272
use AOI21X1  _929_
timestamp 1727487319
transform -1 0 810 0 1 5470
box -6 -8 106 272
use NAND3X1  _930_
timestamp 1727494898
transform -1 0 490 0 -1 5990
box -6 -8 106 272
use OAI21X1  _931_
timestamp 1727498925
transform -1 0 970 0 -1 5990
box -6 -8 106 272
use AOI21X1  _932_
timestamp 1727487319
transform 1 0 230 0 -1 5990
box -6 -8 106 272
use NAND2X1  _933_
timestamp 1727494699
transform 1 0 2130 0 -1 4950
box -6 -8 86 272
use INVX2  _934_
timestamp 1727493898
transform -1 0 3370 0 1 4430
box -6 -8 66 272
use NAND2X1  _935_
timestamp 1727494699
transform 1 0 1590 0 1 4430
box -6 -8 86 272
use OAI21X1  _936_
timestamp 1727498925
transform 1 0 1430 0 1 4430
box -6 -8 106 272
use OAI21X1  _937_
timestamp 1727498925
transform -1 0 1770 0 -1 4950
box -6 -8 106 272
use OAI21X1  _938_
timestamp 1727498925
transform -1 0 330 0 -1 5470
box -6 -8 106 272
use NAND3X1  _939_
timestamp 1727494898
transform -1 0 170 0 -1 5990
box -6 -8 106 272
use NAND3X1  _940_
timestamp 1727494898
transform -1 0 490 0 1 5470
box -6 -8 106 272
use INVX1  _941_
timestamp 1727493700
transform -1 0 130 0 1 4950
box -6 -8 66 272
use NAND3X1  _942_
timestamp 1727494898
transform -1 0 170 0 1 5470
box -6 -8 106 272
use NAND3X1  _943_
timestamp 1727494898
transform 1 0 190 0 1 4950
box -6 -8 106 272
use INVX1  _944_
timestamp 1727493700
transform -1 0 570 0 -1 4950
box -6 -8 66 272
use AOI21X1  _945_
timestamp 1727487319
transform 1 0 350 0 -1 4950
box -6 -8 106 272
use AOI21X1  _946_
timestamp 1727487319
transform -1 0 170 0 -1 5470
box -6 -8 106 272
use INVX1  _947_
timestamp 1727493700
transform -1 0 130 0 -1 4950
box -6 -8 66 272
use OAI21X1  _948_
timestamp 1727498925
transform 1 0 190 0 -1 4950
box -6 -8 106 272
use AOI21X1  _949_
timestamp 1727487319
transform -1 0 170 0 -1 3390
box -6 -8 106 272
use NAND3X1  _950_
timestamp 1727494898
transform 1 0 230 0 -1 3390
box -6 -8 106 272
use NAND2X1  _951_
timestamp 1727494699
transform 1 0 250 0 1 2870
box -6 -8 86 272
use OAI22X1  _952_
timestamp 1727495774
transform -1 0 190 0 1 2870
box -6 -8 126 272
use INVX1  _953_
timestamp 1727493700
transform 1 0 950 0 1 1830
box -6 -8 66 272
use AND2X2  _954_
timestamp 1727487319
transform 1 0 1890 0 1 3910
box -6 -8 106 273
use NAND2X1  _955_
timestamp 1727494699
transform -1 0 150 0 1 3910
box -6 -8 86 272
use INVX1  _956_
timestamp 1727493700
transform -1 0 130 0 1 3390
box -6 -8 66 272
use AOI21X1  _957_
timestamp 1727487319
transform 1 0 230 0 1 5470
box -6 -8 106 272
use NAND2X1  _958_
timestamp 1727494699
transform 1 0 2470 0 1 4430
box -6 -8 86 272
use INVX1  _959_
timestamp 1727493700
transform -1 0 1550 0 -1 4430
box -6 -8 66 272
use AND2X2  _960_
timestamp 1727487319
transform 1 0 1770 0 -1 4430
box -6 -8 106 273
use OAI21X1  _961_
timestamp 1727498925
transform -1 0 1710 0 -1 4430
box -6 -8 106 272
use INVX2  _962_
timestamp 1727493898
transform 1 0 4030 0 1 4430
box -6 -8 66 272
use OAI21X1  _963_
timestamp 1727498925
transform -1 0 2170 0 -1 4430
box -6 -8 106 272
use NAND3X1  _964_
timestamp 1727494898
transform 1 0 1850 0 1 4430
box -6 -8 106 272
use INVX1  _965_
timestamp 1727493700
transform -1 0 1790 0 1 4430
box -6 -8 66 272
use NAND2X1  _966_
timestamp 1727494699
transform -1 0 2010 0 -1 4430
box -6 -8 86 272
use OAI21X1  _967_
timestamp 1727498925
transform -1 0 2070 0 -1 4950
box -6 -8 106 272
use NAND3X1  _968_
timestamp 1727494898
transform 1 0 2010 0 1 4430
box -6 -8 106 272
use NAND2X1  _969_
timestamp 1727494699
transform 1 0 2270 0 -1 4950
box -6 -8 86 272
use AOI21X1  _970_
timestamp 1727487319
transform 1 0 1270 0 -1 5990
box -6 -8 106 272
use NAND2X1  _971_
timestamp 1727494699
transform 1 0 3310 0 1 5470
box -6 -8 86 272
use AND2X2  _972_
timestamp 1727487319
transform -1 0 3250 0 -1 5990
box -6 -8 106 273
use NAND2X1  _973_
timestamp 1727494699
transform 1 0 2710 0 1 5470
box -6 -8 86 272
use NAND2X1  _974_
timestamp 1727494699
transform 1 0 2870 0 -1 5990
box -6 -8 86 272
use NAND2X1  _975_
timestamp 1727494699
transform -1 0 2530 0 -1 5990
box -6 -8 86 272
use NAND3X1  _976_
timestamp 1727494898
transform -1 0 2650 0 1 5470
box -6 -8 106 272
use INVX1  _977_
timestamp 1727493700
transform -1 0 2590 0 -1 5470
box -6 -8 66 272
use NAND2X1  _978_
timestamp 1727494699
transform 1 0 2590 0 -1 5990
box -6 -8 86 272
use OAI21X1  _979_
timestamp 1727498925
transform -1 0 2950 0 1 5470
box -6 -8 106 272
use NAND3X1  _980_
timestamp 1727494898
transform -1 0 2470 0 -1 5470
box -6 -8 106 272
use NAND3X1  _981_
timestamp 1727494898
transform -1 0 1830 0 -1 5470
box -6 -8 106 272
use OAI21X1  _982_
timestamp 1727498925
transform 1 0 1570 0 -1 5990
box -6 -8 106 272
use AOI21X1  _983_
timestamp 1727487319
transform -1 0 2310 0 -1 5470
box -6 -8 106 272
use AOI21X1  _984_
timestamp 1727487319
transform -1 0 2490 0 1 5470
box -6 -8 106 272
use OAI21X1  _985_
timestamp 1727498925
transform -1 0 1990 0 -1 5470
box -6 -8 106 272
use NAND3X1  _986_
timestamp 1727494898
transform -1 0 1830 0 1 4950
box -6 -8 106 272
use AND2X2  _987_
timestamp 1727487319
transform 1 0 2410 0 -1 4950
box -6 -8 106 273
use NAND3X1  _988_
timestamp 1727494898
transform 1 0 2050 0 1 4950
box -6 -8 106 272
use OAI21X1  _989_
timestamp 1727498925
transform -1 0 2150 0 -1 5470
box -6 -8 106 272
use NAND3X1  _990_
timestamp 1727494898
transform 1 0 2570 0 -1 4950
box -6 -8 106 272
use NAND3X1  _991_
timestamp 1727494898
transform -1 0 310 0 1 3910
box -6 -8 106 272
use OAI21X1  _992_
timestamp 1727498925
transform -1 0 490 0 -1 5470
box -6 -8 106 272
use NAND2X1  _993_
timestamp 1727494699
transform -1 0 590 0 -1 3910
box -6 -8 86 272
use NAND2X1  _994_
timestamp 1727494699
transform -1 0 450 0 -1 3910
box -6 -8 86 272
use NAND3X1  _995_
timestamp 1727494898
transform 1 0 210 0 -1 3910
box -6 -8 106 272
use NAND3X1  _996_
timestamp 1727494898
transform -1 0 910 0 -1 3910
box -6 -8 106 272
use NAND2X1  _997_
timestamp 1727494699
transform -1 0 150 0 -1 3910
box -6 -8 86 272
use NAND3X1  _998_
timestamp 1727494898
transform 1 0 470 0 1 3390
box -6 -8 106 272
use NAND2X1  _999_
timestamp 1727494699
transform 1 0 810 0 -1 3390
box -6 -8 86 272
use NAND2X1  _1000_
timestamp 1727494699
transform -1 0 590 0 -1 3390
box -6 -8 86 272
use OR2X2  _1001_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727496117
transform 1 0 950 0 -1 3390
box -6 -8 106 272
use AOI22X1  _1002_
timestamp 1727487144
transform -1 0 770 0 -1 3390
box -6 -8 126 272
use INVX1  _1003_
timestamp 1727493700
transform -1 0 1430 0 -1 3390
box -6 -8 66 272
use NAND3X1  _1004_
timestamp 1727494898
transform -1 0 1350 0 1 2870
box -6 -8 106 272
use OAI21X1  _1005_
timestamp 1727498925
transform 1 0 1310 0 1 1830
box -6 -8 106 272
use INVX1  _1006_
timestamp 1727493700
transform 1 0 1390 0 -1 1830
box -6 -8 66 272
use AOI21X1  _1007_
timestamp 1727487319
transform -1 0 750 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1008_
timestamp 1727498925
transform 1 0 630 0 1 3390
box -6 -8 106 272
use NAND2X1  _1009_
timestamp 1727494699
transform 1 0 2330 0 1 4430
box -6 -8 86 272
use OAI21X1  _1010_
timestamp 1727498925
transform 1 0 2170 0 1 4430
box -6 -8 106 272
use INVX1  _1011_
timestamp 1727493700
transform -1 0 2190 0 -1 3910
box -6 -8 66 272
use INVX1  _1012_
timestamp 1727493700
transform 1 0 2890 0 -1 4950
box -6 -8 66 272
use AOI21X1  _1013_
timestamp 1727487319
transform 1 0 2730 0 -1 4950
box -6 -8 106 272
use NAND2X1  _1014_
timestamp 1727494699
transform 1 0 2890 0 1 4430
box -6 -8 86 272
use AND2X2  _1015_
timestamp 1727487319
transform -1 0 3690 0 -1 4950
box -6 -8 106 273
use OAI21X1  _1016_
timestamp 1727498925
transform 1 0 2610 0 1 4430
box -6 -8 106 272
use AND2X2  _1017_
timestamp 1727487319
transform -1 0 3850 0 -1 4950
box -6 -8 106 273
use OAI21X1  _1018_
timestamp 1727498925
transform 1 0 3430 0 -1 4950
box -6 -8 106 272
use NAND3X1  _1019_
timestamp 1727494898
transform 1 0 3030 0 1 4430
box -6 -8 106 272
use INVX1  _1020_
timestamp 1727493700
transform -1 0 2830 0 1 4430
box -6 -8 66 272
use NAND2X1  _1021_
timestamp 1727494699
transform 1 0 3290 0 -1 4950
box -6 -8 86 272
use OAI21X1  _1022_
timestamp 1727498925
transform 1 0 2230 0 -1 4430
box -6 -8 106 272
use NAND3X1  _1023_
timestamp 1727494898
transform 1 0 2790 0 -1 4430
box -6 -8 106 272
use NAND2X1  _1024_
timestamp 1727494699
transform 1 0 3110 0 -1 4430
box -6 -8 86 272
use NOR2X1  _1025_
timestamp 1727495070
transform -1 0 2810 0 -1 5990
box -6 -8 86 272
use AOI21X1  _1026_
timestamp 1727487319
transform 1 0 2650 0 -1 5470
box -6 -8 106 272
use NAND2X1  _1027_
timestamp 1727494699
transform 1 0 3630 0 -1 5990
box -6 -8 86 272
use AND2X2  _1028_
timestamp 1727487319
transform -1 0 4290 0 1 5470
box -6 -8 106 273
use OAI21X1  _1029_
timestamp 1727498925
transform 1 0 4030 0 1 5470
box -6 -8 106 272
use NAND2X1  _1030_
timestamp 1727494699
transform -1 0 4010 0 -1 5990
box -6 -8 86 272
use NAND3X1  _1031_
timestamp 1727494898
transform -1 0 3870 0 -1 5990
box -6 -8 106 272
use NAND3X1  _1032_
timestamp 1727494898
transform -1 0 3570 0 -1 5990
box -6 -8 106 272
use INVX1  _1033_
timestamp 1727493700
transform -1 0 3670 0 1 5470
box -6 -8 66 272
use AND2X2  _1034_
timestamp 1727487319
transform 1 0 5130 0 -1 5990
box -6 -8 106 273
use NAND2X1  _1035_
timestamp 1727494699
transform 1 0 3730 0 1 5470
box -6 -8 86 272
use OAI21X1  _1036_
timestamp 1727498925
transform 1 0 3870 0 1 5470
box -6 -8 106 272
use NAND3X1  _1037_
timestamp 1727494898
transform -1 0 3230 0 -1 5470
box -6 -8 106 272
use NAND3X1  _1038_
timestamp 1727494898
transform -1 0 2790 0 1 4950
box -6 -8 106 272
use AOI22X1  _1039_
timestamp 1727487144
transform 1 0 3010 0 1 5470
box -6 -8 126 272
use OAI21X1  _1040_
timestamp 1727498925
transform -1 0 2910 0 -1 5470
box -6 -8 106 272
use AOI21X1  _1041_
timestamp 1727487319
transform -1 0 3550 0 1 5470
box -6 -8 106 272
use AOI21X1  _1042_
timestamp 1727487319
transform -1 0 3410 0 -1 5990
box -6 -8 106 272
use OAI21X1  _1043_
timestamp 1727498925
transform -1 0 3070 0 -1 5470
box -6 -8 106 272
use NAND3X1  _1044_
timestamp 1727494898
transform -1 0 2630 0 1 4950
box -6 -8 106 272
use AND2X2  _1045_
timestamp 1727487319
transform -1 0 3050 0 -1 4430
box -6 -8 106 273
use NAND3X1  _1046_
timestamp 1727494898
transform 1 0 2850 0 1 4950
box -6 -8 106 272
use OAI21X1  _1047_
timestamp 1727498925
transform 1 0 3010 0 1 4950
box -6 -8 106 272
use NAND3X1  _1048_
timestamp 1727494898
transform -1 0 2630 0 1 3910
box -6 -8 106 272
use NAND3X1  _1049_
timestamp 1727494898
transform -1 0 2150 0 1 3910
box -6 -8 106 272
use AOI21X1  _1050_
timestamp 1727487319
transform 1 0 1890 0 1 4950
box -6 -8 106 272
use OAI21X1  _1051_
timestamp 1727498925
transform -1 0 2310 0 1 4950
box -6 -8 106 272
use AOI21X1  _1052_
timestamp 1727487319
transform -1 0 2790 0 1 3910
box -6 -8 106 272
use AOI21X1  _1053_
timestamp 1727487319
transform -1 0 2470 0 1 4950
box -6 -8 106 272
use OAI21X1  _1054_
timestamp 1727498925
transform 1 0 2370 0 1 3910
box -6 -8 106 272
use NAND3X1  _1055_
timestamp 1727494898
transform -1 0 2070 0 -1 3910
box -6 -8 106 272
use NAND3X1  _1056_
timestamp 1727494898
transform -1 0 2510 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1057_
timestamp 1727498925
transform -1 0 2310 0 1 3910
box -6 -8 106 272
use NAND3X1  _1058_
timestamp 1727494898
transform 1 0 2110 0 1 3390
box -6 -8 106 272
use NAND3X1  _1059_
timestamp 1727494898
transform -1 0 2050 0 1 3390
box -6 -8 106 272
use INVX1  _1060_
timestamp 1727493700
transform -1 0 410 0 1 3390
box -6 -8 66 272
use AOI21X1  _1061_
timestamp 1727487319
transform 1 0 190 0 1 3390
box -6 -8 106 272
use AOI21X1  _1062_
timestamp 1727487319
transform -1 0 1890 0 1 3390
box -6 -8 106 272
use AOI21X1  _1063_
timestamp 1727487319
transform -1 0 1910 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1064_
timestamp 1727498925
transform -1 0 1730 0 1 3390
box -6 -8 106 272
use AND2X2  _1065_
timestamp 1727487319
transform -1 0 2310 0 -1 3390
box -6 -8 106 273
use NOR2X1  _1066_
timestamp 1727495070
transform 1 0 1890 0 1 2870
box -6 -8 86 272
use INVX1  _1067_
timestamp 1727493700
transform 1 0 2490 0 1 2870
box -6 -8 66 272
use OAI21X1  _1068_
timestamp 1727498925
transform -1 0 2430 0 1 2870
box -6 -8 106 272
use OAI22X1  _1069_
timestamp 1727495774
transform 1 0 1710 0 1 2870
box -6 -8 126 272
use INVX1  _1070_
timestamp 1727493700
transform 1 0 890 0 -1 1310
box -6 -8 66 272
use NAND3X1  _1071_
timestamp 1727494898
transform 1 0 2370 0 -1 3390
box -6 -8 106 272
use AOI21X1  _1072_
timestamp 1727487319
transform -1 0 2350 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1073_
timestamp 1727498925
transform 1 0 2270 0 1 3390
box -6 -8 106 272
use NAND2X1  _1074_
timestamp 1727494699
transform -1 0 3090 0 -1 3910
box -6 -8 86 272
use AOI21X1  _1075_
timestamp 1727487319
transform 1 0 3170 0 1 4950
box -6 -8 106 272
use OAI21X1  _1076_
timestamp 1727498925
transform 1 0 3130 0 -1 4950
box -6 -8 106 272
use NAND2X1  _1077_
timestamp 1727494699
transform 1 0 4150 0 1 4430
box -6 -8 86 272
use AND2X2  _1078_
timestamp 1727487319
transform 1 0 4530 0 -1 4430
box -6 -8 106 273
use OAI21X1  _1079_
timestamp 1727498925
transform 1 0 4370 0 -1 4430
box -6 -8 106 272
use AND2X2  _1080_
timestamp 1727487319
transform 1 0 3770 0 -1 4430
box -6 -8 106 273
use OAI21X1  _1081_
timestamp 1727498925
transform -1 0 4030 0 -1 4430
box -6 -8 106 272
use NAND3X1  _1082_
timestamp 1727494898
transform -1 0 4190 0 -1 4430
box -6 -8 106 272
use INVX1  _1083_
timestamp 1727493700
transform 1 0 4250 0 -1 4430
box -6 -8 66 272
use NAND2X1  _1084_
timestamp 1727494699
transform 1 0 4430 0 1 3910
box -6 -8 86 272
use NAND2X1  _1085_
timestamp 1727494699
transform 1 0 4450 0 1 4430
box -6 -8 86 272
use OAI21X1  _1086_
timestamp 1727498925
transform 1 0 4290 0 1 4430
box -6 -8 106 272
use NAND3X1  _1087_
timestamp 1727494898
transform -1 0 4370 0 1 3910
box -6 -8 106 272
use NAND2X1  _1088_
timestamp 1727494699
transform -1 0 4210 0 1 3910
box -6 -8 86 272
use AOI22X1  _1089_
timestamp 1727487144
transform -1 0 3410 0 -1 5470
box -6 -8 126 272
use NAND2X1  _1090_
timestamp 1727494699
transform -1 0 4710 0 1 5470
box -6 -8 86 272
use AND2X2  _1091_
timestamp 1727487319
transform 1 0 3810 0 -1 5470
box -6 -8 106 273
use OAI21X1  _1092_
timestamp 1727498925
transform -1 0 4030 0 1 4950
box -6 -8 106 272
use OAI21X1  _1093_
timestamp 1727498925
transform -1 0 3430 0 1 4950
box -6 -8 106 272
use NAND3X1  _1094_
timestamp 1727494898
transform -1 0 3710 0 1 4950
box -6 -8 106 272
use INVX1  _1095_
timestamp 1727493700
transform -1 0 4490 0 -1 5470
box -6 -8 66 272
use NAND2X1  _1096_
timestamp 1727494699
transform -1 0 4050 0 -1 5470
box -6 -8 86 272
use AOI22X1  _1097_
timestamp 1727487144
transform -1 0 4330 0 -1 5990
box -6 -8 126 272
use INVX1  _1098_
timestamp 1727493700
transform -1 0 4590 0 -1 5990
box -6 -8 66 272
use NAND3X1  _1099_
timestamp 1727494898
transform -1 0 4210 0 -1 5470
box -6 -8 106 272
use NAND3X1  _1100_
timestamp 1727494898
transform 1 0 3710 0 1 4430
box -6 -8 106 272
use AOI22X1  _1101_
timestamp 1727487144
transform -1 0 3750 0 -1 5470
box -6 -8 126 272
use OAI21X1  _1102_
timestamp 1727498925
transform -1 0 3570 0 -1 5470
box -6 -8 106 272
use AOI21X1  _1103_
timestamp 1727487319
transform -1 0 4370 0 -1 5470
box -6 -8 106 272
use AOI21X1  _1104_
timestamp 1727487319
transform 1 0 3770 0 1 4950
box -6 -8 106 272
use OAI21X1  _1105_
timestamp 1727498925
transform -1 0 4010 0 -1 4950
box -6 -8 106 272
use NAND3X1  _1106_
timestamp 1727494898
transform -1 0 3910 0 1 3910
box -6 -8 106 272
use AND2X2  _1107_
timestamp 1727487319
transform -1 0 4170 0 -1 3910
box -6 -8 106 273
use NAND3X1  _1108_
timestamp 1727494898
transform -1 0 3650 0 1 4430
box -6 -8 106 272
use OAI21X1  _1109_
timestamp 1727498925
transform 1 0 4070 0 -1 4950
box -6 -8 106 272
use NAND3X1  _1110_
timestamp 1727494898
transform -1 0 3730 0 -1 3910
box -6 -8 106 272
use NAND3X1  _1111_
timestamp 1727494898
transform -1 0 3330 0 1 3390
box -6 -8 106 272
use INVX1  _1112_
timestamp 1727493700
transform -1 0 3310 0 -1 4430
box -6 -8 66 272
use AOI21X1  _1113_
timestamp 1727487319
transform 1 0 3090 0 1 3910
box -6 -8 106 272
use AOI21X1  _1114_
timestamp 1727487319
transform -1 0 3570 0 -1 3910
box -6 -8 106 272
use AOI21X1  _1115_
timestamp 1727487319
transform -1 0 3750 0 1 3910
box -6 -8 106 272
use OAI21X1  _1116_
timestamp 1727498925
transform -1 0 3250 0 -1 3910
box -6 -8 106 272
use NAND3X1  _1117_
timestamp 1727494898
transform -1 0 2850 0 1 3390
box -6 -8 106 272
use INVX1  _1118_
timestamp 1727493700
transform 1 0 3590 0 -1 3390
box -6 -8 66 272
use NAND3X1  _1119_
timestamp 1727494898
transform -1 0 3170 0 1 3390
box -6 -8 106 272
use OAI21X1  _1120_
timestamp 1727498925
transform 1 0 3310 0 -1 3910
box -6 -8 106 272
use NAND3X1  _1121_
timestamp 1727494898
transform -1 0 3370 0 -1 3390
box -6 -8 106 272
use AOI21X1  _1122_
timestamp 1727487319
transform -1 0 2770 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1123_
timestamp 1727494898
transform -1 0 3010 0 1 3390
box -6 -8 106 272
use NAND3X1  _1124_
timestamp 1727494898
transform -1 0 3530 0 -1 3390
box -6 -8 106 272
use AOI22X1  _1125_
timestamp 1727487144
transform 1 0 2430 0 1 3390
box -6 -8 126 272
use NOR2X1  _1126_
timestamp 1727495070
transform -1 0 2610 0 -1 3390
box -6 -8 86 272
use AOI21X1  _1127_
timestamp 1727487319
transform -1 0 2850 0 1 2870
box -6 -8 106 272
use OAI21X1  _1128_
timestamp 1727498925
transform 1 0 2610 0 1 2870
box -6 -8 106 272
use INVX1  _1129_
timestamp 1727493700
transform -1 0 3050 0 -1 3390
box -6 -8 66 272
use NAND3X1  _1130_
timestamp 1727494898
transform 1 0 3110 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1131_
timestamp 1727494898
transform 1 0 2830 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1132_
timestamp 1727494699
transform 1 0 3210 0 1 2870
box -6 -8 86 272
use NOR2X1  _1133_
timestamp 1727495070
transform -1 0 2730 0 -1 2870
box -6 -8 86 272
use OAI21X1  _1134_
timestamp 1727498925
transform 1 0 2790 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1135_
timestamp 1727498925
transform 1 0 1250 0 -1 1310
box -6 -8 106 272
use INVX1  _1136_
timestamp 1727493700
transform 1 0 4150 0 -1 2350
box -6 -8 66 272
use NAND2X1  _1137_
timestamp 1727494699
transform -1 0 3150 0 1 2870
box -6 -8 86 272
use NAND2X1  _1138_
timestamp 1727494699
transform 1 0 3350 0 1 2870
box -6 -8 86 272
use OAI21X1  _1139_
timestamp 1727498925
transform 1 0 3230 0 -1 2870
box -6 -8 106 272
use AOI21X1  _1140_
timestamp 1727487319
transform 1 0 3390 0 1 3390
box -6 -8 106 272
use OAI21X1  _1141_
timestamp 1727498925
transform 1 0 3710 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1142_
timestamp 1727494699
transform 1 0 4230 0 -1 3910
box -6 -8 86 272
use INVX1  _1143_
timestamp 1727493700
transform 1 0 4030 0 1 3390
box -6 -8 66 272
use INVX1  _1144_
timestamp 1727493700
transform -1 0 3850 0 -1 3910
box -6 -8 66 272
use AOI21X1  _1145_
timestamp 1727487319
transform 1 0 3910 0 -1 3910
box -6 -8 106 272
use INVX2  _1146_
timestamp 1727493898
transform -1 0 5050 0 1 4950
box -6 -8 66 272
use NOR2X1  _1147_
timestamp 1727495070
transform 1 0 4390 0 1 4950
box -6 -8 86 272
use AND2X2  _1148_
timestamp 1727487319
transform 1 0 5110 0 1 5470
box -6 -8 106 273
use NAND3X1  _1149_
timestamp 1727494898
transform 1 0 4950 0 1 5470
box -6 -8 106 272
use AOI22X1  _1150_
timestamp 1727487144
transform 1 0 4950 0 -1 5990
box -6 -8 126 272
use INVX1  _1151_
timestamp 1727493700
transform -1 0 4770 0 1 4950
box -6 -8 66 272
use NAND3X1  _1152_
timestamp 1727494898
transform -1 0 4810 0 -1 5470
box -6 -8 106 272
use NAND2X1  _1153_
timestamp 1727494699
transform 1 0 5130 0 -1 4950
box -6 -8 86 272
use NOR2X1  _1154_
timestamp 1727495070
transform 1 0 4830 0 -1 4950
box -6 -8 86 272
use OAI22X1  _1155_
timestamp 1727495774
transform 1 0 4530 0 1 4950
box -6 -8 126 272
use NAND2X1  _1156_
timestamp 1727494699
transform 1 0 4870 0 -1 5470
box -6 -8 86 272
use AND2X2  _1157_
timestamp 1727487319
transform -1 0 4890 0 -1 5990
box -6 -8 106 273
use AOI22X1  _1158_
timestamp 1727487144
transform 1 0 4770 0 1 5470
box -6 -8 126 272
use NAND2X1  _1159_
timestamp 1727494699
transform 1 0 5470 0 -1 5990
box -6 -8 86 272
use NAND2X1  _1160_
timestamp 1727494699
transform -1 0 5350 0 1 5470
box -6 -8 86 272
use AOI22X1  _1161_
timestamp 1727487144
transform -1 0 5410 0 -1 5990
box -6 -8 126 272
use INVX1  _1162_
timestamp 1727493700
transform 1 0 5770 0 -1 5990
box -6 -8 66 272
use OAI21X1  _1163_
timestamp 1727498925
transform 1 0 5610 0 -1 5990
box -6 -8 106 272
use NOR2X1  _1164_
timestamp 1727495070
transform -1 0 5830 0 -1 5470
box -6 -8 86 272
use OAI21X1  _1165_
timestamp 1727498925
transform -1 0 4570 0 1 5470
box -6 -8 106 272
use INVX1  _1166_
timestamp 1727493700
transform -1 0 5370 0 -1 5470
box -6 -8 66 272
use AOI21X1  _1167_
timestamp 1727487319
transform 1 0 5410 0 1 5470
box -6 -8 106 272
use NOR2X1  _1168_
timestamp 1727495070
transform 1 0 5570 0 1 5470
box -6 -8 86 272
use OAI21X1  _1169_
timestamp 1727498925
transform 1 0 5430 0 -1 5470
box -6 -8 106 272
use AND2X2  _1170_
timestamp 1727487319
transform 1 0 4550 0 -1 5470
box -6 -8 106 273
use NAND2X1  _1171_
timestamp 1727494699
transform 1 0 5850 0 1 5470
box -6 -8 86 272
use NAND2X1  _1172_
timestamp 1727494699
transform -1 0 5250 0 -1 5470
box -6 -8 86 272
use NAND2X1  _1173_
timestamp 1727494699
transform 1 0 5110 0 1 4950
box -6 -8 86 272
use NAND2X1  _1174_
timestamp 1727494699
transform 1 0 4890 0 1 3910
box -6 -8 86 272
use NAND3X1  _1175_
timestamp 1727494898
transform -1 0 4630 0 -1 3910
box -6 -8 106 272
use AOI21X1  _1176_
timestamp 1727487319
transform 1 0 3870 0 1 4430
box -6 -8 106 272
use OAI21X1  _1177_
timestamp 1727498925
transform -1 0 4070 0 1 3910
box -6 -8 106 272
use NOR2X1  _1178_
timestamp 1727495070
transform 1 0 4690 0 -1 4430
box -6 -8 86 272
use AOI21X1  _1179_
timestamp 1727487319
transform -1 0 5110 0 -1 5470
box -6 -8 106 272
use OAI21X1  _1180_
timestamp 1727498925
transform 1 0 4730 0 1 3910
box -6 -8 106 272
use NAND3X1  _1181_
timestamp 1727494898
transform -1 0 4410 0 1 3390
box -6 -8 106 272
use NAND3X1  _1182_
timestamp 1727494898
transform 1 0 4850 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1183_
timestamp 1727498925
transform -1 0 4670 0 1 3910
box -6 -8 106 272
use NAND3X1  _1184_
timestamp 1727494898
transform 1 0 3870 0 1 3390
box -6 -8 106 272
use NAND3X1  _1185_
timestamp 1727494898
transform 1 0 3990 0 -1 3390
box -6 -8 106 272
use INVX1  _1186_
timestamp 1727493700
transform -1 0 3930 0 -1 3390
box -6 -8 66 272
use AOI21X1  _1187_
timestamp 1727487319
transform -1 0 3810 0 1 3390
box -6 -8 106 272
use AOI21X1  _1188_
timestamp 1727487319
transform -1 0 4250 0 1 3390
box -6 -8 106 272
use OAI21X1  _1189_
timestamp 1727498925
transform -1 0 3650 0 1 3390
box -6 -8 106 272
use NAND2X1  _1190_
timestamp 1727494699
transform -1 0 4230 0 -1 3390
box -6 -8 86 272
use INVX1  _1191_
timestamp 1727493700
transform 1 0 4390 0 -1 2870
box -6 -8 66 272
use NOR2X1  _1192_
timestamp 1727495070
transform 1 0 4510 0 1 2350
box -6 -8 86 272
use INVX1  _1193_
timestamp 1727493700
transform -1 0 4170 0 -1 2870
box -6 -8 66 272
use OAI21X1  _1194_
timestamp 1727498925
transform 1 0 4230 0 -1 2870
box -6 -8 106 272
use OAI22X1  _1195_
timestamp 1727495774
transform 1 0 4330 0 1 2350
box -6 -8 126 272
use INVX1  _1196_
timestamp 1727493700
transform 1 0 4550 0 -1 1830
box -6 -8 66 272
use INVX8  _1197_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727494223
transform -1 0 2370 0 -1 790
box -6 -8 126 272
use INVX1  _1198_
timestamp 1727493700
transform -1 0 4570 0 -1 2870
box -6 -8 66 272
use AOI21X1  _1199_
timestamp 1727487319
transform 1 0 4650 0 1 2350
box -6 -8 106 272
use AOI21X1  _1200_
timestamp 1727487319
transform -1 0 4790 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1201_
timestamp 1727498925
transform 1 0 4630 0 1 3390
box -6 -8 106 272
use AOI21X1  _1202_
timestamp 1727487319
transform 1 0 4830 0 1 4950
box -6 -8 106 272
use INVX1  _1203_
timestamp 1727493700
transform -1 0 5330 0 1 3390
box -6 -8 66 272
use NAND2X1  _1204_
timestamp 1727494699
transform -1 0 5790 0 1 5470
box -6 -8 86 272
use OAI21X1  _1205_
timestamp 1727498925
transform 1 0 5590 0 -1 5470
box -6 -8 106 272
use NOR2X1  _1206_
timestamp 1727495070
transform -1 0 4670 0 1 4430
box -6 -8 86 272
use NAND2X1  _1207_
timestamp 1727494699
transform 1 0 5030 0 1 3910
box -6 -8 86 272
use INVX1  _1208_
timestamp 1727493700
transform 1 0 5150 0 -1 3910
box -6 -8 66 272
use NAND2X1  _1209_
timestamp 1727494699
transform 1 0 5270 0 -1 4950
box -6 -8 86 272
use OAI21X1  _1210_
timestamp 1727498925
transform 1 0 4970 0 -1 4950
box -6 -8 106 272
use NAND3X1  _1211_
timestamp 1727494898
transform 1 0 5190 0 1 4430
box -6 -8 106 272
use NAND2X1  _1212_
timestamp 1727494699
transform -1 0 4970 0 1 4430
box -6 -8 86 272
use OAI21X1  _1213_
timestamp 1727498925
transform -1 0 5130 0 1 4430
box -6 -8 106 272
use OAI21X1  _1214_
timestamp 1727498925
transform 1 0 4730 0 1 4430
box -6 -8 106 272
use NAND2X1  _1215_
timestamp 1727494699
transform 1 0 5790 0 -1 4950
box -6 -8 86 272
use OAI21X1  _1216_
timestamp 1727498925
transform 1 0 5690 0 1 4950
box -6 -8 106 272
use OAI21X1  _1217_
timestamp 1727498925
transform 1 0 5250 0 1 4950
box -6 -8 106 272
use INVX1  _1218_
timestamp 1727493700
transform 1 0 5530 0 -1 4950
box -6 -8 66 272
use NAND3X1  _1219_
timestamp 1727494898
transform 1 0 5930 0 -1 4950
box -6 -8 106 272
use NAND3X1  _1220_
timestamp 1727494898
transform -1 0 5850 0 -1 4430
box -6 -8 106 272
use NAND2X1  _1221_
timestamp 1727494699
transform 1 0 5990 0 1 5470
box -6 -8 86 272
use AOI21X1  _1222_
timestamp 1727487319
transform 1 0 5890 0 -1 5470
box -6 -8 106 272
use AOI21X1  _1223_
timestamp 1727487319
transform 1 0 5490 0 1 4430
box -6 -8 106 272
use INVX1  _1224_
timestamp 1727493700
transform 1 0 5970 0 1 4430
box -6 -8 66 272
use OAI21X1  _1225_
timestamp 1727498925
transform 1 0 5810 0 1 4430
box -6 -8 106 272
use NAND3X1  _1226_
timestamp 1727494898
transform 1 0 5390 0 1 3390
box -6 -8 106 272
use NAND3X1  _1227_
timestamp 1727494898
transform 1 0 5910 0 -1 4430
box -6 -8 106 272
use OAI21X1  _1228_
timestamp 1727498925
transform -1 0 5750 0 1 4430
box -6 -8 106 272
use NAND3X1  _1229_
timestamp 1727494898
transform -1 0 5370 0 -1 3910
box -6 -8 106 272
use AOI21X1  _1230_
timestamp 1727487319
transform -1 0 5130 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1231_
timestamp 1727494898
transform 1 0 5430 0 -1 3910
box -6 -8 106 272
use NAND3X1  _1232_
timestamp 1727494898
transform -1 0 5210 0 1 3390
box -6 -8 106 272
use AOI22X1  _1233_
timestamp 1727487144
transform -1 0 5050 0 1 3390
box -6 -8 126 272
use NOR2X1  _1234_
timestamp 1727495070
transform 1 0 4890 0 -1 3390
box -6 -8 86 272
use OR2X2  _1235_
timestamp 1727496117
transform 1 0 4750 0 -1 2350
box -6 -8 106 272
use AOI21X1  _1236_
timestamp 1727487319
transform 1 0 4410 0 -1 2350
box -6 -8 106 272
use AOI22X1  _1237_
timestamp 1727487144
transform 1 0 4570 0 -1 2350
box -6 -8 126 272
use INVX1  _1238_
timestamp 1727493700
transform -1 0 3110 0 1 1830
box -6 -8 66 272
use NAND2X1  _1239_
timestamp 1727494699
transform 1 0 4790 0 1 3390
box -6 -8 86 272
use NAND3X1  _1240_
timestamp 1727494898
transform -1 0 4570 0 1 3390
box -6 -8 106 272
use NAND3X1  _1241_
timestamp 1727494898
transform -1 0 4830 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1242_
timestamp 1727494699
transform -1 0 4510 0 -1 3390
box -6 -8 86 272
use NOR2X1  _1243_
timestamp 1727495070
transform -1 0 4370 0 -1 3390
box -6 -8 86 272
use OAI21X1  _1244_
timestamp 1727498925
transform 1 0 4570 0 -1 3390
box -6 -8 106 272
use AOI21X1  _1245_
timestamp 1727487319
transform -1 0 4330 0 1 2870
box -6 -8 106 272
use NAND2X1  _1246_
timestamp 1727494699
transform -1 0 5730 0 -1 3390
box -6 -8 86 272
use OAI21X1  _1247_
timestamp 1727498925
transform 1 0 5170 0 1 3910
box -6 -8 106 272
use INVX1  _1248_
timestamp 1727493700
transform -1 0 5650 0 -1 3910
box -6 -8 66 272
use NAND2X1  _1249_
timestamp 1727494699
transform -1 0 5490 0 1 4950
box -6 -8 86 272
use NAND2X1  _1250_
timestamp 1727494699
transform 1 0 5350 0 1 4430
box -6 -8 86 272
use NAND2X1  _1251_
timestamp 1727494699
transform 1 0 5310 0 -1 4430
box -6 -8 86 272
use OAI21X1  _1252_
timestamp 1727498925
transform 1 0 4990 0 -1 4430
box -6 -8 106 272
use NAND2X1  _1253_
timestamp 1727494699
transform -1 0 5530 0 -1 4430
box -6 -8 86 272
use OAI21X1  _1254_
timestamp 1727498925
transform -1 0 5250 0 -1 4430
box -6 -8 106 272
use OR2X2  _1255_
timestamp 1727496117
transform 1 0 5590 0 -1 4430
box -6 -8 106 272
use OAI21X1  _1256_
timestamp 1727498925
transform 1 0 4830 0 -1 4430
box -6 -8 106 272
use NAND2X1  _1257_
timestamp 1727494699
transform 1 0 5650 0 1 3910
box -6 -8 86 272
use AOI21X1  _1258_
timestamp 1727487319
transform -1 0 5890 0 1 3910
box -6 -8 106 272
use NAND3X1  _1259_
timestamp 1727494898
transform 1 0 5950 0 1 3910
box -6 -8 106 272
use INVX1  _1260_
timestamp 1727493700
transform 1 0 5870 0 -1 3910
box -6 -8 66 272
use OAI21X1  _1261_
timestamp 1727498925
transform -1 0 5810 0 -1 3910
box -6 -8 106 272
use INVX1  _1262_
timestamp 1727493700
transform -1 0 5610 0 1 3390
box -6 -8 66 272
use NAND3X1  _1263_
timestamp 1727494898
transform -1 0 5770 0 1 3390
box -6 -8 106 272
use NAND3X1  _1264_
timestamp 1727494898
transform -1 0 5890 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1265_
timestamp 1727494699
transform 1 0 5950 0 -1 3390
box -6 -8 86 272
use NAND3X1  _1266_
timestamp 1727494898
transform -1 0 5590 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1267_
timestamp 1727494699
transform 1 0 4970 0 1 2870
box -6 -8 86 272
use NAND2X1  _1268_
timestamp 1727494699
transform -1 0 3730 0 1 2870
box -6 -8 86 272
use NAND3X1  _1269_
timestamp 1727494898
transform 1 0 2910 0 1 2870
box -6 -8 106 272
use NAND3X1  _1270_
timestamp 1727494898
transform 1 0 4390 0 1 2870
box -6 -8 106 272
use AOI21X1  _1271_
timestamp 1727487319
transform 1 0 3490 0 1 2870
box -6 -8 106 272
use INVX1  _1272_
timestamp 1727493700
transform 1 0 4110 0 1 2870
box -6 -8 66 272
use OAI21X1  _1273_
timestamp 1727498925
transform 1 0 3950 0 1 2870
box -6 -8 106 272
use NAND3X1  _1274_
timestamp 1727494898
transform -1 0 3490 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1275_
timestamp 1727498925
transform 1 0 2970 0 1 2350
box -6 -8 106 272
use NAND2X1  _1276_
timestamp 1727494699
transform -1 0 3350 0 -1 1310
box -6 -8 86 272
use AOI21X1  _1277_
timestamp 1727487319
transform 1 0 5830 0 1 3390
box -6 -8 106 272
use OAI21X1  _1278_
timestamp 1727498925
transform 1 0 5490 0 1 3910
box -6 -8 106 272
use OAI21X1  _1279_
timestamp 1727498925
transform 1 0 5330 0 1 3910
box -6 -8 106 272
use NOR2X1  _1280_
timestamp 1727495070
transform 1 0 5010 0 -1 3910
box -6 -8 86 272
use NAND2X1  _1281_
timestamp 1727494699
transform -1 0 5270 0 -1 3390
box -6 -8 86 272
use AND2X2  _1282_
timestamp 1727487319
transform 1 0 5330 0 -1 3390
box -6 -8 106 273
use OR2X2  _1283_
timestamp 1727496117
transform 1 0 5810 0 1 2870
box -6 -8 106 272
use NAND2X1  _1284_
timestamp 1727494699
transform 1 0 5670 0 1 2870
box -6 -8 86 272
use NAND2X1  _1285_
timestamp 1727494699
transform 1 0 5970 0 1 2870
box -6 -8 86 272
use NOR2X1  _1286_
timestamp 1727495070
transform 1 0 5930 0 -1 2870
box -6 -8 86 272
use AND2X2  _1287_
timestamp 1727487319
transform -1 0 5870 0 -1 2870
box -6 -8 106 273
use NOR2X1  _1288_
timestamp 1727495070
transform -1 0 5270 0 -1 2870
box -6 -8 86 272
use INVX1  _1289_
timestamp 1727493700
transform -1 0 4050 0 -1 2870
box -6 -8 66 272
use NAND3X1  _1290_
timestamp 1727494898
transform -1 0 3950 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1291_
timestamp 1727498925
transform 1 0 3790 0 1 2870
box -6 -8 106 272
use NAND2X1  _1292_
timestamp 1727494699
transform -1 0 3790 0 -1 2870
box -6 -8 86 272
use NAND3X1  _1293_
timestamp 1727494898
transform -1 0 3650 0 -1 2870
box -6 -8 106 272
use NAND2X1  _1294_
timestamp 1727494699
transform 1 0 3410 0 -1 1310
box -6 -8 86 272
use INVX1  _1295_
timestamp 1727493700
transform -1 0 6030 0 -1 2350
box -6 -8 66 272
use NAND3X1  _1296_
timestamp 1727494898
transform -1 0 4910 0 1 2870
box -6 -8 106 272
use NOR2X1  _1297_
timestamp 1727495070
transform -1 0 4710 0 -1 2870
box -6 -8 86 272
use INVX1  _1298_
timestamp 1727493700
transform 1 0 4690 0 1 2870
box -6 -8 66 272
use NOR2X1  _1299_
timestamp 1727495070
transform 1 0 5630 0 -1 2870
box -6 -8 86 272
use NOR2X1  _1300_
timestamp 1727495070
transform 1 0 5490 0 -1 2870
box -6 -8 86 272
use OAI21X1  _1301_
timestamp 1727498925
transform 1 0 4770 0 -1 2870
box -6 -8 106 272
use AOI21X1  _1302_
timestamp 1727487319
transform 1 0 4810 0 1 2350
box -6 -8 106 272
use INVX1  _1303_
timestamp 1727493700
transform 1 0 5550 0 1 2870
box -6 -8 66 272
use NAND3X1  _1304_
timestamp 1727494898
transform -1 0 5490 0 1 2870
box -6 -8 106 272
use INVX1  _1305_
timestamp 1727493700
transform 1 0 5270 0 1 2870
box -6 -8 66 272
use OAI21X1  _1306_
timestamp 1727498925
transform 1 0 5330 0 -1 2870
box -6 -8 106 272
use NAND2X1  _1307_
timestamp 1727494699
transform 1 0 5390 0 1 2350
box -6 -8 86 272
use NAND2X1  _1308_
timestamp 1727494699
transform -1 0 5610 0 -1 2350
box -6 -8 86 272
use INVX1  _1309_
timestamp 1727493700
transform 1 0 5670 0 -1 2350
box -6 -8 66 272
use OAI21X1  _1310_
timestamp 1727498925
transform 1 0 5690 0 1 2350
box -6 -8 106 272
use OAI22X1  _1311_
timestamp 1727495774
transform -1 0 5910 0 -1 2350
box -6 -8 126 272
use INVX1  _1312_
timestamp 1727493700
transform 1 0 5150 0 -1 2350
box -6 -8 66 272
use OR2X2  _1313_
timestamp 1727496117
transform -1 0 5630 0 1 2350
box -6 -8 106 272
use INVX1  _1314_
timestamp 1727493700
transform -1 0 4990 0 -1 2870
box -6 -8 66 272
use OAI21X1  _1315_
timestamp 1727498925
transform -1 0 5210 0 1 2870
box -6 -8 106 272
use NOR2X1  _1316_
timestamp 1727495070
transform -1 0 5130 0 -1 2870
box -6 -8 86 272
use AOI22X1  _1317_
timestamp 1727487144
transform 1 0 5210 0 1 2350
box -6 -8 126 272
use NOR2X1  _1318_
timestamp 1727495070
transform -1 0 2050 0 -1 2870
box -6 -8 86 272
use INVX1  _1319_
timestamp 1727493700
transform 1 0 2110 0 -1 2870
box -6 -8 66 272
use NAND2X1  _1320_
timestamp 1727494699
transform -1 0 2110 0 1 2870
box -6 -8 86 272
use NAND2X1  _1321_
timestamp 1727494699
transform 1 0 2150 0 1 2350
box -6 -8 86 272
use NAND2X1  _1322_
timestamp 1727494699
transform 1 0 2350 0 -1 1310
box -6 -8 86 272
use OAI21X1  _1323_
timestamp 1727498925
transform 1 0 2190 0 -1 1310
box -6 -8 106 272
use NOR2X1  _1324_
timestamp 1727495070
transform 1 0 1570 0 1 2350
box -6 -8 86 272
use NOR2X1  _1325_
timestamp 1727495070
transform 1 0 1830 0 -1 2870
box -6 -8 86 272
use NOR2X1  _1326_
timestamp 1727495070
transform -1 0 1790 0 1 2350
box -6 -8 86 272
use NAND2X1  _1327_
timestamp 1727494699
transform -1 0 1930 0 1 2350
box -6 -8 86 272
use OAI21X1  _1328_
timestamp 1727498925
transform 1 0 1990 0 1 2350
box -6 -8 106 272
use NAND2X1  _1329_
timestamp 1727494699
transform -1 0 2370 0 1 2350
box -6 -8 86 272
use NAND2X1  _1330_
timestamp 1727494699
transform -1 0 2430 0 -1 270
box -6 -8 86 272
use OAI21X1  _1331_
timestamp 1727498925
transform -1 0 2590 0 -1 270
box -6 -8 106 272
use OAI21X1  _1332_
timestamp 1727498925
transform -1 0 1510 0 1 2350
box -6 -8 106 272
use NOR2X1  _1333_
timestamp 1727495070
transform -1 0 930 0 -1 2870
box -6 -8 86 272
use NOR2X1  _1334_
timestamp 1727495070
transform -1 0 910 0 1 2870
box -6 -8 86 272
use NOR2X1  _1335_
timestamp 1727495070
transform -1 0 910 0 1 2350
box -6 -8 86 272
use NAND2X1  _1336_
timestamp 1727494699
transform 1 0 1130 0 1 2350
box -6 -8 86 272
use OR2X2  _1337_
timestamp 1727496117
transform 1 0 970 0 1 2350
box -6 -8 106 272
use NAND2X1  _1338_
timestamp 1727494699
transform 1 0 1270 0 1 2350
box -6 -8 86 272
use NAND2X1  _1339_
timestamp 1727494699
transform 1 0 1790 0 -1 790
box -6 -8 86 272
use OAI21X1  _1340_
timestamp 1727498925
transform 1 0 1630 0 -1 790
box -6 -8 106 272
use AOI21X1  _1341_
timestamp 1727487319
transform -1 0 770 0 1 2350
box -6 -8 106 272
use NOR2X1  _1342_
timestamp 1727495070
transform -1 0 650 0 -1 2350
box -6 -8 86 272
use NOR2X1  _1343_
timestamp 1727495070
transform -1 0 510 0 -1 2350
box -6 -8 86 272
use OAI21X1  _1344_
timestamp 1727498925
transform 1 0 650 0 1 1830
box -6 -8 106 272
use INVX1  _1345_
timestamp 1727493700
transform -1 0 250 0 -1 2350
box -6 -8 66 272
use INVX1  _1346_
timestamp 1727493700
transform -1 0 590 0 1 1830
box -6 -8 66 272
use INVX1  _1347_
timestamp 1727493700
transform -1 0 370 0 -1 2350
box -6 -8 66 272
use NAND3X1  _1348_
timestamp 1727494898
transform -1 0 310 0 1 1830
box -6 -8 106 272
use NAND2X1  _1349_
timestamp 1727494699
transform 1 0 810 0 1 1830
box -6 -8 86 272
use NAND2X1  _1350_
timestamp 1727494699
transform 1 0 1770 0 1 270
box -6 -8 86 272
use OAI21X1  _1351_
timestamp 1727498925
transform 1 0 1370 0 1 270
box -6 -8 106 272
use NAND2X1  _1352_
timestamp 1727494699
transform -1 0 1570 0 -1 790
box -6 -8 86 272
use NOR2X1  _1353_
timestamp 1727495070
transform -1 0 150 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1354_
timestamp 1727495070
transform -1 0 150 0 1 1830
box -6 -8 86 272
use OAI21X1  _1355_
timestamp 1727498925
transform -1 0 470 0 1 1830
box -6 -8 106 272
use INVX1  _1356_
timestamp 1727493700
transform 1 0 370 0 -1 1310
box -6 -8 66 272
use OAI21X1  _1357_
timestamp 1727498925
transform 1 0 210 0 -1 1310
box -6 -8 106 272
use NOR2X1  _1358_
timestamp 1727495070
transform -1 0 150 0 -1 1310
box -6 -8 86 272
use NAND2X1  _1359_
timestamp 1727494699
transform 1 0 230 0 1 790
box -6 -8 86 272
use NAND2X1  _1360_
timestamp 1727494699
transform 1 0 490 0 -1 1310
box -6 -8 86 272
use OAI21X1  _1361_
timestamp 1727498925
transform 1 0 1410 0 1 790
box -6 -8 106 272
use INVX1  _1362_
timestamp 1727493700
transform -1 0 130 0 -1 270
box -6 -8 66 272
use AOI21X1  _1363_
timestamp 1727487319
transform -1 0 170 0 1 790
box -6 -8 106 272
use NOR2X1  _1364_
timestamp 1727495070
transform -1 0 810 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1365_
timestamp 1727495070
transform -1 0 450 0 1 1310
box -6 -8 86 272
use NOR2X1  _1366_
timestamp 1727495070
transform -1 0 590 0 1 1310
box -6 -8 86 272
use AND2X2  _1367_
timestamp 1727487319
transform 1 0 370 0 1 270
box -6 -8 106 273
use NOR2X1  _1368_
timestamp 1727495070
transform -1 0 150 0 1 270
box -6 -8 86 272
use OAI21X1  _1369_
timestamp 1727498925
transform 1 0 210 0 1 270
box -6 -8 106 272
use OAI21X1  _1370_
timestamp 1727498925
transform 1 0 190 0 -1 270
box -6 -8 106 272
use NAND2X1  _1371_
timestamp 1727494699
transform 1 0 1310 0 -1 270
box -6 -8 86 272
use NAND2X1  _1372_
timestamp 1727494699
transform -1 0 150 0 1 1310
box -6 -8 86 272
use OAI21X1  _1373_
timestamp 1727498925
transform -1 0 310 0 1 1310
box -6 -8 106 272
use AND2X2  _1374_
timestamp 1727487319
transform 1 0 70 0 -1 790
box -6 -8 106 273
use AOI21X1  _1375_
timestamp 1727487319
transform 1 0 230 0 -1 790
box -6 -8 106 272
use NOR2X1  _1376_
timestamp 1727495070
transform -1 0 1070 0 1 790
box -6 -8 86 272
use NOR2X1  _1377_
timestamp 1727495070
transform 1 0 1350 0 -1 790
box -6 -8 86 272
use NOR2X1  _1378_
timestamp 1727495070
transform 1 0 970 0 -1 790
box -6 -8 86 272
use INVX1  _1379_
timestamp 1727493700
transform -1 0 870 0 1 270
box -6 -8 66 272
use AND2X2  _1380_
timestamp 1727487319
transform 1 0 750 0 -1 270
box -6 -8 106 273
use OAI21X1  _1381_
timestamp 1727498925
transform -1 0 690 0 -1 270
box -6 -8 106 272
use OAI21X1  _1382_
timestamp 1727498925
transform 1 0 910 0 -1 270
box -6 -8 106 272
use INVX1  _1383_
timestamp 1727493700
transform -1 0 750 0 -1 790
box -6 -8 66 272
use OAI21X1  _1384_
timestamp 1727498925
transform -1 0 910 0 -1 790
box -6 -8 106 272
use NOR2X1  _1385_
timestamp 1727495070
transform 1 0 630 0 -1 1310
box -6 -8 86 272
use NOR2X1  _1386_
timestamp 1727495070
transform 1 0 850 0 1 790
box -6 -8 86 272
use NOR2X1  _1387_
timestamp 1727495070
transform -1 0 470 0 -1 790
box -6 -8 86 272
use OR2X2  _1388_
timestamp 1727496117
transform 1 0 1070 0 1 270
box -6 -8 106 272
use NAND2X1  _1389_
timestamp 1727494699
transform -1 0 1010 0 1 270
box -6 -8 86 272
use NAND2X1  _1390_
timestamp 1727494699
transform 1 0 1230 0 1 270
box -6 -8 86 272
use NAND2X1  _1391_
timestamp 1727494699
transform 1 0 1850 0 -1 270
box -6 -8 86 272
use OAI21X1  _1392_
timestamp 1727498925
transform 1 0 1450 0 -1 270
box -6 -8 106 272
use NAND2X1  _1393_
timestamp 1727494699
transform -1 0 4370 0 1 790
box -6 -8 86 272
use INVX1  _1394_
timestamp 1727493700
transform -1 0 590 0 1 270
box -6 -8 66 272
use OAI21X1  _1395_
timestamp 1727498925
transform -1 0 630 0 -1 790
box -6 -8 106 272
use AND2X2  _1396_
timestamp 1727487319
transform -1 0 750 0 1 270
box -6 -8 106 273
use AOI21X1  _1397_
timestamp 1727487319
transform 1 0 530 0 1 790
box -6 -8 106 272
use NAND3X1  _1398_
timestamp 1727494898
transform 1 0 370 0 1 790
box -6 -8 106 272
use AND2X2  _1399_
timestamp 1727487319
transform 1 0 690 0 1 790
box -6 -8 106 273
use INVX1  _1400_
timestamp 1727493700
transform -1 0 4070 0 1 790
box -6 -8 66 272
use NOR2X1  _1401_
timestamp 1727495070
transform 1 0 4010 0 -1 2350
box -6 -8 86 272
use NOR2X1  _1402_
timestamp 1727495070
transform 1 0 4270 0 -1 2350
box -6 -8 86 272
use NOR2X1  _1403_
timestamp 1727495070
transform 1 0 4150 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1404_
timestamp 1727495070
transform -1 0 4150 0 -1 1310
box -6 -8 86 272
use INVX1  _1405_
timestamp 1727493700
transform -1 0 3850 0 -1 1310
box -6 -8 66 272
use OAI21X1  _1406_
timestamp 1727498925
transform -1 0 3810 0 1 790
box -6 -8 106 272
use OAI21X1  _1407_
timestamp 1727498925
transform 1 0 4130 0 1 790
box -6 -8 106 272
use AOI21X1  _1408_
timestamp 1727487319
transform 1 0 4370 0 -1 1310
box -6 -8 106 272
use NOR2X1  _1409_
timestamp 1727495070
transform 1 0 4510 0 1 1310
box -6 -8 86 272
use NOR2X1  _1410_
timestamp 1727495070
transform 1 0 4650 0 1 1310
box -6 -8 86 272
use NOR2X1  _1411_
timestamp 1727495070
transform 1 0 4530 0 -1 1310
box -6 -8 86 272
use AND2X2  _1412_
timestamp 1727487319
transform 1 0 4810 0 -1 1310
box -6 -8 106 273
use NOR2X1  _1413_
timestamp 1727495070
transform -1 0 4750 0 -1 1310
box -6 -8 86 272
use OAI21X1  _1414_
timestamp 1727498925
transform 1 0 4810 0 1 790
box -6 -8 106 272
use OAI21X1  _1415_
timestamp 1727498925
transform -1 0 4930 0 -1 790
box -6 -8 106 272
use NAND2X1  _1416_
timestamp 1727494699
transform -1 0 3370 0 -1 790
box -6 -8 86 272
use AND2X2  _1417_
timestamp 1727487319
transform -1 0 4310 0 -1 1310
box -6 -8 106 273
use OAI21X1  _1418_
timestamp 1727498925
transform -1 0 4450 0 1 1310
box -6 -8 106 272
use OAI21X1  _1419_
timestamp 1727498925
transform 1 0 4190 0 1 1310
box -6 -8 106 272
use AOI21X1  _1420_
timestamp 1727487319
transform -1 0 4010 0 -1 1310
box -6 -8 106 272
use NOR2X1  _1421_
timestamp 1727495070
transform -1 0 3130 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1422_
timestamp 1727495070
transform -1 0 2990 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1423_
timestamp 1727495070
transform -1 0 2790 0 -1 790
box -6 -8 86 272
use INVX1  _1424_
timestamp 1727493700
transform 1 0 2850 0 -1 790
box -6 -8 66 272
use AND2X2  _1425_
timestamp 1727487319
transform 1 0 2970 0 -1 790
box -6 -8 106 273
use OAI21X1  _1426_
timestamp 1727498925
transform -1 0 3230 0 1 790
box -6 -8 106 272
use OAI21X1  _1427_
timestamp 1727498925
transform 1 0 3130 0 -1 790
box -6 -8 106 272
use INVX1  _1428_
timestamp 1727493700
transform -1 0 2490 0 -1 790
box -6 -8 66 272
use OAI21X1  _1429_
timestamp 1727498925
transform -1 0 2650 0 -1 790
box -6 -8 106 272
use NOR2X1  _1430_
timestamp 1727495070
transform -1 0 2770 0 1 790
box -6 -8 86 272
use NAND2X1  _1431_
timestamp 1727494699
transform 1 0 2750 0 -1 1310
box -6 -8 86 272
use INVX1  _1432_
timestamp 1727493700
transform 1 0 2890 0 -1 1310
box -6 -8 66 272
use NOR2X1  _1433_
timestamp 1727495070
transform 1 0 2830 0 1 790
box -6 -8 86 272
use INVX1  _1434_
timestamp 1727493700
transform -1 0 2630 0 1 790
box -6 -8 66 272
use OR2X2  _1435_
timestamp 1727496117
transform 1 0 2770 0 1 270
box -6 -8 106 272
use AOI21X1  _1436_
timestamp 1727487319
transform 1 0 2610 0 1 270
box -6 -8 106 272
use AOI22X1  _1437_
timestamp 1727487144
transform -1 0 3130 0 -1 270
box -6 -8 126 272
use NAND2X1  _1438_
timestamp 1727494699
transform -1 0 5390 0 1 270
box -6 -8 86 272
use AOI21X1  _1439_
timestamp 1727487319
transform 1 0 2970 0 1 790
box -6 -8 106 272
use NOR2X1  _1440_
timestamp 1727495070
transform 1 0 3290 0 1 790
box -6 -8 86 272
use NAND2X1  _1441_
timestamp 1727494699
transform -1 0 3650 0 1 790
box -6 -8 86 272
use NAND2X1  _1442_
timestamp 1727494699
transform 1 0 3430 0 1 790
box -6 -8 86 272
use NAND2X1  _1443_
timestamp 1727494699
transform -1 0 3950 0 1 790
box -6 -8 86 272
use NOR2X1  _1444_
timestamp 1727495070
transform 1 0 4070 0 -1 790
box -6 -8 86 272
use OR2X2  _1445_
timestamp 1727496117
transform 1 0 4670 0 -1 790
box -6 -8 106 272
use NOR2X1  _1446_
timestamp 1727495070
transform 1 0 5830 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1447_
timestamp 1727495070
transform 1 0 5690 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1448_
timestamp 1727495070
transform -1 0 5870 0 -1 1310
box -6 -8 86 272
use NOR2X1  _1449_
timestamp 1727495070
transform -1 0 5750 0 -1 790
box -6 -8 86 272
use NOR2X1  _1450_
timestamp 1727495070
transform -1 0 4610 0 -1 790
box -6 -8 86 272
use INVX1  _1451_
timestamp 1727493700
transform 1 0 5990 0 1 270
box -6 -8 66 272
use OAI21X1  _1452_
timestamp 1727498925
transform -1 0 5910 0 -1 790
box -6 -8 106 272
use OAI21X1  _1453_
timestamp 1727498925
transform 1 0 5690 0 1 270
box -6 -8 106 272
use INVX1  _1454_
timestamp 1727493700
transform 1 0 5770 0 -1 270
box -6 -8 66 272
use INVX1  _1455_
timestamp 1727493700
transform -1 0 5990 0 -1 1310
box -6 -8 66 272
use OAI21X1  _1456_
timestamp 1727498925
transform 1 0 5870 0 1 790
box -6 -8 106 272
use NOR2X1  _1457_
timestamp 1727495070
transform -1 0 5350 0 -1 2350
box -6 -8 86 272
use NOR2X1  _1458_
timestamp 1727495070
transform -1 0 5450 0 1 1830
box -6 -8 86 272
use NOR2X1  _1459_
timestamp 1727495070
transform 1 0 5990 0 1 4950
box -6 -8 86 272
use INVX1  _1460_
timestamp 1727493700
transform 1 0 5990 0 1 3390
box -6 -8 66 272
use OR2X2  _1461_
timestamp 1727496117
transform 1 0 5890 0 -1 5990
box -6 -8 106 272
use AOI21X1  _1462_
timestamp 1727487319
transform -1 0 5950 0 1 270
box -6 -8 106 272
use AOI22X1  _1463_
timestamp 1727487144
transform 1 0 5890 0 -1 270
box -6 -8 126 272
use NAND2X1  _1464_
timestamp 1727494699
transform -1 0 5050 0 1 790
box -6 -8 86 272
use AOI21X1  _1465_
timestamp 1727487319
transform -1 0 6050 0 1 1310
box -6 -8 106 272
use NOR2X1  _1466_
timestamp 1727495070
transform 1 0 5970 0 -1 790
box -6 -8 86 272
use INVX1  _1467_
timestamp 1727493700
transform 1 0 5750 0 1 790
box -6 -8 66 272
use OAI21X1  _1468_
timestamp 1727498925
transform -1 0 5690 0 1 790
box -6 -8 106 272
use NOR2X1  _1469_
timestamp 1727495070
transform 1 0 5250 0 -1 1310
box -6 -8 86 272
use INVX1  _1470_
timestamp 1727493700
transform 1 0 5670 0 -1 1310
box -6 -8 66 272
use AOI21X1  _1471_
timestamp 1727487319
transform -1 0 5610 0 -1 790
box -6 -8 106 272
use OAI21X1  _1472_
timestamp 1727498925
transform -1 0 5370 0 1 790
box -6 -8 106 272
use OAI21X1  _1473_
timestamp 1727498925
transform -1 0 5210 0 1 790
box -6 -8 106 272
use NAND2X1  _1474_
timestamp 1727494699
transform 1 0 5150 0 -1 270
box -6 -8 86 272
use NAND3X1  _1475_
timestamp 1727494898
transform -1 0 5490 0 -1 1310
box -6 -8 106 272
use OAI21X1  _1476_
timestamp 1727498925
transform 1 0 5430 0 1 790
box -6 -8 106 272
use NAND2X1  _1477_
timestamp 1727494699
transform 1 0 5370 0 -1 790
box -6 -8 86 272
use OAI21X1  _1478_
timestamp 1727498925
transform -1 0 5250 0 1 270
box -6 -8 106 272
use INVX1  _1479_
timestamp 1727493700
transform 1 0 2670 0 -1 1830
box -6 -8 66 272
use NAND3X1  _1480_
timestamp 1727494898
transform 1 0 4210 0 -1 790
box -6 -8 106 272
use NAND2X1  _1481_
timestamp 1727494699
transform 1 0 4010 0 -1 1830
box -6 -8 86 272
use OAI21X1  _1482_
timestamp 1727498925
transform 1 0 3850 0 -1 1830
box -6 -8 106 272
use INVX1  _1483_
timestamp 1727493700
transform 1 0 2890 0 -1 270
box -6 -8 66 272
use NAND2X1  _1484_
timestamp 1727494699
transform 1 0 4450 0 1 1830
box -6 -8 86 272
use OAI21X1  _1485_
timestamp 1727498925
transform 1 0 4050 0 1 1830
box -6 -8 106 272
use INVX1  _1486_
timestamp 1727493700
transform -1 0 3370 0 1 270
box -6 -8 66 272
use NAND2X1  _1487_
timestamp 1727494699
transform -1 0 5030 0 1 1310
box -6 -8 86 272
use OAI21X1  _1488_
timestamp 1727498925
transform 1 0 4790 0 1 1310
box -6 -8 106 272
use INVX1  _1489_
timestamp 1727493700
transform -1 0 3490 0 1 270
box -6 -8 66 272
use NAND2X1  _1490_
timestamp 1727494699
transform -1 0 4910 0 -1 1830
box -6 -8 86 272
use OAI21X1  _1491_
timestamp 1727498925
transform 1 0 4670 0 -1 1830
box -6 -8 106 272
use NOR2X1  _1492_
timestamp 1727495070
transform -1 0 3630 0 1 270
box -6 -8 86 272
use NOR2X1  _1493_
timestamp 1727495070
transform 1 0 3530 0 1 2350
box -6 -8 86 272
use AOI21X1  _1494_
timestamp 1727487319
transform 1 0 3130 0 1 2350
box -6 -8 106 272
use NOR2X1  _1495_
timestamp 1727495070
transform 1 0 3390 0 1 1310
box -6 -8 86 272
use AOI21X1  _1496_
timestamp 1727487319
transform 1 0 2990 0 1 1310
box -6 -8 106 272
use NOR2X1  _1497_
timestamp 1727495070
transform -1 0 3470 0 -1 2350
box -6 -8 86 272
use AOI21X1  _1498_
timestamp 1727487319
transform 1 0 3230 0 -1 2350
box -6 -8 106 272
use NOR2X1  _1499_
timestamp 1727495070
transform 1 0 2850 0 1 1310
box -6 -8 86 272
use AOI21X1  _1500_
timestamp 1727487319
transform -1 0 2790 0 1 1310
box -6 -8 106 272
use INVX1  _1501_
timestamp 1727493700
transform -1 0 2270 0 1 1310
box -6 -8 66 272
use OAI21X1  _1502_
timestamp 1727498925
transform 1 0 2350 0 -1 1830
box -6 -8 106 272
use OAI21X1  _1503_
timestamp 1727498925
transform -1 0 2610 0 -1 1830
box -6 -8 106 272
use OAI21X1  _1504_
timestamp 1727498925
transform -1 0 1890 0 -1 1830
box -6 -8 106 272
use OAI21X1  _1505_
timestamp 1727498925
transform -1 0 2290 0 -1 1830
box -6 -8 106 272
use OAI21X1  _1506_
timestamp 1727498925
transform 1 0 1750 0 1 1310
box -6 -8 106 272
use OAI21X1  _1507_
timestamp 1727498925
transform -1 0 2150 0 1 1310
box -6 -8 106 272
use OAI21X1  _1508_
timestamp 1727498925
transform -1 0 1530 0 1 1310
box -6 -8 106 272
use OAI21X1  _1509_
timestamp 1727498925
transform -1 0 1690 0 1 1310
box -6 -8 106 272
use NOR2X1  _1510_
timestamp 1727495070
transform -1 0 2510 0 1 2350
box -6 -8 86 272
use AOI21X1  _1511_
timestamp 1727487319
transform -1 0 2670 0 1 2350
box -6 -8 106 272
use NOR2X1  _1512_
timestamp 1727495070
transform -1 0 2390 0 -1 2350
box -6 -8 86 272
use AOI21X1  _1513_
timestamp 1727487319
transform 1 0 2410 0 1 1830
box -6 -8 106 272
use NOR2X1  _1514_
timestamp 1727495070
transform -1 0 2770 0 -1 2350
box -6 -8 86 272
use AOI21X1  _1515_
timestamp 1727487319
transform -1 0 2930 0 -1 2350
box -6 -8 106 272
use NOR2X1  _1516_
timestamp 1727495070
transform -1 0 1690 0 1 1830
box -6 -8 86 272
use AOI21X1  _1517_
timestamp 1727487319
transform -1 0 2090 0 1 1830
box -6 -8 106 272
use NAND2X1  _1518_
timestamp 1727494699
transform -1 0 1410 0 1 3390
box -6 -8 86 272
use OAI21X1  _1519_
timestamp 1727498925
transform 1 0 1170 0 1 3390
box -6 -8 106 272
use NAND2X1  _1520_
timestamp 1727494699
transform 1 0 970 0 -1 3910
box -6 -8 86 272
use OAI21X1  _1521_
timestamp 1727498925
transform -1 0 1010 0 1 3910
box -6 -8 106 272
use NAND2X1  _1522_
timestamp 1727494699
transform -1 0 450 0 1 3910
box -6 -8 86 272
use OAI21X1  _1523_
timestamp 1727498925
transform -1 0 610 0 1 3910
box -6 -8 106 272
use NAND2X1  _1524_
timestamp 1727494699
transform 1 0 1470 0 1 3910
box -6 -8 86 272
use OAI21X1  _1525_
timestamp 1727498925
transform -1 0 1410 0 1 3910
box -6 -8 106 272
use DFFPOSX1  _1526_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727503886
transform 1 0 2790 0 1 3910
box -6 -8 246 272
use DFFPOSX1  _1527_
timestamp 1727503886
transform 1 0 2490 0 -1 4430
box -6 -8 246 272
use DFFPOSX1  _1528_
timestamp 1727503886
transform 1 0 3350 0 1 3910
box -6 -8 246 272
use DFFPOSX1  _1529_
timestamp 1727503886
transform 1 0 3470 0 -1 4430
box -6 -8 246 272
use DFFPOSX1  _1530_
timestamp 1727503886
transform -1 0 2150 0 -1 3390
box -6 -8 246 272
use DFFPOSX1  _1531_
timestamp 1727503886
transform 1 0 1170 0 -1 2350
box -6 -8 246 272
use DFFPOSX1  _1532_
timestamp 1727503886
transform -1 0 1170 0 -1 2870
box -6 -8 246 272
use DFFPOSX1  _1533_
timestamp 1727503886
transform -1 0 1010 0 -1 2350
box -6 -8 246 272
use DFFPOSX1  _1534_
timestamp 1727503886
transform -1 0 510 0 -1 1830
box -6 -8 246 272
use DFFPOSX1  _1535_
timestamp 1727503886
transform -1 0 1170 0 -1 1830
box -6 -8 246 272
use DFFPOSX1  _1536_
timestamp 1727503886
transform -1 0 1290 0 -1 790
box -6 -8 246 272
use DFFPOSX1  _1537_
timestamp 1727503886
transform -1 0 830 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1538_
timestamp 1727503886
transform 1 0 3710 0 -1 2350
box -6 -8 246 272
use DFFPOSX1  _1539_
timestamp 1727503886
transform 1 0 3770 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1540_
timestamp 1727503886
transform -1 0 3730 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1541_
timestamp 1727503886
transform 1 0 1990 0 1 790
box -6 -8 246 272
use DFFPOSX1  _1542_
timestamp 1727503886
transform 1 0 5450 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1543_
timestamp 1727503886
transform 1 0 4850 0 -1 2350
box -6 -8 246 272
use DFFPOSX1  _1544_
timestamp 1727503886
transform 1 0 5650 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1545_
timestamp 1727503886
transform -1 0 5650 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1546_
timestamp 1727503886
transform 1 0 1430 0 -1 3390
box -6 -8 246 272
use DFFPOSX1  _1547_
timestamp 1727503886
transform 1 0 1410 0 -1 2870
box -6 -8 246 272
use DFFPOSX1  _1548_
timestamp 1727503886
transform 1 0 430 0 -1 2870
box -6 -8 246 272
use DFFPOSX1  _1549_
timestamp 1727503886
transform 1 0 250 0 1 2350
box -6 -8 246 272
use DFFPOSX1  _1550_
timestamp 1727503886
transform -1 0 250 0 1 2350
box -6 -8 246 272
use DFFPOSX1  _1551_
timestamp 1727503886
transform -1 0 1250 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1552_
timestamp 1727503886
transform -1 0 1410 0 -1 2870
box -6 -8 246 272
use DFFPOSX1  _1553_
timestamp 1727503886
transform -1 0 1190 0 -1 1310
box -6 -8 246 272
use DFFPOSX1  _1554_
timestamp 1727503886
transform -1 0 4270 0 1 2350
box -6 -8 246 272
use DFFPOSX1  _1555_
timestamp 1727503886
transform -1 0 4770 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1556_
timestamp 1727503886
transform 1 0 2930 0 -1 2350
box -6 -8 246 272
use DFFPOSX1  _1557_
timestamp 1727503886
transform -1 0 3730 0 -1 1310
box -6 -8 246 272
use DFFPOSX1  _1558_
timestamp 1727503886
transform 1 0 5790 0 1 2350
box -6 -8 246 272
use DFFPOSX1  _1559_
timestamp 1727503886
transform 1 0 4910 0 1 2350
box -6 -8 246 272
use DFFPOSX1  _1560_
timestamp 1727503886
transform 1 0 1750 0 1 790
box -6 -8 246 272
use DFFPOSX1  _1561_
timestamp 1727503886
transform -1 0 2830 0 -1 270
box -6 -8 246 272
use DFFPOSX1  _1562_
timestamp 1727503886
transform 1 0 1850 0 1 270
box -6 -8 246 272
use DFFPOSX1  _1563_
timestamp 1727503886
transform 1 0 1470 0 1 270
box -6 -8 246 272
use DFFPOSX1  _1564_
timestamp 1727503886
transform 1 0 1510 0 1 790
box -6 -8 246 272
use DFFPOSX1  _1565_
timestamp 1727503886
transform -1 0 530 0 -1 270
box -6 -8 246 272
use DFFPOSX1  _1566_
timestamp 1727503886
transform 1 0 1010 0 -1 270
box -6 -8 246 272
use DFFPOSX1  _1567_
timestamp 1727503886
transform 1 0 1550 0 -1 270
box -6 -8 246 272
use DFFPOSX1  _1568_
timestamp 1727503886
transform -1 0 4610 0 1 790
box -6 -8 246 272
use DFFPOSX1  _1569_
timestamp 1727503886
transform 1 0 4450 0 1 270
box -6 -8 246 272
use DFFPOSX1  _1570_
timestamp 1727503886
transform 1 0 3370 0 -1 790
box -6 -8 246 272
use DFFPOSX1  _1571_
timestamp 1727503886
transform 1 0 3130 0 -1 270
box -6 -8 246 272
use DFFPOSX1  _1572_
timestamp 1727503886
transform -1 0 5630 0 1 270
box -6 -8 246 272
use DFFPOSX1  _1573_
timestamp 1727503886
transform -1 0 5710 0 -1 270
box -6 -8 246 272
use DFFPOSX1  _1574_
timestamp 1727503886
transform -1 0 5310 0 -1 790
box -6 -8 246 272
use DFFPOSX1  _1575_
timestamp 1727503886
transform -1 0 5470 0 -1 270
box -6 -8 246 272
use DFFPOSX1  _1576_
timestamp 1727503886
transform 1 0 3550 0 -1 1830
box -6 -8 246 272
use DFFPOSX1  _1577_
timestamp 1727503886
transform 1 0 4150 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1578_
timestamp 1727503886
transform -1 0 5410 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1579_
timestamp 1727503886
transform 1 0 4910 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1580_
timestamp 1727503886
transform 1 0 3230 0 1 2350
box -6 -8 246 272
use DFFPOSX1  _1581_
timestamp 1727503886
transform 1 0 3090 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1582_
timestamp 1727503886
transform -1 0 3710 0 -1 2350
box -6 -8 246 272
use DFFPOSX1  _1583_
timestamp 1727503886
transform -1 0 2630 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1584_
timestamp 1727503886
transform -1 0 2990 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1585_
timestamp 1727503886
transform -1 0 2130 0 -1 1830
box -6 -8 246 272
use DFFPOSX1  _1586_
timestamp 1727503886
transform -1 0 2130 0 -1 1310
box -6 -8 246 272
use DFFPOSX1  _1587_
timestamp 1727503886
transform -1 0 1370 0 1 1310
box -6 -8 246 272
use DFFPOSX1  _1588_
timestamp 1727503886
transform -1 0 2630 0 -1 2350
box -6 -8 246 272
use DFFPOSX1  _1589_
timestamp 1727503886
transform 1 0 2510 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1590_
timestamp 1727503886
transform -1 0 2910 0 1 2350
box -6 -8 246 272
use DFFPOSX1  _1591_
timestamp 1727503886
transform -1 0 1930 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1592_
timestamp 1727503886
transform 1 0 870 0 1 3390
box -6 -8 246 272
use DFFPOSX1  _1593_
timestamp 1727503886
transform -1 0 850 0 1 3910
box -6 -8 246 272
use DFFPOSX1  _1594_
timestamp 1727503886
transform 1 0 910 0 -1 4430
box -6 -8 246 272
use DFFPOSX1  _1595_
timestamp 1727503886
transform 1 0 1010 0 1 3910
box -6 -8 246 272
use DFFPOSX1  _1596_
timestamp 1727503886
transform 1 0 10 0 -1 2870
box -6 -8 246 272
use DFFPOSX1  _1597_
timestamp 1727503886
transform -1 0 3350 0 1 1830
box -6 -8 246 272
use DFFPOSX1  _1598_
timestamp 1727503886
transform 1 0 2870 0 1 270
box -6 -8 246 272
use DFFPOSX1  _1599_
timestamp 1727503886
transform 1 0 3750 0 1 270
box -6 -8 246 272
use DFFPOSX1  _1600_
timestamp 1727503886
transform 1 0 3770 0 -1 790
box -6 -8 246 272
use BUFX2  _1601_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487319
transform 1 0 5970 0 -1 1830
box -6 -8 86 272
use BUFX2  _1602_
timestamp 1727487319
transform 1 0 5990 0 -1 3910
box -6 -8 86 272
use BUFX2  _1603_
timestamp 1727487319
transform 1 0 5650 0 -1 4950
box -6 -8 86 272
use BUFX2  _1604_
timestamp 1727487319
transform 1 0 5550 0 1 4950
box -6 -8 86 272
use BUFX2  _1605_
timestamp 1727487319
transform 1 0 5850 0 1 4950
box -6 -8 86 272
use BUFX2  _1606_
timestamp 1727487319
transform 1 0 4430 0 -1 270
box -6 -8 86 272
use BUFX2  _1607_
timestamp 1727487319
transform 1 0 4570 0 -1 270
box -6 -8 86 272
use BUFX2  _1608_
timestamp 1727487319
transform 1 0 4710 0 -1 270
box -6 -8 86 272
use BUFX2  _1609_
timestamp 1727487319
transform 1 0 4290 0 -1 270
box -6 -8 86 272
use BUFX2  BUFX2_insert0
timestamp 1727487319
transform -1 0 1890 0 -1 1310
box -6 -8 86 272
use BUFX2  BUFX2_insert1
timestamp 1727487319
transform -1 0 1650 0 1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert2
timestamp 1727487319
transform 1 0 4990 0 -1 790
box -6 -8 86 272
use BUFX2  BUFX2_insert3
timestamp 1727487319
transform 1 0 3470 0 -1 1830
box -6 -8 86 272
use BUFX2  BUFX2_insert4
timestamp 1727487319
transform 1 0 2230 0 -1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert5
timestamp 1727487319
transform 1 0 1750 0 -1 2350
box -6 -8 86 272
use BUFX2  BUFX2_insert6
timestamp 1727487319
transform -1 0 3170 0 -1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert7
timestamp 1727487319
transform -1 0 4630 0 1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert16
timestamp 1727487319
transform -1 0 2190 0 -1 790
box -6 -8 86 272
use BUFX2  BUFX2_insert17
timestamp 1727487319
transform 1 0 2330 0 1 270
box -6 -8 86 272
use BUFX2  BUFX2_insert18
timestamp 1727487319
transform 1 0 2470 0 1 270
box -6 -8 86 272
use BUFX2  BUFX2_insert19
timestamp 1727487319
transform 1 0 5010 0 1 270
box -6 -8 86 272
use BUFX2  BUFX2_insert20
timestamp 1727487319
transform -1 0 4750 0 1 790
box -6 -8 86 272
use BUFX2  BUFX2_insert21
timestamp 1727487319
transform 1 0 4070 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert22
timestamp 1727487319
transform -1 0 1670 0 -1 5470
box -6 -8 86 272
use BUFX2  BUFX2_insert23
timestamp 1727487319
transform 1 0 3010 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert24
timestamp 1727487319
transform -1 0 2330 0 1 5470
box -6 -8 86 272
use BUFX2  BUFX2_insert25
timestamp 1727487319
transform 1 0 2950 0 -1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert26
timestamp 1727487319
transform -1 0 2690 0 1 3390
box -6 -8 86 272
use BUFX2  BUFX2_insert27
timestamp 1727487319
transform 1 0 790 0 1 3390
box -6 -8 86 272
use BUFX2  BUFX2_insert28
timestamp 1727487319
transform -1 0 2110 0 -1 2350
box -6 -8 86 272
use BUFX2  BUFX2_insert29
timestamp 1727487319
transform -1 0 2250 0 -1 2350
box -6 -8 86 272
use BUFX2  BUFX2_insert30
timestamp 1727487319
transform -1 0 1950 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert31
timestamp 1727487319
transform 1 0 2010 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert32
timestamp 1727487319
transform 1 0 4650 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert33
timestamp 1727487319
transform -1 0 4470 0 -1 5990
box -6 -8 86 272
use CLKBUF1  CLKBUF1_insert8 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727490190
transform 1 0 3010 0 -1 1310
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert9
timestamp 1727490190
transform -1 0 1310 0 -1 3390
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert10
timestamp 1727490190
transform -1 0 2690 0 -1 1310
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert11
timestamp 1727490190
transform 1 0 5750 0 1 1830
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert12
timestamp 1727490190
transform -1 0 3990 0 1 1830
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert13
timestamp 1727490190
transform 1 0 4290 0 -1 1830
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert14
timestamp 1727490190
transform -1 0 2350 0 1 1830
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert15
timestamp 1727490190
transform -1 0 1610 0 -1 1310
box -6 -8 206 272
use FILL  FILL89250x27450 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727493435
transform 1 0 5950 0 1 1830
box -6 -8 26 272
use FILL  FILL89550x11850
timestamp 1727493435
transform 1 0 5970 0 1 790
box -6 -8 26 272
use FILL  FILL89550x27450
timestamp 1727493435
transform 1 0 5970 0 1 1830
box -6 -8 26 272
use FILL  FILL89850x11850
timestamp 1727493435
transform 1 0 5990 0 1 790
box -6 -8 26 272
use FILL  FILL89850x15750
timestamp 1727493435
transform -1 0 6010 0 -1 1310
box -6 -8 26 272
use FILL  FILL89850x27450
timestamp 1727493435
transform 1 0 5990 0 1 1830
box -6 -8 26 272
use FILL  FILL89850x78150
timestamp 1727493435
transform -1 0 6010 0 -1 5470
box -6 -8 26 272
use FILL  FILL89850x85950
timestamp 1727493435
transform -1 0 6010 0 -1 5990
box -6 -8 26 272
use FILL  FILL90150x150
timestamp 1727493435
transform -1 0 6030 0 -1 270
box -6 -8 26 272
use FILL  FILL90150x11850
timestamp 1727493435
transform 1 0 6010 0 1 790
box -6 -8 26 272
use FILL  FILL90150x15750
timestamp 1727493435
transform -1 0 6030 0 -1 1310
box -6 -8 26 272
use FILL  FILL90150x27450
timestamp 1727493435
transform 1 0 6010 0 1 1830
box -6 -8 26 272
use FILL  FILL90150x39150
timestamp 1727493435
transform -1 0 6030 0 -1 2870
box -6 -8 26 272
use FILL  FILL90150x62550
timestamp 1727493435
transform -1 0 6030 0 -1 4430
box -6 -8 26 272
use FILL  FILL90150x78150
timestamp 1727493435
transform -1 0 6030 0 -1 5470
box -6 -8 26 272
use FILL  FILL90150x85950
timestamp 1727493435
transform -1 0 6030 0 -1 5990
box -6 -8 26 272
use FILL  FILL90450x150
timestamp 1727493435
transform -1 0 6050 0 -1 270
box -6 -8 26 272
use FILL  FILL90450x11850
timestamp 1727493435
transform 1 0 6030 0 1 790
box -6 -8 26 272
use FILL  FILL90450x15750
timestamp 1727493435
transform -1 0 6050 0 -1 1310
box -6 -8 26 272
use FILL  FILL90450x27450
timestamp 1727493435
transform 1 0 6030 0 1 1830
box -6 -8 26 272
use FILL  FILL90450x31350
timestamp 1727493435
transform -1 0 6050 0 -1 2350
box -6 -8 26 272
use FILL  FILL90450x35250
timestamp 1727493435
transform 1 0 6030 0 1 2350
box -6 -8 26 272
use FILL  FILL90450x39150
timestamp 1727493435
transform -1 0 6050 0 -1 2870
box -6 -8 26 272
use FILL  FILL90450x46950
timestamp 1727493435
transform -1 0 6050 0 -1 3390
box -6 -8 26 272
use FILL  FILL90450x62550
timestamp 1727493435
transform -1 0 6050 0 -1 4430
box -6 -8 26 272
use FILL  FILL90450x66450
timestamp 1727493435
transform 1 0 6030 0 1 4430
box -6 -8 26 272
use FILL  FILL90450x70350
timestamp 1727493435
transform -1 0 6050 0 -1 4950
box -6 -8 26 272
use FILL  FILL90450x78150
timestamp 1727493435
transform -1 0 6050 0 -1 5470
box -6 -8 26 272
use FILL  FILL90450x85950
timestamp 1727493435
transform -1 0 6050 0 -1 5990
box -6 -8 26 272
use FILL  FILL90750x150
timestamp 1727493435
transform -1 0 6070 0 -1 270
box -6 -8 26 272
use FILL  FILL90750x4050
timestamp 1727493435
transform 1 0 6050 0 1 270
box -6 -8 26 272
use FILL  FILL90750x7950
timestamp 1727493435
transform -1 0 6070 0 -1 790
box -6 -8 26 272
use FILL  FILL90750x11850
timestamp 1727493435
transform 1 0 6050 0 1 790
box -6 -8 26 272
use FILL  FILL90750x15750
timestamp 1727493435
transform -1 0 6070 0 -1 1310
box -6 -8 26 272
use FILL  FILL90750x19650
timestamp 1727493435
transform 1 0 6050 0 1 1310
box -6 -8 26 272
use FILL  FILL90750x23550
timestamp 1727493435
transform -1 0 6070 0 -1 1830
box -6 -8 26 272
use FILL  FILL90750x27450
timestamp 1727493435
transform 1 0 6050 0 1 1830
box -6 -8 26 272
use FILL  FILL90750x31350
timestamp 1727493435
transform -1 0 6070 0 -1 2350
box -6 -8 26 272
use FILL  FILL90750x35250
timestamp 1727493435
transform 1 0 6050 0 1 2350
box -6 -8 26 272
use FILL  FILL90750x39150
timestamp 1727493435
transform -1 0 6070 0 -1 2870
box -6 -8 26 272
use FILL  FILL90750x43050
timestamp 1727493435
transform 1 0 6050 0 1 2870
box -6 -8 26 272
use FILL  FILL90750x46950
timestamp 1727493435
transform -1 0 6070 0 -1 3390
box -6 -8 26 272
use FILL  FILL90750x50850
timestamp 1727493435
transform 1 0 6050 0 1 3390
box -6 -8 26 272
use FILL  FILL90750x58650
timestamp 1727493435
transform 1 0 6050 0 1 3910
box -6 -8 26 272
use FILL  FILL90750x62550
timestamp 1727493435
transform -1 0 6070 0 -1 4430
box -6 -8 26 272
use FILL  FILL90750x66450
timestamp 1727493435
transform 1 0 6050 0 1 4430
box -6 -8 26 272
use FILL  FILL90750x70350
timestamp 1727493435
transform -1 0 6070 0 -1 4950
box -6 -8 26 272
use FILL  FILL90750x78150
timestamp 1727493435
transform -1 0 6070 0 -1 5470
box -6 -8 26 272
use FILL  FILL90750x85950
timestamp 1727493435
transform -1 0 6070 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__760_
timestamp 1727493435
transform 1 0 4810 0 1 270
box -6 -8 26 272
use FILL  FILL_0__761_
timestamp 1727493435
transform 1 0 3630 0 1 270
box -6 -8 26 272
use FILL  FILL_0__762_
timestamp 1727493435
transform 1 0 3110 0 1 270
box -6 -8 26 272
use FILL  FILL_0__763_
timestamp 1727493435
transform 1 0 4310 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__764_
timestamp 1727493435
transform -1 0 2750 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__765_
timestamp 1727493435
transform -1 0 1870 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__766_
timestamp 1727493435
transform -1 0 1890 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__767_
timestamp 1727493435
transform -1 0 4310 0 1 270
box -6 -8 26 272
use FILL  FILL_0__768_
timestamp 1727493435
transform 1 0 3950 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__769_
timestamp 1727493435
transform 1 0 4690 0 1 270
box -6 -8 26 272
use FILL  FILL_0__770_
timestamp 1727493435
transform -1 0 4810 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__771_
timestamp 1727493435
transform -1 0 4950 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__772_
timestamp 1727493435
transform -1 0 2130 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__773_
timestamp 1727493435
transform -1 0 4090 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__774_
timestamp 1727493435
transform 1 0 4150 0 1 270
box -6 -8 26 272
use FILL  FILL_0__775_
timestamp 1727493435
transform 1 0 3610 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__776_
timestamp 1727493435
transform 1 0 2090 0 1 270
box -6 -8 26 272
use FILL  FILL_0__777_
timestamp 1727493435
transform -1 0 4010 0 1 270
box -6 -8 26 272
use FILL  FILL_0__778_
timestamp 1727493435
transform 1 0 3370 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__779_
timestamp 1727493435
transform -1 0 3510 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__780_
timestamp 1727493435
transform -1 0 3810 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__781_
timestamp 1727493435
transform 1 0 1930 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__782_
timestamp 1727493435
transform -1 0 3650 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__783_
timestamp 1727493435
transform -1 0 3390 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__784_
timestamp 1727493435
transform -1 0 2530 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__785_
timestamp 1727493435
transform -1 0 4330 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__786_
timestamp 1727493435
transform -1 0 3150 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__787_
timestamp 1727493435
transform -1 0 4490 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__788_
timestamp 1727493435
transform 1 0 4610 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__789_
timestamp 1727493435
transform -1 0 3450 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__790_
timestamp 1727493435
transform -1 0 4050 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__791_
timestamp 1727493435
transform -1 0 4190 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__792_
timestamp 1727493435
transform -1 0 5370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__793_
timestamp 1727493435
transform -1 0 4190 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__794_
timestamp 1727493435
transform -1 0 4330 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__795_
timestamp 1727493435
transform 1 0 2650 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__796_
timestamp 1727493435
transform -1 0 2810 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__797_
timestamp 1727493435
transform 1 0 1610 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__798_
timestamp 1727493435
transform -1 0 2350 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__799_
timestamp 1727493435
transform 1 0 1690 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__800_
timestamp 1727493435
transform -1 0 3210 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__801_
timestamp 1727493435
transform 1 0 1550 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__802_
timestamp 1727493435
transform -1 0 3330 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__803_
timestamp 1727493435
transform -1 0 1810 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__804_
timestamp 1727493435
transform -1 0 2330 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__805_
timestamp 1727493435
transform 1 0 2110 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__806_
timestamp 1727493435
transform 1 0 1410 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__807_
timestamp 1727493435
transform 1 0 1830 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__808_
timestamp 1727493435
transform 1 0 1530 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__809_
timestamp 1727493435
transform 1 0 910 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__810_
timestamp 1727493435
transform 1 0 2450 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__811_
timestamp 1727493435
transform 1 0 1030 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__812_
timestamp 1727493435
transform -1 0 670 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__813_
timestamp 1727493435
transform 1 0 1410 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__814_
timestamp 1727493435
transform -1 0 1030 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__815_
timestamp 1727493435
transform -1 0 170 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__816_
timestamp 1727493435
transform -1 0 1470 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__817_
timestamp 1727493435
transform 1 0 510 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__818_
timestamp 1727493435
transform -1 0 830 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__819_
timestamp 1727493435
transform 1 0 1590 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__820_
timestamp 1727493435
transform 1 0 1170 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__821_
timestamp 1727493435
transform 1 0 1070 0 1 790
box -6 -8 26 272
use FILL  FILL_0__822_
timestamp 1727493435
transform -1 0 1630 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__823_
timestamp 1727493435
transform 1 0 1190 0 1 790
box -6 -8 26 272
use FILL  FILL_0__824_
timestamp 1727493435
transform 1 0 710 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__825_
timestamp 1727493435
transform 1 0 990 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__826_
timestamp 1727493435
transform 1 0 830 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__827_
timestamp 1727493435
transform 1 0 3910 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__828_
timestamp 1727493435
transform -1 0 3630 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__829_
timestamp 1727493435
transform -1 0 3770 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__830_
timestamp 1727493435
transform 1 0 4010 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__831_
timestamp 1727493435
transform -1 0 3490 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__832_
timestamp 1727493435
transform -1 0 3630 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__833_
timestamp 1727493435
transform 1 0 3130 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__834_
timestamp 1727493435
transform 1 0 3350 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__835_
timestamp 1727493435
transform 1 0 3250 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__836_
timestamp 1727493435
transform 1 0 2390 0 1 790
box -6 -8 26 272
use FILL  FILL_0__837_
timestamp 1727493435
transform 1 0 2270 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__838_
timestamp 1727493435
transform -1 0 2250 0 1 790
box -6 -8 26 272
use FILL  FILL_0__839_
timestamp 1727493435
transform -1 0 5530 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__840_
timestamp 1727493435
transform -1 0 4930 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__841_
timestamp 1727493435
transform -1 0 5370 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__842_
timestamp 1727493435
transform 1 0 5350 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__843_
timestamp 1727493435
transform 1 0 4770 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__844_
timestamp 1727493435
transform -1 0 5170 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__845_
timestamp 1727493435
transform -1 0 4930 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__846_
timestamp 1727493435
transform 1 0 5030 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__847_
timestamp 1727493435
transform -1 0 5050 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__848_
timestamp 1727493435
transform 1 0 5490 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__849_
timestamp 1727493435
transform -1 0 5070 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__850_
timestamp 1727493435
transform 1 0 5190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__851_
timestamp 1727493435
transform 1 0 1670 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__852_
timestamp 1727493435
transform -1 0 1470 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__853_
timestamp 1727493435
transform -1 0 1430 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__854_
timestamp 1727493435
transform 1 0 1650 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__855_
timestamp 1727493435
transform -1 0 1090 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__856_
timestamp 1727493435
transform 1 0 1290 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__857_
timestamp 1727493435
transform 1 0 1150 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__858_
timestamp 1727493435
transform 1 0 1170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__859_
timestamp 1727493435
transform -1 0 1070 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__860_
timestamp 1727493435
transform -1 0 4310 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__861_
timestamp 1727493435
transform -1 0 1230 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__862_
timestamp 1727493435
transform -1 0 1310 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__863_
timestamp 1727493435
transform -1 0 1370 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__864_
timestamp 1727493435
transform -1 0 690 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__865_
timestamp 1727493435
transform 1 0 1470 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__866_
timestamp 1727493435
transform -1 0 1250 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__867_
timestamp 1727493435
transform 1 0 1210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__868_
timestamp 1727493435
transform 1 0 890 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__869_
timestamp 1727493435
transform 1 0 730 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__870_
timestamp 1727493435
transform 1 0 1350 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__871_
timestamp 1727493435
transform -1 0 1390 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__872_
timestamp 1727493435
transform -1 0 950 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__873_
timestamp 1727493435
transform -1 0 470 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__874_
timestamp 1727493435
transform -1 0 590 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__875_
timestamp 1727493435
transform 1 0 750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__876_
timestamp 1727493435
transform -1 0 350 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__877_
timestamp 1727493435
transform -1 0 610 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__878_
timestamp 1727493435
transform -1 0 470 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__879_
timestamp 1727493435
transform -1 0 490 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__880_
timestamp 1727493435
transform -1 0 630 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__881_
timestamp 1727493435
transform -1 0 510 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__882_
timestamp 1727493435
transform 1 0 1770 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__883_
timestamp 1727493435
transform 1 0 1050 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__884_
timestamp 1727493435
transform 1 0 1250 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__885_
timestamp 1727493435
transform 1 0 1530 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__886_
timestamp 1727493435
transform 1 0 1250 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__887_
timestamp 1727493435
transform 1 0 1670 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__888_
timestamp 1727493435
transform -1 0 1110 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__889_
timestamp 1727493435
transform -1 0 830 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__890_
timestamp 1727493435
transform -1 0 1870 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__891_
timestamp 1727493435
transform -1 0 950 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__892_
timestamp 1727493435
transform -1 0 830 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__893_
timestamp 1727493435
transform -1 0 510 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__894_
timestamp 1727493435
transform -1 0 470 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__895_
timestamp 1727493435
transform 1 0 890 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__896_
timestamp 1727493435
transform -1 0 670 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__897_
timestamp 1727493435
transform -1 0 1570 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__898_
timestamp 1727493435
transform -1 0 1090 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__899_
timestamp 1727493435
transform 1 0 2950 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__900_
timestamp 1727493435
transform 1 0 3130 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__901_
timestamp 1727493435
transform -1 0 1410 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__902_
timestamp 1727493435
transform -1 0 1110 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__903_
timestamp 1727493435
transform 1 0 730 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__904_
timestamp 1727493435
transform -1 0 310 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__905_
timestamp 1727493435
transform -1 0 30 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__906_
timestamp 1727493435
transform -1 0 630 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__907_
timestamp 1727493435
transform -1 0 590 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__908_
timestamp 1727493435
transform -1 0 150 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__909_
timestamp 1727493435
transform 1 0 170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__910_
timestamp 1727493435
transform -1 0 30 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__911_
timestamp 1727493435
transform -1 0 350 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__912_
timestamp 1727493435
transform -1 0 270 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__913_
timestamp 1727493435
transform 1 0 10 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__914_
timestamp 1727493435
transform 1 0 330 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__915_
timestamp 1727493435
transform 1 0 770 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__916_
timestamp 1727493435
transform -1 0 310 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__917_
timestamp 1727493435
transform 1 0 930 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__918_
timestamp 1727493435
transform 1 0 2230 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__919_
timestamp 1727493435
transform 1 0 1670 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__920_
timestamp 1727493435
transform -1 0 2030 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__921_
timestamp 1727493435
transform 1 0 1090 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__922_
timestamp 1727493435
transform -1 0 1390 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__923_
timestamp 1727493435
transform 1 0 970 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__924_
timestamp 1727493435
transform -1 0 510 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__925_
timestamp 1727493435
transform -1 0 2110 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__926_
timestamp 1727493435
transform 1 0 1390 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__927_
timestamp 1727493435
transform -1 0 670 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__928_
timestamp 1727493435
transform 1 0 490 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__929_
timestamp 1727493435
transform -1 0 670 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__930_
timestamp 1727493435
transform -1 0 350 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__931_
timestamp 1727493435
transform -1 0 830 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__932_
timestamp 1727493435
transform 1 0 170 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__933_
timestamp 1727493435
transform 1 0 2070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__934_
timestamp 1727493435
transform -1 0 3270 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__935_
timestamp 1727493435
transform 1 0 1530 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__936_
timestamp 1727493435
transform 1 0 1370 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__937_
timestamp 1727493435
transform -1 0 1630 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__938_
timestamp 1727493435
transform -1 0 190 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__939_
timestamp 1727493435
transform -1 0 30 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__940_
timestamp 1727493435
transform -1 0 350 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__941_
timestamp 1727493435
transform -1 0 30 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__942_
timestamp 1727493435
transform -1 0 30 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__943_
timestamp 1727493435
transform 1 0 130 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__944_
timestamp 1727493435
transform -1 0 470 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__945_
timestamp 1727493435
transform 1 0 290 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__946_
timestamp 1727493435
transform -1 0 30 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__947_
timestamp 1727493435
transform -1 0 30 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__948_
timestamp 1727493435
transform 1 0 130 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__949_
timestamp 1727493435
transform -1 0 30 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__950_
timestamp 1727493435
transform 1 0 170 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__951_
timestamp 1727493435
transform 1 0 190 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__952_
timestamp 1727493435
transform -1 0 30 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__953_
timestamp 1727493435
transform 1 0 890 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__954_
timestamp 1727493435
transform 1 0 1830 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__955_
timestamp 1727493435
transform -1 0 30 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__956_
timestamp 1727493435
transform -1 0 30 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__957_
timestamp 1727493435
transform 1 0 170 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__958_
timestamp 1727493435
transform 1 0 2410 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__959_
timestamp 1727493435
transform -1 0 1450 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__960_
timestamp 1727493435
transform 1 0 1710 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__961_
timestamp 1727493435
transform -1 0 1570 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__962_
timestamp 1727493435
transform 1 0 3970 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__963_
timestamp 1727493435
transform -1 0 2030 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__964_
timestamp 1727493435
transform 1 0 1790 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__965_
timestamp 1727493435
transform -1 0 1690 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__966_
timestamp 1727493435
transform -1 0 1890 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__967_
timestamp 1727493435
transform -1 0 1930 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__968_
timestamp 1727493435
transform 1 0 1950 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__969_
timestamp 1727493435
transform 1 0 2210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__970_
timestamp 1727493435
transform 1 0 1210 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__971_
timestamp 1727493435
transform 1 0 3250 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__972_
timestamp 1727493435
transform -1 0 3110 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__973_
timestamp 1727493435
transform 1 0 2650 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__974_
timestamp 1727493435
transform 1 0 2810 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__975_
timestamp 1727493435
transform -1 0 2410 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__976_
timestamp 1727493435
transform -1 0 2510 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__977_
timestamp 1727493435
transform -1 0 2490 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__978_
timestamp 1727493435
transform 1 0 2530 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__979_
timestamp 1727493435
transform -1 0 2810 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__980_
timestamp 1727493435
transform -1 0 2330 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__981_
timestamp 1727493435
transform -1 0 1690 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__982_
timestamp 1727493435
transform 1 0 1510 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__983_
timestamp 1727493435
transform -1 0 2170 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__984_
timestamp 1727493435
transform -1 0 2350 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__985_
timestamp 1727493435
transform -1 0 1850 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__986_
timestamp 1727493435
transform -1 0 1690 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__987_
timestamp 1727493435
transform 1 0 2350 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__988_
timestamp 1727493435
transform 1 0 1990 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__989_
timestamp 1727493435
transform -1 0 2010 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__990_
timestamp 1727493435
transform 1 0 2510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__991_
timestamp 1727493435
transform -1 0 170 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__992_
timestamp 1727493435
transform -1 0 350 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__993_
timestamp 1727493435
transform -1 0 470 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__994_
timestamp 1727493435
transform -1 0 330 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__995_
timestamp 1727493435
transform 1 0 150 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__996_
timestamp 1727493435
transform -1 0 770 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__997_
timestamp 1727493435
transform -1 0 30 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__998_
timestamp 1727493435
transform 1 0 410 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__999_
timestamp 1727493435
transform 1 0 770 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1000_
timestamp 1727493435
transform -1 0 470 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1001_
timestamp 1727493435
transform 1 0 890 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1002_
timestamp 1727493435
transform -1 0 610 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1003_
timestamp 1727493435
transform -1 0 1330 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1004_
timestamp 1727493435
transform -1 0 1210 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1005_
timestamp 1727493435
transform 1 0 1250 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1006_
timestamp 1727493435
transform 1 0 1330 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1007_
timestamp 1727493435
transform -1 0 610 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1008_
timestamp 1727493435
transform 1 0 570 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1009_
timestamp 1727493435
transform 1 0 2270 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1010_
timestamp 1727493435
transform 1 0 2110 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1011_
timestamp 1727493435
transform -1 0 2090 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1012_
timestamp 1727493435
transform 1 0 2830 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1013_
timestamp 1727493435
transform 1 0 2670 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1014_
timestamp 1727493435
transform 1 0 2830 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1015_
timestamp 1727493435
transform -1 0 3550 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1016_
timestamp 1727493435
transform 1 0 2550 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1017_
timestamp 1727493435
transform -1 0 3710 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1018_
timestamp 1727493435
transform 1 0 3370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1019_
timestamp 1727493435
transform 1 0 2970 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1020_
timestamp 1727493435
transform -1 0 2730 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1021_
timestamp 1727493435
transform 1 0 3230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1022_
timestamp 1727493435
transform 1 0 2170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1023_
timestamp 1727493435
transform 1 0 2730 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1024_
timestamp 1727493435
transform 1 0 3050 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1025_
timestamp 1727493435
transform -1 0 2690 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1026_
timestamp 1727493435
transform 1 0 2590 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1027_
timestamp 1727493435
transform 1 0 3570 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1028_
timestamp 1727493435
transform -1 0 4150 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1029_
timestamp 1727493435
transform 1 0 3970 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1030_
timestamp 1727493435
transform -1 0 3890 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1031_
timestamp 1727493435
transform -1 0 3730 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1032_
timestamp 1727493435
transform -1 0 3430 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1033_
timestamp 1727493435
transform -1 0 3570 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1034_
timestamp 1727493435
transform 1 0 5070 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1035_
timestamp 1727493435
transform 1 0 3670 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1036_
timestamp 1727493435
transform 1 0 3810 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1037_
timestamp 1727493435
transform -1 0 3090 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1038_
timestamp 1727493435
transform -1 0 2650 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1039_
timestamp 1727493435
transform 1 0 2950 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1040_
timestamp 1727493435
transform -1 0 2770 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1041_
timestamp 1727493435
transform -1 0 3410 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1042_
timestamp 1727493435
transform -1 0 3270 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1043_
timestamp 1727493435
transform -1 0 2930 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1044_
timestamp 1727493435
transform -1 0 2490 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1045_
timestamp 1727493435
transform -1 0 2910 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1046_
timestamp 1727493435
transform 1 0 2790 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1047_
timestamp 1727493435
transform 1 0 2950 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1048_
timestamp 1727493435
transform -1 0 2490 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1049_
timestamp 1727493435
transform -1 0 2010 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1050_
timestamp 1727493435
transform 1 0 1830 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1051_
timestamp 1727493435
transform -1 0 2170 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1052_
timestamp 1727493435
transform -1 0 2650 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1053_
timestamp 1727493435
transform -1 0 2330 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1054_
timestamp 1727493435
transform 1 0 2310 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1055_
timestamp 1727493435
transform -1 0 1930 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1056_
timestamp 1727493435
transform -1 0 2370 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1057_
timestamp 1727493435
transform -1 0 2170 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1058_
timestamp 1727493435
transform 1 0 2050 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1059_
timestamp 1727493435
transform -1 0 1910 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1060_
timestamp 1727493435
transform -1 0 310 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1061_
timestamp 1727493435
transform 1 0 130 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1062_
timestamp 1727493435
transform -1 0 1750 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1063_
timestamp 1727493435
transform -1 0 1770 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1064_
timestamp 1727493435
transform -1 0 1590 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1065_
timestamp 1727493435
transform -1 0 2170 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1066_
timestamp 1727493435
transform 1 0 1830 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1067_
timestamp 1727493435
transform 1 0 2430 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1068_
timestamp 1727493435
transform -1 0 2290 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1069_
timestamp 1727493435
transform 1 0 1650 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1070_
timestamp 1727493435
transform 1 0 830 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1071_
timestamp 1727493435
transform 1 0 2310 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1072_
timestamp 1727493435
transform -1 0 2210 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1073_
timestamp 1727493435
transform 1 0 2210 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1074_
timestamp 1727493435
transform -1 0 2970 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1075_
timestamp 1727493435
transform 1 0 3110 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1076_
timestamp 1727493435
transform 1 0 3070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1077_
timestamp 1727493435
transform 1 0 4090 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1078_
timestamp 1727493435
transform 1 0 4470 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1079_
timestamp 1727493435
transform 1 0 4310 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1080_
timestamp 1727493435
transform 1 0 3710 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1081_
timestamp 1727493435
transform -1 0 3890 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1082_
timestamp 1727493435
transform -1 0 4050 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1083_
timestamp 1727493435
transform 1 0 4190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1084_
timestamp 1727493435
transform 1 0 4370 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1085_
timestamp 1727493435
transform 1 0 4390 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1086_
timestamp 1727493435
transform 1 0 4230 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1087_
timestamp 1727493435
transform -1 0 4230 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1088_
timestamp 1727493435
transform -1 0 4090 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1089_
timestamp 1727493435
transform -1 0 3250 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1090_
timestamp 1727493435
transform -1 0 4590 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1091_
timestamp 1727493435
transform 1 0 3750 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1092_
timestamp 1727493435
transform -1 0 3890 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1093_
timestamp 1727493435
transform -1 0 3290 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1094_
timestamp 1727493435
transform -1 0 3570 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1095_
timestamp 1727493435
transform -1 0 4390 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1096_
timestamp 1727493435
transform -1 0 3930 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1097_
timestamp 1727493435
transform -1 0 4170 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1098_
timestamp 1727493435
transform -1 0 4490 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1099_
timestamp 1727493435
transform -1 0 4070 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1100_
timestamp 1727493435
transform 1 0 3650 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1101_
timestamp 1727493435
transform -1 0 3590 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1102_
timestamp 1727493435
transform -1 0 3430 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1103_
timestamp 1727493435
transform -1 0 4230 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1104_
timestamp 1727493435
transform 1 0 3710 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1105_
timestamp 1727493435
transform -1 0 3870 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1106_
timestamp 1727493435
transform -1 0 3770 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1107_
timestamp 1727493435
transform -1 0 4030 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1108_
timestamp 1727493435
transform -1 0 3510 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1109_
timestamp 1727493435
transform 1 0 4010 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1110_
timestamp 1727493435
transform -1 0 3590 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1111_
timestamp 1727493435
transform -1 0 3190 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1112_
timestamp 1727493435
transform -1 0 3210 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1113_
timestamp 1727493435
transform 1 0 3030 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1114_
timestamp 1727493435
transform -1 0 3430 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1115_
timestamp 1727493435
transform -1 0 3610 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1116_
timestamp 1727493435
transform -1 0 3110 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1117_
timestamp 1727493435
transform -1 0 2710 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1118_
timestamp 1727493435
transform 1 0 3530 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1119_
timestamp 1727493435
transform -1 0 3030 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1120_
timestamp 1727493435
transform 1 0 3250 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1121_
timestamp 1727493435
transform -1 0 3230 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1122_
timestamp 1727493435
transform -1 0 2630 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1123_
timestamp 1727493435
transform -1 0 2870 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1124_
timestamp 1727493435
transform -1 0 3390 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1125_
timestamp 1727493435
transform 1 0 2370 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1126_
timestamp 1727493435
transform -1 0 2490 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1127_
timestamp 1727493435
transform -1 0 2730 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1128_
timestamp 1727493435
transform 1 0 2550 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1129_
timestamp 1727493435
transform -1 0 2950 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1130_
timestamp 1727493435
transform 1 0 3050 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1131_
timestamp 1727493435
transform 1 0 2770 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1132_
timestamp 1727493435
transform 1 0 3150 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1133_
timestamp 1727493435
transform -1 0 2610 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1134_
timestamp 1727493435
transform 1 0 2730 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1135_
timestamp 1727493435
transform 1 0 1190 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1136_
timestamp 1727493435
transform 1 0 4090 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1137_
timestamp 1727493435
transform -1 0 3030 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1138_
timestamp 1727493435
transform 1 0 3290 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1139_
timestamp 1727493435
transform 1 0 3170 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1140_
timestamp 1727493435
transform 1 0 3330 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1141_
timestamp 1727493435
transform 1 0 3650 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1142_
timestamp 1727493435
transform 1 0 4170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1143_
timestamp 1727493435
transform 1 0 3970 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1144_
timestamp 1727493435
transform -1 0 3750 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1145_
timestamp 1727493435
transform 1 0 3850 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1146_
timestamp 1727493435
transform -1 0 4950 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1147_
timestamp 1727493435
transform 1 0 4330 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1148_
timestamp 1727493435
transform 1 0 5050 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1149_
timestamp 1727493435
transform 1 0 4890 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1150_
timestamp 1727493435
transform 1 0 4890 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1151_
timestamp 1727493435
transform -1 0 4670 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1152_
timestamp 1727493435
transform -1 0 4670 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1153_
timestamp 1727493435
transform 1 0 5070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1154_
timestamp 1727493435
transform 1 0 4770 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1155_
timestamp 1727493435
transform 1 0 4470 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1156_
timestamp 1727493435
transform 1 0 4810 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1157_
timestamp 1727493435
transform -1 0 4750 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1158_
timestamp 1727493435
transform 1 0 4710 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1159_
timestamp 1727493435
transform 1 0 5410 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1160_
timestamp 1727493435
transform -1 0 5230 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1161_
timestamp 1727493435
transform -1 0 5250 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1162_
timestamp 1727493435
transform 1 0 5710 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1163_
timestamp 1727493435
transform 1 0 5550 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1164_
timestamp 1727493435
transform -1 0 5710 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1165_
timestamp 1727493435
transform -1 0 4430 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1166_
timestamp 1727493435
transform -1 0 5270 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1167_
timestamp 1727493435
transform 1 0 5350 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1168_
timestamp 1727493435
transform 1 0 5510 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1169_
timestamp 1727493435
transform 1 0 5370 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1170_
timestamp 1727493435
transform 1 0 4490 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1171_
timestamp 1727493435
transform 1 0 5790 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1172_
timestamp 1727493435
transform -1 0 5130 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1173_
timestamp 1727493435
transform 1 0 5050 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1174_
timestamp 1727493435
transform 1 0 4830 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1175_
timestamp 1727493435
transform -1 0 4490 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1176_
timestamp 1727493435
transform 1 0 3810 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1177_
timestamp 1727493435
transform -1 0 3930 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1178_
timestamp 1727493435
transform 1 0 4630 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1179_
timestamp 1727493435
transform -1 0 4970 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1180_
timestamp 1727493435
transform 1 0 4670 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1181_
timestamp 1727493435
transform -1 0 4270 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1182_
timestamp 1727493435
transform 1 0 4790 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1183_
timestamp 1727493435
transform -1 0 4530 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1184_
timestamp 1727493435
transform 1 0 3810 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1185_
timestamp 1727493435
transform 1 0 3930 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1186_
timestamp 1727493435
transform -1 0 3830 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1187_
timestamp 1727493435
transform -1 0 3670 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1188_
timestamp 1727493435
transform -1 0 4110 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1189_
timestamp 1727493435
transform -1 0 3510 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1190_
timestamp 1727493435
transform -1 0 4110 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1191_
timestamp 1727493435
transform 1 0 4330 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1192_
timestamp 1727493435
transform 1 0 4450 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1193_
timestamp 1727493435
transform -1 0 4070 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1194_
timestamp 1727493435
transform 1 0 4170 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1195_
timestamp 1727493435
transform 1 0 4270 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1196_
timestamp 1727493435
transform 1 0 4490 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1197_
timestamp 1727493435
transform -1 0 2210 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1198_
timestamp 1727493435
transform -1 0 4470 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1199_
timestamp 1727493435
transform 1 0 4590 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1200_
timestamp 1727493435
transform -1 0 4650 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1201_
timestamp 1727493435
transform 1 0 4570 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1202_
timestamp 1727493435
transform 1 0 4770 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1203_
timestamp 1727493435
transform -1 0 5230 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1204_
timestamp 1727493435
transform -1 0 5670 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1205_
timestamp 1727493435
transform 1 0 5530 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1206_
timestamp 1727493435
transform -1 0 4550 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1207_
timestamp 1727493435
transform 1 0 4970 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1208_
timestamp 1727493435
transform 1 0 5090 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1209_
timestamp 1727493435
transform 1 0 5210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1210_
timestamp 1727493435
transform 1 0 4910 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1211_
timestamp 1727493435
transform 1 0 5130 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1212_
timestamp 1727493435
transform -1 0 4850 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1213_
timestamp 1727493435
transform -1 0 4990 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1214_
timestamp 1727493435
transform 1 0 4670 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1215_
timestamp 1727493435
transform 1 0 5730 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1216_
timestamp 1727493435
transform 1 0 5630 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1217_
timestamp 1727493435
transform 1 0 5190 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1218_
timestamp 1727493435
transform 1 0 5470 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1219_
timestamp 1727493435
transform 1 0 5870 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1220_
timestamp 1727493435
transform -1 0 5710 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1221_
timestamp 1727493435
transform 1 0 5930 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1222_
timestamp 1727493435
transform 1 0 5830 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1223_
timestamp 1727493435
transform 1 0 5430 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1224_
timestamp 1727493435
transform 1 0 5910 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1225_
timestamp 1727493435
transform 1 0 5750 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1226_
timestamp 1727493435
transform 1 0 5330 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1227_
timestamp 1727493435
transform 1 0 5850 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1228_
timestamp 1727493435
transform -1 0 5610 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1229_
timestamp 1727493435
transform -1 0 5230 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1230_
timestamp 1727493435
transform -1 0 4990 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1231_
timestamp 1727493435
transform 1 0 5370 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1232_
timestamp 1727493435
transform -1 0 5070 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1233_
timestamp 1727493435
transform -1 0 4890 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1234_
timestamp 1727493435
transform 1 0 4830 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1235_
timestamp 1727493435
transform 1 0 4690 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1236_
timestamp 1727493435
transform 1 0 4350 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1237_
timestamp 1727493435
transform 1 0 4510 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1238_
timestamp 1727493435
transform -1 0 3010 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1239_
timestamp 1727493435
transform 1 0 4730 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1240_
timestamp 1727493435
transform -1 0 4430 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1241_
timestamp 1727493435
transform -1 0 4690 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1242_
timestamp 1727493435
transform -1 0 4390 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1243_
timestamp 1727493435
transform -1 0 4250 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1244_
timestamp 1727493435
transform 1 0 4510 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1245_
timestamp 1727493435
transform -1 0 4190 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1246_
timestamp 1727493435
transform -1 0 5610 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1247_
timestamp 1727493435
transform 1 0 5110 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1248_
timestamp 1727493435
transform -1 0 5550 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1249_
timestamp 1727493435
transform -1 0 5370 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1250_
timestamp 1727493435
transform 1 0 5290 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1251_
timestamp 1727493435
transform 1 0 5250 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1252_
timestamp 1727493435
transform 1 0 4930 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1253_
timestamp 1727493435
transform -1 0 5410 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1254_
timestamp 1727493435
transform -1 0 5110 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1255_
timestamp 1727493435
transform 1 0 5530 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1256_
timestamp 1727493435
transform 1 0 4770 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1257_
timestamp 1727493435
transform 1 0 5590 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1258_
timestamp 1727493435
transform -1 0 5750 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1259_
timestamp 1727493435
transform 1 0 5890 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1260_
timestamp 1727493435
transform 1 0 5810 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1261_
timestamp 1727493435
transform -1 0 5670 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1262_
timestamp 1727493435
transform -1 0 5510 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1263_
timestamp 1727493435
transform -1 0 5630 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1264_
timestamp 1727493435
transform -1 0 5750 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1265_
timestamp 1727493435
transform 1 0 5890 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1266_
timestamp 1727493435
transform -1 0 5450 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1267_
timestamp 1727493435
transform 1 0 4910 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1268_
timestamp 1727493435
transform -1 0 3610 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1269_
timestamp 1727493435
transform 1 0 2850 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1270_
timestamp 1727493435
transform 1 0 4330 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1271_
timestamp 1727493435
transform 1 0 3430 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1272_
timestamp 1727493435
transform 1 0 4050 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1273_
timestamp 1727493435
transform 1 0 3890 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1274_
timestamp 1727493435
transform -1 0 3350 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1275_
timestamp 1727493435
transform 1 0 2910 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1276_
timestamp 1727493435
transform -1 0 3230 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1277_
timestamp 1727493435
transform 1 0 5770 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1278_
timestamp 1727493435
transform 1 0 5430 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1279_
timestamp 1727493435
transform 1 0 5270 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1280_
timestamp 1727493435
transform 1 0 4950 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1281_
timestamp 1727493435
transform -1 0 5150 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1282_
timestamp 1727493435
transform 1 0 5270 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1283_
timestamp 1727493435
transform 1 0 5750 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1284_
timestamp 1727493435
transform 1 0 5610 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1285_
timestamp 1727493435
transform 1 0 5910 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1286_
timestamp 1727493435
transform 1 0 5870 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1287_
timestamp 1727493435
transform -1 0 5730 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1288_
timestamp 1727493435
transform -1 0 5150 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1289_
timestamp 1727493435
transform -1 0 3970 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1290_
timestamp 1727493435
transform -1 0 3810 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1291_
timestamp 1727493435
transform 1 0 3730 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1292_
timestamp 1727493435
transform -1 0 3670 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1293_
timestamp 1727493435
transform -1 0 3510 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1294_
timestamp 1727493435
transform 1 0 3350 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1295_
timestamp 1727493435
transform -1 0 5930 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1296_
timestamp 1727493435
transform -1 0 4770 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1297_
timestamp 1727493435
transform -1 0 4590 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1298_
timestamp 1727493435
transform 1 0 4630 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1299_
timestamp 1727493435
transform 1 0 5570 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1300_
timestamp 1727493435
transform 1 0 5430 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1301_
timestamp 1727493435
transform 1 0 4710 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1302_
timestamp 1727493435
transform 1 0 4750 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1303_
timestamp 1727493435
transform 1 0 5490 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1304_
timestamp 1727493435
transform -1 0 5350 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1305_
timestamp 1727493435
transform 1 0 5210 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1306_
timestamp 1727493435
transform 1 0 5270 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1307_
timestamp 1727493435
transform 1 0 5330 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1308_
timestamp 1727493435
transform -1 0 5490 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1309_
timestamp 1727493435
transform 1 0 5610 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1310_
timestamp 1727493435
transform 1 0 5630 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1311_
timestamp 1727493435
transform -1 0 5750 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1312_
timestamp 1727493435
transform 1 0 5090 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1313_
timestamp 1727493435
transform -1 0 5490 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1314_
timestamp 1727493435
transform -1 0 4890 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1315_
timestamp 1727493435
transform -1 0 5070 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1316_
timestamp 1727493435
transform -1 0 5010 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1317_
timestamp 1727493435
transform 1 0 5150 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1318_
timestamp 1727493435
transform -1 0 1930 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1319_
timestamp 1727493435
transform 1 0 2050 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1320_
timestamp 1727493435
transform -1 0 1990 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1321_
timestamp 1727493435
transform 1 0 2090 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1322_
timestamp 1727493435
transform 1 0 2290 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1323_
timestamp 1727493435
transform 1 0 2130 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1324_
timestamp 1727493435
transform 1 0 1510 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1325_
timestamp 1727493435
transform 1 0 1770 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1326_
timestamp 1727493435
transform -1 0 1670 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1327_
timestamp 1727493435
transform -1 0 1810 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1328_
timestamp 1727493435
transform 1 0 1930 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1329_
timestamp 1727493435
transform -1 0 2250 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1330_
timestamp 1727493435
transform -1 0 2310 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1331_
timestamp 1727493435
transform -1 0 2450 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1332_
timestamp 1727493435
transform -1 0 1370 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1333_
timestamp 1727493435
transform -1 0 810 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1334_
timestamp 1727493435
transform -1 0 790 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1335_
timestamp 1727493435
transform -1 0 790 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1336_
timestamp 1727493435
transform 1 0 1070 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1337_
timestamp 1727493435
transform 1 0 910 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1338_
timestamp 1727493435
transform 1 0 1210 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1339_
timestamp 1727493435
transform 1 0 1730 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1340_
timestamp 1727493435
transform 1 0 1570 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1341_
timestamp 1727493435
transform -1 0 630 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1342_
timestamp 1727493435
transform -1 0 530 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1343_
timestamp 1727493435
transform -1 0 390 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1344_
timestamp 1727493435
transform 1 0 590 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1345_
timestamp 1727493435
transform -1 0 150 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1346_
timestamp 1727493435
transform -1 0 490 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1347_
timestamp 1727493435
transform -1 0 270 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1348_
timestamp 1727493435
transform -1 0 170 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1349_
timestamp 1727493435
transform 1 0 750 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1350_
timestamp 1727493435
transform 1 0 1710 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1351_
timestamp 1727493435
transform 1 0 1310 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1352_
timestamp 1727493435
transform -1 0 1450 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1353_
timestamp 1727493435
transform -1 0 30 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1354_
timestamp 1727493435
transform -1 0 30 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1355_
timestamp 1727493435
transform -1 0 330 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1356_
timestamp 1727493435
transform 1 0 310 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1357_
timestamp 1727493435
transform 1 0 150 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1358_
timestamp 1727493435
transform -1 0 30 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1359_
timestamp 1727493435
transform 1 0 170 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1360_
timestamp 1727493435
transform 1 0 430 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1361_
timestamp 1727493435
transform 1 0 1350 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1362_
timestamp 1727493435
transform -1 0 30 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1363_
timestamp 1727493435
transform -1 0 30 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1364_
timestamp 1727493435
transform -1 0 690 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1365_
timestamp 1727493435
transform -1 0 330 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1366_
timestamp 1727493435
transform -1 0 470 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1367_
timestamp 1727493435
transform 1 0 310 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1368_
timestamp 1727493435
transform -1 0 30 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1369_
timestamp 1727493435
transform 1 0 150 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1370_
timestamp 1727493435
transform 1 0 130 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1371_
timestamp 1727493435
transform 1 0 1250 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1372_
timestamp 1727493435
transform -1 0 30 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1373_
timestamp 1727493435
transform -1 0 170 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1374_
timestamp 1727493435
transform 1 0 10 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1375_
timestamp 1727493435
transform 1 0 170 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1376_
timestamp 1727493435
transform -1 0 950 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1377_
timestamp 1727493435
transform 1 0 1290 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1378_
timestamp 1727493435
transform 1 0 910 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1379_
timestamp 1727493435
transform -1 0 770 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1380_
timestamp 1727493435
transform 1 0 690 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1381_
timestamp 1727493435
transform -1 0 550 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1382_
timestamp 1727493435
transform 1 0 850 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1383_
timestamp 1727493435
transform -1 0 650 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1384_
timestamp 1727493435
transform -1 0 770 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1385_
timestamp 1727493435
transform 1 0 570 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1386_
timestamp 1727493435
transform 1 0 790 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1387_
timestamp 1727493435
transform -1 0 350 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1388_
timestamp 1727493435
transform 1 0 1010 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1389_
timestamp 1727493435
transform -1 0 890 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1390_
timestamp 1727493435
transform 1 0 1170 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1391_
timestamp 1727493435
transform 1 0 1790 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1392_
timestamp 1727493435
transform 1 0 1390 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1393_
timestamp 1727493435
transform -1 0 4250 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1394_
timestamp 1727493435
transform -1 0 490 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1395_
timestamp 1727493435
transform -1 0 490 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1396_
timestamp 1727493435
transform -1 0 610 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1397_
timestamp 1727493435
transform 1 0 470 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1398_
timestamp 1727493435
transform 1 0 310 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1399_
timestamp 1727493435
transform 1 0 630 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1400_
timestamp 1727493435
transform -1 0 3970 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1401_
timestamp 1727493435
transform 1 0 3950 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1402_
timestamp 1727493435
transform 1 0 4210 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1403_
timestamp 1727493435
transform 1 0 4090 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1404_
timestamp 1727493435
transform -1 0 4030 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1405_
timestamp 1727493435
transform -1 0 3750 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1406_
timestamp 1727493435
transform -1 0 3670 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1407_
timestamp 1727493435
transform 1 0 4070 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1408_
timestamp 1727493435
transform 1 0 4310 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1409_
timestamp 1727493435
transform 1 0 4450 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1410_
timestamp 1727493435
transform 1 0 4590 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1411_
timestamp 1727493435
transform 1 0 4470 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1412_
timestamp 1727493435
transform 1 0 4750 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1413_
timestamp 1727493435
transform -1 0 4630 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1414_
timestamp 1727493435
transform 1 0 4750 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1415_
timestamp 1727493435
transform -1 0 4790 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1416_
timestamp 1727493435
transform -1 0 3250 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1417_
timestamp 1727493435
transform -1 0 4170 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1418_
timestamp 1727493435
transform -1 0 4310 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1419_
timestamp 1727493435
transform 1 0 4130 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1420_
timestamp 1727493435
transform -1 0 3870 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1421_
timestamp 1727493435
transform -1 0 3010 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1422_
timestamp 1727493435
transform -1 0 2870 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1423_
timestamp 1727493435
transform -1 0 2670 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1424_
timestamp 1727493435
transform 1 0 2790 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1425_
timestamp 1727493435
transform 1 0 2910 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1426_
timestamp 1727493435
transform -1 0 3090 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1427_
timestamp 1727493435
transform 1 0 3070 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1428_
timestamp 1727493435
transform -1 0 2390 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1429_
timestamp 1727493435
transform -1 0 2510 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1430_
timestamp 1727493435
transform -1 0 2650 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1431_
timestamp 1727493435
transform 1 0 2690 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1432_
timestamp 1727493435
transform 1 0 2830 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1433_
timestamp 1727493435
transform 1 0 2770 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1434_
timestamp 1727493435
transform -1 0 2530 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1435_
timestamp 1727493435
transform 1 0 2710 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1436_
timestamp 1727493435
transform 1 0 2550 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1437_
timestamp 1727493435
transform -1 0 2970 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1438_
timestamp 1727493435
transform -1 0 5270 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1439_
timestamp 1727493435
transform 1 0 2910 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1440_
timestamp 1727493435
transform 1 0 3230 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1441_
timestamp 1727493435
transform -1 0 3530 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1442_
timestamp 1727493435
transform 1 0 3370 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1443_
timestamp 1727493435
transform -1 0 3830 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1444_
timestamp 1727493435
transform 1 0 4010 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1445_
timestamp 1727493435
transform 1 0 4610 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1446_
timestamp 1727493435
transform 1 0 5770 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1447_
timestamp 1727493435
transform 1 0 5630 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1448_
timestamp 1727493435
transform -1 0 5750 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1449_
timestamp 1727493435
transform -1 0 5630 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1450_
timestamp 1727493435
transform -1 0 4490 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1451_
timestamp 1727493435
transform 1 0 5950 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1452_
timestamp 1727493435
transform -1 0 5770 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1453_
timestamp 1727493435
transform 1 0 5630 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1454_
timestamp 1727493435
transform 1 0 5710 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1455_
timestamp 1727493435
transform -1 0 5890 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1456_
timestamp 1727493435
transform 1 0 5810 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1457_
timestamp 1727493435
transform -1 0 5230 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1458_
timestamp 1727493435
transform -1 0 5330 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1459_
timestamp 1727493435
transform 1 0 5930 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1460_
timestamp 1727493435
transform 1 0 5930 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1461_
timestamp 1727493435
transform 1 0 5830 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1462_
timestamp 1727493435
transform -1 0 5810 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1463_
timestamp 1727493435
transform 1 0 5830 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1464_
timestamp 1727493435
transform -1 0 4930 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1465_
timestamp 1727493435
transform -1 0 5910 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1466_
timestamp 1727493435
transform 1 0 5910 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1467_
timestamp 1727493435
transform 1 0 5690 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1468_
timestamp 1727493435
transform -1 0 5550 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1469_
timestamp 1727493435
transform 1 0 5190 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1470_
timestamp 1727493435
transform 1 0 5610 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1471_
timestamp 1727493435
transform -1 0 5470 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1472_
timestamp 1727493435
transform -1 0 5230 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1473_
timestamp 1727493435
transform -1 0 5070 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1474_
timestamp 1727493435
transform 1 0 5090 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1475_
timestamp 1727493435
transform -1 0 5350 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1476_
timestamp 1727493435
transform 1 0 5370 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1477_
timestamp 1727493435
transform 1 0 5310 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1478_
timestamp 1727493435
transform -1 0 5110 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1479_
timestamp 1727493435
transform 1 0 2610 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1480_
timestamp 1727493435
transform 1 0 4150 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1481_
timestamp 1727493435
transform 1 0 3950 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1482_
timestamp 1727493435
transform 1 0 3790 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1483_
timestamp 1727493435
transform 1 0 2830 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1484_
timestamp 1727493435
transform 1 0 4390 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1485_
timestamp 1727493435
transform 1 0 3990 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1486_
timestamp 1727493435
transform -1 0 3270 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1487_
timestamp 1727493435
transform -1 0 4910 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1488_
timestamp 1727493435
transform 1 0 4730 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1489_
timestamp 1727493435
transform -1 0 3390 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1490_
timestamp 1727493435
transform -1 0 4790 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1491_
timestamp 1727493435
transform 1 0 4610 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1492_
timestamp 1727493435
transform -1 0 3510 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1493_
timestamp 1727493435
transform 1 0 3470 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1494_
timestamp 1727493435
transform 1 0 3070 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1495_
timestamp 1727493435
transform 1 0 3330 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1496_
timestamp 1727493435
transform 1 0 2930 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1497_
timestamp 1727493435
transform -1 0 3350 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1498_
timestamp 1727493435
transform 1 0 3170 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1499_
timestamp 1727493435
transform 1 0 2790 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1500_
timestamp 1727493435
transform -1 0 2650 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1501_
timestamp 1727493435
transform -1 0 2170 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1502_
timestamp 1727493435
transform 1 0 2290 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1503_
timestamp 1727493435
transform -1 0 2470 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1504_
timestamp 1727493435
transform -1 0 1750 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1505_
timestamp 1727493435
transform -1 0 2150 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1506_
timestamp 1727493435
transform 1 0 1690 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1507_
timestamp 1727493435
transform -1 0 2010 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1508_
timestamp 1727493435
transform -1 0 1390 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1509_
timestamp 1727493435
transform -1 0 1550 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1510_
timestamp 1727493435
transform -1 0 2390 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1511_
timestamp 1727493435
transform -1 0 2530 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1512_
timestamp 1727493435
transform -1 0 2270 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1513_
timestamp 1727493435
transform 1 0 2350 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1514_
timestamp 1727493435
transform -1 0 2650 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1515_
timestamp 1727493435
transform -1 0 2790 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1516_
timestamp 1727493435
transform -1 0 1570 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1517_
timestamp 1727493435
transform -1 0 1950 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1518_
timestamp 1727493435
transform -1 0 1290 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1519_
timestamp 1727493435
transform 1 0 1110 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1520_
timestamp 1727493435
transform 1 0 910 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1521_
timestamp 1727493435
transform -1 0 870 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1522_
timestamp 1727493435
transform -1 0 330 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1523_
timestamp 1727493435
transform -1 0 470 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1524_
timestamp 1727493435
transform 1 0 1410 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1525_
timestamp 1727493435
transform -1 0 1270 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1601_
timestamp 1727493435
transform 1 0 5910 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1602_
timestamp 1727493435
transform 1 0 5930 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1603_
timestamp 1727493435
transform 1 0 5590 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1604_
timestamp 1727493435
transform 1 0 5490 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1605_
timestamp 1727493435
transform 1 0 5790 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1606_
timestamp 1727493435
transform 1 0 4370 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1607_
timestamp 1727493435
transform 1 0 4510 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1608_
timestamp 1727493435
transform 1 0 4650 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1609_
timestamp 1727493435
transform 1 0 4230 0 -1 270
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1727493435
transform -1 0 1770 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1727493435
transform -1 0 1530 0 1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1727493435
transform 1 0 4930 0 -1 790
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1727493435
transform 1 0 3410 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1727493435
transform 1 0 2170 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1727493435
transform 1 0 1690 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1727493435
transform -1 0 3050 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert7
timestamp 1727493435
transform -1 0 4510 0 1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1727493435
transform -1 0 2070 0 -1 790
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1727493435
transform 1 0 2270 0 1 270
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1727493435
transform 1 0 2410 0 1 270
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1727493435
transform 1 0 4950 0 1 270
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1727493435
transform -1 0 4630 0 1 790
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1727493435
transform 1 0 4010 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1727493435
transform -1 0 1550 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1727493435
transform 1 0 2950 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1727493435
transform -1 0 2210 0 1 5470
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1727493435
transform 1 0 2890 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1727493435
transform -1 0 2570 0 1 3390
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1727493435
transform 1 0 730 0 1 3390
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1727493435
transform -1 0 1990 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1727493435
transform -1 0 2130 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1727493435
transform -1 0 1830 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1727493435
transform 1 0 1950 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1727493435
transform 1 0 4590 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert33
timestamp 1727493435
transform -1 0 4350 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1727493435
transform 1 0 2950 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1727493435
transform -1 0 1070 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1727493435
transform -1 0 2450 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1727493435
transform 1 0 5690 0 1 1830
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1727493435
transform -1 0 3750 0 1 1830
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert13
timestamp 1727493435
transform 1 0 4230 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert14
timestamp 1727493435
transform -1 0 2110 0 1 1830
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert15
timestamp 1727493435
transform -1 0 1370 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__760_
timestamp 1727493435
transform 1 0 4830 0 1 270
box -6 -8 26 272
use FILL  FILL_1__761_
timestamp 1727493435
transform 1 0 3650 0 1 270
box -6 -8 26 272
use FILL  FILL_1__762_
timestamp 1727493435
transform 1 0 3130 0 1 270
box -6 -8 26 272
use FILL  FILL_1__763_
timestamp 1727493435
transform 1 0 4330 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__764_
timestamp 1727493435
transform -1 0 2770 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__765_
timestamp 1727493435
transform -1 0 1890 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__766_
timestamp 1727493435
transform -1 0 1910 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__767_
timestamp 1727493435
transform -1 0 4330 0 1 270
box -6 -8 26 272
use FILL  FILL_1__768_
timestamp 1727493435
transform 1 0 3970 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__769_
timestamp 1727493435
transform 1 0 4710 0 1 270
box -6 -8 26 272
use FILL  FILL_1__770_
timestamp 1727493435
transform -1 0 4830 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__771_
timestamp 1727493435
transform -1 0 4970 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__772_
timestamp 1727493435
transform -1 0 2150 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__773_
timestamp 1727493435
transform -1 0 4110 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__774_
timestamp 1727493435
transform 1 0 4170 0 1 270
box -6 -8 26 272
use FILL  FILL_1__775_
timestamp 1727493435
transform 1 0 3630 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__776_
timestamp 1727493435
transform 1 0 2110 0 1 270
box -6 -8 26 272
use FILL  FILL_1__777_
timestamp 1727493435
transform -1 0 4030 0 1 270
box -6 -8 26 272
use FILL  FILL_1__778_
timestamp 1727493435
transform 1 0 3390 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__779_
timestamp 1727493435
transform -1 0 3530 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__780_
timestamp 1727493435
transform -1 0 3830 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__781_
timestamp 1727493435
transform 1 0 1950 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__782_
timestamp 1727493435
transform -1 0 3670 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__783_
timestamp 1727493435
transform -1 0 3410 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__784_
timestamp 1727493435
transform -1 0 2550 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__785_
timestamp 1727493435
transform -1 0 4350 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__786_
timestamp 1727493435
transform -1 0 3170 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__787_
timestamp 1727493435
transform -1 0 4510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__788_
timestamp 1727493435
transform 1 0 4630 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__789_
timestamp 1727493435
transform -1 0 3470 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__790_
timestamp 1727493435
transform -1 0 4070 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__791_
timestamp 1727493435
transform -1 0 4210 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__792_
timestamp 1727493435
transform -1 0 5390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__793_
timestamp 1727493435
transform -1 0 4210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__794_
timestamp 1727493435
transform -1 0 4350 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__795_
timestamp 1727493435
transform 1 0 2670 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__796_
timestamp 1727493435
transform -1 0 2830 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__797_
timestamp 1727493435
transform 1 0 1630 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__798_
timestamp 1727493435
transform -1 0 2370 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__799_
timestamp 1727493435
transform 1 0 1710 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__800_
timestamp 1727493435
transform -1 0 3230 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__801_
timestamp 1727493435
transform 1 0 1570 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__802_
timestamp 1727493435
transform -1 0 3350 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__803_
timestamp 1727493435
transform -1 0 1830 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__804_
timestamp 1727493435
transform -1 0 2350 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__805_
timestamp 1727493435
transform 1 0 2130 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__806_
timestamp 1727493435
transform 1 0 1430 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__807_
timestamp 1727493435
transform 1 0 1850 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__808_
timestamp 1727493435
transform 1 0 1550 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__809_
timestamp 1727493435
transform 1 0 930 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__810_
timestamp 1727493435
transform 1 0 2470 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__811_
timestamp 1727493435
transform 1 0 1050 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__812_
timestamp 1727493435
transform -1 0 690 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__813_
timestamp 1727493435
transform 1 0 1430 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__814_
timestamp 1727493435
transform -1 0 1050 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__815_
timestamp 1727493435
transform -1 0 190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__816_
timestamp 1727493435
transform -1 0 1490 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__817_
timestamp 1727493435
transform 1 0 530 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__818_
timestamp 1727493435
transform -1 0 850 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__819_
timestamp 1727493435
transform 1 0 1610 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__820_
timestamp 1727493435
transform 1 0 1190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__821_
timestamp 1727493435
transform 1 0 1090 0 1 790
box -6 -8 26 272
use FILL  FILL_1__822_
timestamp 1727493435
transform -1 0 1650 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__823_
timestamp 1727493435
transform 1 0 1210 0 1 790
box -6 -8 26 272
use FILL  FILL_1__824_
timestamp 1727493435
transform 1 0 730 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__825_
timestamp 1727493435
transform 1 0 1010 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__826_
timestamp 1727493435
transform 1 0 850 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__827_
timestamp 1727493435
transform 1 0 3930 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__828_
timestamp 1727493435
transform -1 0 3650 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__829_
timestamp 1727493435
transform -1 0 3790 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__830_
timestamp 1727493435
transform 1 0 4030 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__831_
timestamp 1727493435
transform -1 0 3510 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__832_
timestamp 1727493435
transform -1 0 3650 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__833_
timestamp 1727493435
transform 1 0 3150 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__834_
timestamp 1727493435
transform 1 0 3370 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__835_
timestamp 1727493435
transform 1 0 3270 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__836_
timestamp 1727493435
transform 1 0 2410 0 1 790
box -6 -8 26 272
use FILL  FILL_1__837_
timestamp 1727493435
transform 1 0 2290 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__838_
timestamp 1727493435
transform -1 0 2270 0 1 790
box -6 -8 26 272
use FILL  FILL_1__839_
timestamp 1727493435
transform -1 0 5550 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__840_
timestamp 1727493435
transform -1 0 4950 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__841_
timestamp 1727493435
transform -1 0 5390 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__842_
timestamp 1727493435
transform 1 0 5370 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__843_
timestamp 1727493435
transform 1 0 4790 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__844_
timestamp 1727493435
transform -1 0 5190 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__845_
timestamp 1727493435
transform -1 0 4950 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__846_
timestamp 1727493435
transform 1 0 5050 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__847_
timestamp 1727493435
transform -1 0 5070 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__848_
timestamp 1727493435
transform 1 0 5510 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__849_
timestamp 1727493435
transform -1 0 5090 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__850_
timestamp 1727493435
transform 1 0 5210 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__851_
timestamp 1727493435
transform 1 0 1690 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__852_
timestamp 1727493435
transform -1 0 1490 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__853_
timestamp 1727493435
transform -1 0 1450 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__854_
timestamp 1727493435
transform 1 0 1670 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__855_
timestamp 1727493435
transform -1 0 1110 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__856_
timestamp 1727493435
transform 1 0 1310 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__857_
timestamp 1727493435
transform 1 0 1170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__858_
timestamp 1727493435
transform 1 0 1190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__859_
timestamp 1727493435
transform -1 0 1090 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__860_
timestamp 1727493435
transform -1 0 4330 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__861_
timestamp 1727493435
transform -1 0 1250 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__862_
timestamp 1727493435
transform -1 0 1330 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__863_
timestamp 1727493435
transform -1 0 1390 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__864_
timestamp 1727493435
transform -1 0 710 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__865_
timestamp 1727493435
transform 1 0 1490 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__866_
timestamp 1727493435
transform -1 0 1270 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__867_
timestamp 1727493435
transform 1 0 1230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__868_
timestamp 1727493435
transform 1 0 910 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__869_
timestamp 1727493435
transform 1 0 750 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__870_
timestamp 1727493435
transform 1 0 1370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__871_
timestamp 1727493435
transform -1 0 1410 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__872_
timestamp 1727493435
transform -1 0 970 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__873_
timestamp 1727493435
transform -1 0 490 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__874_
timestamp 1727493435
transform -1 0 610 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__875_
timestamp 1727493435
transform 1 0 770 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__876_
timestamp 1727493435
transform -1 0 370 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__877_
timestamp 1727493435
transform -1 0 630 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__878_
timestamp 1727493435
transform -1 0 490 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__879_
timestamp 1727493435
transform -1 0 510 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__880_
timestamp 1727493435
transform -1 0 650 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__881_
timestamp 1727493435
transform -1 0 530 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__882_
timestamp 1727493435
transform 1 0 1790 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__883_
timestamp 1727493435
transform 1 0 1070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__884_
timestamp 1727493435
transform 1 0 1270 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__885_
timestamp 1727493435
transform 1 0 1550 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__886_
timestamp 1727493435
transform 1 0 1270 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__887_
timestamp 1727493435
transform 1 0 1690 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__888_
timestamp 1727493435
transform -1 0 1130 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__889_
timestamp 1727493435
transform -1 0 850 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__890_
timestamp 1727493435
transform -1 0 1890 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__891_
timestamp 1727493435
transform -1 0 970 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__892_
timestamp 1727493435
transform -1 0 850 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__893_
timestamp 1727493435
transform -1 0 530 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__894_
timestamp 1727493435
transform -1 0 490 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__895_
timestamp 1727493435
transform 1 0 910 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__896_
timestamp 1727493435
transform -1 0 690 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__897_
timestamp 1727493435
transform -1 0 1590 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__898_
timestamp 1727493435
transform -1 0 1110 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__899_
timestamp 1727493435
transform 1 0 2970 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__900_
timestamp 1727493435
transform 1 0 3150 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__901_
timestamp 1727493435
transform -1 0 1430 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__902_
timestamp 1727493435
transform -1 0 1130 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__903_
timestamp 1727493435
transform 1 0 750 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__904_
timestamp 1727493435
transform -1 0 330 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__905_
timestamp 1727493435
transform -1 0 50 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__906_
timestamp 1727493435
transform -1 0 650 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__907_
timestamp 1727493435
transform -1 0 610 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__908_
timestamp 1727493435
transform -1 0 170 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__909_
timestamp 1727493435
transform 1 0 190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__910_
timestamp 1727493435
transform -1 0 50 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__911_
timestamp 1727493435
transform -1 0 370 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__912_
timestamp 1727493435
transform -1 0 290 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__913_
timestamp 1727493435
transform 1 0 30 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__914_
timestamp 1727493435
transform 1 0 350 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__915_
timestamp 1727493435
transform 1 0 790 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__916_
timestamp 1727493435
transform -1 0 330 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__917_
timestamp 1727493435
transform 1 0 950 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__918_
timestamp 1727493435
transform 1 0 2250 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__919_
timestamp 1727493435
transform 1 0 1690 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__920_
timestamp 1727493435
transform -1 0 2050 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__921_
timestamp 1727493435
transform 1 0 1110 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__922_
timestamp 1727493435
transform -1 0 1410 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__923_
timestamp 1727493435
transform 1 0 990 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__924_
timestamp 1727493435
transform -1 0 530 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__925_
timestamp 1727493435
transform -1 0 2130 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__926_
timestamp 1727493435
transform 1 0 1410 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__927_
timestamp 1727493435
transform -1 0 690 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__928_
timestamp 1727493435
transform 1 0 510 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__929_
timestamp 1727493435
transform -1 0 690 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__930_
timestamp 1727493435
transform -1 0 370 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__931_
timestamp 1727493435
transform -1 0 850 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__932_
timestamp 1727493435
transform 1 0 190 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__933_
timestamp 1727493435
transform 1 0 2090 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__934_
timestamp 1727493435
transform -1 0 3290 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__935_
timestamp 1727493435
transform 1 0 1550 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__936_
timestamp 1727493435
transform 1 0 1390 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__937_
timestamp 1727493435
transform -1 0 1650 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__938_
timestamp 1727493435
transform -1 0 210 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__939_
timestamp 1727493435
transform -1 0 50 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__940_
timestamp 1727493435
transform -1 0 370 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__941_
timestamp 1727493435
transform -1 0 50 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__942_
timestamp 1727493435
transform -1 0 50 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__943_
timestamp 1727493435
transform 1 0 150 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__944_
timestamp 1727493435
transform -1 0 490 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__945_
timestamp 1727493435
transform 1 0 310 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__946_
timestamp 1727493435
transform -1 0 50 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__947_
timestamp 1727493435
transform -1 0 50 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__948_
timestamp 1727493435
transform 1 0 150 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__949_
timestamp 1727493435
transform -1 0 50 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__950_
timestamp 1727493435
transform 1 0 190 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__951_
timestamp 1727493435
transform 1 0 210 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__952_
timestamp 1727493435
transform -1 0 50 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__953_
timestamp 1727493435
transform 1 0 910 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__954_
timestamp 1727493435
transform 1 0 1850 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__955_
timestamp 1727493435
transform -1 0 50 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__956_
timestamp 1727493435
transform -1 0 50 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__957_
timestamp 1727493435
transform 1 0 190 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__958_
timestamp 1727493435
transform 1 0 2430 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__959_
timestamp 1727493435
transform -1 0 1470 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__960_
timestamp 1727493435
transform 1 0 1730 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__961_
timestamp 1727493435
transform -1 0 1590 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__962_
timestamp 1727493435
transform 1 0 3990 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__963_
timestamp 1727493435
transform -1 0 2050 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__964_
timestamp 1727493435
transform 1 0 1810 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__965_
timestamp 1727493435
transform -1 0 1710 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__966_
timestamp 1727493435
transform -1 0 1910 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__967_
timestamp 1727493435
transform -1 0 1950 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__968_
timestamp 1727493435
transform 1 0 1970 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__969_
timestamp 1727493435
transform 1 0 2230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__970_
timestamp 1727493435
transform 1 0 1230 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__971_
timestamp 1727493435
transform 1 0 3270 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__972_
timestamp 1727493435
transform -1 0 3130 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__973_
timestamp 1727493435
transform 1 0 2670 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__974_
timestamp 1727493435
transform 1 0 2830 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__975_
timestamp 1727493435
transform -1 0 2430 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__976_
timestamp 1727493435
transform -1 0 2530 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__977_
timestamp 1727493435
transform -1 0 2510 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__978_
timestamp 1727493435
transform 1 0 2550 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__979_
timestamp 1727493435
transform -1 0 2830 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__980_
timestamp 1727493435
transform -1 0 2350 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__981_
timestamp 1727493435
transform -1 0 1710 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__982_
timestamp 1727493435
transform 1 0 1530 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__983_
timestamp 1727493435
transform -1 0 2190 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__984_
timestamp 1727493435
transform -1 0 2370 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__985_
timestamp 1727493435
transform -1 0 1870 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__986_
timestamp 1727493435
transform -1 0 1710 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__987_
timestamp 1727493435
transform 1 0 2370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__988_
timestamp 1727493435
transform 1 0 2010 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__989_
timestamp 1727493435
transform -1 0 2030 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__990_
timestamp 1727493435
transform 1 0 2530 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__991_
timestamp 1727493435
transform -1 0 190 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__992_
timestamp 1727493435
transform -1 0 370 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__993_
timestamp 1727493435
transform -1 0 490 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__994_
timestamp 1727493435
transform -1 0 350 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__995_
timestamp 1727493435
transform 1 0 170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__996_
timestamp 1727493435
transform -1 0 790 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__997_
timestamp 1727493435
transform -1 0 50 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__998_
timestamp 1727493435
transform 1 0 430 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__999_
timestamp 1727493435
transform 1 0 790 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1000_
timestamp 1727493435
transform -1 0 490 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1001_
timestamp 1727493435
transform 1 0 910 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1002_
timestamp 1727493435
transform -1 0 630 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1003_
timestamp 1727493435
transform -1 0 1350 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1004_
timestamp 1727493435
transform -1 0 1230 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1005_
timestamp 1727493435
transform 1 0 1270 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1006_
timestamp 1727493435
transform 1 0 1350 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1007_
timestamp 1727493435
transform -1 0 630 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1008_
timestamp 1727493435
transform 1 0 590 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1009_
timestamp 1727493435
transform 1 0 2290 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1010_
timestamp 1727493435
transform 1 0 2130 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1011_
timestamp 1727493435
transform -1 0 2110 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1012_
timestamp 1727493435
transform 1 0 2850 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1013_
timestamp 1727493435
transform 1 0 2690 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1014_
timestamp 1727493435
transform 1 0 2850 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1015_
timestamp 1727493435
transform -1 0 3570 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1016_
timestamp 1727493435
transform 1 0 2570 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1017_
timestamp 1727493435
transform -1 0 3730 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1018_
timestamp 1727493435
transform 1 0 3390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1019_
timestamp 1727493435
transform 1 0 2990 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1020_
timestamp 1727493435
transform -1 0 2750 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1021_
timestamp 1727493435
transform 1 0 3250 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1022_
timestamp 1727493435
transform 1 0 2190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1023_
timestamp 1727493435
transform 1 0 2750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1024_
timestamp 1727493435
transform 1 0 3070 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1025_
timestamp 1727493435
transform -1 0 2710 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1026_
timestamp 1727493435
transform 1 0 2610 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1027_
timestamp 1727493435
transform 1 0 3590 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1028_
timestamp 1727493435
transform -1 0 4170 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1029_
timestamp 1727493435
transform 1 0 3990 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1030_
timestamp 1727493435
transform -1 0 3910 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1031_
timestamp 1727493435
transform -1 0 3750 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1032_
timestamp 1727493435
transform -1 0 3450 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1033_
timestamp 1727493435
transform -1 0 3590 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1034_
timestamp 1727493435
transform 1 0 5090 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1035_
timestamp 1727493435
transform 1 0 3690 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1036_
timestamp 1727493435
transform 1 0 3830 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1037_
timestamp 1727493435
transform -1 0 3110 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1038_
timestamp 1727493435
transform -1 0 2670 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1039_
timestamp 1727493435
transform 1 0 2970 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1040_
timestamp 1727493435
transform -1 0 2790 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1041_
timestamp 1727493435
transform -1 0 3430 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1042_
timestamp 1727493435
transform -1 0 3290 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1043_
timestamp 1727493435
transform -1 0 2950 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1044_
timestamp 1727493435
transform -1 0 2510 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1045_
timestamp 1727493435
transform -1 0 2930 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1046_
timestamp 1727493435
transform 1 0 2810 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1047_
timestamp 1727493435
transform 1 0 2970 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1048_
timestamp 1727493435
transform -1 0 2510 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1049_
timestamp 1727493435
transform -1 0 2030 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1050_
timestamp 1727493435
transform 1 0 1850 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1051_
timestamp 1727493435
transform -1 0 2190 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1052_
timestamp 1727493435
transform -1 0 2670 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1053_
timestamp 1727493435
transform -1 0 2350 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1054_
timestamp 1727493435
transform 1 0 2330 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1055_
timestamp 1727493435
transform -1 0 1950 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1056_
timestamp 1727493435
transform -1 0 2390 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1057_
timestamp 1727493435
transform -1 0 2190 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1058_
timestamp 1727493435
transform 1 0 2070 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1059_
timestamp 1727493435
transform -1 0 1930 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1060_
timestamp 1727493435
transform -1 0 330 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1061_
timestamp 1727493435
transform 1 0 150 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1062_
timestamp 1727493435
transform -1 0 1770 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1063_
timestamp 1727493435
transform -1 0 1790 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1064_
timestamp 1727493435
transform -1 0 1610 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1065_
timestamp 1727493435
transform -1 0 2190 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1066_
timestamp 1727493435
transform 1 0 1850 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1067_
timestamp 1727493435
transform 1 0 2450 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1068_
timestamp 1727493435
transform -1 0 2310 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1069_
timestamp 1727493435
transform 1 0 1670 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1070_
timestamp 1727493435
transform 1 0 850 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1071_
timestamp 1727493435
transform 1 0 2330 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1072_
timestamp 1727493435
transform -1 0 2230 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1073_
timestamp 1727493435
transform 1 0 2230 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1074_
timestamp 1727493435
transform -1 0 2990 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1075_
timestamp 1727493435
transform 1 0 3130 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1076_
timestamp 1727493435
transform 1 0 3090 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1077_
timestamp 1727493435
transform 1 0 4110 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1078_
timestamp 1727493435
transform 1 0 4490 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1079_
timestamp 1727493435
transform 1 0 4330 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1080_
timestamp 1727493435
transform 1 0 3730 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1081_
timestamp 1727493435
transform -1 0 3910 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1082_
timestamp 1727493435
transform -1 0 4070 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1083_
timestamp 1727493435
transform 1 0 4210 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1084_
timestamp 1727493435
transform 1 0 4390 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1085_
timestamp 1727493435
transform 1 0 4410 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1086_
timestamp 1727493435
transform 1 0 4250 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1087_
timestamp 1727493435
transform -1 0 4250 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1088_
timestamp 1727493435
transform -1 0 4110 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1089_
timestamp 1727493435
transform -1 0 3270 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1090_
timestamp 1727493435
transform -1 0 4610 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1091_
timestamp 1727493435
transform 1 0 3770 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1092_
timestamp 1727493435
transform -1 0 3910 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1093_
timestamp 1727493435
transform -1 0 3310 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1094_
timestamp 1727493435
transform -1 0 3590 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1095_
timestamp 1727493435
transform -1 0 4410 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1096_
timestamp 1727493435
transform -1 0 3950 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1097_
timestamp 1727493435
transform -1 0 4190 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1098_
timestamp 1727493435
transform -1 0 4510 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1099_
timestamp 1727493435
transform -1 0 4090 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1100_
timestamp 1727493435
transform 1 0 3670 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1101_
timestamp 1727493435
transform -1 0 3610 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1102_
timestamp 1727493435
transform -1 0 3450 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1103_
timestamp 1727493435
transform -1 0 4250 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1104_
timestamp 1727493435
transform 1 0 3730 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1105_
timestamp 1727493435
transform -1 0 3890 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1106_
timestamp 1727493435
transform -1 0 3790 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1107_
timestamp 1727493435
transform -1 0 4050 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1108_
timestamp 1727493435
transform -1 0 3530 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1109_
timestamp 1727493435
transform 1 0 4030 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1110_
timestamp 1727493435
transform -1 0 3610 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1111_
timestamp 1727493435
transform -1 0 3210 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1112_
timestamp 1727493435
transform -1 0 3230 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1113_
timestamp 1727493435
transform 1 0 3050 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1114_
timestamp 1727493435
transform -1 0 3450 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1115_
timestamp 1727493435
transform -1 0 3630 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1116_
timestamp 1727493435
transform -1 0 3130 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1117_
timestamp 1727493435
transform -1 0 2730 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1118_
timestamp 1727493435
transform 1 0 3550 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1119_
timestamp 1727493435
transform -1 0 3050 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1120_
timestamp 1727493435
transform 1 0 3270 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1121_
timestamp 1727493435
transform -1 0 3250 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1122_
timestamp 1727493435
transform -1 0 2650 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1123_
timestamp 1727493435
transform -1 0 2890 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1124_
timestamp 1727493435
transform -1 0 3410 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1125_
timestamp 1727493435
transform 1 0 2390 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1126_
timestamp 1727493435
transform -1 0 2510 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1127_
timestamp 1727493435
transform -1 0 2750 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1128_
timestamp 1727493435
transform 1 0 2570 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1129_
timestamp 1727493435
transform -1 0 2970 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1130_
timestamp 1727493435
transform 1 0 3070 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1131_
timestamp 1727493435
transform 1 0 2790 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1132_
timestamp 1727493435
transform 1 0 3170 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1133_
timestamp 1727493435
transform -1 0 2630 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1134_
timestamp 1727493435
transform 1 0 2750 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1135_
timestamp 1727493435
transform 1 0 1210 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1136_
timestamp 1727493435
transform 1 0 4110 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1137_
timestamp 1727493435
transform -1 0 3050 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1138_
timestamp 1727493435
transform 1 0 3310 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1139_
timestamp 1727493435
transform 1 0 3190 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1140_
timestamp 1727493435
transform 1 0 3350 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1141_
timestamp 1727493435
transform 1 0 3670 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1142_
timestamp 1727493435
transform 1 0 4190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1143_
timestamp 1727493435
transform 1 0 3990 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1144_
timestamp 1727493435
transform -1 0 3770 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1145_
timestamp 1727493435
transform 1 0 3870 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1146_
timestamp 1727493435
transform -1 0 4970 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1147_
timestamp 1727493435
transform 1 0 4350 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1148_
timestamp 1727493435
transform 1 0 5070 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1149_
timestamp 1727493435
transform 1 0 4910 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1150_
timestamp 1727493435
transform 1 0 4910 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1151_
timestamp 1727493435
transform -1 0 4690 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1152_
timestamp 1727493435
transform -1 0 4690 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1153_
timestamp 1727493435
transform 1 0 5090 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1154_
timestamp 1727493435
transform 1 0 4790 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1155_
timestamp 1727493435
transform 1 0 4490 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1156_
timestamp 1727493435
transform 1 0 4830 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1157_
timestamp 1727493435
transform -1 0 4770 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1158_
timestamp 1727493435
transform 1 0 4730 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1159_
timestamp 1727493435
transform 1 0 5430 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1160_
timestamp 1727493435
transform -1 0 5250 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1161_
timestamp 1727493435
transform -1 0 5270 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1162_
timestamp 1727493435
transform 1 0 5730 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1163_
timestamp 1727493435
transform 1 0 5570 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1164_
timestamp 1727493435
transform -1 0 5730 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1165_
timestamp 1727493435
transform -1 0 4450 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1166_
timestamp 1727493435
transform -1 0 5290 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1167_
timestamp 1727493435
transform 1 0 5370 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1168_
timestamp 1727493435
transform 1 0 5530 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1169_
timestamp 1727493435
transform 1 0 5390 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1170_
timestamp 1727493435
transform 1 0 4510 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1171_
timestamp 1727493435
transform 1 0 5810 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1172_
timestamp 1727493435
transform -1 0 5150 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1173_
timestamp 1727493435
transform 1 0 5070 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1174_
timestamp 1727493435
transform 1 0 4850 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1175_
timestamp 1727493435
transform -1 0 4510 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1176_
timestamp 1727493435
transform 1 0 3830 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1177_
timestamp 1727493435
transform -1 0 3950 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1178_
timestamp 1727493435
transform 1 0 4650 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1179_
timestamp 1727493435
transform -1 0 4990 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1180_
timestamp 1727493435
transform 1 0 4690 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1181_
timestamp 1727493435
transform -1 0 4290 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1182_
timestamp 1727493435
transform 1 0 4810 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1183_
timestamp 1727493435
transform -1 0 4550 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1184_
timestamp 1727493435
transform 1 0 3830 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1185_
timestamp 1727493435
transform 1 0 3950 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1186_
timestamp 1727493435
transform -1 0 3850 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1187_
timestamp 1727493435
transform -1 0 3690 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1188_
timestamp 1727493435
transform -1 0 4130 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1189_
timestamp 1727493435
transform -1 0 3530 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1190_
timestamp 1727493435
transform -1 0 4130 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1191_
timestamp 1727493435
transform 1 0 4350 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1192_
timestamp 1727493435
transform 1 0 4470 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1193_
timestamp 1727493435
transform -1 0 4090 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1194_
timestamp 1727493435
transform 1 0 4190 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1195_
timestamp 1727493435
transform 1 0 4290 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1196_
timestamp 1727493435
transform 1 0 4510 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1197_
timestamp 1727493435
transform -1 0 2230 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1198_
timestamp 1727493435
transform -1 0 4490 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1199_
timestamp 1727493435
transform 1 0 4610 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1200_
timestamp 1727493435
transform -1 0 4670 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1201_
timestamp 1727493435
transform 1 0 4590 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1202_
timestamp 1727493435
transform 1 0 4790 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1203_
timestamp 1727493435
transform -1 0 5250 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1204_
timestamp 1727493435
transform -1 0 5690 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1205_
timestamp 1727493435
transform 1 0 5550 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1206_
timestamp 1727493435
transform -1 0 4570 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1207_
timestamp 1727493435
transform 1 0 4990 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1208_
timestamp 1727493435
transform 1 0 5110 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1209_
timestamp 1727493435
transform 1 0 5230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1210_
timestamp 1727493435
transform 1 0 4930 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1211_
timestamp 1727493435
transform 1 0 5150 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1212_
timestamp 1727493435
transform -1 0 4870 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1213_
timestamp 1727493435
transform -1 0 5010 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1214_
timestamp 1727493435
transform 1 0 4690 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1215_
timestamp 1727493435
transform 1 0 5750 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1216_
timestamp 1727493435
transform 1 0 5650 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1217_
timestamp 1727493435
transform 1 0 5210 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1218_
timestamp 1727493435
transform 1 0 5490 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1219_
timestamp 1727493435
transform 1 0 5890 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1220_
timestamp 1727493435
transform -1 0 5730 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1221_
timestamp 1727493435
transform 1 0 5950 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1222_
timestamp 1727493435
transform 1 0 5850 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1223_
timestamp 1727493435
transform 1 0 5450 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1224_
timestamp 1727493435
transform 1 0 5930 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1225_
timestamp 1727493435
transform 1 0 5770 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1226_
timestamp 1727493435
transform 1 0 5350 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1227_
timestamp 1727493435
transform 1 0 5870 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1228_
timestamp 1727493435
transform -1 0 5630 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1229_
timestamp 1727493435
transform -1 0 5250 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1230_
timestamp 1727493435
transform -1 0 5010 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1231_
timestamp 1727493435
transform 1 0 5390 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1232_
timestamp 1727493435
transform -1 0 5090 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1233_
timestamp 1727493435
transform -1 0 4910 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1234_
timestamp 1727493435
transform 1 0 4850 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1235_
timestamp 1727493435
transform 1 0 4710 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1236_
timestamp 1727493435
transform 1 0 4370 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1237_
timestamp 1727493435
transform 1 0 4530 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1238_
timestamp 1727493435
transform -1 0 3030 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1239_
timestamp 1727493435
transform 1 0 4750 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1240_
timestamp 1727493435
transform -1 0 4450 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1241_
timestamp 1727493435
transform -1 0 4710 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1242_
timestamp 1727493435
transform -1 0 4410 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1243_
timestamp 1727493435
transform -1 0 4270 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1244_
timestamp 1727493435
transform 1 0 4530 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1245_
timestamp 1727493435
transform -1 0 4210 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1246_
timestamp 1727493435
transform -1 0 5630 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1247_
timestamp 1727493435
transform 1 0 5130 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1248_
timestamp 1727493435
transform -1 0 5570 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1249_
timestamp 1727493435
transform -1 0 5390 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1250_
timestamp 1727493435
transform 1 0 5310 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1251_
timestamp 1727493435
transform 1 0 5270 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1252_
timestamp 1727493435
transform 1 0 4950 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1253_
timestamp 1727493435
transform -1 0 5430 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1254_
timestamp 1727493435
transform -1 0 5130 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1255_
timestamp 1727493435
transform 1 0 5550 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1256_
timestamp 1727493435
transform 1 0 4790 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1257_
timestamp 1727493435
transform 1 0 5610 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1258_
timestamp 1727493435
transform -1 0 5770 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1259_
timestamp 1727493435
transform 1 0 5910 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1260_
timestamp 1727493435
transform 1 0 5830 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1261_
timestamp 1727493435
transform -1 0 5690 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1262_
timestamp 1727493435
transform -1 0 5530 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1263_
timestamp 1727493435
transform -1 0 5650 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1264_
timestamp 1727493435
transform -1 0 5770 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1265_
timestamp 1727493435
transform 1 0 5910 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1266_
timestamp 1727493435
transform -1 0 5470 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1267_
timestamp 1727493435
transform 1 0 4930 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1268_
timestamp 1727493435
transform -1 0 3630 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1269_
timestamp 1727493435
transform 1 0 2870 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1270_
timestamp 1727493435
transform 1 0 4350 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1271_
timestamp 1727493435
transform 1 0 3450 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1272_
timestamp 1727493435
transform 1 0 4070 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1273_
timestamp 1727493435
transform 1 0 3910 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1274_
timestamp 1727493435
transform -1 0 3370 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1275_
timestamp 1727493435
transform 1 0 2930 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1276_
timestamp 1727493435
transform -1 0 3250 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1277_
timestamp 1727493435
transform 1 0 5790 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1278_
timestamp 1727493435
transform 1 0 5450 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1279_
timestamp 1727493435
transform 1 0 5290 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1280_
timestamp 1727493435
transform 1 0 4970 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1281_
timestamp 1727493435
transform -1 0 5170 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1282_
timestamp 1727493435
transform 1 0 5290 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1283_
timestamp 1727493435
transform 1 0 5770 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1284_
timestamp 1727493435
transform 1 0 5630 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1285_
timestamp 1727493435
transform 1 0 5930 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1286_
timestamp 1727493435
transform 1 0 5890 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1287_
timestamp 1727493435
transform -1 0 5750 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1288_
timestamp 1727493435
transform -1 0 5170 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1289_
timestamp 1727493435
transform -1 0 3990 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1290_
timestamp 1727493435
transform -1 0 3830 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1291_
timestamp 1727493435
transform 1 0 3750 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1292_
timestamp 1727493435
transform -1 0 3690 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1293_
timestamp 1727493435
transform -1 0 3530 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1294_
timestamp 1727493435
transform 1 0 3370 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1295_
timestamp 1727493435
transform -1 0 5950 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1296_
timestamp 1727493435
transform -1 0 4790 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1297_
timestamp 1727493435
transform -1 0 4610 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1298_
timestamp 1727493435
transform 1 0 4650 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1299_
timestamp 1727493435
transform 1 0 5590 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1300_
timestamp 1727493435
transform 1 0 5450 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1301_
timestamp 1727493435
transform 1 0 4730 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1302_
timestamp 1727493435
transform 1 0 4770 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1303_
timestamp 1727493435
transform 1 0 5510 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1304_
timestamp 1727493435
transform -1 0 5370 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1305_
timestamp 1727493435
transform 1 0 5230 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1306_
timestamp 1727493435
transform 1 0 5290 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1307_
timestamp 1727493435
transform 1 0 5350 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1308_
timestamp 1727493435
transform -1 0 5510 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1309_
timestamp 1727493435
transform 1 0 5630 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1310_
timestamp 1727493435
transform 1 0 5650 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1311_
timestamp 1727493435
transform -1 0 5770 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1312_
timestamp 1727493435
transform 1 0 5110 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1313_
timestamp 1727493435
transform -1 0 5510 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1314_
timestamp 1727493435
transform -1 0 4910 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1315_
timestamp 1727493435
transform -1 0 5090 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1316_
timestamp 1727493435
transform -1 0 5030 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1317_
timestamp 1727493435
transform 1 0 5170 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1318_
timestamp 1727493435
transform -1 0 1950 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1319_
timestamp 1727493435
transform 1 0 2070 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1320_
timestamp 1727493435
transform -1 0 2010 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1321_
timestamp 1727493435
transform 1 0 2110 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1322_
timestamp 1727493435
transform 1 0 2310 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1323_
timestamp 1727493435
transform 1 0 2150 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1324_
timestamp 1727493435
transform 1 0 1530 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1325_
timestamp 1727493435
transform 1 0 1790 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1326_
timestamp 1727493435
transform -1 0 1690 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1327_
timestamp 1727493435
transform -1 0 1830 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1328_
timestamp 1727493435
transform 1 0 1950 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1329_
timestamp 1727493435
transform -1 0 2270 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1330_
timestamp 1727493435
transform -1 0 2330 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1331_
timestamp 1727493435
transform -1 0 2470 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1332_
timestamp 1727493435
transform -1 0 1390 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1333_
timestamp 1727493435
transform -1 0 830 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1334_
timestamp 1727493435
transform -1 0 810 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1335_
timestamp 1727493435
transform -1 0 810 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1336_
timestamp 1727493435
transform 1 0 1090 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1337_
timestamp 1727493435
transform 1 0 930 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1338_
timestamp 1727493435
transform 1 0 1230 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1339_
timestamp 1727493435
transform 1 0 1750 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1340_
timestamp 1727493435
transform 1 0 1590 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1341_
timestamp 1727493435
transform -1 0 650 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1342_
timestamp 1727493435
transform -1 0 550 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1343_
timestamp 1727493435
transform -1 0 410 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1344_
timestamp 1727493435
transform 1 0 610 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1345_
timestamp 1727493435
transform -1 0 170 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1346_
timestamp 1727493435
transform -1 0 510 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1347_
timestamp 1727493435
transform -1 0 290 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1348_
timestamp 1727493435
transform -1 0 190 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1349_
timestamp 1727493435
transform 1 0 770 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1350_
timestamp 1727493435
transform 1 0 1730 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1351_
timestamp 1727493435
transform 1 0 1330 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1352_
timestamp 1727493435
transform -1 0 1470 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1353_
timestamp 1727493435
transform -1 0 50 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1354_
timestamp 1727493435
transform -1 0 50 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1355_
timestamp 1727493435
transform -1 0 350 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1356_
timestamp 1727493435
transform 1 0 330 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1357_
timestamp 1727493435
transform 1 0 170 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1358_
timestamp 1727493435
transform -1 0 50 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1359_
timestamp 1727493435
transform 1 0 190 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1360_
timestamp 1727493435
transform 1 0 450 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1361_
timestamp 1727493435
transform 1 0 1370 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1362_
timestamp 1727493435
transform -1 0 50 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1363_
timestamp 1727493435
transform -1 0 50 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1364_
timestamp 1727493435
transform -1 0 710 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1365_
timestamp 1727493435
transform -1 0 350 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1366_
timestamp 1727493435
transform -1 0 490 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1367_
timestamp 1727493435
transform 1 0 330 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1368_
timestamp 1727493435
transform -1 0 50 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1369_
timestamp 1727493435
transform 1 0 170 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1370_
timestamp 1727493435
transform 1 0 150 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1371_
timestamp 1727493435
transform 1 0 1270 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1372_
timestamp 1727493435
transform -1 0 50 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1373_
timestamp 1727493435
transform -1 0 190 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1374_
timestamp 1727493435
transform 1 0 30 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1375_
timestamp 1727493435
transform 1 0 190 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1376_
timestamp 1727493435
transform -1 0 970 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1377_
timestamp 1727493435
transform 1 0 1310 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1378_
timestamp 1727493435
transform 1 0 930 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1379_
timestamp 1727493435
transform -1 0 790 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1380_
timestamp 1727493435
transform 1 0 710 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1381_
timestamp 1727493435
transform -1 0 570 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1382_
timestamp 1727493435
transform 1 0 870 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1383_
timestamp 1727493435
transform -1 0 670 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1384_
timestamp 1727493435
transform -1 0 790 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1385_
timestamp 1727493435
transform 1 0 590 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1386_
timestamp 1727493435
transform 1 0 810 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1387_
timestamp 1727493435
transform -1 0 370 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1388_
timestamp 1727493435
transform 1 0 1030 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1389_
timestamp 1727493435
transform -1 0 910 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1390_
timestamp 1727493435
transform 1 0 1190 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1391_
timestamp 1727493435
transform 1 0 1810 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1392_
timestamp 1727493435
transform 1 0 1410 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1393_
timestamp 1727493435
transform -1 0 4270 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1394_
timestamp 1727493435
transform -1 0 510 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1395_
timestamp 1727493435
transform -1 0 510 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1396_
timestamp 1727493435
transform -1 0 630 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1397_
timestamp 1727493435
transform 1 0 490 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1398_
timestamp 1727493435
transform 1 0 330 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1399_
timestamp 1727493435
transform 1 0 650 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1400_
timestamp 1727493435
transform -1 0 3990 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1401_
timestamp 1727493435
transform 1 0 3970 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1402_
timestamp 1727493435
transform 1 0 4230 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1403_
timestamp 1727493435
transform 1 0 4110 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1404_
timestamp 1727493435
transform -1 0 4050 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1405_
timestamp 1727493435
transform -1 0 3770 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1406_
timestamp 1727493435
transform -1 0 3690 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1407_
timestamp 1727493435
transform 1 0 4090 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1408_
timestamp 1727493435
transform 1 0 4330 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1409_
timestamp 1727493435
transform 1 0 4470 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1410_
timestamp 1727493435
transform 1 0 4610 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1411_
timestamp 1727493435
transform 1 0 4490 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1412_
timestamp 1727493435
transform 1 0 4770 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1413_
timestamp 1727493435
transform -1 0 4650 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1414_
timestamp 1727493435
transform 1 0 4770 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1415_
timestamp 1727493435
transform -1 0 4810 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1416_
timestamp 1727493435
transform -1 0 3270 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1417_
timestamp 1727493435
transform -1 0 4190 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1418_
timestamp 1727493435
transform -1 0 4330 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1419_
timestamp 1727493435
transform 1 0 4150 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1420_
timestamp 1727493435
transform -1 0 3890 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1421_
timestamp 1727493435
transform -1 0 3030 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1422_
timestamp 1727493435
transform -1 0 2890 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1423_
timestamp 1727493435
transform -1 0 2690 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1424_
timestamp 1727493435
transform 1 0 2810 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1425_
timestamp 1727493435
transform 1 0 2930 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1426_
timestamp 1727493435
transform -1 0 3110 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1427_
timestamp 1727493435
transform 1 0 3090 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1428_
timestamp 1727493435
transform -1 0 2410 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1429_
timestamp 1727493435
transform -1 0 2530 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1430_
timestamp 1727493435
transform -1 0 2670 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1431_
timestamp 1727493435
transform 1 0 2710 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1432_
timestamp 1727493435
transform 1 0 2850 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1433_
timestamp 1727493435
transform 1 0 2790 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1434_
timestamp 1727493435
transform -1 0 2550 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1435_
timestamp 1727493435
transform 1 0 2730 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1436_
timestamp 1727493435
transform 1 0 2570 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1437_
timestamp 1727493435
transform -1 0 2990 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1438_
timestamp 1727493435
transform -1 0 5290 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1439_
timestamp 1727493435
transform 1 0 2930 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1440_
timestamp 1727493435
transform 1 0 3250 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1441_
timestamp 1727493435
transform -1 0 3550 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1442_
timestamp 1727493435
transform 1 0 3390 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1443_
timestamp 1727493435
transform -1 0 3850 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1444_
timestamp 1727493435
transform 1 0 4030 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1445_
timestamp 1727493435
transform 1 0 4630 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1446_
timestamp 1727493435
transform 1 0 5790 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1447_
timestamp 1727493435
transform 1 0 5650 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1448_
timestamp 1727493435
transform -1 0 5770 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1449_
timestamp 1727493435
transform -1 0 5650 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1450_
timestamp 1727493435
transform -1 0 4510 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1451_
timestamp 1727493435
transform 1 0 5970 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1452_
timestamp 1727493435
transform -1 0 5790 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1453_
timestamp 1727493435
transform 1 0 5650 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1454_
timestamp 1727493435
transform 1 0 5730 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1455_
timestamp 1727493435
transform -1 0 5910 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1456_
timestamp 1727493435
transform 1 0 5830 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1457_
timestamp 1727493435
transform -1 0 5250 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1458_
timestamp 1727493435
transform -1 0 5350 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1459_
timestamp 1727493435
transform 1 0 5950 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1460_
timestamp 1727493435
transform 1 0 5950 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1461_
timestamp 1727493435
transform 1 0 5850 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1462_
timestamp 1727493435
transform -1 0 5830 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1463_
timestamp 1727493435
transform 1 0 5850 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1464_
timestamp 1727493435
transform -1 0 4950 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1465_
timestamp 1727493435
transform -1 0 5930 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1466_
timestamp 1727493435
transform 1 0 5930 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1467_
timestamp 1727493435
transform 1 0 5710 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1468_
timestamp 1727493435
transform -1 0 5570 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1469_
timestamp 1727493435
transform 1 0 5210 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1470_
timestamp 1727493435
transform 1 0 5630 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1471_
timestamp 1727493435
transform -1 0 5490 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1472_
timestamp 1727493435
transform -1 0 5250 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1473_
timestamp 1727493435
transform -1 0 5090 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1474_
timestamp 1727493435
transform 1 0 5110 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1475_
timestamp 1727493435
transform -1 0 5370 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1476_
timestamp 1727493435
transform 1 0 5390 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1477_
timestamp 1727493435
transform 1 0 5330 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1478_
timestamp 1727493435
transform -1 0 5130 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1479_
timestamp 1727493435
transform 1 0 2630 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1480_
timestamp 1727493435
transform 1 0 4170 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1481_
timestamp 1727493435
transform 1 0 3970 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1482_
timestamp 1727493435
transform 1 0 3810 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1483_
timestamp 1727493435
transform 1 0 2850 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1484_
timestamp 1727493435
transform 1 0 4410 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1485_
timestamp 1727493435
transform 1 0 4010 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1486_
timestamp 1727493435
transform -1 0 3290 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1487_
timestamp 1727493435
transform -1 0 4930 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1488_
timestamp 1727493435
transform 1 0 4750 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1489_
timestamp 1727493435
transform -1 0 3410 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1490_
timestamp 1727493435
transform -1 0 4810 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1491_
timestamp 1727493435
transform 1 0 4630 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1492_
timestamp 1727493435
transform -1 0 3530 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1493_
timestamp 1727493435
transform 1 0 3490 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1494_
timestamp 1727493435
transform 1 0 3090 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1495_
timestamp 1727493435
transform 1 0 3350 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1496_
timestamp 1727493435
transform 1 0 2950 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1497_
timestamp 1727493435
transform -1 0 3370 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1498_
timestamp 1727493435
transform 1 0 3190 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1499_
timestamp 1727493435
transform 1 0 2810 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1500_
timestamp 1727493435
transform -1 0 2670 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1501_
timestamp 1727493435
transform -1 0 2190 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1502_
timestamp 1727493435
transform 1 0 2310 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1503_
timestamp 1727493435
transform -1 0 2490 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1504_
timestamp 1727493435
transform -1 0 1770 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1505_
timestamp 1727493435
transform -1 0 2170 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1506_
timestamp 1727493435
transform 1 0 1710 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1507_
timestamp 1727493435
transform -1 0 2030 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1508_
timestamp 1727493435
transform -1 0 1410 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1509_
timestamp 1727493435
transform -1 0 1570 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1510_
timestamp 1727493435
transform -1 0 2410 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1511_
timestamp 1727493435
transform -1 0 2550 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1512_
timestamp 1727493435
transform -1 0 2290 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1513_
timestamp 1727493435
transform 1 0 2370 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1514_
timestamp 1727493435
transform -1 0 2670 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1515_
timestamp 1727493435
transform -1 0 2810 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1516_
timestamp 1727493435
transform -1 0 1590 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1517_
timestamp 1727493435
transform -1 0 1970 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1518_
timestamp 1727493435
transform -1 0 1310 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1519_
timestamp 1727493435
transform 1 0 1130 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1520_
timestamp 1727493435
transform 1 0 930 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1521_
timestamp 1727493435
transform -1 0 890 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1522_
timestamp 1727493435
transform -1 0 350 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1523_
timestamp 1727493435
transform -1 0 490 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1524_
timestamp 1727493435
transform 1 0 1430 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1525_
timestamp 1727493435
transform -1 0 1290 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1601_
timestamp 1727493435
transform 1 0 5930 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1602_
timestamp 1727493435
transform 1 0 5950 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1603_
timestamp 1727493435
transform 1 0 5610 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1604_
timestamp 1727493435
transform 1 0 5510 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1605_
timestamp 1727493435
transform 1 0 5810 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1606_
timestamp 1727493435
transform 1 0 4390 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1607_
timestamp 1727493435
transform 1 0 4530 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1608_
timestamp 1727493435
transform 1 0 4670 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1609_
timestamp 1727493435
transform 1 0 4250 0 -1 270
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1727493435
transform -1 0 1790 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1727493435
transform -1 0 1550 0 1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1727493435
transform 1 0 4950 0 -1 790
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1727493435
transform 1 0 3430 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1727493435
transform 1 0 2190 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1727493435
transform 1 0 1710 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert6
timestamp 1727493435
transform -1 0 3070 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert7
timestamp 1727493435
transform -1 0 4530 0 1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1727493435
transform -1 0 2090 0 -1 790
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1727493435
transform 1 0 2290 0 1 270
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1727493435
transform 1 0 2430 0 1 270
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1727493435
transform 1 0 4970 0 1 270
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1727493435
transform -1 0 4650 0 1 790
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1727493435
transform 1 0 4030 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1727493435
transform -1 0 1570 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1727493435
transform 1 0 2970 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1727493435
transform -1 0 2230 0 1 5470
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1727493435
transform 1 0 2910 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1727493435
transform -1 0 2590 0 1 3390
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert27
timestamp 1727493435
transform 1 0 750 0 1 3390
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1727493435
transform -1 0 2010 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert29
timestamp 1727493435
transform -1 0 2150 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1727493435
transform -1 0 1850 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert31
timestamp 1727493435
transform 1 0 1970 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1727493435
transform 1 0 4610 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert33
timestamp 1727493435
transform -1 0 4370 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1727493435
transform 1 0 2970 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1727493435
transform -1 0 1090 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1727493435
transform -1 0 2470 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1727493435
transform 1 0 5710 0 1 1830
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1727493435
transform -1 0 3770 0 1 1830
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert13
timestamp 1727493435
transform 1 0 4250 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert14
timestamp 1727493435
transform -1 0 2130 0 1 1830
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert15
timestamp 1727493435
transform -1 0 1390 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__760_
timestamp 1727493435
transform 1 0 4850 0 1 270
box -6 -8 26 272
use FILL  FILL_2__761_
timestamp 1727493435
transform 1 0 3670 0 1 270
box -6 -8 26 272
use FILL  FILL_2__762_
timestamp 1727493435
transform 1 0 3150 0 1 270
box -6 -8 26 272
use FILL  FILL_2__763_
timestamp 1727493435
transform 1 0 4350 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__764_
timestamp 1727493435
transform -1 0 2790 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__765_
timestamp 1727493435
transform -1 0 1910 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__766_
timestamp 1727493435
transform -1 0 1930 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__767_
timestamp 1727493435
transform -1 0 4350 0 1 270
box -6 -8 26 272
use FILL  FILL_2__768_
timestamp 1727493435
transform 1 0 3990 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__769_
timestamp 1727493435
transform 1 0 4730 0 1 270
box -6 -8 26 272
use FILL  FILL_2__770_
timestamp 1727493435
transform -1 0 4850 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__771_
timestamp 1727493435
transform -1 0 4990 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__772_
timestamp 1727493435
transform -1 0 2170 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__773_
timestamp 1727493435
transform -1 0 4130 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__774_
timestamp 1727493435
transform 1 0 4190 0 1 270
box -6 -8 26 272
use FILL  FILL_2__775_
timestamp 1727493435
transform 1 0 3650 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__776_
timestamp 1727493435
transform 1 0 2130 0 1 270
box -6 -8 26 272
use FILL  FILL_2__777_
timestamp 1727493435
transform -1 0 4050 0 1 270
box -6 -8 26 272
use FILL  FILL_2__778_
timestamp 1727493435
transform 1 0 3410 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__779_
timestamp 1727493435
transform -1 0 3550 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__780_
timestamp 1727493435
transform -1 0 3850 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__781_
timestamp 1727493435
transform 1 0 1970 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__782_
timestamp 1727493435
transform -1 0 3690 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__783_
timestamp 1727493435
transform -1 0 3430 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__784_
timestamp 1727493435
transform -1 0 2570 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__785_
timestamp 1727493435
transform -1 0 4370 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__786_
timestamp 1727493435
transform -1 0 3190 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__787_
timestamp 1727493435
transform -1 0 4530 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__788_
timestamp 1727493435
transform 1 0 4650 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__789_
timestamp 1727493435
transform -1 0 3490 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__790_
timestamp 1727493435
transform -1 0 4090 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__791_
timestamp 1727493435
transform -1 0 4230 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__792_
timestamp 1727493435
transform -1 0 5410 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__793_
timestamp 1727493435
transform -1 0 4230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__794_
timestamp 1727493435
transform -1 0 4370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__795_
timestamp 1727493435
transform 1 0 2690 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__796_
timestamp 1727493435
transform -1 0 2850 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__797_
timestamp 1727493435
transform 1 0 1650 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__798_
timestamp 1727493435
transform -1 0 2390 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__799_
timestamp 1727493435
transform 1 0 1730 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__800_
timestamp 1727493435
transform -1 0 3250 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__801_
timestamp 1727493435
transform 1 0 1590 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__802_
timestamp 1727493435
transform -1 0 3370 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__803_
timestamp 1727493435
transform -1 0 1850 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__804_
timestamp 1727493435
transform -1 0 2370 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__805_
timestamp 1727493435
transform 1 0 2150 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__806_
timestamp 1727493435
transform 1 0 1450 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__807_
timestamp 1727493435
transform 1 0 1870 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__808_
timestamp 1727493435
transform 1 0 1570 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__809_
timestamp 1727493435
transform 1 0 950 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__810_
timestamp 1727493435
transform 1 0 2490 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__811_
timestamp 1727493435
transform 1 0 1070 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__812_
timestamp 1727493435
transform -1 0 710 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__813_
timestamp 1727493435
transform 1 0 1450 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__814_
timestamp 1727493435
transform -1 0 1070 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__815_
timestamp 1727493435
transform -1 0 210 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__816_
timestamp 1727493435
transform -1 0 1510 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__817_
timestamp 1727493435
transform 1 0 550 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__818_
timestamp 1727493435
transform -1 0 870 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__819_
timestamp 1727493435
transform 1 0 1630 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__820_
timestamp 1727493435
transform 1 0 1210 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__821_
timestamp 1727493435
transform 1 0 1110 0 1 790
box -6 -8 26 272
use FILL  FILL_2__822_
timestamp 1727493435
transform -1 0 1670 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__823_
timestamp 1727493435
transform 1 0 1230 0 1 790
box -6 -8 26 272
use FILL  FILL_2__824_
timestamp 1727493435
transform 1 0 750 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__825_
timestamp 1727493435
transform 1 0 1030 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__826_
timestamp 1727493435
transform 1 0 870 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__827_
timestamp 1727493435
transform 1 0 3950 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__828_
timestamp 1727493435
transform -1 0 3670 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__829_
timestamp 1727493435
transform -1 0 3810 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__830_
timestamp 1727493435
transform 1 0 4050 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__831_
timestamp 1727493435
transform -1 0 3530 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__832_
timestamp 1727493435
transform -1 0 3670 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__833_
timestamp 1727493435
transform 1 0 3170 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__834_
timestamp 1727493435
transform 1 0 3390 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__835_
timestamp 1727493435
transform 1 0 3290 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__836_
timestamp 1727493435
transform 1 0 2430 0 1 790
box -6 -8 26 272
use FILL  FILL_2__838_
timestamp 1727493435
transform -1 0 2290 0 1 790
box -6 -8 26 272
use FILL  FILL_2__839_
timestamp 1727493435
transform -1 0 5570 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__840_
timestamp 1727493435
transform -1 0 4970 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__841_
timestamp 1727493435
transform -1 0 5410 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__842_
timestamp 1727493435
transform 1 0 5390 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__843_
timestamp 1727493435
transform 1 0 4810 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__844_
timestamp 1727493435
transform -1 0 5210 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__845_
timestamp 1727493435
transform -1 0 4970 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__846_
timestamp 1727493435
transform 1 0 5070 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__847_
timestamp 1727493435
transform -1 0 5090 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__848_
timestamp 1727493435
transform 1 0 5530 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__849_
timestamp 1727493435
transform -1 0 5110 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__850_
timestamp 1727493435
transform 1 0 5230 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__851_
timestamp 1727493435
transform 1 0 1710 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__852_
timestamp 1727493435
transform -1 0 1510 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__853_
timestamp 1727493435
transform -1 0 1470 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__854_
timestamp 1727493435
transform 1 0 1690 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__855_
timestamp 1727493435
transform -1 0 1130 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__856_
timestamp 1727493435
transform 1 0 1330 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__857_
timestamp 1727493435
transform 1 0 1190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__858_
timestamp 1727493435
transform 1 0 1210 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__859_
timestamp 1727493435
transform -1 0 1110 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__860_
timestamp 1727493435
transform -1 0 4350 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__861_
timestamp 1727493435
transform -1 0 1270 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__862_
timestamp 1727493435
transform -1 0 1350 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__863_
timestamp 1727493435
transform -1 0 1410 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__864_
timestamp 1727493435
transform -1 0 730 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__865_
timestamp 1727493435
transform 1 0 1510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__866_
timestamp 1727493435
transform -1 0 1290 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__867_
timestamp 1727493435
transform 1 0 1250 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__868_
timestamp 1727493435
transform 1 0 930 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__869_
timestamp 1727493435
transform 1 0 770 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__870_
timestamp 1727493435
transform 1 0 1390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__871_
timestamp 1727493435
transform -1 0 1430 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__872_
timestamp 1727493435
transform -1 0 990 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__873_
timestamp 1727493435
transform -1 0 510 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__874_
timestamp 1727493435
transform -1 0 630 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__875_
timestamp 1727493435
transform 1 0 790 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__876_
timestamp 1727493435
transform -1 0 390 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__877_
timestamp 1727493435
transform -1 0 650 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__878_
timestamp 1727493435
transform -1 0 510 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__879_
timestamp 1727493435
transform -1 0 530 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__880_
timestamp 1727493435
transform -1 0 670 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__881_
timestamp 1727493435
transform -1 0 550 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__882_
timestamp 1727493435
transform 1 0 1810 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__883_
timestamp 1727493435
transform 1 0 1090 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__884_
timestamp 1727493435
transform 1 0 1290 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__885_
timestamp 1727493435
transform 1 0 1570 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__886_
timestamp 1727493435
transform 1 0 1290 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__887_
timestamp 1727493435
transform 1 0 1710 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__888_
timestamp 1727493435
transform -1 0 1150 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__889_
timestamp 1727493435
transform -1 0 870 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__890_
timestamp 1727493435
transform -1 0 1910 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__891_
timestamp 1727493435
transform -1 0 990 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__892_
timestamp 1727493435
transform -1 0 870 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__893_
timestamp 1727493435
transform -1 0 550 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__894_
timestamp 1727493435
transform -1 0 510 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__895_
timestamp 1727493435
transform 1 0 930 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__896_
timestamp 1727493435
transform -1 0 710 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__897_
timestamp 1727493435
transform -1 0 1610 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__898_
timestamp 1727493435
transform -1 0 1130 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__899_
timestamp 1727493435
transform 1 0 2990 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__900_
timestamp 1727493435
transform 1 0 3170 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__901_
timestamp 1727493435
transform -1 0 1450 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__902_
timestamp 1727493435
transform -1 0 1150 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__903_
timestamp 1727493435
transform 1 0 770 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__904_
timestamp 1727493435
transform -1 0 350 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__905_
timestamp 1727493435
transform -1 0 70 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__906_
timestamp 1727493435
transform -1 0 670 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__907_
timestamp 1727493435
transform -1 0 630 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__908_
timestamp 1727493435
transform -1 0 190 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__909_
timestamp 1727493435
transform 1 0 210 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__910_
timestamp 1727493435
transform -1 0 70 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__911_
timestamp 1727493435
transform -1 0 390 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__912_
timestamp 1727493435
transform -1 0 310 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__913_
timestamp 1727493435
transform 1 0 50 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__914_
timestamp 1727493435
transform 1 0 370 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__915_
timestamp 1727493435
transform 1 0 810 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__916_
timestamp 1727493435
transform -1 0 350 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__917_
timestamp 1727493435
transform 1 0 970 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__918_
timestamp 1727493435
transform 1 0 2270 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__919_
timestamp 1727493435
transform 1 0 1710 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__920_
timestamp 1727493435
transform -1 0 2070 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__921_
timestamp 1727493435
transform 1 0 1130 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__922_
timestamp 1727493435
transform -1 0 1430 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__923_
timestamp 1727493435
transform 1 0 1010 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__924_
timestamp 1727493435
transform -1 0 550 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__925_
timestamp 1727493435
transform -1 0 2150 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__926_
timestamp 1727493435
transform 1 0 1430 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__927_
timestamp 1727493435
transform -1 0 710 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__928_
timestamp 1727493435
transform 1 0 530 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__929_
timestamp 1727493435
transform -1 0 710 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__930_
timestamp 1727493435
transform -1 0 390 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__931_
timestamp 1727493435
transform -1 0 870 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__932_
timestamp 1727493435
transform 1 0 210 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__933_
timestamp 1727493435
transform 1 0 2110 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__934_
timestamp 1727493435
transform -1 0 3310 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__935_
timestamp 1727493435
transform 1 0 1570 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__936_
timestamp 1727493435
transform 1 0 1410 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__937_
timestamp 1727493435
transform -1 0 1670 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__938_
timestamp 1727493435
transform -1 0 230 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__939_
timestamp 1727493435
transform -1 0 70 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__940_
timestamp 1727493435
transform -1 0 390 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__941_
timestamp 1727493435
transform -1 0 70 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__942_
timestamp 1727493435
transform -1 0 70 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__943_
timestamp 1727493435
transform 1 0 170 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__944_
timestamp 1727493435
transform -1 0 510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__945_
timestamp 1727493435
transform 1 0 330 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__946_
timestamp 1727493435
transform -1 0 70 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__947_
timestamp 1727493435
transform -1 0 70 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__948_
timestamp 1727493435
transform 1 0 170 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__949_
timestamp 1727493435
transform -1 0 70 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__950_
timestamp 1727493435
transform 1 0 210 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__951_
timestamp 1727493435
transform 1 0 230 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__952_
timestamp 1727493435
transform -1 0 70 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__953_
timestamp 1727493435
transform 1 0 930 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__954_
timestamp 1727493435
transform 1 0 1870 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__955_
timestamp 1727493435
transform -1 0 70 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__956_
timestamp 1727493435
transform -1 0 70 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__957_
timestamp 1727493435
transform 1 0 210 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__958_
timestamp 1727493435
transform 1 0 2450 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__959_
timestamp 1727493435
transform -1 0 1490 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__960_
timestamp 1727493435
transform 1 0 1750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__961_
timestamp 1727493435
transform -1 0 1610 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__962_
timestamp 1727493435
transform 1 0 4010 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__963_
timestamp 1727493435
transform -1 0 2070 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__964_
timestamp 1727493435
transform 1 0 1830 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__965_
timestamp 1727493435
transform -1 0 1730 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__966_
timestamp 1727493435
transform -1 0 1930 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__967_
timestamp 1727493435
transform -1 0 1970 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__968_
timestamp 1727493435
transform 1 0 1990 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__969_
timestamp 1727493435
transform 1 0 2250 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__970_
timestamp 1727493435
transform 1 0 1250 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__971_
timestamp 1727493435
transform 1 0 3290 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__972_
timestamp 1727493435
transform -1 0 3150 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__973_
timestamp 1727493435
transform 1 0 2690 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__974_
timestamp 1727493435
transform 1 0 2850 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__975_
timestamp 1727493435
transform -1 0 2450 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__976_
timestamp 1727493435
transform -1 0 2550 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__977_
timestamp 1727493435
transform -1 0 2530 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__978_
timestamp 1727493435
transform 1 0 2570 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__979_
timestamp 1727493435
transform -1 0 2850 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__980_
timestamp 1727493435
transform -1 0 2370 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__981_
timestamp 1727493435
transform -1 0 1730 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__982_
timestamp 1727493435
transform 1 0 1550 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__983_
timestamp 1727493435
transform -1 0 2210 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__984_
timestamp 1727493435
transform -1 0 2390 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__985_
timestamp 1727493435
transform -1 0 1890 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__986_
timestamp 1727493435
transform -1 0 1730 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__987_
timestamp 1727493435
transform 1 0 2390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__988_
timestamp 1727493435
transform 1 0 2030 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__989_
timestamp 1727493435
transform -1 0 2050 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__990_
timestamp 1727493435
transform 1 0 2550 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__991_
timestamp 1727493435
transform -1 0 210 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__992_
timestamp 1727493435
transform -1 0 390 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__993_
timestamp 1727493435
transform -1 0 510 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__994_
timestamp 1727493435
transform -1 0 370 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__995_
timestamp 1727493435
transform 1 0 190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__996_
timestamp 1727493435
transform -1 0 810 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__997_
timestamp 1727493435
transform -1 0 70 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__998_
timestamp 1727493435
transform 1 0 450 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1000_
timestamp 1727493435
transform -1 0 510 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1001_
timestamp 1727493435
transform 1 0 930 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1002_
timestamp 1727493435
transform -1 0 650 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1003_
timestamp 1727493435
transform -1 0 1370 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1004_
timestamp 1727493435
transform -1 0 1250 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1005_
timestamp 1727493435
transform 1 0 1290 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1006_
timestamp 1727493435
transform 1 0 1370 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1007_
timestamp 1727493435
transform -1 0 650 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1008_
timestamp 1727493435
transform 1 0 610 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1009_
timestamp 1727493435
transform 1 0 2310 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1010_
timestamp 1727493435
transform 1 0 2150 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1011_
timestamp 1727493435
transform -1 0 2130 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1012_
timestamp 1727493435
transform 1 0 2870 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1013_
timestamp 1727493435
transform 1 0 2710 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1014_
timestamp 1727493435
transform 1 0 2870 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1015_
timestamp 1727493435
transform -1 0 3590 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1016_
timestamp 1727493435
transform 1 0 2590 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1017_
timestamp 1727493435
transform -1 0 3750 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1018_
timestamp 1727493435
transform 1 0 3410 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1019_
timestamp 1727493435
transform 1 0 3010 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1020_
timestamp 1727493435
transform -1 0 2770 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1021_
timestamp 1727493435
transform 1 0 3270 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1022_
timestamp 1727493435
transform 1 0 2210 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1023_
timestamp 1727493435
transform 1 0 2770 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1024_
timestamp 1727493435
transform 1 0 3090 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1025_
timestamp 1727493435
transform -1 0 2730 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1026_
timestamp 1727493435
transform 1 0 2630 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1027_
timestamp 1727493435
transform 1 0 3610 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1028_
timestamp 1727493435
transform -1 0 4190 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1029_
timestamp 1727493435
transform 1 0 4010 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1030_
timestamp 1727493435
transform -1 0 3930 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1031_
timestamp 1727493435
transform -1 0 3770 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1032_
timestamp 1727493435
transform -1 0 3470 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1033_
timestamp 1727493435
transform -1 0 3610 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1034_
timestamp 1727493435
transform 1 0 5110 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1035_
timestamp 1727493435
transform 1 0 3710 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1036_
timestamp 1727493435
transform 1 0 3850 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1037_
timestamp 1727493435
transform -1 0 3130 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1038_
timestamp 1727493435
transform -1 0 2690 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1039_
timestamp 1727493435
transform 1 0 2990 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1040_
timestamp 1727493435
transform -1 0 2810 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1041_
timestamp 1727493435
transform -1 0 3450 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1042_
timestamp 1727493435
transform -1 0 3310 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1043_
timestamp 1727493435
transform -1 0 2970 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1044_
timestamp 1727493435
transform -1 0 2530 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1045_
timestamp 1727493435
transform -1 0 2950 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1046_
timestamp 1727493435
transform 1 0 2830 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1047_
timestamp 1727493435
transform 1 0 2990 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1048_
timestamp 1727493435
transform -1 0 2530 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1049_
timestamp 1727493435
transform -1 0 2050 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1050_
timestamp 1727493435
transform 1 0 1870 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1051_
timestamp 1727493435
transform -1 0 2210 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1052_
timestamp 1727493435
transform -1 0 2690 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1053_
timestamp 1727493435
transform -1 0 2370 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1054_
timestamp 1727493435
transform 1 0 2350 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1055_
timestamp 1727493435
transform -1 0 1970 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1056_
timestamp 1727493435
transform -1 0 2410 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1057_
timestamp 1727493435
transform -1 0 2210 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1058_
timestamp 1727493435
transform 1 0 2090 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1059_
timestamp 1727493435
transform -1 0 1950 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1060_
timestamp 1727493435
transform -1 0 350 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1061_
timestamp 1727493435
transform 1 0 170 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1062_
timestamp 1727493435
transform -1 0 1790 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1063_
timestamp 1727493435
transform -1 0 1810 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1064_
timestamp 1727493435
transform -1 0 1630 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1065_
timestamp 1727493435
transform -1 0 2210 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1066_
timestamp 1727493435
transform 1 0 1870 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1067_
timestamp 1727493435
transform 1 0 2470 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1068_
timestamp 1727493435
transform -1 0 2330 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1069_
timestamp 1727493435
transform 1 0 1690 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1070_
timestamp 1727493435
transform 1 0 870 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1071_
timestamp 1727493435
transform 1 0 2350 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1072_
timestamp 1727493435
transform -1 0 2250 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1073_
timestamp 1727493435
transform 1 0 2250 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1074_
timestamp 1727493435
transform -1 0 3010 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1075_
timestamp 1727493435
transform 1 0 3150 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1076_
timestamp 1727493435
transform 1 0 3110 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1077_
timestamp 1727493435
transform 1 0 4130 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1078_
timestamp 1727493435
transform 1 0 4510 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1079_
timestamp 1727493435
transform 1 0 4350 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1080_
timestamp 1727493435
transform 1 0 3750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1081_
timestamp 1727493435
transform -1 0 3930 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1082_
timestamp 1727493435
transform -1 0 4090 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1083_
timestamp 1727493435
transform 1 0 4230 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1084_
timestamp 1727493435
transform 1 0 4410 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1085_
timestamp 1727493435
transform 1 0 4430 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1086_
timestamp 1727493435
transform 1 0 4270 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1087_
timestamp 1727493435
transform -1 0 4270 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1088_
timestamp 1727493435
transform -1 0 4130 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1089_
timestamp 1727493435
transform -1 0 3290 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1090_
timestamp 1727493435
transform -1 0 4630 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1091_
timestamp 1727493435
transform 1 0 3790 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1092_
timestamp 1727493435
transform -1 0 3930 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1093_
timestamp 1727493435
transform -1 0 3330 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1094_
timestamp 1727493435
transform -1 0 3610 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1095_
timestamp 1727493435
transform -1 0 4430 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1096_
timestamp 1727493435
transform -1 0 3970 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1097_
timestamp 1727493435
transform -1 0 4210 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1098_
timestamp 1727493435
transform -1 0 4530 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1099_
timestamp 1727493435
transform -1 0 4110 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1100_
timestamp 1727493435
transform 1 0 3690 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1101_
timestamp 1727493435
transform -1 0 3630 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1102_
timestamp 1727493435
transform -1 0 3470 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1103_
timestamp 1727493435
transform -1 0 4270 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1104_
timestamp 1727493435
transform 1 0 3750 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1105_
timestamp 1727493435
transform -1 0 3910 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1106_
timestamp 1727493435
transform -1 0 3810 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1107_
timestamp 1727493435
transform -1 0 4070 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1108_
timestamp 1727493435
transform -1 0 3550 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1109_
timestamp 1727493435
transform 1 0 4050 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1110_
timestamp 1727493435
transform -1 0 3630 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1111_
timestamp 1727493435
transform -1 0 3230 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1112_
timestamp 1727493435
transform -1 0 3250 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1113_
timestamp 1727493435
transform 1 0 3070 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1114_
timestamp 1727493435
transform -1 0 3470 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1115_
timestamp 1727493435
transform -1 0 3650 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1116_
timestamp 1727493435
transform -1 0 3150 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1117_
timestamp 1727493435
transform -1 0 2750 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1118_
timestamp 1727493435
transform 1 0 3570 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1119_
timestamp 1727493435
transform -1 0 3070 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1120_
timestamp 1727493435
transform 1 0 3290 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1121_
timestamp 1727493435
transform -1 0 3270 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1122_
timestamp 1727493435
transform -1 0 2670 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1123_
timestamp 1727493435
transform -1 0 2910 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1124_
timestamp 1727493435
transform -1 0 3430 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1125_
timestamp 1727493435
transform 1 0 2410 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1126_
timestamp 1727493435
transform -1 0 2530 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1128_
timestamp 1727493435
transform 1 0 2590 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1129_
timestamp 1727493435
transform -1 0 2990 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1130_
timestamp 1727493435
transform 1 0 3090 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1131_
timestamp 1727493435
transform 1 0 2810 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1132_
timestamp 1727493435
transform 1 0 3190 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1133_
timestamp 1727493435
transform -1 0 2650 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1134_
timestamp 1727493435
transform 1 0 2770 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1135_
timestamp 1727493435
transform 1 0 1230 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1136_
timestamp 1727493435
transform 1 0 4130 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1137_
timestamp 1727493435
transform -1 0 3070 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1138_
timestamp 1727493435
transform 1 0 3330 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1139_
timestamp 1727493435
transform 1 0 3210 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1140_
timestamp 1727493435
transform 1 0 3370 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1141_
timestamp 1727493435
transform 1 0 3690 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1142_
timestamp 1727493435
transform 1 0 4210 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1143_
timestamp 1727493435
transform 1 0 4010 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1144_
timestamp 1727493435
transform -1 0 3790 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1145_
timestamp 1727493435
transform 1 0 3890 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1146_
timestamp 1727493435
transform -1 0 4990 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1147_
timestamp 1727493435
transform 1 0 4370 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1148_
timestamp 1727493435
transform 1 0 5090 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1149_
timestamp 1727493435
transform 1 0 4930 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1150_
timestamp 1727493435
transform 1 0 4930 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1151_
timestamp 1727493435
transform -1 0 4710 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1152_
timestamp 1727493435
transform -1 0 4710 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1153_
timestamp 1727493435
transform 1 0 5110 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1154_
timestamp 1727493435
transform 1 0 4810 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1155_
timestamp 1727493435
transform 1 0 4510 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1156_
timestamp 1727493435
transform 1 0 4850 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1157_
timestamp 1727493435
transform -1 0 4790 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1158_
timestamp 1727493435
transform 1 0 4750 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1159_
timestamp 1727493435
transform 1 0 5450 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1160_
timestamp 1727493435
transform -1 0 5270 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1161_
timestamp 1727493435
transform -1 0 5290 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1162_
timestamp 1727493435
transform 1 0 5750 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1163_
timestamp 1727493435
transform 1 0 5590 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1164_
timestamp 1727493435
transform -1 0 5750 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1165_
timestamp 1727493435
transform -1 0 4470 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1166_
timestamp 1727493435
transform -1 0 5310 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1167_
timestamp 1727493435
transform 1 0 5390 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1168_
timestamp 1727493435
transform 1 0 5550 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1169_
timestamp 1727493435
transform 1 0 5410 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1170_
timestamp 1727493435
transform 1 0 4530 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1171_
timestamp 1727493435
transform 1 0 5830 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1172_
timestamp 1727493435
transform -1 0 5170 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1173_
timestamp 1727493435
transform 1 0 5090 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1174_
timestamp 1727493435
transform 1 0 4870 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1175_
timestamp 1727493435
transform -1 0 4530 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1176_
timestamp 1727493435
transform 1 0 3850 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1177_
timestamp 1727493435
transform -1 0 3970 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1178_
timestamp 1727493435
transform 1 0 4670 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1179_
timestamp 1727493435
transform -1 0 5010 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1180_
timestamp 1727493435
transform 1 0 4710 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1181_
timestamp 1727493435
transform -1 0 4310 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1182_
timestamp 1727493435
transform 1 0 4830 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1183_
timestamp 1727493435
transform -1 0 4570 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1184_
timestamp 1727493435
transform 1 0 3850 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1185_
timestamp 1727493435
transform 1 0 3970 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1186_
timestamp 1727493435
transform -1 0 3870 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1187_
timestamp 1727493435
transform -1 0 3710 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1188_
timestamp 1727493435
transform -1 0 4150 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1189_
timestamp 1727493435
transform -1 0 3550 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1190_
timestamp 1727493435
transform -1 0 4150 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1191_
timestamp 1727493435
transform 1 0 4370 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1192_
timestamp 1727493435
transform 1 0 4490 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1193_
timestamp 1727493435
transform -1 0 4110 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1194_
timestamp 1727493435
transform 1 0 4210 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1195_
timestamp 1727493435
transform 1 0 4310 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1196_
timestamp 1727493435
transform 1 0 4530 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1197_
timestamp 1727493435
transform -1 0 2250 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1198_
timestamp 1727493435
transform -1 0 4510 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1199_
timestamp 1727493435
transform 1 0 4630 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1200_
timestamp 1727493435
transform -1 0 4690 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1201_
timestamp 1727493435
transform 1 0 4610 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1202_
timestamp 1727493435
transform 1 0 4810 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1203_
timestamp 1727493435
transform -1 0 5270 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1204_
timestamp 1727493435
transform -1 0 5710 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1205_
timestamp 1727493435
transform 1 0 5570 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1206_
timestamp 1727493435
transform -1 0 4590 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1207_
timestamp 1727493435
transform 1 0 5010 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1208_
timestamp 1727493435
transform 1 0 5130 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1209_
timestamp 1727493435
transform 1 0 5250 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1210_
timestamp 1727493435
transform 1 0 4950 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1211_
timestamp 1727493435
transform 1 0 5170 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1212_
timestamp 1727493435
transform -1 0 4890 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1213_
timestamp 1727493435
transform -1 0 5030 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1214_
timestamp 1727493435
transform 1 0 4710 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1215_
timestamp 1727493435
transform 1 0 5770 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1216_
timestamp 1727493435
transform 1 0 5670 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1217_
timestamp 1727493435
transform 1 0 5230 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1218_
timestamp 1727493435
transform 1 0 5510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1219_
timestamp 1727493435
transform 1 0 5910 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1220_
timestamp 1727493435
transform -1 0 5750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1221_
timestamp 1727493435
transform 1 0 5970 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1222_
timestamp 1727493435
transform 1 0 5870 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1223_
timestamp 1727493435
transform 1 0 5470 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1224_
timestamp 1727493435
transform 1 0 5950 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1225_
timestamp 1727493435
transform 1 0 5790 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1226_
timestamp 1727493435
transform 1 0 5370 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1227_
timestamp 1727493435
transform 1 0 5890 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1228_
timestamp 1727493435
transform -1 0 5650 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1229_
timestamp 1727493435
transform -1 0 5270 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1230_
timestamp 1727493435
transform -1 0 5030 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1231_
timestamp 1727493435
transform 1 0 5410 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1232_
timestamp 1727493435
transform -1 0 5110 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1233_
timestamp 1727493435
transform -1 0 4930 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1234_
timestamp 1727493435
transform 1 0 4870 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1235_
timestamp 1727493435
transform 1 0 4730 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1236_
timestamp 1727493435
transform 1 0 4390 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1237_
timestamp 1727493435
transform 1 0 4550 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1238_
timestamp 1727493435
transform -1 0 3050 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1239_
timestamp 1727493435
transform 1 0 4770 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1240_
timestamp 1727493435
transform -1 0 4470 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1241_
timestamp 1727493435
transform -1 0 4730 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1242_
timestamp 1727493435
transform -1 0 4430 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1243_
timestamp 1727493435
transform -1 0 4290 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1244_
timestamp 1727493435
transform 1 0 4550 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1245_
timestamp 1727493435
transform -1 0 4230 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1246_
timestamp 1727493435
transform -1 0 5650 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1247_
timestamp 1727493435
transform 1 0 5150 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1248_
timestamp 1727493435
transform -1 0 5590 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1249_
timestamp 1727493435
transform -1 0 5410 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1250_
timestamp 1727493435
transform 1 0 5330 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1251_
timestamp 1727493435
transform 1 0 5290 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1252_
timestamp 1727493435
transform 1 0 4970 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1253_
timestamp 1727493435
transform -1 0 5450 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1254_
timestamp 1727493435
transform -1 0 5150 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1255_
timestamp 1727493435
transform 1 0 5570 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1256_
timestamp 1727493435
transform 1 0 4810 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1257_
timestamp 1727493435
transform 1 0 5630 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1258_
timestamp 1727493435
transform -1 0 5790 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1259_
timestamp 1727493435
transform 1 0 5930 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1260_
timestamp 1727493435
transform 1 0 5850 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1261_
timestamp 1727493435
transform -1 0 5710 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1262_
timestamp 1727493435
transform -1 0 5550 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1263_
timestamp 1727493435
transform -1 0 5670 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1264_
timestamp 1727493435
transform -1 0 5790 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1265_
timestamp 1727493435
transform 1 0 5930 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1266_
timestamp 1727493435
transform -1 0 5490 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1267_
timestamp 1727493435
transform 1 0 4950 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1268_
timestamp 1727493435
transform -1 0 3650 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1269_
timestamp 1727493435
transform 1 0 2890 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1270_
timestamp 1727493435
transform 1 0 4370 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1271_
timestamp 1727493435
transform 1 0 3470 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1272_
timestamp 1727493435
transform 1 0 4090 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1273_
timestamp 1727493435
transform 1 0 3930 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1274_
timestamp 1727493435
transform -1 0 3390 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1275_
timestamp 1727493435
transform 1 0 2950 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1276_
timestamp 1727493435
transform -1 0 3270 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1277_
timestamp 1727493435
transform 1 0 5810 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1278_
timestamp 1727493435
transform 1 0 5470 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1279_
timestamp 1727493435
transform 1 0 5310 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1280_
timestamp 1727493435
transform 1 0 4990 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1281_
timestamp 1727493435
transform -1 0 5190 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1282_
timestamp 1727493435
transform 1 0 5310 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1283_
timestamp 1727493435
transform 1 0 5790 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1284_
timestamp 1727493435
transform 1 0 5650 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1285_
timestamp 1727493435
transform 1 0 5950 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1286_
timestamp 1727493435
transform 1 0 5910 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1287_
timestamp 1727493435
transform -1 0 5770 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1288_
timestamp 1727493435
transform -1 0 5190 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1290_
timestamp 1727493435
transform -1 0 3850 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1291_
timestamp 1727493435
transform 1 0 3770 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1292_
timestamp 1727493435
transform -1 0 3710 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1293_
timestamp 1727493435
transform -1 0 3550 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1294_
timestamp 1727493435
transform 1 0 3390 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1295_
timestamp 1727493435
transform -1 0 5970 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1296_
timestamp 1727493435
transform -1 0 4810 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1297_
timestamp 1727493435
transform -1 0 4630 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1298_
timestamp 1727493435
transform 1 0 4670 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1299_
timestamp 1727493435
transform 1 0 5610 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1300_
timestamp 1727493435
transform 1 0 5470 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1301_
timestamp 1727493435
transform 1 0 4750 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1302_
timestamp 1727493435
transform 1 0 4790 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1303_
timestamp 1727493435
transform 1 0 5530 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1304_
timestamp 1727493435
transform -1 0 5390 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1305_
timestamp 1727493435
transform 1 0 5250 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1306_
timestamp 1727493435
transform 1 0 5310 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1307_
timestamp 1727493435
transform 1 0 5370 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1308_
timestamp 1727493435
transform -1 0 5530 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1309_
timestamp 1727493435
transform 1 0 5650 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1310_
timestamp 1727493435
transform 1 0 5670 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1311_
timestamp 1727493435
transform -1 0 5790 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1312_
timestamp 1727493435
transform 1 0 5130 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1313_
timestamp 1727493435
transform -1 0 5530 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1314_
timestamp 1727493435
transform -1 0 4930 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1315_
timestamp 1727493435
transform -1 0 5110 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1316_
timestamp 1727493435
transform -1 0 5050 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1317_
timestamp 1727493435
transform 1 0 5190 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1318_
timestamp 1727493435
transform -1 0 1970 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1319_
timestamp 1727493435
transform 1 0 2090 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1320_
timestamp 1727493435
transform -1 0 2030 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1321_
timestamp 1727493435
transform 1 0 2130 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1322_
timestamp 1727493435
transform 1 0 2330 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1323_
timestamp 1727493435
transform 1 0 2170 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1324_
timestamp 1727493435
transform 1 0 1550 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1325_
timestamp 1727493435
transform 1 0 1810 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1326_
timestamp 1727493435
transform -1 0 1710 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1327_
timestamp 1727493435
transform -1 0 1850 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1328_
timestamp 1727493435
transform 1 0 1970 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1329_
timestamp 1727493435
transform -1 0 2290 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1330_
timestamp 1727493435
transform -1 0 2350 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1331_
timestamp 1727493435
transform -1 0 2490 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1332_
timestamp 1727493435
transform -1 0 1410 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1333_
timestamp 1727493435
transform -1 0 850 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1334_
timestamp 1727493435
transform -1 0 830 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1335_
timestamp 1727493435
transform -1 0 830 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1336_
timestamp 1727493435
transform 1 0 1110 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1337_
timestamp 1727493435
transform 1 0 950 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1338_
timestamp 1727493435
transform 1 0 1250 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1339_
timestamp 1727493435
transform 1 0 1770 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1340_
timestamp 1727493435
transform 1 0 1610 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1341_
timestamp 1727493435
transform -1 0 670 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1342_
timestamp 1727493435
transform -1 0 570 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1343_
timestamp 1727493435
transform -1 0 430 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1344_
timestamp 1727493435
transform 1 0 630 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1345_
timestamp 1727493435
transform -1 0 190 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1346_
timestamp 1727493435
transform -1 0 530 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1347_
timestamp 1727493435
transform -1 0 310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1348_
timestamp 1727493435
transform -1 0 210 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1349_
timestamp 1727493435
transform 1 0 790 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1350_
timestamp 1727493435
transform 1 0 1750 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1351_
timestamp 1727493435
transform 1 0 1350 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1352_
timestamp 1727493435
transform -1 0 1490 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1353_
timestamp 1727493435
transform -1 0 70 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1354_
timestamp 1727493435
transform -1 0 70 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1355_
timestamp 1727493435
transform -1 0 370 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1356_
timestamp 1727493435
transform 1 0 350 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1357_
timestamp 1727493435
transform 1 0 190 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1358_
timestamp 1727493435
transform -1 0 70 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1359_
timestamp 1727493435
transform 1 0 210 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1360_
timestamp 1727493435
transform 1 0 470 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1361_
timestamp 1727493435
transform 1 0 1390 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1362_
timestamp 1727493435
transform -1 0 70 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1363_
timestamp 1727493435
transform -1 0 70 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1364_
timestamp 1727493435
transform -1 0 730 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1365_
timestamp 1727493435
transform -1 0 370 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1366_
timestamp 1727493435
transform -1 0 510 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1367_
timestamp 1727493435
transform 1 0 350 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1368_
timestamp 1727493435
transform -1 0 70 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1369_
timestamp 1727493435
transform 1 0 190 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1370_
timestamp 1727493435
transform 1 0 170 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1371_
timestamp 1727493435
transform 1 0 1290 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1372_
timestamp 1727493435
transform -1 0 70 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1373_
timestamp 1727493435
transform -1 0 210 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1374_
timestamp 1727493435
transform 1 0 50 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1375_
timestamp 1727493435
transform 1 0 210 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1376_
timestamp 1727493435
transform -1 0 990 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1377_
timestamp 1727493435
transform 1 0 1330 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1378_
timestamp 1727493435
transform 1 0 950 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1379_
timestamp 1727493435
transform -1 0 810 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1380_
timestamp 1727493435
transform 1 0 730 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1381_
timestamp 1727493435
transform -1 0 590 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1382_
timestamp 1727493435
transform 1 0 890 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1383_
timestamp 1727493435
transform -1 0 690 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1384_
timestamp 1727493435
transform -1 0 810 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1385_
timestamp 1727493435
transform 1 0 610 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1386_
timestamp 1727493435
transform 1 0 830 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1387_
timestamp 1727493435
transform -1 0 390 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1388_
timestamp 1727493435
transform 1 0 1050 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1389_
timestamp 1727493435
transform -1 0 930 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1390_
timestamp 1727493435
transform 1 0 1210 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1391_
timestamp 1727493435
transform 1 0 1830 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1392_
timestamp 1727493435
transform 1 0 1430 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1393_
timestamp 1727493435
transform -1 0 4290 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1394_
timestamp 1727493435
transform -1 0 530 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1395_
timestamp 1727493435
transform -1 0 530 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1396_
timestamp 1727493435
transform -1 0 650 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1397_
timestamp 1727493435
transform 1 0 510 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1398_
timestamp 1727493435
transform 1 0 350 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1399_
timestamp 1727493435
transform 1 0 670 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1400_
timestamp 1727493435
transform -1 0 4010 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1401_
timestamp 1727493435
transform 1 0 3990 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1402_
timestamp 1727493435
transform 1 0 4250 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1403_
timestamp 1727493435
transform 1 0 4130 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1404_
timestamp 1727493435
transform -1 0 4070 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1405_
timestamp 1727493435
transform -1 0 3790 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1406_
timestamp 1727493435
transform -1 0 3710 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1407_
timestamp 1727493435
transform 1 0 4110 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1408_
timestamp 1727493435
transform 1 0 4350 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1409_
timestamp 1727493435
transform 1 0 4490 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1410_
timestamp 1727493435
transform 1 0 4630 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1411_
timestamp 1727493435
transform 1 0 4510 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1412_
timestamp 1727493435
transform 1 0 4790 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1413_
timestamp 1727493435
transform -1 0 4670 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1414_
timestamp 1727493435
transform 1 0 4790 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1415_
timestamp 1727493435
transform -1 0 4830 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1416_
timestamp 1727493435
transform -1 0 3290 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1417_
timestamp 1727493435
transform -1 0 4210 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1418_
timestamp 1727493435
transform -1 0 4350 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1419_
timestamp 1727493435
transform 1 0 4170 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1420_
timestamp 1727493435
transform -1 0 3910 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1421_
timestamp 1727493435
transform -1 0 3050 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1422_
timestamp 1727493435
transform -1 0 2910 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1423_
timestamp 1727493435
transform -1 0 2710 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1424_
timestamp 1727493435
transform 1 0 2830 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1425_
timestamp 1727493435
transform 1 0 2950 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1426_
timestamp 1727493435
transform -1 0 3130 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1427_
timestamp 1727493435
transform 1 0 3110 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1428_
timestamp 1727493435
transform -1 0 2430 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1429_
timestamp 1727493435
transform -1 0 2550 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1430_
timestamp 1727493435
transform -1 0 2690 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1431_
timestamp 1727493435
transform 1 0 2730 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1432_
timestamp 1727493435
transform 1 0 2870 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1433_
timestamp 1727493435
transform 1 0 2810 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1434_
timestamp 1727493435
transform -1 0 2570 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1435_
timestamp 1727493435
transform 1 0 2750 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1436_
timestamp 1727493435
transform 1 0 2590 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1437_
timestamp 1727493435
transform -1 0 3010 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1438_
timestamp 1727493435
transform -1 0 5310 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1439_
timestamp 1727493435
transform 1 0 2950 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1440_
timestamp 1727493435
transform 1 0 3270 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1441_
timestamp 1727493435
transform -1 0 3570 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1442_
timestamp 1727493435
transform 1 0 3410 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1443_
timestamp 1727493435
transform -1 0 3870 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1444_
timestamp 1727493435
transform 1 0 4050 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1445_
timestamp 1727493435
transform 1 0 4650 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1446_
timestamp 1727493435
transform 1 0 5810 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1447_
timestamp 1727493435
transform 1 0 5670 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1448_
timestamp 1727493435
transform -1 0 5790 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1449_
timestamp 1727493435
transform -1 0 5670 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1450_
timestamp 1727493435
transform -1 0 4530 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1452_
timestamp 1727493435
transform -1 0 5810 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1453_
timestamp 1727493435
transform 1 0 5670 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1454_
timestamp 1727493435
transform 1 0 5750 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1455_
timestamp 1727493435
transform -1 0 5930 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1456_
timestamp 1727493435
transform 1 0 5850 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1457_
timestamp 1727493435
transform -1 0 5270 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1458_
timestamp 1727493435
transform -1 0 5370 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1459_
timestamp 1727493435
transform 1 0 5970 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1460_
timestamp 1727493435
transform 1 0 5970 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1461_
timestamp 1727493435
transform 1 0 5870 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1462_
timestamp 1727493435
transform -1 0 5850 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1463_
timestamp 1727493435
transform 1 0 5870 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1464_
timestamp 1727493435
transform -1 0 4970 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1465_
timestamp 1727493435
transform -1 0 5950 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1466_
timestamp 1727493435
transform 1 0 5950 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1467_
timestamp 1727493435
transform 1 0 5730 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1468_
timestamp 1727493435
transform -1 0 5590 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1469_
timestamp 1727493435
transform 1 0 5230 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1470_
timestamp 1727493435
transform 1 0 5650 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1471_
timestamp 1727493435
transform -1 0 5510 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1472_
timestamp 1727493435
transform -1 0 5270 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1473_
timestamp 1727493435
transform -1 0 5110 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1474_
timestamp 1727493435
transform 1 0 5130 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1475_
timestamp 1727493435
transform -1 0 5390 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1476_
timestamp 1727493435
transform 1 0 5410 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1477_
timestamp 1727493435
transform 1 0 5350 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1478_
timestamp 1727493435
transform -1 0 5150 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1479_
timestamp 1727493435
transform 1 0 2650 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1480_
timestamp 1727493435
transform 1 0 4190 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1481_
timestamp 1727493435
transform 1 0 3990 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1482_
timestamp 1727493435
transform 1 0 3830 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1483_
timestamp 1727493435
transform 1 0 2870 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1484_
timestamp 1727493435
transform 1 0 4430 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1485_
timestamp 1727493435
transform 1 0 4030 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1486_
timestamp 1727493435
transform -1 0 3310 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1487_
timestamp 1727493435
transform -1 0 4950 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1488_
timestamp 1727493435
transform 1 0 4770 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1489_
timestamp 1727493435
transform -1 0 3430 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1490_
timestamp 1727493435
transform -1 0 4830 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1491_
timestamp 1727493435
transform 1 0 4650 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1492_
timestamp 1727493435
transform -1 0 3550 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1493_
timestamp 1727493435
transform 1 0 3510 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1494_
timestamp 1727493435
transform 1 0 3110 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1495_
timestamp 1727493435
transform 1 0 3370 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1496_
timestamp 1727493435
transform 1 0 2970 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1497_
timestamp 1727493435
transform -1 0 3390 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1498_
timestamp 1727493435
transform 1 0 3210 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1499_
timestamp 1727493435
transform 1 0 2830 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1500_
timestamp 1727493435
transform -1 0 2690 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1501_
timestamp 1727493435
transform -1 0 2210 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1502_
timestamp 1727493435
transform 1 0 2330 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1503_
timestamp 1727493435
transform -1 0 2510 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1504_
timestamp 1727493435
transform -1 0 1790 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1505_
timestamp 1727493435
transform -1 0 2190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1506_
timestamp 1727493435
transform 1 0 1730 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1507_
timestamp 1727493435
transform -1 0 2050 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1508_
timestamp 1727493435
transform -1 0 1430 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1509_
timestamp 1727493435
transform -1 0 1590 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1510_
timestamp 1727493435
transform -1 0 2430 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1511_
timestamp 1727493435
transform -1 0 2570 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1512_
timestamp 1727493435
transform -1 0 2310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1513_
timestamp 1727493435
transform 1 0 2390 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1514_
timestamp 1727493435
transform -1 0 2690 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1515_
timestamp 1727493435
transform -1 0 2830 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1516_
timestamp 1727493435
transform -1 0 1610 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1517_
timestamp 1727493435
transform -1 0 1990 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1518_
timestamp 1727493435
transform -1 0 1330 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1519_
timestamp 1727493435
transform 1 0 1150 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1520_
timestamp 1727493435
transform 1 0 950 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1521_
timestamp 1727493435
transform -1 0 910 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1522_
timestamp 1727493435
transform -1 0 370 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1523_
timestamp 1727493435
transform -1 0 510 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1524_
timestamp 1727493435
transform 1 0 1450 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1525_
timestamp 1727493435
transform -1 0 1310 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1601_
timestamp 1727493435
transform 1 0 5950 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1602_
timestamp 1727493435
transform 1 0 5970 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1603_
timestamp 1727493435
transform 1 0 5630 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1604_
timestamp 1727493435
transform 1 0 5530 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1605_
timestamp 1727493435
transform 1 0 5830 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1606_
timestamp 1727493435
transform 1 0 4410 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1607_
timestamp 1727493435
transform 1 0 4550 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1608_
timestamp 1727493435
transform 1 0 4690 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1609_
timestamp 1727493435
transform 1 0 4270 0 -1 270
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert0
timestamp 1727493435
transform -1 0 1810 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert1
timestamp 1727493435
transform -1 0 1570 0 1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert2
timestamp 1727493435
transform 1 0 4970 0 -1 790
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert3
timestamp 1727493435
transform 1 0 3450 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert4
timestamp 1727493435
transform 1 0 2210 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert5
timestamp 1727493435
transform 1 0 1730 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert6
timestamp 1727493435
transform -1 0 3090 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert7
timestamp 1727493435
transform -1 0 4550 0 1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert16
timestamp 1727493435
transform -1 0 2110 0 -1 790
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert17
timestamp 1727493435
transform 1 0 2310 0 1 270
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert18
timestamp 1727493435
transform 1 0 2450 0 1 270
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert19
timestamp 1727493435
transform 1 0 4990 0 1 270
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert20
timestamp 1727493435
transform -1 0 4670 0 1 790
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert21
timestamp 1727493435
transform 1 0 4050 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert22
timestamp 1727493435
transform -1 0 1590 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert23
timestamp 1727493435
transform 1 0 2990 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert24
timestamp 1727493435
transform -1 0 2250 0 1 5470
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert25
timestamp 1727493435
transform 1 0 2930 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert26
timestamp 1727493435
transform -1 0 2610 0 1 3390
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert27
timestamp 1727493435
transform 1 0 770 0 1 3390
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert28
timestamp 1727493435
transform -1 0 2030 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert29
timestamp 1727493435
transform -1 0 2170 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert30
timestamp 1727493435
transform -1 0 1870 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert31
timestamp 1727493435
transform 1 0 1990 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert32
timestamp 1727493435
transform 1 0 4630 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert33
timestamp 1727493435
transform -1 0 4390 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert8
timestamp 1727493435
transform 1 0 2990 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert9
timestamp 1727493435
transform -1 0 1110 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert10
timestamp 1727493435
transform -1 0 2490 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert11
timestamp 1727493435
transform 1 0 5730 0 1 1830
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert12
timestamp 1727493435
transform -1 0 3790 0 1 1830
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert13
timestamp 1727493435
transform 1 0 4270 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert14
timestamp 1727493435
transform -1 0 2150 0 1 1830
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert15
timestamp 1727493435
transform -1 0 1410 0 -1 1310
box -6 -8 26 272
<< labels >>
flabel metal1 s 6077 2 6137 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -57 2 3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s 5476 6036 5484 6044 3 FreeSans 16 90 0 0 Cin[5]
port 2 nsew
flabel metal3 s 5436 6036 5444 6044 3 FreeSans 16 90 0 0 Cin[4]
port 3 nsew
flabel metal3 s 5376 6036 5384 6044 3 FreeSans 16 90 0 0 Cin[3]
port 4 nsew
flabel metal3 s 5336 6036 5344 6044 3 FreeSans 16 90 0 0 Cin[2]
port 5 nsew
flabel metal3 s 4096 6036 4104 6044 3 FreeSans 16 90 0 0 Cin[1]
port 6 nsew
flabel metal3 s 4056 6036 4064 6044 3 FreeSans 16 90 0 0 Cin[0]
port 7 nsew
flabel metal2 s -23 2737 -17 2743 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal2 s 6117 1697 6123 1703 3 FreeSans 16 0 0 0 Vld
port 9 nsew
flabel metal2 s -23 4077 -17 4083 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal2 s -23 4037 -17 4043 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal2 s -23 3777 -17 3783 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal2 s -23 3537 -17 3543 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal2 s 6117 5117 6123 5123 3 FreeSans 16 0 0 0 Xout[3]
port 14 nsew
flabel metal2 s 6117 5077 6123 5083 3 FreeSans 16 0 0 0 Xout[2]
port 15 nsew
flabel metal2 s 6117 4817 6123 4823 3 FreeSans 16 0 0 0 Xout[1]
port 16 nsew
flabel metal2 s 6117 3777 6123 3783 3 FreeSans 16 0 0 0 Xout[0]
port 17 nsew
flabel metal3 s 3456 -24 3464 -16 7 FreeSans 16 270 0 0 Yin[3]
port 18 nsew
flabel metal3 s 3336 -24 3344 -16 7 FreeSans 16 270 0 0 Yin[2]
port 19 nsew
flabel metal3 s 2916 -24 2924 -16 7 FreeSans 16 270 0 0 Yin[1]
port 20 nsew
flabel metal3 s 2696 -24 2704 -16 7 FreeSans 16 270 0 0 Yin[0]
port 21 nsew
flabel metal3 s 4776 -24 4784 -16 7 FreeSans 16 270 0 0 Yout[3]
port 22 nsew
flabel metal3 s 4736 -24 4744 -16 7 FreeSans 16 270 0 0 Yout[2]
port 23 nsew
flabel metal3 s 4596 -24 4604 -16 7 FreeSans 16 270 0 0 Yout[1]
port 24 nsew
flabel metal3 s 4456 -24 4464 -16 7 FreeSans 16 270 0 0 Yout[0]
port 25 nsew
flabel metal3 s 1316 6036 1324 6044 3 FreeSans 16 90 0 0 clk
port 26 nsew
<< properties >>
string FIXED_BBOX -40 -40 6120 6040
<< end >>
