magic
tech scmos
magscale 1 2
timestamp 1727399082
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
<< ptransistor >>
rect 26 166 30 246
rect 34 166 38 246
rect 56 206 60 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 42 40 54
rect 24 14 26 42
rect 38 14 40 42
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
<< pdiffusion >>
rect 24 166 26 246
rect 30 166 34 246
rect 38 166 40 246
rect 52 206 56 246
rect 60 206 62 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 42
rect 46 14 58 54
rect 66 14 78 54
<< pdcontact >>
rect 12 166 24 246
rect 40 166 52 246
rect 62 206 74 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 26 246 30 250
rect 34 246 38 250
rect 56 246 60 250
rect 26 162 30 166
rect 12 154 30 162
rect 12 109 16 154
rect 34 123 38 166
rect 56 162 60 206
rect 56 154 66 162
rect 60 123 66 154
rect 36 111 44 123
rect 12 66 16 97
rect 12 59 24 66
rect 20 54 24 59
rect 40 54 44 111
rect 60 54 64 123
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
<< polycontact >>
rect 24 111 36 123
rect 4 97 16 109
rect 64 111 76 123
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 12 246 24 252
rect 62 246 74 252
rect 23 123 37 137
rect 43 97 51 166
rect 63 123 77 137
rect 3 83 17 97
rect 43 83 57 97
rect 49 75 57 83
rect 49 68 74 75
rect 6 54 58 57
rect 18 48 46 54
rect 66 54 74 68
rect 26 8 38 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect 23 123 37 137
rect 63 123 77 137
rect 3 83 17 97
rect 43 83 57 97
<< labels >>
rlabel metal1 23 123 37 137 0 B
port 1 nsew signal input
rlabel metal1 -6 252 106 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal1 43 83 57 97 0 Y
port 3 nsew signal output
rlabel metal1 63 123 77 137 0 C
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
