magic
tech scmos
magscale 1 2
timestamp 1749781196
<< checkpaint >>
rect -40 -40 331 707
<< metal1 >>
rect 0 0 32 667
rect 257 0 291 667
<< metal2 >>
rect 87 622 101 667
rect 127 591 141 616
rect 87 579 141 591
rect 87 552 101 579
rect 127 520 141 546
rect 87 508 141 520
rect 87 482 101 508
rect 127 451 141 476
rect 87 439 141 451
rect 87 413 101 439
rect 127 381 141 406
rect 87 369 141 381
rect 87 342 101 369
rect 127 310 141 336
rect 87 298 141 310
rect 87 272 101 298
rect 127 240 141 266
rect 87 228 141 240
rect 87 202 101 228
rect 127 171 141 196
rect 87 159 141 171
rect 87 132 101 159
rect 127 103 141 126
rect 87 91 141 103
rect 87 62 101 91
rect 127 0 141 56
<< m2p >>
rect 87 622 101 667
rect 87 579 141 591
rect 87 508 141 520
rect 127 0 141 56
use INVX1  INVX1_0 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1749781103
transform 0 1 24 -1 0 79
box -12 -8 72 252
use INVX1  INVX1_1
timestamp 1749781103
transform 0 1 24 -1 0 149
box -12 -8 72 252
use INVX1  INVX1_2
timestamp 1749781103
transform 0 1 24 -1 0 219
box -12 -8 72 252
use INVX1  INVX1_3
timestamp 1749781103
transform 0 1 24 -1 0 289
box -12 -8 72 252
use INVX1  INVX1_4
timestamp 1749781103
transform 0 1 24 -1 0 359
box -12 -8 72 252
use INVX1  INVX1_5
timestamp 1749781103
transform 0 1 24 -1 0 429
box -12 -8 72 252
use INVX1  INVX1_6
timestamp 1749781103
transform 0 1 24 -1 0 499
box -12 -8 72 252
use INVX1  INVX1_7
timestamp 1749781103
transform 0 1 24 -1 0 569
box -12 -8 72 252
use INVX1  INVX1_8
timestamp 1749781103
transform 0 1 24 -1 0 639
box -12 -8 72 252
<< labels >>
rlabel metal1 0 0 32 32 0 gnd
port 2 nsew ground bidirectional abutment
rlabel metal2 87 622 101 667 0 In
port 3 nsew signal input
rlabel metal2 87 579 141 591 0 Out1
port 4 nsew signal output
rlabel metal2 87 508 141 520 0 Out2
port 5 nsew signal output
rlabel metal2 127 0 141 56 0 Out3
port 6 nsew signal output
rlabel metal1 257 0 291 34 0 vdd
port 1 nsew power bidirectional abutment
<< end >>
