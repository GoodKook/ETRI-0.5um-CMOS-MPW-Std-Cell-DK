magic
tech scmos
magscale 1 6
timestamp 1555589239
<< checkpaint >>
rect -122 -178 218 530
<< ntransistor >>
rect 43 0 53 400
<< ndiffusion >>
rect 0 0 43 400
rect 53 0 96 400
<< polysilicon >>
rect 43 400 53 410
rect 43 -24 53 0
<< metal1 >>
rect -2 -2 40 402
rect 56 -2 98 402
use CONT  CONT_0
array 0 0 0 0 6 56
timestamp 1555589239
transform 1 0 78 0 1 20
box -6 -6 6 6
use CONT  CONT_1
array 0 0 0 0 6 56
timestamp 1555589239
transform 1 0 18 0 1 20
box -6 -6 6 6
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_0
timestamp 1555589239
transform -1 0 66 0 -1 -22
box 0 0 36 36
<< end >>
