magic
tech scmos
magscale 1 2
timestamp 1702345906
<< nwell >>
rect -13 194 474 272
<< ntransistor >>
rect 24 14 28 54
rect 36 14 40 54
rect 60 14 64 54
rect 72 14 76 54
rect 122 14 126 34
rect 142 14 146 34
rect 162 14 166 34
rect 213 14 217 34
rect 233 14 237 34
rect 273 14 277 34
rect 293 14 297 34
rect 342 14 346 54
rect 354 14 358 54
rect 377 14 381 54
rect 389 14 393 54
rect 434 14 438 34
<< ptransistor >>
rect 22 206 26 246
rect 42 206 46 246
rect 62 206 66 246
rect 82 206 86 246
rect 126 226 130 246
rect 146 226 150 246
rect 166 206 170 246
rect 213 206 217 246
rect 233 206 237 246
rect 273 226 277 246
rect 293 226 297 246
rect 333 206 337 246
rect 353 206 357 246
rect 373 206 377 246
rect 393 206 397 246
rect 434 206 438 246
<< ndiffusion >>
rect 20 14 24 54
rect 28 14 36 54
rect 40 14 44 54
rect 56 14 60 54
rect 64 14 72 54
rect 76 14 80 54
rect 120 14 122 34
rect 126 14 128 34
rect 140 14 142 34
rect 146 14 148 34
rect 160 14 162 34
rect 166 14 168 34
rect 211 14 213 34
rect 217 14 219 34
rect 231 14 233 34
rect 237 14 239 34
rect 271 14 273 34
rect 277 14 279 34
rect 291 14 293 34
rect 297 14 299 34
rect 338 14 342 54
rect 346 14 354 54
rect 358 14 361 54
rect 373 14 377 54
rect 381 14 389 54
rect 393 14 397 54
rect 432 14 434 34
rect 438 14 440 34
<< pdiffusion >>
rect 20 206 22 246
rect 26 206 28 246
rect 40 206 42 246
rect 46 206 48 246
rect 60 206 62 246
rect 66 206 68 246
rect 80 206 82 246
rect 86 206 88 246
rect 124 227 126 246
rect 112 226 126 227
rect 130 226 132 246
rect 144 226 146 246
rect 150 226 152 246
rect 164 206 166 246
rect 170 206 172 246
rect 211 206 213 246
rect 217 206 219 246
rect 231 206 233 246
rect 237 206 239 246
rect 271 226 273 246
rect 277 226 279 246
rect 291 226 293 246
rect 297 226 299 246
rect 331 206 333 246
rect 337 206 339 246
rect 351 206 353 246
rect 357 206 359 246
rect 371 206 373 246
rect 377 206 379 246
rect 391 206 393 246
rect 397 206 399 246
rect 432 206 434 246
rect 438 206 440 246
<< ndcontact >>
rect 8 14 20 54
rect 44 14 56 54
rect 80 14 92 54
rect 108 14 120 34
rect 128 14 140 34
rect 148 14 160 34
rect 168 14 180 34
rect 199 14 211 34
rect 219 14 231 34
rect 239 14 251 34
rect 259 14 271 34
rect 279 14 291 34
rect 299 14 311 34
rect 326 14 338 54
rect 361 14 373 54
rect 397 14 409 54
rect 420 14 432 34
rect 440 14 452 34
<< pdcontact >>
rect 8 206 20 246
rect 28 206 40 246
rect 48 206 60 246
rect 68 206 80 246
rect 88 206 100 246
rect 112 227 124 246
rect 132 226 144 246
rect 152 206 164 246
rect 172 206 184 246
rect 199 206 211 246
rect 219 206 231 246
rect 239 206 251 246
rect 259 226 271 246
rect 279 226 291 246
rect 299 226 311 246
rect 319 206 331 246
rect 339 206 351 246
rect 359 206 371 246
rect 379 206 391 246
rect 399 206 411 246
rect 420 206 432 246
rect 440 206 452 246
<< psubstratepcontact >>
rect -6 -6 466 6
<< nsubstratencontact >>
rect -6 254 466 266
<< polysilicon >>
rect 22 246 26 250
rect 42 246 46 250
rect 62 246 66 250
rect 82 246 86 250
rect 126 246 130 250
rect 146 246 150 250
rect 166 246 170 250
rect 213 246 217 250
rect 233 246 237 250
rect 273 246 277 250
rect 293 246 297 250
rect 333 246 337 250
rect 353 246 357 250
rect 373 246 377 250
rect 393 246 397 250
rect 434 246 438 250
rect 22 115 26 206
rect 42 188 46 206
rect 22 103 24 115
rect 24 54 28 103
rect 44 72 48 176
rect 62 172 66 206
rect 36 54 40 60
rect 60 54 64 160
rect 82 118 86 206
rect 84 106 86 118
rect 82 85 86 106
rect 126 99 130 226
rect 146 133 150 226
rect 72 81 86 85
rect 72 54 76 81
rect 146 79 150 121
rect 122 75 150 79
rect 122 34 126 75
rect 166 74 170 206
rect 213 147 217 206
rect 233 166 237 206
rect 273 192 277 226
rect 257 180 277 192
rect 233 159 252 166
rect 213 135 225 147
rect 166 73 182 74
rect 162 62 182 73
rect 142 34 146 54
rect 162 34 166 62
rect 213 54 217 135
rect 245 119 252 159
rect 233 112 252 119
rect 233 74 237 112
rect 273 111 277 180
rect 293 144 297 226
rect 333 194 337 206
rect 297 132 311 138
rect 273 105 297 111
rect 186 47 217 54
rect 213 34 217 47
rect 233 34 237 62
rect 273 34 277 54
rect 293 34 297 105
rect 305 66 311 132
rect 325 60 331 188
rect 353 166 357 206
rect 373 195 377 206
rect 372 192 377 195
rect 337 161 357 166
rect 337 147 342 161
rect 337 135 339 147
rect 372 137 377 180
rect 393 161 397 206
rect 337 68 342 135
rect 363 131 377 137
rect 363 88 368 131
rect 392 116 397 149
rect 364 76 368 88
rect 337 64 358 68
rect 325 56 346 60
rect 342 54 346 56
rect 354 54 358 64
rect 363 60 368 76
rect 372 111 397 116
rect 372 68 377 111
rect 434 88 438 206
rect 397 76 438 88
rect 372 64 393 68
rect 363 56 381 60
rect 377 54 381 56
rect 389 54 393 64
rect 434 34 438 76
rect 24 10 28 14
rect 36 10 40 14
rect 60 10 64 14
rect 72 10 76 14
rect 122 10 126 14
rect 142 10 146 14
rect 162 10 166 14
rect 213 10 217 14
rect 233 10 237 14
rect 273 10 277 14
rect 293 10 297 14
rect 342 10 346 14
rect 354 10 358 14
rect 377 10 381 14
rect 389 10 393 14
rect 434 10 438 14
<< polycontact >>
rect 38 176 50 188
rect 24 103 36 115
rect 36 60 48 72
rect 60 160 72 172
rect 72 106 84 118
rect 146 121 158 133
rect 126 87 138 99
rect 245 180 257 192
rect 225 135 237 147
rect 142 54 154 66
rect 182 62 194 74
rect 321 188 333 200
rect 285 132 297 144
rect 225 62 237 74
rect 174 41 186 54
rect 273 54 285 66
rect 305 54 317 66
rect 365 180 377 192
rect 339 135 351 147
rect 385 149 397 161
rect 352 76 364 88
rect 385 76 397 88
<< metal1 >>
rect -6 266 466 268
rect -6 252 466 254
rect 8 246 20 252
rect 48 246 60 252
rect 88 246 100 252
rect 172 246 184 252
rect 219 246 231 252
rect 319 246 331 252
rect 359 246 370 252
rect 399 246 411 252
rect 440 246 452 252
rect 26 206 28 212
rect 26 200 32 206
rect 8 194 32 200
rect 8 87 16 194
rect 68 186 80 206
rect 199 197 211 206
rect 50 179 166 186
rect 199 183 203 197
rect 239 180 245 206
rect 293 192 321 200
rect 339 187 346 206
rect 383 200 391 206
rect 383 194 409 200
rect 420 194 432 206
rect 159 174 166 179
rect 72 160 126 168
rect 159 167 263 174
rect 339 180 365 187
rect 403 174 409 194
rect 313 167 409 174
rect 159 154 385 161
rect 159 149 166 154
rect 93 142 166 149
rect 23 123 37 137
rect 63 123 77 137
rect 24 115 36 123
rect 68 118 77 123
rect 93 118 100 142
rect 158 125 203 129
rect 285 128 297 132
rect 217 125 297 128
rect 158 121 297 125
rect 315 135 339 147
rect 68 106 72 118
rect 84 111 100 118
rect 315 115 321 135
rect 113 108 321 115
rect 29 100 36 103
rect 113 100 120 108
rect 29 93 120 100
rect 8 78 106 87
rect 8 54 16 78
rect 48 60 92 68
rect 82 54 92 60
rect 126 66 132 87
rect 183 83 197 97
rect 223 83 237 97
rect 183 74 194 83
rect 126 59 142 66
rect 154 59 174 66
rect 225 74 237 83
rect 345 76 352 88
rect 364 76 385 88
rect 168 47 174 59
rect 285 54 305 66
rect 345 54 355 76
rect 403 54 409 167
rect 199 40 203 54
rect 199 34 211 40
rect 338 46 355 54
rect 423 137 432 194
rect 423 123 437 137
rect 423 34 432 123
rect 44 8 56 14
rect 168 8 180 14
rect 219 8 231 14
rect 361 8 373 14
rect 440 8 452 14
rect -6 6 466 8
rect -6 -8 466 -6
<< m2contact >>
rect 112 213 126 227
rect 132 212 146 226
rect 259 212 273 226
rect 279 212 293 226
rect 299 212 313 226
rect 148 192 162 206
rect 203 183 217 197
rect 245 192 259 206
rect 279 192 293 206
rect 126 158 140 172
rect 263 167 277 181
rect 299 167 313 181
rect 203 125 217 139
rect 237 134 251 148
rect 106 73 120 87
rect 108 34 122 48
rect 128 34 142 48
rect 148 34 162 48
rect 203 40 217 54
rect 239 34 253 48
rect 259 34 273 48
rect 279 34 293 48
rect 299 34 313 48
<< metal2 >>
rect 106 213 112 227
rect 106 87 116 213
rect 132 172 140 212
rect 108 48 117 73
rect 132 48 140 158
rect 148 48 156 192
rect 206 139 213 183
rect 245 148 253 192
rect 265 181 273 212
rect 279 206 293 212
rect 251 134 253 148
rect 206 54 213 125
rect 245 48 253 134
rect 265 48 273 167
rect 285 48 293 192
rect 299 181 308 212
rect 299 48 308 167
<< m1p >>
rect -6 252 466 268
rect 23 123 37 137
rect 63 123 77 137
rect 423 123 437 137
rect 183 83 197 97
rect 223 83 237 97
rect -6 -8 466 8
<< labels >>
rlabel nsubstratencontact 230 260 230 260 0 vdd
port 6 nsew power bidirectional abutment
rlabel psubstratepcontact 230 0 230 0 0 gnd
port 7 nsew ground bidirectional abutment
rlabel metal1 430 131 430 131 0 Q
port 5 nsew signal output
rlabel metal1 30 130 30 130 0 R
port 3 nsew signal input
rlabel metal1 69 131 69 131 0 S
port 2 nsew signal input
rlabel metal1 231 91 231 91 0 CLK
port 4 nsew clock input
rlabel metal1 190 91 190 91 0 D
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 460 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
