magic
tech scmos
magscale 1 2
timestamp 1726639203
<< checkpaint >>
rect 3015 5567 3106 5576
rect 3192 5567 3296 5568
rect -103 -64 5863 5567
<< nwell >>
rect 655 5113 727 5127
<< metal1 >>
rect -63 5218 -3 5478
rect 5730 5462 5823 5478
rect 2807 5397 2873 5403
rect 3787 5397 3813 5403
rect 297 5377 333 5383
rect 297 5343 303 5377
rect 3627 5383 3640 5387
rect 3627 5373 3643 5383
rect 3637 5347 3643 5373
rect 277 5340 303 5343
rect 273 5337 303 5340
rect 273 5327 287 5337
rect 687 5337 733 5343
rect 3627 5337 3643 5347
rect 3627 5333 3640 5337
rect 3947 5337 3973 5343
rect 127 5317 233 5323
rect 3067 5317 3153 5323
rect 3307 5317 3433 5323
rect 3787 5317 3833 5323
rect 4967 5317 5013 5323
rect 3307 5297 3333 5303
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 2787 5137 2853 5143
rect 3227 5137 3253 5143
rect 2407 5117 2493 5123
rect 627 5097 673 5103
rect 1917 5097 1953 5103
rect 547 5083 560 5087
rect 920 5083 933 5087
rect 547 5073 563 5083
rect 557 5047 563 5073
rect 917 5073 933 5083
rect 1917 5083 1923 5097
rect 2107 5097 2173 5103
rect 2387 5097 2423 5103
rect 1877 5077 1923 5083
rect 2417 5083 2423 5097
rect 2647 5097 2693 5103
rect 3047 5097 3113 5103
rect 3947 5097 3993 5103
rect 4707 5100 4743 5103
rect 4707 5097 4747 5100
rect 2417 5077 2463 5083
rect 917 5047 923 5073
rect 1877 5047 1883 5077
rect 547 5037 563 5047
rect 547 5033 560 5037
rect 907 5037 923 5047
rect 907 5033 920 5037
rect 1867 5037 1883 5047
rect 2457 5047 2463 5077
rect 2547 5077 2573 5083
rect 2817 5077 2853 5083
rect 2817 5047 2823 5077
rect 3397 5047 3403 5093
rect 2457 5037 2473 5047
rect 1867 5033 1880 5037
rect 2460 5033 2473 5037
rect 2817 5037 2833 5047
rect 2820 5033 2833 5037
rect 3387 5037 3403 5047
rect 3387 5033 3400 5037
rect 3677 5043 3683 5093
rect 3817 5077 3839 5083
rect 3817 5047 3823 5077
rect 3947 5077 3973 5083
rect 4227 5077 4253 5083
rect 4327 5083 4340 5087
rect 4327 5073 4343 5083
rect 4733 5086 4747 5097
rect 5487 5097 5573 5103
rect 4567 5077 4603 5083
rect 3647 5037 3683 5043
rect 3807 5037 3823 5047
rect 3807 5033 3820 5037
rect 3347 5017 3413 5023
rect 4337 5023 4343 5073
rect 4597 5047 4603 5077
rect 4960 5083 4973 5087
rect 4957 5073 4973 5083
rect 5500 5083 5513 5087
rect 5497 5073 5513 5083
rect 4957 5047 4963 5073
rect 5497 5047 5503 5073
rect 4597 5037 4613 5047
rect 4600 5033 4613 5037
rect 4947 5037 4963 5047
rect 4947 5033 4960 5037
rect 5227 5037 5253 5043
rect 5497 5037 5513 5047
rect 5500 5033 5513 5037
rect 4307 5017 4343 5023
rect 4827 5017 4853 5023
rect 5763 4958 5823 5462
rect 5730 4942 5823 4958
rect 1527 4877 1573 4883
rect 460 4863 473 4867
rect 457 4853 473 4863
rect 707 4857 743 4863
rect 457 4823 463 4853
rect 427 4817 463 4823
rect 737 4827 743 4857
rect 1107 4863 1120 4867
rect 1107 4853 1123 4863
rect 2727 4863 2740 4867
rect 2727 4853 2743 4863
rect 3407 4857 3433 4863
rect 3767 4863 3780 4867
rect 4640 4863 4653 4867
rect 3767 4853 3783 4863
rect 1117 4827 1123 4853
rect 1667 4843 1680 4847
rect 1667 4833 1683 4843
rect 1677 4827 1683 4833
rect 737 4817 753 4827
rect 740 4813 753 4817
rect 1117 4817 1133 4827
rect 1120 4813 1133 4817
rect 1677 4817 1693 4827
rect 1680 4813 1693 4817
rect 2737 4823 2743 4853
rect 3777 4827 3783 4853
rect 4637 4853 4653 4863
rect 4637 4827 4643 4853
rect 2737 4817 2773 4823
rect 3147 4817 3213 4823
rect 3777 4817 3793 4827
rect 3780 4813 3793 4817
rect 3947 4817 3973 4823
rect 4347 4817 4383 4823
rect 4627 4817 4643 4827
rect 4627 4813 4640 4817
rect 5207 4817 5233 4823
rect 581 4797 653 4803
rect 1467 4797 1553 4803
rect 1947 4797 1973 4803
rect 2447 4803 2460 4807
rect 2447 4793 2463 4803
rect 3767 4797 3853 4803
rect 2457 4783 2463 4793
rect 4287 4797 4353 4803
rect 5567 4797 5633 4803
rect 2457 4777 2513 4783
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 647 4577 693 4583
rect 2607 4577 2693 4583
rect 3547 4577 3573 4583
rect 627 4563 640 4567
rect 627 4553 643 4563
rect 637 4543 643 4553
rect 887 4557 933 4563
rect 1167 4557 1213 4563
rect 2280 4563 2293 4567
rect 2277 4553 2293 4563
rect 2787 4563 2800 4567
rect 2787 4553 2803 4563
rect 3167 4563 3180 4567
rect 3320 4563 3333 4567
rect 3167 4553 3183 4563
rect 637 4537 663 4543
rect 657 4527 663 4537
rect 2277 4527 2283 4553
rect 2797 4527 2803 4553
rect 657 4517 673 4527
rect 660 4513 673 4517
rect 2277 4517 2293 4527
rect 2280 4513 2293 4517
rect 2787 4517 2803 4527
rect 3177 4527 3183 4553
rect 3317 4553 3333 4563
rect 3407 4557 3443 4563
rect 3317 4527 3323 4553
rect 3177 4517 3193 4527
rect 2787 4513 2800 4517
rect 3180 4513 3193 4517
rect 3307 4517 3323 4527
rect 3437 4527 3443 4557
rect 3567 4557 3593 4563
rect 4257 4557 4303 4563
rect 4577 4557 4613 4563
rect 4297 4527 4303 4557
rect 3437 4517 3453 4527
rect 3307 4513 3320 4517
rect 3440 4513 3453 4517
rect 4297 4517 4313 4527
rect 4300 4513 4313 4517
rect 367 4497 393 4503
rect 3667 4497 3713 4503
rect 5763 4438 5823 4942
rect 5730 4422 5823 4438
rect 107 4357 153 4363
rect 687 4357 713 4363
rect 3997 4357 4019 4363
rect 527 4343 540 4347
rect 527 4333 543 4343
rect 667 4337 693 4343
rect 1280 4343 1293 4347
rect 1277 4333 1293 4343
rect 2200 4343 2213 4347
rect 2197 4333 2213 4343
rect 2400 4343 2413 4347
rect 2397 4333 2413 4343
rect 2880 4343 2893 4347
rect 2877 4333 2893 4343
rect 3407 4343 3420 4347
rect 3407 4333 3423 4343
rect 3827 4343 3840 4347
rect 3997 4343 4003 4357
rect 4100 4363 4113 4367
rect 4097 4357 4113 4363
rect 4100 4353 4113 4357
rect 4127 4357 4153 4363
rect 3827 4333 3843 4343
rect 537 4307 543 4333
rect 1277 4307 1283 4333
rect 527 4297 543 4307
rect 527 4293 540 4297
rect 1127 4297 1153 4303
rect 1267 4297 1283 4307
rect 2197 4307 2203 4333
rect 2397 4307 2403 4333
rect 2197 4297 2213 4307
rect 1267 4293 1280 4297
rect 2200 4293 2213 4297
rect 2387 4297 2403 4307
rect 2877 4307 2883 4333
rect 2877 4297 2893 4307
rect 2387 4293 2400 4297
rect 2880 4293 2893 4297
rect 1347 4277 1433 4283
rect 1627 4277 1713 4283
rect 3417 4286 3423 4333
rect 3517 4300 3573 4303
rect 3513 4297 3573 4300
rect 3513 4287 3527 4297
rect 3837 4303 3843 4333
rect 3977 4337 4003 4343
rect 3977 4307 3983 4337
rect 5027 4343 5040 4347
rect 5027 4333 5043 4343
rect 5167 4343 5180 4347
rect 5167 4333 5183 4343
rect 3807 4297 3873 4303
rect 3967 4297 3983 4307
rect 3967 4293 3980 4297
rect 4107 4297 4153 4303
rect 4247 4297 4273 4303
rect 4507 4297 4553 4303
rect 5037 4303 5043 4333
rect 5017 4300 5043 4303
rect 5013 4297 5043 4300
rect 5177 4303 5183 4333
rect 5177 4297 5213 4303
rect 5013 4287 5027 4297
rect 5067 4277 5113 4283
rect 1367 4257 1393 4263
rect 5307 4257 5333 4263
rect 5267 4237 5313 4243
rect 5327 4237 5353 4243
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 587 4077 633 4083
rect 107 4057 233 4063
rect 617 4057 653 4063
rect 617 4043 623 4057
rect 967 4057 1013 4063
rect 1867 4057 1953 4063
rect 2987 4057 3033 4063
rect 3347 4057 3373 4063
rect 740 4043 753 4047
rect 577 4037 623 4043
rect 577 4007 583 4037
rect 567 3997 583 4007
rect 737 4033 753 4043
rect 2007 4043 2020 4047
rect 2040 4043 2053 4047
rect 2007 4033 2023 4043
rect 737 4006 743 4033
rect 2017 4007 2023 4033
rect 567 3993 580 3997
rect 2007 3997 2023 4007
rect 2037 4033 2053 4043
rect 2180 4043 2193 4047
rect 2177 4033 2193 4043
rect 2460 4043 2473 4047
rect 2457 4033 2473 4043
rect 2587 4037 2613 4043
rect 3140 4043 3153 4047
rect 3137 4033 3153 4043
rect 3257 4037 3293 4043
rect 2037 4007 2043 4033
rect 2177 4007 2183 4033
rect 2037 3997 2053 4007
rect 2007 3993 2020 3997
rect 2040 3993 2053 3997
rect 2177 3997 2193 4007
rect 2180 3993 2193 3997
rect 2457 3987 2463 4033
rect 3137 4007 3143 4033
rect 3257 4007 3263 4037
rect 3397 4043 3403 4073
rect 3607 4057 3633 4063
rect 3727 4057 3793 4063
rect 4067 4057 4113 4063
rect 3860 4043 3873 4047
rect 3377 4037 3403 4043
rect 3377 4007 3383 4037
rect 3857 4033 3873 4043
rect 3977 4037 4013 4043
rect 3857 4007 3863 4033
rect 3137 3997 3153 4007
rect 3140 3993 3153 3997
rect 3257 3997 3273 4007
rect 3260 3993 3273 3997
rect 3367 3997 3383 4007
rect 3367 3993 3380 3997
rect 3847 3997 3863 4007
rect 3977 4007 3983 4037
rect 4327 4043 4340 4047
rect 4360 4043 4373 4047
rect 4327 4033 4343 4043
rect 4337 4007 4343 4033
rect 3977 3997 3993 4007
rect 3847 3993 3860 3997
rect 3980 3993 3993 3997
rect 4327 3997 4343 4007
rect 4357 4033 4373 4043
rect 5007 4037 5033 4043
rect 5247 4037 5283 4043
rect 4357 4007 4363 4033
rect 5277 4007 5283 4037
rect 4357 3997 4373 4007
rect 4327 3993 4340 3997
rect 4360 3993 4373 3997
rect 5277 3997 5293 4007
rect 5280 3993 5293 3997
rect 4607 3977 4633 3983
rect 5763 3918 5823 4422
rect 5730 3902 5823 3918
rect 967 3837 1033 3843
rect 2387 3837 2433 3843
rect 3647 3837 3673 3843
rect 667 3823 680 3827
rect 820 3823 833 3827
rect 667 3813 683 3823
rect 677 3787 683 3813
rect 817 3813 833 3823
rect 1780 3823 1793 3827
rect 1087 3817 1123 3823
rect 817 3787 823 3813
rect 1117 3787 1123 3817
rect 1777 3813 1793 3823
rect 1880 3823 1893 3827
rect 1877 3813 1893 3823
rect 2127 3823 2140 3827
rect 2640 3823 2653 3827
rect 2127 3813 2143 3823
rect 677 3777 693 3787
rect 680 3773 693 3777
rect 817 3777 833 3787
rect 820 3773 833 3777
rect 967 3777 993 3783
rect 1117 3777 1133 3787
rect 1120 3773 1133 3777
rect 1513 3783 1527 3793
rect 1777 3787 1783 3813
rect 1877 3787 1883 3813
rect 1487 3780 1527 3783
rect 1487 3777 1523 3780
rect 1627 3777 1659 3783
rect 1727 3777 1753 3783
rect 1777 3777 1793 3787
rect 1780 3773 1793 3777
rect 1877 3777 1893 3787
rect 1880 3773 1893 3777
rect 1187 3757 1253 3763
rect 2137 3763 2143 3813
rect 2637 3813 2653 3823
rect 3747 3823 3760 3827
rect 3747 3813 3763 3823
rect 2637 3787 2643 3813
rect 2627 3777 2643 3787
rect 2627 3773 2640 3777
rect 3757 3783 3763 3813
rect 3727 3777 3763 3783
rect 3873 3783 3887 3793
rect 3873 3780 3913 3783
rect 3877 3777 3913 3780
rect 3997 3783 4003 3833
rect 3967 3777 4003 3783
rect 4157 3787 4163 3813
rect 4397 3787 4403 3833
rect 5540 3823 5553 3827
rect 4157 3777 4173 3787
rect 4160 3773 4173 3777
rect 4387 3777 4403 3787
rect 5537 3813 5553 3823
rect 5537 3787 5543 3813
rect 5537 3777 5553 3787
rect 4387 3773 4400 3777
rect 5540 3773 5553 3777
rect 2137 3757 2173 3763
rect 4407 3737 4473 3743
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 2827 3557 2873 3563
rect 107 3537 193 3543
rect 807 3537 833 3543
rect 2467 3537 2493 3543
rect 2720 3546 2740 3547
rect 2697 3537 2713 3543
rect 40 3523 53 3527
rect 37 3513 53 3523
rect 307 3517 333 3523
rect 947 3523 960 3527
rect 947 3513 963 3523
rect 1397 3517 1433 3523
rect 37 3487 43 3513
rect 957 3487 963 3513
rect 1097 3487 1103 3513
rect 1397 3487 1403 3517
rect 1820 3523 1833 3527
rect 1817 3513 1833 3523
rect 2027 3517 2073 3523
rect 2173 3523 2187 3533
rect 2173 3520 2203 3523
rect 2177 3517 2203 3520
rect 1817 3487 1823 3513
rect 37 3477 53 3487
rect 40 3473 53 3477
rect 957 3477 973 3487
rect 960 3473 973 3477
rect 1087 3477 1103 3487
rect 1087 3473 1100 3477
rect 1387 3477 1403 3487
rect 1387 3473 1400 3477
rect 1807 3477 1823 3487
rect 2197 3483 2203 3517
rect 2447 3523 2460 3527
rect 2447 3513 2463 3523
rect 2457 3487 2463 3513
rect 2197 3477 2233 3483
rect 1807 3473 1820 3477
rect 2447 3477 2463 3487
rect 2697 3487 2703 3537
rect 2727 3543 2740 3546
rect 2727 3537 2743 3543
rect 2727 3533 2740 3537
rect 2847 3517 2873 3523
rect 3237 3487 3243 3533
rect 3467 3523 3480 3527
rect 3467 3513 3483 3523
rect 2697 3477 2713 3487
rect 2447 3473 2460 3477
rect 2700 3473 2713 3477
rect 3237 3477 3253 3487
rect 3240 3473 3253 3477
rect 547 3457 593 3463
rect 667 3457 753 3463
rect 3477 3463 3483 3513
rect 4337 3487 4343 3533
rect 4460 3523 4473 3527
rect 4457 3513 4473 3523
rect 4900 3523 4913 3527
rect 4897 3513 4913 3523
rect 5040 3523 5053 3527
rect 5037 3517 5053 3523
rect 5040 3513 5053 3517
rect 5537 3517 5593 3523
rect 4457 3487 4463 3513
rect 4897 3487 4903 3513
rect 3607 3477 3633 3483
rect 4337 3477 4353 3487
rect 4340 3473 4353 3477
rect 4457 3477 4473 3487
rect 4460 3473 4473 3477
rect 4887 3477 4903 3487
rect 4887 3473 4900 3477
rect 3477 3457 3513 3463
rect 4587 3457 4613 3463
rect 5717 3446 5723 3533
rect 2207 3417 2233 3423
rect 5763 3398 5823 3902
rect 5730 3382 5823 3398
rect 1827 3337 1873 3343
rect 3847 3337 3893 3343
rect 207 3317 233 3323
rect 1847 3317 1893 3323
rect 4827 3317 4873 3323
rect 4980 3323 4993 3327
rect 4977 3313 4993 3323
rect 647 3303 660 3307
rect 1280 3303 1293 3307
rect 647 3293 663 3303
rect 657 3267 663 3293
rect 1277 3293 1293 3303
rect 1387 3303 1400 3307
rect 1700 3303 1713 3307
rect 1387 3293 1403 3303
rect 647 3257 663 3267
rect 647 3253 660 3257
rect 1107 3257 1133 3263
rect 1277 3266 1283 3293
rect 1397 3267 1403 3293
rect 1387 3257 1403 3267
rect 1697 3293 1713 3303
rect 1697 3263 1703 3293
rect 2257 3267 2263 3313
rect 2367 3303 2380 3307
rect 3680 3303 3693 3307
rect 2367 3293 2383 3303
rect 1697 3257 1743 3263
rect 1387 3253 1400 3257
rect 627 3237 693 3243
rect 1737 3243 1743 3257
rect 2247 3257 2263 3267
rect 2377 3267 2383 3293
rect 3677 3293 3693 3303
rect 4597 3297 4633 3303
rect 3677 3267 3683 3293
rect 2377 3257 2393 3267
rect 2247 3253 2260 3257
rect 2380 3253 2393 3257
rect 3677 3257 3693 3267
rect 3680 3253 3693 3257
rect 4597 3263 4603 3297
rect 4977 3263 4983 3313
rect 5400 3303 5413 3307
rect 5397 3293 5413 3303
rect 5527 3303 5540 3307
rect 5527 3293 5543 3303
rect 5397 3267 5403 3293
rect 5537 3267 5543 3293
rect 4557 3257 4603 3263
rect 4957 3257 4983 3263
rect 5117 3257 5153 3263
rect 4957 3247 4963 3257
rect 5387 3257 5403 3267
rect 5387 3253 5400 3257
rect 5527 3257 5543 3267
rect 5527 3253 5540 3257
rect 1737 3237 1773 3243
rect 1967 3237 2033 3243
rect 2847 3237 2933 3243
rect 4407 3237 4453 3243
rect 4947 3237 4963 3247
rect 4947 3233 4960 3237
rect 1967 3217 2013 3223
rect 2127 3223 2140 3227
rect 2127 3220 2143 3223
rect 2127 3213 2147 3220
rect 2133 3206 2147 3213
rect 2087 3197 2112 3203
rect 3857 3200 3893 3203
rect 3853 3197 3893 3200
rect 3853 3187 3867 3197
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 387 3037 453 3043
rect 547 3017 573 3023
rect 1887 3017 1913 3023
rect 2207 3017 2233 3023
rect 2967 3017 3013 3023
rect 4187 3017 4253 3023
rect 4761 3017 4813 3023
rect 4867 3017 4933 3023
rect 5087 3017 5153 3023
rect 877 2997 913 3003
rect 877 2967 883 2997
rect 1120 3003 1133 3007
rect 1117 2997 1133 3003
rect 1120 2993 1133 2997
rect 1440 3003 1453 3007
rect 1437 2993 1453 3003
rect 1527 2997 1573 3003
rect 1687 2997 1713 3003
rect 1847 2997 1913 3003
rect 867 2957 883 2967
rect 1437 2967 1443 2993
rect 3347 2997 3373 3003
rect 4087 2997 4113 3003
rect 4747 2997 4793 3003
rect 4897 2997 4933 3003
rect 4897 2967 4903 2997
rect 5547 3003 5560 3007
rect 5547 2997 5563 3003
rect 5547 2993 5560 2997
rect 5667 2997 5693 3003
rect 1437 2957 1453 2967
rect 867 2953 880 2957
rect 1440 2953 1453 2957
rect 4897 2957 4913 2967
rect 4900 2953 4913 2957
rect 5763 2878 5823 3382
rect 5730 2862 5823 2878
rect 107 2797 193 2803
rect 280 2783 293 2787
rect 277 2773 293 2783
rect 547 2783 560 2787
rect 547 2773 563 2783
rect 1707 2783 1720 2787
rect 1940 2783 1953 2787
rect 1707 2773 1723 2783
rect 277 2747 283 2773
rect 557 2747 563 2773
rect 1717 2747 1723 2773
rect 1937 2773 1953 2783
rect 4000 2783 4013 2787
rect 3997 2773 4013 2783
rect 4780 2783 4793 2787
rect 4777 2773 4793 2783
rect 5160 2783 5173 2787
rect 5157 2773 5173 2783
rect 5427 2783 5440 2787
rect 5427 2773 5443 2783
rect 5527 2783 5540 2787
rect 5527 2773 5543 2783
rect 1937 2747 1943 2773
rect 3997 2747 4003 2773
rect 4777 2747 4783 2773
rect 277 2737 293 2747
rect 280 2733 293 2737
rect 547 2737 563 2747
rect 547 2733 560 2737
rect 807 2737 833 2743
rect 1717 2737 1733 2747
rect 1720 2733 1733 2737
rect 1937 2737 1953 2747
rect 1940 2733 1953 2737
rect 3997 2737 4013 2747
rect 4000 2733 4013 2737
rect 4777 2737 4793 2747
rect 4780 2733 4793 2737
rect 5157 2743 5163 2773
rect 5437 2747 5443 2773
rect 5537 2747 5543 2773
rect 5137 2740 5203 2743
rect 5133 2737 5203 2740
rect 5437 2737 5453 2747
rect 5133 2727 5147 2737
rect 127 2717 193 2723
rect 5197 2723 5203 2737
rect 5440 2733 5453 2737
rect 5527 2737 5543 2747
rect 5527 2733 5540 2737
rect 5197 2717 5233 2723
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 107 2497 233 2503
rect 967 2477 1003 2483
rect 2867 2477 2913 2483
rect 3027 2477 3053 2483
rect 3160 2483 3173 2487
rect 3157 2473 3173 2483
rect 3157 2447 3163 2473
rect 3157 2437 3173 2447
rect 3160 2433 3173 2437
rect 5763 2358 5823 2862
rect 5730 2342 5823 2358
rect 5007 2277 5053 2283
rect 1867 2263 1880 2267
rect 1867 2253 1883 2263
rect 1877 2227 1883 2253
rect 1977 2257 2013 2263
rect 1977 2227 1983 2257
rect 3427 2257 3453 2263
rect 1867 2217 1883 2227
rect 1867 2213 1880 2217
rect 1967 2217 1983 2227
rect 4297 2227 4303 2273
rect 4297 2217 4313 2227
rect 1967 2213 1980 2217
rect 4300 2213 4313 2217
rect 5507 2217 5553 2223
rect 3907 2157 3933 2163
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 1147 1977 1193 1983
rect 1127 1957 1163 1963
rect 1157 1927 1163 1957
rect 1387 1957 1413 1963
rect 2360 1963 2373 1967
rect 2357 1953 2373 1963
rect 2587 1963 2600 1967
rect 2587 1953 2603 1963
rect 4487 1963 4500 1967
rect 4487 1957 4503 1963
rect 4487 1953 4500 1957
rect 4707 1963 4720 1967
rect 4707 1953 4723 1963
rect 5347 1963 5360 1967
rect 5347 1953 5363 1963
rect 2357 1927 2363 1953
rect 2597 1927 2603 1953
rect 4717 1927 4723 1953
rect 5357 1927 5363 1953
rect 1157 1917 1173 1927
rect 1160 1913 1173 1917
rect 2357 1917 2373 1927
rect 2360 1913 2373 1917
rect 2597 1917 2613 1927
rect 2600 1913 2613 1917
rect 4717 1917 4733 1927
rect 4720 1913 4733 1917
rect 5357 1917 5373 1927
rect 5360 1913 5373 1917
rect 1787 1897 1853 1903
rect 5763 1838 5823 2342
rect 5730 1822 5823 1838
rect 2237 1757 2273 1763
rect 607 1737 643 1743
rect 637 1707 643 1737
rect 1837 1737 1873 1743
rect 1837 1707 1843 1737
rect 637 1697 653 1707
rect 640 1693 653 1697
rect 1827 1697 1843 1707
rect 1827 1693 1840 1697
rect 2237 1703 2243 1757
rect 2820 1763 2833 1767
rect 2817 1753 2833 1763
rect 2207 1697 2243 1703
rect 2817 1703 2823 1753
rect 4720 1743 4733 1747
rect 4717 1740 4733 1743
rect 4713 1733 4733 1740
rect 4807 1743 4820 1747
rect 4807 1733 4823 1743
rect 5047 1743 5060 1747
rect 5047 1733 5063 1743
rect 4713 1726 4727 1733
rect 4817 1707 4823 1733
rect 5057 1707 5063 1733
rect 2787 1697 2823 1703
rect 3447 1697 3473 1703
rect 4807 1697 4823 1707
rect 4807 1693 4820 1697
rect 5047 1697 5063 1707
rect 5047 1693 5060 1697
rect 2087 1677 2153 1683
rect 4467 1677 4493 1683
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 707 1457 753 1463
rect 1767 1443 1780 1447
rect 4520 1443 4533 1447
rect 1767 1437 1783 1443
rect 1767 1433 1780 1437
rect 4517 1433 4533 1443
rect 4900 1443 4913 1447
rect 4897 1437 4913 1443
rect 4900 1433 4913 1437
rect 4517 1407 4523 1433
rect 4517 1397 4533 1407
rect 4520 1393 4533 1397
rect 5763 1318 5823 1822
rect 5730 1302 5823 1318
rect 720 1223 733 1227
rect 717 1213 733 1223
rect 1947 1223 1960 1227
rect 4660 1223 4673 1227
rect 1947 1213 1963 1223
rect 717 1187 723 1213
rect 1957 1187 1963 1213
rect 707 1177 723 1187
rect 707 1173 720 1177
rect 1207 1177 1233 1183
rect 1947 1177 1963 1187
rect 4657 1213 4673 1223
rect 5200 1223 5213 1227
rect 5197 1213 5213 1223
rect 4657 1183 4663 1213
rect 4773 1187 4787 1193
rect 5197 1187 5203 1213
rect 4657 1177 4693 1183
rect 1947 1173 1960 1177
rect 4773 1180 4793 1187
rect 4777 1177 4793 1180
rect 4780 1173 4793 1177
rect 5197 1177 5213 1187
rect 5200 1173 5213 1177
rect 2087 1157 2133 1163
rect 5167 1157 5233 1163
rect 2107 1137 2133 1143
rect 4913 1143 4927 1153
rect 4913 1140 4953 1143
rect 4917 1137 4953 1140
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 4487 957 4533 963
rect 787 943 800 947
rect 787 933 803 943
rect 607 923 620 927
rect 760 926 780 927
rect 760 923 773 926
rect 607 913 623 923
rect 757 917 773 923
rect 760 913 773 917
rect 617 887 623 913
rect 607 877 623 887
rect 797 887 803 933
rect 3927 937 3973 943
rect 933 923 947 933
rect 917 920 947 923
rect 917 917 943 920
rect 797 877 813 887
rect 607 873 620 877
rect 800 873 813 877
rect 917 867 923 917
rect 1407 923 1420 927
rect 1407 913 1423 923
rect 2087 917 2113 923
rect 2167 917 2193 923
rect 2347 923 2360 927
rect 2347 913 2363 923
rect 2487 923 2500 927
rect 2487 913 2503 923
rect 4207 917 4233 923
rect 1417 887 1423 913
rect 1407 877 1423 887
rect 1407 873 1420 877
rect 2357 866 2363 913
rect 2497 887 2503 913
rect 2487 877 2503 887
rect 2487 873 2500 877
rect 5763 798 5823 1302
rect 5730 782 5823 798
rect 2707 717 2743 723
rect 2337 697 2373 703
rect 27 677 74 683
rect 2337 667 2343 697
rect 587 657 623 663
rect 2327 657 2343 667
rect 2327 653 2340 657
rect 2737 663 2743 717
rect 3707 703 3720 707
rect 4180 703 4193 707
rect 3707 693 3723 703
rect 3717 667 3723 693
rect 2707 657 2743 663
rect 3587 657 3613 663
rect 3707 657 3723 667
rect 4177 693 4193 703
rect 4320 703 4333 707
rect 4317 693 4333 703
rect 4177 667 4183 693
rect 4317 667 4323 693
rect 4177 657 4193 667
rect 3707 653 3720 657
rect 4180 653 4193 657
rect 4317 657 4333 667
rect 4320 653 4333 657
rect 407 637 453 643
rect 3607 617 3653 623
rect -63 522 30 538
rect -63 18 -3 522
rect 1747 417 1773 423
rect 3567 417 3593 423
rect 4097 417 4133 423
rect 1867 403 1880 407
rect 1867 393 1883 403
rect 1877 367 1883 393
rect 2637 397 2673 403
rect 2637 367 2643 397
rect 2727 397 2753 403
rect 1867 357 1883 367
rect 1867 353 1880 357
rect 2627 357 2643 367
rect 2627 353 2640 357
rect 2777 363 2783 413
rect 2747 357 2783 363
rect 4097 367 4103 417
rect 4217 417 4253 423
rect 4097 357 4113 367
rect 4100 353 4113 357
rect 4217 363 4223 417
rect 4527 417 4573 423
rect 4217 357 4243 363
rect 867 337 913 343
rect 2107 337 2133 343
rect 2847 337 2893 343
rect 4237 343 4243 357
rect 4237 340 4263 343
rect 4237 337 4267 340
rect 2967 317 2993 323
rect 4253 326 4267 337
rect 5763 278 5823 782
rect 5730 262 5823 278
rect 5027 217 5053 223
rect 5027 197 5073 203
rect 2700 183 2713 187
rect 2697 173 2713 183
rect 3267 183 3280 187
rect 3267 173 3283 183
rect 3887 183 3900 187
rect 3887 173 3903 183
rect 4927 183 4940 187
rect 4927 173 4943 183
rect 5467 183 5480 187
rect 5467 173 5483 183
rect 2697 147 2703 173
rect 3277 147 3283 173
rect 3897 147 3903 173
rect 4937 147 4943 173
rect 5477 147 5483 173
rect 1707 137 1733 143
rect 2697 137 2713 147
rect 2700 133 2713 137
rect 3277 137 3293 147
rect 3280 133 3293 137
rect 3787 137 3813 143
rect 3897 137 3913 147
rect 3900 133 3913 137
rect 4937 137 4953 147
rect 4940 133 4953 137
rect 5477 137 5493 147
rect 5480 133 5493 137
rect 967 117 1013 123
rect 2447 97 2473 103
rect 3367 77 3433 83
rect -63 2 30 18
rect 5763 2 5823 262
<< m2contact >>
rect 2793 5393 2807 5407
rect 2873 5393 2887 5407
rect 3773 5393 3787 5407
rect 3813 5393 3827 5407
rect 333 5373 347 5387
rect 3613 5373 3627 5387
rect 673 5333 687 5347
rect 733 5333 747 5347
rect 3613 5333 3627 5347
rect 3933 5333 3947 5347
rect 3973 5333 3987 5347
rect 113 5313 127 5327
rect 233 5313 247 5327
rect 273 5313 287 5327
rect 3053 5313 3067 5327
rect 3153 5313 3167 5327
rect 3293 5313 3307 5327
rect 3433 5313 3447 5327
rect 3773 5313 3787 5327
rect 3833 5313 3847 5327
rect 4953 5313 4967 5327
rect 5013 5313 5027 5327
rect 3293 5292 3307 5306
rect 3333 5293 3347 5307
rect 2773 5133 2787 5147
rect 2853 5133 2867 5147
rect 3213 5133 3227 5147
rect 3253 5133 3267 5147
rect 2393 5113 2407 5127
rect 2493 5113 2507 5127
rect 613 5093 627 5107
rect 673 5093 687 5107
rect 533 5073 547 5087
rect 933 5073 947 5087
rect 1953 5093 1967 5107
rect 2093 5093 2107 5107
rect 2173 5093 2187 5107
rect 2373 5093 2387 5107
rect 2633 5093 2647 5107
rect 2693 5093 2707 5107
rect 3033 5093 3047 5107
rect 3113 5093 3127 5107
rect 3393 5093 3407 5107
rect 3673 5093 3687 5107
rect 3933 5093 3947 5107
rect 3993 5093 4007 5107
rect 4693 5093 4707 5107
rect 533 5033 547 5047
rect 893 5033 907 5047
rect 1853 5033 1867 5047
rect 2533 5073 2547 5087
rect 2573 5073 2587 5087
rect 2853 5073 2867 5087
rect 2473 5033 2487 5047
rect 2833 5033 2847 5047
rect 3373 5033 3387 5047
rect 3633 5033 3647 5047
rect 3839 5073 3853 5087
rect 3933 5072 3947 5086
rect 3973 5073 3987 5087
rect 4213 5073 4227 5087
rect 4253 5073 4267 5087
rect 4313 5073 4327 5087
rect 4553 5073 4567 5087
rect 5473 5093 5487 5107
rect 5573 5093 5587 5107
rect 3793 5033 3807 5047
rect 3333 5010 3347 5024
rect 3413 5013 3427 5027
rect 4293 5013 4307 5027
rect 4733 5072 4747 5086
rect 4973 5073 4987 5087
rect 5513 5073 5527 5087
rect 4613 5033 4627 5047
rect 4933 5033 4947 5047
rect 5213 5033 5227 5047
rect 5253 5033 5267 5047
rect 5513 5033 5527 5047
rect 4813 5013 4827 5027
rect 4853 5013 4867 5027
rect 1513 4873 1527 4887
rect 1573 4873 1587 4887
rect 473 4853 487 4867
rect 693 4853 707 4867
rect 413 4813 427 4827
rect 1093 4853 1107 4867
rect 2713 4853 2727 4867
rect 3393 4853 3407 4867
rect 3433 4853 3447 4867
rect 3753 4853 3767 4867
rect 1653 4833 1667 4847
rect 753 4813 767 4827
rect 1133 4813 1147 4827
rect 1693 4813 1707 4827
rect 4653 4853 4667 4867
rect 2773 4813 2787 4827
rect 3133 4813 3147 4827
rect 3213 4813 3227 4827
rect 3793 4813 3807 4827
rect 3933 4813 3947 4827
rect 3973 4813 3987 4827
rect 4333 4813 4347 4827
rect 4613 4813 4627 4827
rect 5193 4813 5207 4827
rect 5233 4813 5247 4827
rect 567 4793 581 4807
rect 653 4793 667 4807
rect 1453 4793 1467 4807
rect 1553 4793 1567 4807
rect 1933 4793 1947 4807
rect 1973 4793 1987 4807
rect 2433 4793 2447 4807
rect 3753 4793 3767 4807
rect 3853 4792 3867 4806
rect 4273 4791 4287 4805
rect 4353 4793 4367 4807
rect 5553 4793 5567 4807
rect 5633 4793 5647 4807
rect 2513 4773 2527 4787
rect 4533 4633 4547 4647
rect 633 4573 647 4587
rect 693 4573 707 4587
rect 2593 4573 2607 4587
rect 2693 4573 2707 4587
rect 3533 4573 3547 4587
rect 3573 4573 3587 4587
rect 613 4553 627 4567
rect 873 4552 887 4566
rect 933 4553 947 4567
rect 1153 4553 1167 4567
rect 1213 4553 1227 4567
rect 2293 4553 2307 4567
rect 2773 4553 2787 4567
rect 3153 4553 3167 4567
rect 673 4513 687 4527
rect 2293 4513 2307 4527
rect 2773 4513 2787 4527
rect 3333 4553 3347 4567
rect 3393 4553 3407 4567
rect 3193 4513 3207 4527
rect 3293 4513 3307 4527
rect 3553 4553 3567 4567
rect 3593 4552 3607 4566
rect 4613 4553 4627 4567
rect 3453 4513 3467 4527
rect 4313 4513 4327 4527
rect 353 4493 367 4507
rect 393 4493 407 4507
rect 3653 4493 3667 4507
rect 3713 4493 3727 4507
rect 93 4352 107 4366
rect 153 4353 167 4367
rect 673 4353 687 4367
rect 713 4353 727 4367
rect 513 4333 527 4347
rect 653 4333 667 4347
rect 693 4333 707 4347
rect 1293 4333 1307 4347
rect 2213 4333 2227 4347
rect 2413 4333 2427 4347
rect 2893 4333 2907 4347
rect 3393 4333 3407 4347
rect 3813 4333 3827 4347
rect 4019 4353 4033 4367
rect 4113 4353 4127 4367
rect 4153 4353 4167 4367
rect 513 4293 527 4307
rect 1113 4293 1127 4307
rect 1153 4293 1167 4307
rect 1253 4293 1267 4307
rect 2213 4293 2227 4307
rect 2373 4293 2387 4307
rect 2893 4293 2907 4307
rect 1333 4273 1347 4287
rect 1433 4273 1447 4287
rect 1613 4273 1627 4287
rect 1713 4273 1727 4287
rect 3573 4293 3587 4307
rect 3793 4293 3807 4307
rect 5013 4333 5027 4347
rect 5153 4333 5167 4347
rect 3873 4293 3887 4307
rect 3953 4293 3967 4307
rect 4093 4293 4107 4307
rect 4153 4293 4167 4307
rect 4233 4293 4247 4307
rect 4273 4293 4287 4307
rect 4493 4293 4507 4307
rect 4553 4293 4567 4307
rect 3413 4272 3427 4286
rect 3513 4273 3527 4287
rect 5213 4293 5227 4307
rect 5013 4273 5027 4287
rect 5053 4273 5067 4287
rect 5113 4273 5127 4287
rect 1353 4253 1367 4267
rect 1393 4253 1407 4267
rect 5293 4253 5307 4267
rect 5333 4253 5347 4267
rect 5253 4232 5267 4246
rect 5313 4233 5327 4247
rect 5353 4233 5367 4247
rect 573 4073 587 4087
rect 633 4073 647 4087
rect 3393 4073 3407 4087
rect 93 4053 107 4067
rect 233 4053 247 4067
rect 653 4053 667 4067
rect 953 4054 967 4068
rect 1013 4053 1027 4067
rect 1853 4053 1867 4067
rect 1953 4053 1967 4067
rect 2973 4053 2987 4067
rect 3033 4053 3047 4067
rect 3333 4053 3347 4067
rect 3373 4053 3387 4067
rect 553 3993 567 4007
rect 753 4033 767 4047
rect 1993 4033 2007 4047
rect 733 3992 747 4006
rect 1993 3993 2007 4007
rect 2053 4033 2067 4047
rect 2193 4033 2207 4047
rect 2473 4033 2487 4047
rect 2573 4033 2587 4047
rect 2613 4033 2627 4047
rect 3153 4033 3167 4047
rect 2053 3993 2067 4007
rect 2193 3993 2207 4007
rect 3293 4033 3307 4047
rect 3593 4053 3607 4067
rect 3633 4052 3647 4066
rect 3713 4053 3727 4067
rect 3793 4053 3807 4067
rect 4053 4053 4067 4067
rect 4113 4053 4127 4067
rect 3873 4033 3887 4047
rect 3153 3993 3167 4007
rect 3273 3993 3287 4007
rect 3353 3993 3367 4007
rect 3833 3993 3847 4007
rect 4013 4033 4027 4047
rect 4313 4033 4327 4047
rect 3993 3993 4007 4007
rect 4313 3993 4327 4007
rect 4373 4033 4387 4047
rect 4993 4033 5007 4047
rect 5033 4033 5047 4047
rect 5233 4033 5247 4047
rect 4373 3993 4387 4007
rect 5293 3993 5307 4007
rect 2453 3973 2467 3987
rect 4593 3973 4607 3987
rect 4633 3973 4647 3987
rect 953 3833 967 3847
rect 1033 3833 1047 3847
rect 2373 3833 2387 3847
rect 2433 3833 2447 3847
rect 3633 3833 3647 3847
rect 3673 3832 3687 3846
rect 3993 3833 4007 3847
rect 4393 3833 4407 3847
rect 653 3813 667 3827
rect 833 3813 847 3827
rect 1073 3813 1087 3827
rect 1793 3813 1807 3827
rect 1893 3813 1907 3827
rect 2113 3813 2127 3827
rect 1513 3793 1527 3807
rect 693 3773 707 3787
rect 833 3773 847 3787
rect 953 3772 967 3786
rect 993 3773 1007 3787
rect 1133 3773 1147 3787
rect 1473 3773 1487 3787
rect 1613 3773 1627 3787
rect 1659 3773 1673 3787
rect 1713 3773 1727 3787
rect 1753 3773 1767 3787
rect 1793 3773 1807 3787
rect 1893 3773 1907 3787
rect 1173 3753 1187 3767
rect 1253 3753 1267 3767
rect 2653 3813 2667 3827
rect 3733 3813 3747 3827
rect 2613 3773 2627 3787
rect 3713 3773 3727 3787
rect 3873 3793 3887 3807
rect 3913 3773 3927 3787
rect 3953 3773 3967 3787
rect 4153 3813 4167 3827
rect 4173 3773 4187 3787
rect 4373 3773 4387 3787
rect 5553 3813 5567 3827
rect 5553 3773 5567 3787
rect 2173 3753 2187 3767
rect 4393 3733 4407 3747
rect 4473 3732 4487 3746
rect 4993 3613 5007 3627
rect 2813 3553 2827 3567
rect 2873 3553 2887 3567
rect 93 3533 107 3547
rect 193 3533 207 3547
rect 793 3533 807 3547
rect 833 3533 847 3547
rect 2173 3533 2187 3547
rect 2453 3533 2467 3547
rect 2493 3533 2507 3547
rect 53 3513 67 3527
rect 293 3513 307 3527
rect 333 3513 347 3527
rect 933 3513 947 3527
rect 1093 3513 1107 3527
rect 1433 3513 1447 3527
rect 1833 3513 1847 3527
rect 2013 3513 2027 3527
rect 2073 3513 2087 3527
rect 53 3473 67 3487
rect 973 3473 987 3487
rect 1073 3473 1087 3487
rect 1373 3473 1387 3487
rect 1793 3473 1807 3487
rect 2433 3513 2447 3527
rect 2233 3473 2247 3487
rect 2433 3473 2447 3487
rect 2713 3532 2727 3546
rect 3233 3533 3247 3547
rect 4333 3533 4347 3547
rect 5713 3533 5727 3547
rect 2833 3513 2847 3527
rect 2873 3513 2887 3527
rect 3453 3513 3467 3527
rect 2713 3473 2727 3487
rect 3253 3473 3267 3487
rect 533 3453 547 3467
rect 593 3453 607 3467
rect 653 3453 667 3467
rect 753 3453 767 3467
rect 4473 3513 4487 3527
rect 4913 3513 4927 3527
rect 5053 3513 5067 3527
rect 5593 3513 5607 3527
rect 3593 3473 3607 3487
rect 3633 3473 3647 3487
rect 4353 3473 4367 3487
rect 4473 3473 4487 3487
rect 4873 3473 4887 3487
rect 3513 3453 3527 3467
rect 4573 3453 4587 3467
rect 4613 3452 4627 3466
rect 5713 3432 5727 3446
rect 2193 3413 2207 3427
rect 2233 3413 2247 3427
rect 1813 3332 1827 3346
rect 1873 3333 1887 3347
rect 3833 3333 3847 3347
rect 3893 3333 3907 3347
rect 193 3313 207 3327
rect 233 3313 247 3327
rect 1833 3313 1847 3327
rect 1893 3312 1907 3326
rect 2253 3313 2267 3327
rect 4813 3315 4827 3329
rect 4873 3313 4887 3327
rect 4993 3313 5007 3327
rect 633 3293 647 3307
rect 1293 3293 1307 3307
rect 1373 3293 1387 3307
rect 633 3253 647 3267
rect 1093 3253 1107 3267
rect 1133 3253 1147 3267
rect 1273 3252 1287 3266
rect 1373 3253 1387 3267
rect 1713 3293 1727 3307
rect 2353 3293 2367 3307
rect 613 3233 627 3247
rect 693 3233 707 3247
rect 2233 3253 2247 3267
rect 3693 3293 3707 3307
rect 2393 3253 2407 3267
rect 3693 3253 3707 3267
rect 4633 3293 4647 3307
rect 5413 3293 5427 3307
rect 5513 3293 5527 3307
rect 5153 3253 5167 3267
rect 5373 3253 5387 3267
rect 5513 3253 5527 3267
rect 1773 3233 1787 3247
rect 1953 3233 1967 3247
rect 2033 3233 2047 3247
rect 2833 3233 2847 3247
rect 2933 3233 2947 3247
rect 4393 3232 4407 3246
rect 4453 3233 4467 3247
rect 4933 3233 4947 3247
rect 1953 3212 1967 3226
rect 2013 3213 2027 3227
rect 2113 3213 2127 3227
rect 2073 3193 2087 3207
rect 2112 3192 2126 3206
rect 2133 3192 2147 3206
rect 3893 3192 3907 3206
rect 3853 3173 3867 3187
rect 5073 3173 5087 3187
rect 373 3033 387 3047
rect 453 3033 467 3047
rect 533 3013 547 3027
rect 573 3013 587 3027
rect 1873 3013 1887 3027
rect 1913 3013 1927 3027
rect 2193 3013 2207 3027
rect 2233 3013 2247 3027
rect 2953 3013 2967 3027
rect 3013 3013 3027 3027
rect 4173 3013 4187 3027
rect 4253 3013 4267 3027
rect 4747 3013 4761 3027
rect 4813 3013 4827 3027
rect 4853 3013 4867 3027
rect 4933 3013 4947 3027
rect 5073 3013 5087 3027
rect 5153 3013 5167 3027
rect 913 2993 927 3007
rect 1133 2993 1147 3007
rect 1453 2993 1467 3007
rect 1513 2993 1527 3007
rect 1573 2993 1587 3007
rect 1673 2993 1687 3007
rect 1713 2993 1727 3007
rect 1833 2993 1847 3007
rect 853 2953 867 2967
rect 1913 2992 1927 3006
rect 3333 2993 3347 3007
rect 3373 2992 3387 3006
rect 4073 2993 4087 3007
rect 4113 2993 4127 3007
rect 4733 2992 4747 3006
rect 4793 2993 4807 3007
rect 4933 2992 4947 3006
rect 5533 2993 5547 3007
rect 5653 2993 5667 3007
rect 5693 2993 5707 3007
rect 1453 2953 1467 2967
rect 4913 2953 4927 2967
rect 93 2792 107 2806
rect 193 2793 207 2807
rect 293 2773 307 2787
rect 533 2773 547 2787
rect 1693 2773 1707 2787
rect 1953 2773 1967 2787
rect 4013 2773 4027 2787
rect 4793 2773 4807 2787
rect 5173 2773 5187 2787
rect 5413 2773 5427 2787
rect 5513 2773 5527 2787
rect 293 2733 307 2747
rect 533 2733 547 2747
rect 793 2733 807 2747
rect 833 2733 847 2747
rect 1733 2733 1747 2747
rect 1953 2733 1967 2747
rect 4013 2733 4027 2747
rect 4793 2733 4807 2747
rect 113 2713 127 2727
rect 193 2713 207 2727
rect 5133 2713 5147 2727
rect 5453 2733 5467 2747
rect 5513 2733 5527 2747
rect 5233 2713 5247 2727
rect 93 2493 107 2507
rect 233 2493 247 2507
rect 953 2473 967 2487
rect 2853 2473 2867 2487
rect 2913 2473 2927 2487
rect 3013 2473 3027 2487
rect 3053 2473 3067 2487
rect 3173 2473 3187 2487
rect 3173 2433 3187 2447
rect 4293 2273 4307 2287
rect 4993 2273 5007 2287
rect 5053 2273 5067 2287
rect 1853 2253 1867 2267
rect 2013 2253 2027 2267
rect 3413 2253 3427 2267
rect 3453 2253 3467 2267
rect 1853 2213 1867 2227
rect 1953 2213 1967 2227
rect 4313 2213 4327 2227
rect 5493 2213 5507 2227
rect 5553 2213 5567 2227
rect 3893 2153 3907 2167
rect 3933 2152 3947 2166
rect 4533 2053 4547 2067
rect 1133 1973 1147 1987
rect 1193 1973 1207 1987
rect 1113 1953 1127 1967
rect 1373 1953 1387 1967
rect 1413 1953 1427 1967
rect 2373 1953 2387 1967
rect 2573 1953 2587 1967
rect 4473 1953 4487 1967
rect 4693 1953 4707 1967
rect 5333 1953 5347 1967
rect 1173 1913 1187 1927
rect 2373 1913 2387 1927
rect 2613 1913 2627 1927
rect 4733 1913 4747 1927
rect 5373 1913 5387 1927
rect 1773 1893 1787 1907
rect 1853 1893 1867 1907
rect 593 1733 607 1747
rect 1873 1733 1887 1747
rect 653 1693 667 1707
rect 1813 1693 1827 1707
rect 2193 1693 2207 1707
rect 2273 1753 2287 1767
rect 2833 1753 2847 1767
rect 2773 1693 2787 1707
rect 4733 1733 4747 1747
rect 4793 1733 4807 1747
rect 5033 1733 5047 1747
rect 4713 1712 4727 1726
rect 3433 1693 3447 1707
rect 3473 1693 3487 1707
rect 4793 1693 4807 1707
rect 5033 1693 5047 1707
rect 2073 1673 2087 1687
rect 2153 1672 2167 1686
rect 4453 1673 4467 1687
rect 4493 1673 4507 1687
rect 693 1453 707 1467
rect 753 1453 767 1467
rect 1753 1433 1767 1447
rect 4533 1433 4547 1447
rect 4913 1433 4927 1447
rect 4533 1393 4547 1407
rect 733 1213 747 1227
rect 1933 1213 1947 1227
rect 693 1173 707 1187
rect 1193 1173 1207 1187
rect 1233 1173 1247 1187
rect 1933 1173 1947 1187
rect 4673 1213 4687 1227
rect 5213 1213 5227 1227
rect 4773 1193 4787 1207
rect 4693 1173 4707 1187
rect 4793 1173 4807 1187
rect 5213 1173 5227 1187
rect 2073 1153 2087 1167
rect 2133 1153 2147 1167
rect 4913 1153 4927 1167
rect 5153 1153 5167 1167
rect 5233 1153 5247 1167
rect 2093 1133 2107 1147
rect 2133 1132 2147 1146
rect 4953 1132 4967 1146
rect 4473 952 4487 966
rect 4533 953 4547 967
rect 773 933 787 947
rect 593 913 607 927
rect 773 912 787 926
rect 593 873 607 887
rect 933 933 947 947
rect 3913 933 3927 947
rect 3973 933 3987 947
rect 813 873 827 887
rect 1393 913 1407 927
rect 2073 913 2087 927
rect 2113 913 2127 927
rect 2153 913 2167 927
rect 2193 913 2207 927
rect 2333 913 2347 927
rect 2473 913 2487 927
rect 4193 913 4207 927
rect 4233 913 4247 927
rect 1393 873 1407 887
rect 913 853 927 867
rect 2473 873 2487 887
rect 2353 852 2367 866
rect 2693 713 2707 727
rect 13 673 27 687
rect 2373 693 2387 707
rect 573 653 587 667
rect 2313 653 2327 667
rect 2693 653 2707 667
rect 3693 693 3707 707
rect 3573 653 3587 667
rect 3613 653 3627 667
rect 3693 653 3707 667
rect 4193 693 4207 707
rect 4333 693 4347 707
rect 4193 653 4207 667
rect 4333 653 4347 667
rect 393 633 407 647
rect 453 633 467 647
rect 3593 613 3607 627
rect 3653 613 3667 627
rect 1733 412 1747 426
rect 1773 413 1787 427
rect 2773 413 2787 427
rect 3553 413 3567 427
rect 3593 413 3607 427
rect 1853 393 1867 407
rect 2673 393 2687 407
rect 2713 393 2727 407
rect 2753 393 2767 407
rect 1853 353 1867 367
rect 2613 353 2627 367
rect 2733 353 2747 367
rect 4133 413 4147 427
rect 4113 353 4127 367
rect 4253 413 4267 427
rect 4513 413 4527 427
rect 4573 413 4587 427
rect 853 333 867 347
rect 913 333 927 347
rect 2093 333 2107 347
rect 2133 333 2147 347
rect 2833 333 2847 347
rect 2893 333 2907 347
rect 2953 313 2967 327
rect 2993 313 3007 327
rect 4253 312 4267 326
rect 5013 213 5027 227
rect 5053 213 5067 227
rect 5013 192 5027 206
rect 5073 193 5087 207
rect 2713 173 2727 187
rect 3253 173 3267 187
rect 3873 173 3887 187
rect 4913 173 4927 187
rect 5453 173 5467 187
rect 1693 133 1707 147
rect 1733 133 1747 147
rect 2713 133 2727 147
rect 3293 133 3307 147
rect 3773 133 3787 147
rect 3813 133 3827 147
rect 3913 133 3927 147
rect 4953 133 4967 147
rect 5493 133 5507 147
rect 953 113 967 127
rect 1013 113 1027 127
rect 2433 93 2447 107
rect 2473 93 2487 107
rect 3353 73 3367 87
rect 3433 73 3447 87
<< metal2 >>
rect 2896 5487 2903 5523
rect 216 5389 223 5413
rect 36 5027 43 5373
rect 96 5340 103 5343
rect 93 5327 107 5340
rect 113 5327 127 5333
rect 196 5327 203 5343
rect 233 5327 247 5333
rect 273 5327 287 5333
rect 196 5227 203 5313
rect 296 5167 303 5375
rect 316 5347 323 5473
rect 336 5427 343 5453
rect 347 5383 360 5387
rect 347 5376 363 5383
rect 396 5376 403 5413
rect 347 5373 360 5376
rect 353 5368 360 5373
rect 556 5347 563 5373
rect 116 5076 123 5113
rect 216 5076 223 5113
rect 16 4127 23 4933
rect 36 4827 43 4873
rect 76 4856 83 4933
rect 96 4887 103 5043
rect 136 5040 143 5043
rect 196 5040 203 5043
rect 133 5027 147 5040
rect 193 5027 207 5040
rect 236 4967 243 5043
rect 276 5007 283 5033
rect 116 4856 123 4933
rect 216 4856 223 4933
rect 136 4727 143 4823
rect 36 4526 43 4613
rect 196 4556 203 4613
rect 216 4567 223 4793
rect 236 4727 243 4823
rect 236 4556 243 4653
rect 256 4627 263 4693
rect 276 4607 283 4813
rect 296 4767 303 5073
rect 316 5047 323 5113
rect 376 5007 383 5043
rect 316 4787 323 4893
rect 336 4867 343 4953
rect 356 4856 363 4933
rect 376 4887 383 4993
rect 396 4856 403 4893
rect 416 4887 423 5253
rect 476 5187 483 5333
rect 516 5307 523 5343
rect 556 5267 563 5333
rect 576 5327 583 5413
rect 596 5387 603 5473
rect 616 5376 623 5453
rect 653 5380 667 5393
rect 756 5389 763 5453
rect 656 5376 663 5380
rect 736 5267 743 5333
rect 476 5076 483 5113
rect 536 5087 543 5153
rect 556 5047 563 5213
rect 667 5123 740 5127
rect 667 5113 743 5123
rect 613 5087 627 5093
rect 656 5076 663 5113
rect 687 5093 693 5107
rect 736 5088 743 5113
rect 756 5083 763 5313
rect 776 5307 783 5343
rect 796 5267 803 5313
rect 816 5307 823 5393
rect 896 5376 903 5453
rect 1156 5376 1163 5413
rect 1236 5389 1243 5413
rect 876 5183 883 5343
rect 976 5227 983 5373
rect 1116 5327 1123 5343
rect 1116 5267 1123 5313
rect 1176 5227 1183 5343
rect 1236 5327 1243 5375
rect 1276 5267 1283 5343
rect 856 5176 883 5183
rect 756 5076 783 5083
rect 496 4987 503 5043
rect 536 4907 543 5033
rect 596 4927 603 5043
rect 636 4987 643 5043
rect 707 5036 723 5043
rect 696 4967 703 5033
rect 776 5027 783 5076
rect 856 5076 863 5176
rect 976 5127 983 5173
rect 1056 5167 1063 5213
rect 880 5047 887 5052
rect 916 5047 923 5093
rect 933 5087 947 5093
rect 976 5083 983 5113
rect 956 5076 983 5083
rect 880 5043 893 5047
rect 356 4587 363 4813
rect 376 4767 383 4823
rect 456 4667 463 4873
rect 476 4867 483 4893
rect 536 4869 543 4893
rect 680 4863 693 4867
rect 676 4856 693 4863
rect 680 4853 693 4856
rect 680 4848 687 4853
rect 476 4743 483 4773
rect 496 4767 503 4813
rect 516 4787 523 4823
rect 556 4820 563 4823
rect 553 4807 567 4820
rect 516 4743 523 4773
rect 476 4736 523 4743
rect 596 4667 603 4812
rect 616 4787 623 4823
rect 656 4820 663 4823
rect 653 4807 667 4820
rect 96 4387 103 4512
rect 136 4467 143 4553
rect 156 4516 183 4523
rect 156 4367 163 4516
rect 356 4520 363 4523
rect 316 4447 323 4512
rect 353 4507 367 4520
rect 93 4348 107 4352
rect 236 4336 243 4373
rect 296 4336 303 4373
rect 376 4367 383 4513
rect 396 4507 403 4653
rect 456 4556 463 4613
rect 576 4556 583 4613
rect 616 4567 623 4593
rect 76 4267 83 4303
rect 136 4067 143 4333
rect 176 4267 183 4303
rect 356 4287 363 4303
rect 176 4147 183 4253
rect 356 4247 363 4273
rect 376 4083 383 4293
rect 356 4076 383 4083
rect 93 4040 107 4053
rect 96 4036 103 4040
rect 193 4040 207 4053
rect 233 4047 247 4053
rect 356 4047 363 4076
rect 196 4036 203 4040
rect 373 4040 387 4053
rect 396 4047 403 4453
rect 416 4347 423 4513
rect 436 4387 443 4523
rect 496 4507 503 4553
rect 636 4525 643 4573
rect 456 4349 463 4493
rect 516 4347 523 4373
rect 376 4036 383 4040
rect 416 4036 423 4233
rect 436 4227 443 4303
rect 476 4300 483 4303
rect 473 4287 487 4300
rect 516 4227 523 4293
rect 476 4036 483 4133
rect 516 4036 523 4073
rect 536 4047 543 4433
rect 656 4387 663 4772
rect 716 4607 723 5013
rect 836 4987 843 5043
rect 876 5036 893 5043
rect 880 5033 893 5036
rect 996 5040 1003 5043
rect 993 5027 1007 5040
rect 1036 4987 1043 5033
rect 796 4907 803 4953
rect 836 4947 843 4973
rect 1056 4967 1063 5153
rect 1136 5076 1143 5213
rect 936 4856 943 4933
rect 1056 4856 1063 4893
rect 1076 4883 1083 5033
rect 1116 5007 1123 5043
rect 1076 4880 1103 4883
rect 1076 4876 1107 4880
rect 1093 4867 1107 4876
rect 1156 4856 1163 4953
rect 1176 4867 1183 5133
rect 1196 5107 1203 5193
rect 1276 5187 1283 5253
rect 1316 5127 1323 5343
rect 1336 5267 1343 5333
rect 1356 5147 1363 5343
rect 1236 5076 1243 5113
rect 1396 5107 1403 5413
rect 1476 5388 1483 5453
rect 1556 5427 1563 5473
rect 1556 5376 1563 5413
rect 1436 5340 1443 5343
rect 1433 5327 1447 5340
rect 1216 4907 1223 5043
rect 1316 5007 1323 5073
rect 1336 4887 1343 5093
rect 1416 5076 1423 5233
rect 1516 5088 1523 5193
rect 1536 5147 1543 5343
rect 1576 5247 1583 5343
rect 1576 5103 1583 5233
rect 1556 5096 1583 5103
rect 1556 5076 1563 5096
rect 1596 5083 1603 5333
rect 1656 5287 1663 5375
rect 1756 5376 1763 5433
rect 1856 5389 1863 5413
rect 2016 5389 2023 5433
rect 2036 5407 2043 5473
rect 2396 5407 2403 5453
rect 1676 5107 1683 5373
rect 1776 5287 1783 5343
rect 1836 5247 1843 5343
rect 1596 5076 1623 5083
rect 736 4667 743 4853
rect 756 4767 763 4813
rect 776 4787 783 4823
rect 816 4767 823 4823
rect 876 4727 883 4853
rect 956 4787 963 4823
rect 976 4747 983 4793
rect 756 4647 763 4693
rect 676 4567 683 4593
rect 733 4584 747 4593
rect 707 4580 747 4584
rect 707 4577 743 4580
rect 796 4556 803 4673
rect 836 4556 843 4633
rect 876 4587 883 4713
rect 867 4566 880 4567
rect 867 4553 873 4566
rect 596 4336 603 4373
rect 676 4367 683 4513
rect 716 4447 723 4523
rect 776 4467 783 4513
rect 816 4487 823 4511
rect 856 4467 863 4523
rect 713 4347 727 4353
rect 916 4349 923 4573
rect 936 4567 943 4713
rect 996 4567 1003 4773
rect 1036 4727 1043 4823
rect 1056 4816 1073 4823
rect 936 4423 943 4553
rect 1020 4523 1033 4527
rect 1016 4516 1033 4523
rect 1020 4513 1033 4516
rect 936 4416 963 4423
rect 640 4343 653 4347
rect 636 4336 653 4343
rect 640 4333 653 4336
rect 640 4328 647 4333
rect 576 4300 583 4303
rect 573 4287 587 4300
rect 567 4073 573 4087
rect 616 4067 623 4113
rect 76 3907 83 4003
rect 16 3747 23 3853
rect 36 3787 43 3833
rect 96 3816 103 3853
rect 136 3827 143 3893
rect 173 3820 187 3833
rect 176 3816 183 3820
rect 216 3816 223 3913
rect 256 3787 263 4003
rect 296 3903 303 4033
rect 356 4000 363 4003
rect 276 3896 303 3903
rect 136 3776 153 3783
rect 16 3267 23 3593
rect 56 3527 63 3553
rect 76 3523 83 3772
rect 136 3547 143 3776
rect 93 3523 107 3533
rect 76 3520 107 3523
rect 76 3516 103 3520
rect 136 3516 143 3533
rect 193 3520 207 3533
rect 216 3527 223 3673
rect 276 3667 283 3896
rect 336 3867 343 3993
rect 353 3987 367 4000
rect 496 4000 503 4003
rect 376 3816 383 3893
rect 316 3747 323 3783
rect 196 3516 203 3520
rect 233 3520 247 3533
rect 236 3516 243 3520
rect 376 3516 383 3753
rect 416 3727 423 3853
rect 436 3827 443 3993
rect 493 3987 507 4000
rect 456 3816 463 3893
rect 536 3829 543 4003
rect 556 3927 563 3993
rect 576 3867 583 4052
rect 616 4036 623 4053
rect 636 4047 643 4073
rect 653 4040 667 4053
rect 676 4047 683 4332
rect 696 4147 703 4333
rect 736 4300 743 4303
rect 716 4127 723 4293
rect 733 4287 747 4300
rect 796 4207 803 4303
rect 867 4296 883 4303
rect 656 4036 663 4040
rect 636 4000 643 4003
rect 633 3987 647 4000
rect 676 3967 683 4003
rect 716 3987 723 4033
rect 736 4027 743 4073
rect 767 4043 780 4047
rect 767 4036 783 4043
rect 816 4036 823 4113
rect 856 4047 863 4133
rect 876 4107 883 4296
rect 896 4207 903 4303
rect 936 4287 943 4393
rect 956 4347 963 4416
rect 976 4336 983 4473
rect 996 4407 1003 4513
rect 996 4300 1003 4303
rect 767 4033 780 4036
rect 916 4036 923 4113
rect 956 4068 963 4293
rect 993 4287 1007 4300
rect 1036 4127 1043 4473
rect 1056 4387 1063 4816
rect 1076 4567 1083 4773
rect 1116 4687 1123 4853
rect 1236 4827 1243 4873
rect 1336 4856 1383 4863
rect 1116 4556 1123 4593
rect 1136 4567 1143 4813
rect 1196 4627 1203 4823
rect 1256 4587 1263 4813
rect 1276 4707 1283 4823
rect 1213 4567 1227 4573
rect 1247 4563 1260 4567
rect 1276 4563 1283 4693
rect 1316 4667 1323 4823
rect 1247 4556 1283 4563
rect 1247 4553 1260 4556
rect 1096 4427 1103 4523
rect 1113 4483 1127 4493
rect 1113 4480 1143 4483
rect 1116 4476 1143 4480
rect 1136 4347 1143 4476
rect 1236 4467 1243 4523
rect 1156 4307 1163 4373
rect 1076 4167 1083 4303
rect 1096 4247 1103 4293
rect 1116 4147 1123 4293
rect 1176 4227 1183 4413
rect 736 3927 743 3992
rect 796 3983 803 4003
rect 796 3976 843 3983
rect 656 3827 663 3853
rect 776 3847 783 3973
rect 476 3780 483 3783
rect 36 3367 43 3513
rect 296 3487 303 3513
rect 436 3487 443 3653
rect 56 3447 63 3473
rect 76 3327 83 3483
rect 356 3480 363 3483
rect 16 3047 23 3093
rect 16 2647 23 2993
rect 36 2947 43 3313
rect 96 3296 103 3333
rect 76 3047 83 3263
rect 136 3067 143 3433
rect 256 3347 263 3471
rect 353 3467 367 3480
rect 193 3300 207 3313
rect 233 3308 247 3313
rect 196 3296 203 3300
rect 296 3296 303 3452
rect 176 3043 183 3252
rect 236 3167 243 3294
rect 276 3227 283 3263
rect 156 3036 183 3043
rect 116 2996 123 3033
rect 156 3007 163 3036
rect 36 2747 43 2793
rect 56 2783 63 2953
rect 96 2827 103 2963
rect 136 2960 143 2963
rect 133 2947 147 2960
rect 176 2963 183 3013
rect 233 3000 247 3013
rect 236 2996 243 3000
rect 276 2996 283 3153
rect 296 3107 303 3133
rect 176 2956 203 2963
rect 87 2806 100 2807
rect 87 2793 93 2806
rect 56 2776 83 2783
rect 156 2787 163 2953
rect 196 2907 203 2956
rect 216 2827 223 2963
rect 256 2927 263 2963
rect 126 2733 127 2740
rect 113 2727 127 2733
rect 176 2567 183 2813
rect 193 2787 207 2793
rect 233 2780 247 2793
rect 236 2776 243 2780
rect 253 2723 267 2733
rect 207 2720 267 2723
rect 207 2716 263 2720
rect 36 2367 43 2553
rect 93 2487 107 2493
rect 196 2487 203 2613
rect 276 2527 283 2813
rect 316 2807 323 3213
rect 376 3127 383 3353
rect 396 3347 403 3483
rect 456 3387 463 3773
rect 473 3767 487 3780
rect 516 3727 523 3783
rect 576 3767 583 3783
rect 576 3647 583 3753
rect 616 3727 623 3783
rect 656 3687 663 3773
rect 676 3747 683 3814
rect 816 3786 823 3893
rect 836 3827 843 3976
rect 936 3947 943 4003
rect 896 3903 903 3933
rect 896 3896 933 3903
rect 873 3820 887 3833
rect 876 3816 883 3820
rect 916 3816 923 3873
rect 956 3847 963 3973
rect 976 3887 983 3953
rect 996 3947 1003 4053
rect 1016 3887 1023 4053
rect 1056 4047 1063 4133
rect 1136 4107 1143 4133
rect 1073 4040 1087 4053
rect 1096 4047 1103 4073
rect 1076 4036 1083 4040
rect 1113 4040 1127 4053
rect 1116 4036 1123 4040
rect 1036 3903 1043 3993
rect 1056 3927 1063 4003
rect 1096 3907 1103 4003
rect 1036 3896 1063 3903
rect 1016 3876 1033 3887
rect 1020 3873 1033 3876
rect 1056 3864 1063 3896
rect 1027 3857 1063 3864
rect 956 3807 963 3833
rect 976 3827 983 3852
rect 1026 3832 1027 3840
rect 1047 3833 1053 3847
rect 1013 3820 1027 3832
rect 1060 3823 1073 3827
rect 1016 3816 1023 3820
rect 1056 3816 1073 3823
rect 1060 3813 1073 3816
rect 1060 3808 1067 3813
rect 693 3767 707 3773
rect 687 3740 703 3743
rect 687 3736 707 3740
rect 693 3727 707 3736
rect 776 3687 783 3783
rect 856 3780 863 3783
rect 776 3567 783 3633
rect 796 3607 803 3653
rect 816 3627 823 3713
rect 836 3687 843 3773
rect 853 3767 867 3780
rect 953 3767 967 3772
rect 516 3516 523 3553
rect 556 3517 593 3524
rect 596 3483 603 3513
rect 536 3480 543 3483
rect 533 3467 547 3480
rect 576 3476 603 3483
rect 576 3427 583 3476
rect 593 3447 607 3453
rect 476 3323 483 3393
rect 456 3316 483 3323
rect 456 3309 463 3316
rect 436 3107 443 3263
rect 476 3227 483 3263
rect 373 3047 387 3053
rect 373 3000 387 3012
rect 376 2996 383 3000
rect 416 2996 423 3093
rect 436 3007 443 3053
rect 456 3047 463 3073
rect 476 3027 483 3213
rect 516 3187 523 3333
rect 536 3307 543 3353
rect 556 3347 563 3393
rect 616 3296 623 3453
rect 636 3307 643 3483
rect 656 3347 663 3453
rect 676 3447 683 3471
rect 736 3407 743 3553
rect 836 3547 843 3593
rect 793 3527 807 3533
rect 876 3527 883 3553
rect 913 3520 927 3533
rect 936 3527 943 3633
rect 916 3516 923 3520
rect 776 3467 783 3483
rect 896 3480 903 3483
rect 767 3456 783 3467
rect 816 3463 823 3471
rect 816 3456 843 3463
rect 767 3453 780 3456
rect 696 3296 703 3373
rect 736 3296 743 3333
rect 516 3027 523 3173
rect 536 3067 543 3253
rect 616 3147 623 3233
rect 547 3056 563 3063
rect 456 3016 473 3023
rect 456 2965 463 3016
rect 533 3003 547 3013
rect 516 3000 547 3003
rect 516 2996 543 3000
rect 556 2996 563 3056
rect 596 3047 603 3073
rect 636 3067 643 3253
rect 656 3227 663 3293
rect 776 3267 783 3393
rect 796 3307 803 3433
rect 836 3423 843 3456
rect 856 3447 863 3473
rect 893 3467 907 3480
rect 956 3427 963 3533
rect 976 3527 983 3773
rect 1076 3647 1083 3773
rect 1096 3747 1103 3872
rect 1096 3647 1103 3733
rect 1016 3516 1023 3553
rect 1056 3516 1063 3593
rect 1096 3587 1103 3612
rect 1116 3563 1123 3913
rect 1156 3847 1163 4113
rect 1196 4036 1203 4293
rect 1216 4247 1223 4303
rect 1256 4207 1263 4293
rect 1276 4187 1283 4373
rect 1296 4347 1303 4473
rect 1316 4387 1323 4613
rect 1376 4556 1383 4856
rect 1396 4827 1403 5043
rect 1436 4947 1443 5043
rect 1536 4907 1543 5043
rect 1576 4947 1583 5043
rect 1596 5007 1603 5033
rect 1616 4967 1623 5076
rect 1813 5080 1827 5093
rect 1816 5076 1823 5080
rect 1656 4927 1663 5043
rect 1796 5007 1803 5043
rect 1576 4887 1583 4912
rect 1513 4869 1527 4873
rect 1576 4856 1583 4873
rect 1653 4847 1667 4853
rect 1453 4807 1467 4813
rect 1496 4767 1503 4823
rect 1556 4820 1563 4823
rect 1553 4807 1567 4820
rect 1556 4687 1563 4772
rect 1596 4767 1603 4823
rect 1676 4807 1683 4893
rect 1756 4856 1763 4893
rect 1576 4667 1583 4733
rect 1356 4503 1363 4523
rect 1356 4496 1383 4503
rect 1356 4336 1363 4413
rect 1376 4367 1383 4496
rect 1396 4407 1403 4523
rect 1416 4348 1423 4493
rect 1436 4427 1443 4513
rect 1456 4467 1463 4653
rect 1516 4556 1523 4653
rect 1576 4520 1583 4523
rect 1573 4507 1587 4520
rect 1436 4363 1443 4413
rect 1476 4387 1483 4473
rect 1436 4356 1463 4363
rect 1456 4336 1463 4356
rect 1496 4336 1503 4433
rect 1296 4127 1303 4293
rect 1336 4287 1343 4303
rect 1436 4300 1443 4303
rect 1336 4227 1343 4273
rect 1353 4267 1367 4273
rect 1376 4247 1383 4293
rect 1433 4287 1447 4300
rect 1407 4253 1413 4267
rect 1476 4247 1483 4303
rect 1256 4043 1263 4093
rect 1236 4036 1263 4043
rect 1313 4040 1327 4053
rect 1336 4047 1343 4192
rect 1316 4036 1323 4040
rect 1196 3927 1203 3953
rect 1147 3823 1160 3827
rect 1147 3816 1163 3823
rect 1196 3816 1203 3913
rect 1276 3903 1283 3993
rect 1296 3983 1303 4003
rect 1296 3976 1323 3983
rect 1276 3896 1303 3903
rect 1236 3827 1243 3853
rect 1147 3813 1160 3816
rect 1276 3823 1283 3873
rect 1296 3847 1303 3896
rect 1316 3847 1323 3976
rect 1256 3816 1283 3823
rect 1313 3820 1327 3833
rect 1356 3827 1363 4173
rect 1396 4147 1403 4213
rect 1536 4187 1543 4413
rect 1596 4407 1603 4453
rect 1616 4427 1623 4773
rect 1676 4627 1683 4713
rect 1656 4556 1663 4593
rect 1696 4568 1703 4813
rect 1716 4707 1723 4813
rect 1736 4727 1743 4823
rect 1716 4607 1723 4653
rect 1796 4587 1803 4813
rect 1816 4687 1823 4953
rect 1836 4907 1843 5043
rect 1853 5027 1867 5033
rect 1876 5007 1883 5312
rect 1916 5307 1923 5353
rect 1956 5247 1963 5343
rect 1996 5340 2003 5343
rect 1993 5327 2007 5340
rect 2036 5287 2043 5343
rect 1913 5080 1927 5093
rect 1953 5080 1967 5093
rect 1916 5076 1923 5080
rect 1956 5076 1963 5080
rect 1976 4927 1983 5043
rect 2036 4967 2043 5273
rect 2076 5207 2083 5393
rect 2096 5346 2103 5373
rect 2136 5107 2143 5173
rect 2196 5167 2203 5233
rect 2216 5187 2223 5343
rect 2256 5207 2263 5343
rect 2296 5227 2303 5375
rect 2316 5247 2323 5393
rect 2393 5380 2407 5393
rect 2396 5376 2403 5380
rect 2436 5347 2443 5375
rect 2636 5376 2643 5433
rect 2336 5287 2343 5313
rect 2356 5247 2363 5332
rect 2476 5307 2483 5343
rect 2453 5263 2467 5273
rect 2453 5260 2493 5263
rect 2456 5256 2493 5260
rect 2216 5147 2223 5173
rect 2296 5127 2303 5213
rect 2093 5080 2107 5093
rect 2096 5076 2103 5080
rect 2073 5047 2080 5052
rect 2176 5047 2183 5093
rect 2236 5087 2243 5113
rect 2393 5107 2407 5113
rect 2373 5080 2387 5093
rect 2376 5076 2383 5080
rect 2416 5076 2423 5133
rect 2067 5043 2080 5047
rect 2067 5036 2083 5043
rect 2116 5040 2123 5043
rect 2067 5033 2080 5036
rect 2113 5027 2127 5040
rect 2316 5045 2323 5073
rect 1836 4867 1843 4893
rect 1896 4856 1903 4893
rect 1936 4867 1943 4913
rect 2196 4907 2203 4953
rect 2216 4947 2223 5043
rect 2256 4987 2263 5031
rect 2396 5007 2403 5043
rect 2436 4987 2443 5031
rect 2456 4947 2463 5173
rect 2476 5083 2483 5233
rect 2536 5147 2543 5343
rect 2696 5346 2703 5413
rect 2793 5380 2807 5393
rect 2796 5376 2803 5380
rect 2576 5227 2583 5333
rect 2616 5227 2623 5343
rect 2736 5287 2743 5343
rect 2493 5103 2507 5113
rect 2493 5100 2523 5103
rect 2496 5096 2523 5100
rect 2476 5076 2493 5083
rect 2516 5083 2523 5096
rect 2516 5076 2533 5083
rect 2587 5073 2593 5087
rect 2633 5080 2647 5093
rect 2676 5087 2683 5273
rect 2736 5163 2743 5252
rect 2756 5247 2763 5333
rect 2776 5227 2783 5343
rect 2736 5156 2763 5163
rect 2756 5147 2763 5156
rect 2756 5136 2773 5147
rect 2760 5133 2773 5136
rect 2707 5093 2713 5107
rect 2636 5076 2643 5080
rect 2736 5076 2743 5133
rect 2796 5083 2803 5333
rect 2816 5267 2823 5343
rect 2816 5147 2823 5253
rect 2856 5247 2863 5453
rect 2896 5407 2903 5473
rect 2936 5447 2943 5473
rect 2876 5347 2883 5393
rect 2956 5376 2963 5393
rect 3016 5388 3023 5413
rect 3056 5387 3063 5523
rect 2896 5207 2903 5293
rect 2916 5287 2923 5332
rect 2936 5267 2943 5293
rect 2853 5147 2867 5153
rect 2776 5076 2803 5083
rect 2013 4860 2027 4873
rect 2016 4856 2023 4860
rect 1876 4727 1883 4823
rect 1916 4820 1923 4823
rect 1913 4807 1927 4820
rect 1933 4807 1947 4813
rect 1896 4707 1903 4773
rect 1956 4767 1963 4813
rect 1996 4807 2003 4823
rect 1987 4796 2003 4807
rect 1987 4793 2000 4796
rect 2076 4767 2083 4873
rect 2116 4868 2123 4893
rect 2176 4807 2183 4855
rect 1936 4756 1953 4763
rect 1816 4647 1823 4673
rect 1856 4627 1863 4673
rect 1676 4363 1683 4523
rect 1776 4520 1783 4523
rect 1773 4507 1787 4520
rect 1676 4356 1703 4363
rect 1696 4349 1703 4356
rect 1736 4336 1743 4393
rect 1856 4387 1863 4553
rect 1876 4507 1883 4633
rect 1916 4556 1923 4613
rect 1936 4567 1943 4756
rect 1956 4607 1963 4732
rect 2216 4727 2223 4823
rect 2036 4556 2043 4713
rect 2076 4567 2083 4653
rect 2316 4647 2323 4933
rect 2476 4927 2483 5033
rect 2336 4826 2343 4913
rect 2396 4856 2403 4893
rect 2496 4867 2503 4993
rect 2516 4927 2523 5043
rect 2576 4907 2583 5073
rect 2696 5007 2703 5033
rect 2576 4896 2593 4907
rect 2580 4893 2593 4896
rect 2636 4868 2643 4973
rect 2756 4967 2763 5043
rect 2816 4967 2823 5093
rect 2836 5007 2843 5033
rect 2436 4856 2483 4863
rect 2476 4823 2483 4856
rect 2673 4860 2687 4873
rect 2716 4867 2723 4893
rect 2676 4856 2683 4860
rect 2416 4807 2423 4823
rect 2456 4816 2483 4823
rect 2416 4793 2433 4807
rect 2096 4556 2103 4613
rect 2136 4567 2143 4593
rect 2193 4560 2207 4573
rect 2196 4556 2203 4560
rect 1976 4467 1983 4493
rect 1996 4487 2003 4553
rect 2056 4487 2063 4523
rect 1596 4287 1603 4303
rect 1596 4276 1613 4287
rect 1600 4273 1613 4276
rect 1393 4040 1407 4053
rect 1396 4036 1403 4040
rect 1416 3887 1423 4003
rect 1496 3983 1503 4093
rect 1496 3976 1523 3983
rect 1316 3816 1323 3820
rect 1153 3808 1160 3813
rect 1176 3780 1183 3783
rect 1136 3707 1143 3773
rect 1096 3556 1123 3563
rect 1096 3527 1103 3556
rect 1136 3523 1143 3553
rect 1156 3547 1163 3773
rect 1173 3767 1187 3780
rect 1256 3767 1263 3816
rect 1393 3820 1407 3833
rect 1433 3820 1447 3833
rect 1476 3827 1483 3913
rect 1396 3816 1403 3820
rect 1436 3816 1443 3820
rect 1276 3776 1303 3783
rect 1176 3687 1183 3753
rect 1176 3523 1183 3633
rect 1116 3516 1143 3523
rect 1156 3516 1183 3523
rect 1196 3516 1203 3553
rect 1236 3516 1243 3713
rect 1256 3527 1263 3732
rect 1276 3667 1283 3776
rect 1336 3687 1343 3713
rect 1276 3547 1283 3613
rect 1296 3587 1303 3633
rect 1356 3627 1363 3773
rect 836 3416 873 3423
rect 836 3296 843 3353
rect 976 3347 983 3473
rect 996 3367 1003 3483
rect 1076 3387 1083 3473
rect 1096 3387 1103 3492
rect 1116 3467 1123 3516
rect 1356 3516 1363 3553
rect 1176 3447 1183 3471
rect 976 3296 983 3333
rect 1036 3307 1043 3373
rect 693 3227 707 3233
rect 656 3023 663 3133
rect 716 3127 723 3193
rect 876 3187 883 3295
rect 1136 3267 1143 3333
rect 1216 3327 1223 3471
rect 1336 3447 1343 3483
rect 1373 3463 1387 3473
rect 1356 3460 1387 3463
rect 1356 3456 1383 3460
rect 1256 3267 1263 3373
rect 1276 3287 1283 3413
rect 1356 3407 1363 3456
rect 1396 3427 1403 3733
rect 1416 3707 1423 3783
rect 1416 3527 1423 3672
rect 1456 3527 1463 3593
rect 1476 3567 1483 3773
rect 1496 3747 1503 3833
rect 1516 3807 1523 3976
rect 1536 3927 1543 4003
rect 1596 3867 1603 4113
rect 1616 3927 1623 4133
rect 1636 4067 1643 4333
rect 1656 4247 1663 4293
rect 1676 4267 1683 4303
rect 1716 4300 1723 4303
rect 1713 4287 1727 4300
rect 1656 4047 1663 4233
rect 1676 4067 1683 4093
rect 1716 4067 1723 4252
rect 1673 4040 1687 4053
rect 1676 4036 1683 4040
rect 1716 4036 1723 4053
rect 1636 3947 1643 3993
rect 1616 3843 1623 3913
rect 1596 3836 1623 3843
rect 1596 3816 1603 3836
rect 1636 3827 1643 3853
rect 1656 3827 1663 4003
rect 1736 3947 1743 3993
rect 1756 3947 1763 4173
rect 1776 4127 1783 4373
rect 1916 4307 1923 4335
rect 1816 4300 1843 4303
rect 1816 4296 1847 4300
rect 1793 4283 1807 4293
rect 1833 4287 1847 4296
rect 1793 4280 1823 4283
rect 1796 4276 1823 4280
rect 1816 4247 1823 4276
rect 1796 4187 1803 4233
rect 1836 4167 1843 4273
rect 1856 4227 1863 4253
rect 1876 4227 1883 4303
rect 1936 4147 1943 4433
rect 2076 4347 2083 4513
rect 2116 4336 2123 4513
rect 2176 4447 2183 4523
rect 2216 4487 2223 4511
rect 2156 4336 2163 4393
rect 2176 4347 2183 4373
rect 2056 4306 2063 4333
rect 1956 4147 1963 4193
rect 1836 4036 1843 4132
rect 1853 4067 1867 4073
rect 1916 4036 1923 4093
rect 1976 4067 1983 4293
rect 2016 4287 2023 4303
rect 2016 4107 2023 4273
rect 1987 4060 2003 4063
rect 1987 4056 2007 4060
rect 1953 4047 1967 4053
rect 1993 4047 2007 4056
rect 1736 3827 1743 3933
rect 1756 3787 1763 3912
rect 1516 3607 1523 3772
rect 1476 3516 1483 3553
rect 1293 3307 1307 3313
rect 1336 3296 1343 3353
rect 1356 3327 1363 3393
rect 1376 3307 1383 3333
rect 1416 3323 1423 3473
rect 1496 3387 1503 3473
rect 1516 3363 1523 3572
rect 1556 3523 1563 3773
rect 1576 3747 1583 3783
rect 1596 3587 1603 3753
rect 1616 3527 1623 3733
rect 1736 3687 1743 3773
rect 1536 3516 1563 3523
rect 1536 3367 1543 3516
rect 1640 3523 1653 3527
rect 1636 3516 1653 3523
rect 1640 3513 1653 3516
rect 1576 3383 1583 3483
rect 1556 3376 1583 3383
rect 1496 3356 1523 3363
rect 1396 3316 1423 3323
rect 736 3107 743 3133
rect 573 3007 587 3013
rect 636 3016 663 3023
rect 636 3008 643 3016
rect 676 3008 683 3093
rect 356 2807 363 2963
rect 496 2927 503 2963
rect 616 2960 623 2963
rect 307 2783 320 2787
rect 307 2776 323 2783
rect 356 2776 363 2793
rect 307 2773 320 2776
rect 313 2768 320 2773
rect 376 2740 383 2743
rect 233 2480 247 2493
rect 296 2487 303 2733
rect 373 2727 387 2740
rect 416 2707 423 2873
rect 436 2867 443 2893
rect 516 2776 523 2913
rect 536 2787 543 2893
rect 496 2707 503 2743
rect 236 2476 243 2480
rect 56 2343 63 2433
rect 76 2407 83 2443
rect 116 2367 123 2431
rect 36 2336 63 2343
rect 36 2227 43 2336
rect 136 2227 143 2293
rect 216 2269 223 2353
rect 256 2327 263 2443
rect 296 2307 303 2433
rect 296 2283 303 2293
rect 296 2276 323 2283
rect 316 2256 323 2276
rect 376 2263 383 2413
rect 416 2367 423 2513
rect 436 2287 443 2473
rect 496 2436 523 2443
rect 516 2367 523 2436
rect 536 2423 543 2733
rect 556 2627 563 2933
rect 576 2783 583 2953
rect 613 2947 627 2960
rect 656 2867 663 2963
rect 696 2887 703 2953
rect 716 2947 723 3053
rect 876 3027 883 3173
rect 916 3007 923 3263
rect 956 3260 963 3263
rect 953 3247 967 3260
rect 996 3256 1053 3263
rect 976 3127 983 3193
rect 996 3067 1003 3173
rect 1016 3147 1023 3233
rect 1116 3063 1123 3233
rect 1116 3056 1143 3063
rect 736 2967 743 2994
rect 953 3000 967 3013
rect 1136 3007 1143 3056
rect 956 2996 963 3000
rect 836 2823 843 2963
rect 856 2907 863 2953
rect 876 2947 883 2992
rect 896 2907 903 2953
rect 836 2816 853 2823
rect 576 2776 593 2783
rect 856 2776 863 2813
rect 916 2788 923 2933
rect 1036 2787 1043 2813
rect 616 2740 623 2743
rect 613 2727 627 2740
rect 636 2707 643 2733
rect 656 2476 663 2513
rect 696 2445 703 2773
rect 756 2587 763 2743
rect 796 2707 803 2733
rect 756 2476 763 2513
rect 536 2416 553 2423
rect 376 2256 403 2263
rect 236 2220 243 2223
rect 116 2047 123 2213
rect 233 2203 247 2220
rect 287 2223 300 2227
rect 287 2216 303 2223
rect 336 2220 343 2223
rect 287 2213 300 2216
rect 333 2207 347 2220
rect 233 2197 333 2203
rect 356 2087 363 2213
rect 16 1967 23 1993
rect 36 1927 43 2013
rect 76 1956 83 2033
rect 196 1967 203 2053
rect 236 1956 243 2013
rect 256 1967 263 2073
rect 376 1956 383 1993
rect 396 1967 403 2256
rect 516 2256 523 2313
rect 176 1887 183 1923
rect 216 1903 223 1923
rect 216 1896 243 1903
rect 16 1396 43 1403
rect 16 687 23 1396
rect 56 1228 63 1313
rect 96 1287 103 1873
rect 236 1747 243 1896
rect 116 1327 123 1734
rect 216 1667 223 1703
rect 276 1667 283 1703
rect 227 1656 243 1663
rect 236 1443 243 1656
rect 216 1436 243 1443
rect 376 1436 383 1813
rect 396 1667 403 1893
rect 416 1827 423 2253
rect 456 2220 463 2223
rect 453 2207 467 2220
rect 456 2067 463 2193
rect 556 2167 563 2413
rect 596 2327 603 2443
rect 736 2387 743 2443
rect 836 2387 843 2733
rect 896 2527 903 2733
rect 916 2507 923 2774
rect 976 2707 983 2743
rect 956 2676 1003 2683
rect 956 2647 963 2676
rect 947 2636 963 2647
rect 947 2633 960 2636
rect 956 2487 963 2613
rect 976 2587 983 2653
rect 996 2567 1003 2676
rect 1056 2667 1063 2893
rect 1076 2847 1083 2923
rect 1156 2783 1163 3253
rect 1176 3027 1183 3263
rect 1196 3256 1213 3263
rect 1196 3003 1203 3256
rect 1256 3087 1263 3253
rect 1176 2996 1203 3003
rect 1216 2996 1223 3073
rect 1276 3067 1283 3252
rect 1296 3047 1303 3213
rect 1356 3207 1363 3263
rect 1376 3107 1383 3253
rect 1253 3000 1267 3013
rect 1256 2996 1263 3000
rect 1176 2965 1183 2996
rect 1376 2996 1383 3053
rect 1396 3007 1403 3316
rect 1496 3296 1503 3356
rect 1556 3347 1563 3376
rect 1576 3307 1583 3353
rect 1596 3296 1603 3453
rect 1616 3447 1623 3483
rect 1676 3427 1683 3593
rect 1716 3516 1723 3573
rect 1756 3516 1763 3653
rect 1776 3547 1783 3893
rect 1796 3827 1803 3933
rect 1816 3867 1823 4003
rect 1856 3947 1863 4003
rect 1976 3947 1983 4003
rect 1836 3843 1843 3893
rect 1996 3867 2003 3993
rect 1816 3836 1843 3843
rect 1816 3816 1823 3836
rect 1796 3687 1803 3773
rect 1796 3527 1803 3633
rect 1876 3567 1883 3853
rect 1893 3827 1907 3833
rect 1936 3829 1943 3853
rect 2016 3827 2023 4093
rect 2036 4005 2043 4173
rect 2056 4147 2063 4213
rect 2076 4047 2083 4253
rect 2096 4063 2103 4292
rect 2116 4167 2123 4233
rect 2136 4207 2143 4303
rect 2156 4143 2163 4253
rect 2136 4136 2163 4143
rect 2136 4067 2143 4136
rect 2156 4067 2163 4113
rect 2096 4056 2123 4063
rect 2067 4036 2083 4047
rect 2116 4036 2123 4056
rect 2067 4033 2080 4036
rect 2056 3927 2063 3993
rect 2136 3983 2143 4003
rect 2116 3976 2143 3983
rect 2116 3827 2123 3976
rect 2136 3907 2143 3953
rect 1916 3780 1923 3783
rect 1896 3607 1903 3773
rect 1913 3767 1927 3780
rect 1676 3303 1683 3413
rect 1796 3407 1803 3473
rect 1716 3307 1723 3353
rect 1736 3327 1743 3373
rect 1816 3367 1823 3553
rect 1916 3543 1923 3673
rect 1976 3667 1983 3783
rect 1896 3536 1923 3543
rect 1847 3523 1860 3527
rect 1847 3516 1863 3523
rect 1896 3516 1903 3536
rect 1976 3527 1983 3613
rect 1996 3527 2003 3633
rect 1847 3513 1860 3516
rect 1967 3516 1983 3527
rect 1967 3513 1980 3516
rect 1876 3447 1883 3483
rect 1916 3427 1923 3483
rect 1936 3447 1943 3473
rect 1807 3346 1820 3347
rect 1807 3333 1813 3346
rect 1676 3296 1703 3303
rect 1427 3273 1433 3287
rect 1696 3267 1703 3296
rect 1756 3296 1763 3333
rect 1836 3327 1843 3373
rect 1896 3367 1903 3413
rect 1887 3346 1900 3347
rect 1887 3333 1893 3346
rect 1536 3260 1543 3263
rect 1533 3247 1547 3260
rect 1616 3260 1623 3263
rect 1416 2967 1423 3013
rect 1436 3007 1443 3193
rect 1456 3007 1463 3173
rect 1476 2996 1483 3053
rect 1136 2776 1163 2783
rect 1076 2627 1083 2733
rect 1096 2476 1103 2713
rect 1116 2707 1123 2743
rect 1116 2567 1123 2633
rect 1136 2543 1143 2593
rect 1176 2587 1183 2833
rect 1216 2783 1223 2873
rect 1236 2827 1243 2963
rect 1356 2789 1363 2951
rect 1376 2807 1383 2933
rect 1196 2776 1223 2783
rect 1116 2536 1143 2543
rect 1116 2507 1123 2536
rect 1196 2527 1203 2776
rect 1396 2776 1403 2893
rect 1436 2867 1443 2993
rect 1456 2847 1463 2953
rect 1496 2807 1503 2963
rect 1556 2927 1563 3252
rect 1613 3247 1627 3260
rect 1656 3187 1663 3263
rect 1776 3260 1783 3263
rect 1676 3007 1683 3253
rect 1773 3247 1787 3260
rect 1696 3127 1703 3193
rect 1796 3147 1803 3233
rect 1836 3187 1843 3292
rect 1836 3147 1843 3173
rect 1836 3007 1843 3133
rect 1587 3003 1600 3007
rect 1587 2996 1603 3003
rect 1587 2993 1600 2996
rect 1827 2986 1843 2987
rect 1827 2973 1833 2986
rect 1856 2967 1863 3313
rect 1893 3308 1907 3312
rect 1936 3308 1943 3333
rect 1956 3327 1963 3473
rect 2056 3483 2063 3733
rect 2076 3547 2083 3773
rect 2096 3707 2103 3783
rect 2136 3647 2143 3853
rect 2156 3847 2163 3993
rect 2176 3867 2183 4293
rect 2196 4087 2203 4353
rect 2216 4347 2223 4433
rect 2256 4367 2263 4633
rect 2276 4527 2283 4613
rect 2293 4567 2307 4573
rect 2353 4560 2367 4573
rect 2376 4567 2383 4753
rect 2396 4667 2403 4753
rect 2416 4707 2423 4793
rect 2456 4727 2463 4816
rect 2527 4783 2540 4787
rect 2527 4773 2543 4783
rect 2476 4687 2483 4753
rect 2356 4556 2363 4560
rect 2416 4556 2423 4593
rect 2436 4587 2443 4673
rect 2456 4556 2463 4593
rect 2496 4567 2503 4773
rect 2516 4667 2523 4733
rect 2536 4707 2543 4773
rect 2556 4767 2563 4823
rect 2273 4343 2287 4353
rect 2296 4349 2303 4513
rect 2436 4520 2443 4523
rect 2433 4507 2447 4520
rect 2476 4467 2483 4523
rect 2516 4427 2523 4593
rect 2596 4587 2603 4813
rect 2656 4767 2663 4823
rect 2696 4787 2703 4823
rect 2536 4523 2543 4573
rect 2596 4556 2603 4573
rect 2636 4556 2643 4613
rect 2656 4567 2663 4713
rect 2676 4707 2683 4733
rect 2736 4707 2743 4873
rect 2836 4856 2843 4993
rect 2876 4947 2883 5043
rect 2916 4987 2923 5043
rect 2876 4867 2883 4933
rect 2936 4856 2943 4993
rect 2956 4887 2963 5313
rect 2996 5087 3003 5333
rect 3036 5327 3043 5343
rect 3036 5316 3053 5327
rect 3040 5313 3053 5316
rect 3076 5267 3083 5473
rect 3096 5387 3103 5473
rect 3180 5383 3193 5387
rect 3176 5376 3193 5383
rect 3180 5373 3193 5376
rect 3180 5368 3187 5373
rect 3096 5187 3103 5333
rect 3116 5107 3123 5343
rect 3156 5340 3163 5343
rect 3153 5327 3167 5340
rect 3216 5343 3223 5523
rect 3416 5503 3423 5523
rect 3416 5496 3463 5503
rect 3416 5467 3423 5496
rect 3436 5447 3443 5473
rect 3456 5467 3463 5496
rect 3276 5376 3283 5412
rect 3296 5407 3303 5433
rect 3556 5376 3563 5413
rect 3600 5383 3613 5387
rect 3596 5376 3613 5383
rect 3600 5373 3613 5376
rect 3196 5336 3223 5343
rect 3176 5107 3183 5333
rect 3196 5247 3203 5336
rect 3236 5327 3243 5373
rect 3496 5347 3503 5373
rect 3600 5368 3607 5373
rect 3296 5340 3303 5343
rect 3293 5327 3307 5340
rect 3336 5327 3343 5343
rect 3333 5307 3347 5313
rect 3196 5167 3203 5193
rect 3216 5147 3223 5293
rect 3376 5303 3383 5333
rect 3396 5307 3403 5343
rect 3376 5296 3393 5303
rect 3236 5187 3243 5273
rect 3296 5267 3303 5292
rect 3316 5227 3323 5253
rect 3033 5080 3047 5093
rect 3073 5080 3087 5093
rect 3036 5076 3043 5080
rect 3076 5076 3083 5080
rect 3016 5040 3023 5043
rect 3013 5027 3027 5040
rect 3060 5023 3073 5027
rect 3056 5020 3073 5023
rect 3053 5013 3073 5020
rect 3053 5007 3067 5013
rect 3066 5000 3067 5007
rect 2976 4856 2983 4893
rect 2996 4883 3003 4973
rect 2996 4876 3023 4883
rect 2693 4560 2707 4573
rect 2736 4567 2743 4613
rect 2756 4587 2763 4853
rect 2776 4567 2783 4813
rect 2856 4787 2863 4823
rect 2916 4820 2923 4823
rect 2913 4807 2927 4820
rect 2796 4587 2803 4613
rect 2696 4556 2703 4560
rect 2536 4516 2563 4523
rect 2576 4520 2583 4523
rect 2433 4403 2447 4413
rect 2416 4400 2447 4403
rect 2416 4396 2443 4400
rect 2256 4340 2287 4343
rect 2256 4336 2283 4340
rect 2376 4347 2383 4393
rect 2416 4383 2423 4396
rect 2396 4376 2423 4383
rect 2227 4303 2240 4307
rect 2227 4296 2243 4303
rect 2227 4293 2240 4296
rect 2216 4063 2223 4153
rect 2316 4147 2323 4292
rect 2336 4107 2343 4153
rect 2356 4123 2363 4303
rect 2376 4147 2383 4293
rect 2356 4116 2383 4123
rect 2376 4087 2383 4116
rect 2396 4107 2403 4376
rect 2413 4347 2427 4353
rect 2436 4348 2443 4373
rect 2476 4336 2483 4413
rect 2456 4207 2463 4303
rect 2536 4247 2543 4453
rect 2196 4060 2223 4063
rect 2193 4056 2223 4060
rect 2193 4047 2207 4056
rect 2213 4007 2220 4012
rect 2207 4003 2220 4007
rect 2207 3996 2223 4003
rect 2256 4000 2263 4003
rect 2207 3993 2220 3996
rect 2253 3987 2267 4000
rect 2156 3833 2173 3847
rect 2156 3827 2163 3833
rect 2216 3816 2223 3973
rect 2316 3887 2323 4073
rect 2353 4040 2367 4053
rect 2456 4048 2463 4193
rect 2356 4036 2363 4040
rect 2476 4047 2483 4233
rect 2556 4187 2563 4516
rect 2573 4507 2587 4520
rect 2616 4487 2623 4523
rect 2716 4487 2723 4523
rect 2596 4349 2603 4373
rect 2547 4163 2560 4167
rect 2547 4153 2563 4163
rect 2527 4143 2540 4147
rect 2527 4133 2543 4143
rect 2456 4003 2463 4034
rect 2516 4036 2523 4093
rect 2536 4043 2543 4133
rect 2556 4127 2563 4153
rect 2576 4087 2583 4213
rect 2596 4143 2603 4293
rect 2616 4167 2623 4303
rect 2596 4136 2623 4143
rect 2616 4107 2623 4136
rect 2576 4047 2583 4073
rect 2636 4067 2643 4293
rect 2656 4147 2663 4433
rect 2756 4336 2763 4523
rect 2776 4447 2783 4513
rect 2796 4487 2803 4573
rect 2876 4556 2883 4593
rect 2896 4567 2903 4693
rect 2913 4560 2927 4573
rect 2936 4567 2943 4813
rect 2956 4787 2963 4823
rect 3016 4763 3023 4876
rect 3036 4767 3043 4873
rect 3056 4867 3063 4953
rect 3076 4887 3083 4992
rect 3116 4967 3123 5093
rect 3176 5076 3183 5093
rect 3216 5087 3223 5112
rect 3156 4947 3163 5043
rect 3196 4967 3203 5043
rect 3236 4967 3243 5033
rect 2996 4756 3023 4763
rect 2916 4556 2923 4560
rect 2976 4556 2983 4593
rect 2996 4587 3003 4756
rect 3016 4643 3023 4733
rect 3056 4647 3063 4793
rect 3076 4667 3083 4713
rect 3016 4636 3043 4643
rect 3036 4587 3043 4636
rect 2996 4563 3003 4573
rect 2996 4556 3023 4563
rect 2816 4467 2823 4553
rect 3076 4527 3083 4653
rect 3096 4647 3103 4673
rect 3136 4663 3143 4813
rect 3136 4656 3163 4663
rect 3116 4587 3123 4653
rect 3136 4568 3143 4593
rect 3156 4567 3163 4656
rect 3176 4567 3183 4893
rect 3236 4856 3243 4953
rect 3256 4907 3263 5133
rect 3353 5080 3367 5093
rect 3376 5083 3383 5173
rect 3396 5107 3403 5233
rect 3416 5207 3423 5333
rect 3436 5327 3443 5343
rect 3436 5247 3443 5313
rect 3456 5123 3463 5333
rect 3496 5227 3503 5253
rect 3536 5247 3543 5343
rect 3576 5340 3583 5343
rect 3573 5327 3587 5340
rect 3436 5116 3463 5123
rect 3436 5087 3443 5116
rect 3356 5076 3363 5080
rect 3376 5076 3403 5083
rect 3296 5007 3303 5043
rect 3327 5024 3340 5027
rect 3327 5013 3333 5024
rect 3287 4996 3303 5007
rect 3287 4993 3300 4996
rect 3356 4967 3363 5013
rect 3376 4887 3383 5033
rect 3396 4967 3403 5076
rect 3453 5083 3467 5093
rect 3476 5083 3483 5173
rect 3616 5167 3623 5333
rect 3636 5307 3643 5413
rect 3736 5407 3743 5453
rect 3776 5407 3783 5473
rect 3876 5427 3883 5523
rect 3453 5080 3483 5083
rect 3456 5076 3483 5080
rect 3576 5076 3583 5153
rect 3616 5076 3623 5113
rect 3636 5107 3643 5293
rect 3656 5187 3663 5373
rect 3696 5340 3703 5343
rect 3693 5327 3707 5340
rect 3736 5247 3743 5343
rect 3796 5343 3803 5413
rect 3916 5407 3923 5523
rect 3827 5393 3833 5407
rect 3853 5380 3867 5393
rect 3856 5376 3863 5380
rect 3936 5367 3943 5433
rect 3996 5376 4003 5453
rect 4036 5388 4043 5473
rect 4067 5436 4093 5443
rect 3933 5347 3947 5353
rect 3796 5336 3823 5343
rect 3836 5340 3843 5343
rect 3773 5327 3787 5333
rect 3676 5187 3683 5233
rect 3656 5047 3663 5133
rect 3673 5107 3687 5113
rect 3696 5083 3703 5213
rect 3756 5167 3763 5273
rect 3676 5076 3703 5083
rect 3436 5027 3443 5043
rect 3427 5017 3443 5027
rect 3427 5013 3440 5017
rect 3416 4947 3423 4992
rect 3456 4987 3463 5013
rect 3516 4987 3523 5033
rect 3536 4943 3543 4993
rect 3556 4987 3563 5043
rect 3496 4940 3543 4943
rect 3493 4936 3543 4940
rect 3493 4927 3507 4936
rect 3616 4927 3623 5013
rect 3506 4920 3507 4927
rect 3313 4860 3327 4873
rect 3316 4856 3323 4860
rect 3256 4787 3263 4813
rect 3356 4747 3363 4812
rect 3396 4783 3403 4853
rect 3376 4776 3403 4783
rect 3276 4556 3283 4613
rect 2836 4387 2843 4513
rect 2836 4336 2843 4373
rect 2856 4347 2863 4523
rect 2696 4300 2703 4303
rect 2693 4287 2707 4300
rect 2876 4303 2883 4493
rect 2973 4387 2987 4393
rect 2967 4380 2987 4387
rect 2967 4376 2983 4380
rect 2967 4373 2980 4376
rect 2996 4367 3003 4433
rect 2893 4347 2907 4353
rect 3016 4327 3023 4473
rect 3036 4427 3043 4523
rect 3116 4467 3123 4523
rect 3096 4349 3103 4413
rect 2856 4296 2883 4303
rect 2536 4036 2553 4043
rect 2376 4000 2383 4003
rect 2373 3987 2387 4000
rect 2416 3944 2423 4003
rect 2456 3996 2483 4003
rect 2387 3943 2423 3944
rect 2387 3940 2443 3943
rect 2387 3937 2447 3940
rect 2416 3936 2447 3937
rect 2433 3927 2447 3936
rect 2376 3847 2383 3912
rect 2156 3747 2163 3773
rect 2073 3527 2087 3533
rect 2116 3516 2123 3573
rect 2176 3547 2183 3753
rect 2196 3547 2203 3783
rect 2236 3707 2243 3772
rect 2296 3767 2303 3813
rect 2416 3683 2423 3893
rect 2456 3867 2463 3973
rect 2476 3847 2483 3996
rect 2496 3887 2503 4003
rect 2536 3947 2543 4003
rect 2576 3867 2583 3993
rect 2596 3983 2603 4053
rect 2676 4048 2683 4173
rect 2627 4043 2640 4047
rect 2627 4036 2643 4043
rect 2627 4033 2640 4036
rect 2753 4040 2767 4053
rect 2813 4043 2827 4053
rect 2796 4040 2827 4043
rect 2756 4036 2763 4040
rect 2796 4036 2823 4040
rect 2836 4005 2843 4233
rect 2656 3983 2663 4003
rect 2696 4000 2703 4003
rect 2596 3976 2623 3983
rect 2616 3887 2623 3976
rect 2636 3976 2663 3983
rect 2693 3987 2707 4000
rect 2776 3987 2783 4003
rect 2636 3947 2643 3976
rect 2767 3976 2783 3987
rect 2767 3973 2780 3976
rect 2447 3843 2460 3847
rect 2447 3833 2463 3843
rect 2456 3816 2463 3833
rect 2576 3816 2583 3853
rect 2656 3827 2663 3953
rect 2736 3927 2743 3973
rect 2796 3927 2803 3973
rect 2636 3787 2643 3815
rect 2693 3820 2707 3833
rect 2736 3827 2743 3913
rect 2696 3816 2703 3820
rect 2476 3780 2483 3783
rect 2396 3676 2423 3683
rect 2156 3516 2203 3523
rect 2056 3476 2083 3483
rect 2056 3387 2063 3453
rect 2036 3327 2043 3353
rect 2056 3296 2063 3333
rect 2076 3307 2083 3476
rect 2196 3483 2203 3516
rect 1616 2927 1623 2963
rect 1567 2916 1583 2923
rect 1240 2743 1253 2747
rect 1236 2736 1253 2743
rect 1240 2733 1253 2736
rect 1276 2687 1283 2743
rect 1216 2567 1223 2633
rect 1256 2607 1263 2633
rect 1336 2607 1343 2743
rect 1376 2647 1383 2743
rect 1416 2707 1423 2733
rect 1456 2667 1463 2793
rect 1576 2747 1583 2916
rect 1636 2847 1643 2933
rect 1776 2887 1783 2923
rect 1716 2827 1723 2853
rect 1653 2780 1667 2793
rect 1693 2787 1707 2793
rect 1656 2776 1663 2780
rect 1496 2647 1503 2743
rect 1496 2607 1503 2633
rect 1596 2627 1603 2773
rect 1676 2707 1683 2743
rect 1696 2547 1703 2733
rect 1716 2647 1723 2813
rect 1796 2807 1803 2853
rect 1816 2788 1823 2873
rect 1876 2867 1883 3013
rect 1896 3007 1903 3113
rect 1916 3027 1923 3263
rect 2036 3260 2043 3263
rect 1953 3247 1967 3253
rect 2033 3247 2047 3260
rect 1953 3207 1967 3212
rect 1973 3067 1987 3073
rect 1996 3067 2003 3173
rect 2016 3127 2023 3213
rect 2056 3187 2063 3253
rect 2076 3163 2083 3193
rect 2096 3167 2103 3472
rect 2136 3447 2143 3483
rect 2176 3476 2203 3483
rect 2127 3423 2140 3427
rect 2127 3420 2143 3423
rect 2127 3413 2147 3420
rect 2133 3407 2147 3413
rect 2116 3227 2123 3373
rect 2176 3296 2183 3476
rect 2216 3447 2223 3673
rect 2296 3516 2303 3653
rect 2316 3587 2323 3633
rect 2336 3627 2343 3673
rect 2233 3467 2247 3473
rect 2247 3424 2260 3427
rect 2247 3413 2263 3424
rect 2193 3407 2207 3413
rect 2236 3307 2243 3392
rect 2256 3387 2263 3413
rect 2256 3327 2263 3352
rect 2276 3303 2283 3471
rect 2256 3296 2283 3303
rect 2316 3296 2323 3413
rect 2336 3367 2343 3553
rect 2376 3516 2383 3593
rect 2396 3527 2403 3676
rect 2416 3587 2423 3653
rect 2416 3516 2423 3573
rect 2436 3527 2443 3773
rect 2473 3767 2487 3780
rect 2496 3647 2503 3673
rect 2456 3547 2463 3633
rect 2516 3547 2523 3783
rect 2536 3727 2543 3773
rect 2656 3776 2683 3783
rect 2716 3780 2723 3783
rect 2456 3487 2463 3533
rect 2493 3520 2507 3533
rect 2496 3516 2503 3520
rect 2536 3516 2543 3713
rect 2556 3707 2563 3733
rect 2576 3527 2583 3653
rect 2616 3567 2623 3773
rect 2656 3647 2663 3776
rect 2713 3767 2727 3780
rect 2636 3567 2643 3613
rect 2613 3520 2627 3532
rect 2616 3516 2623 3520
rect 2656 3516 2663 3593
rect 2676 3527 2683 3693
rect 2696 3587 2703 3673
rect 2716 3647 2723 3713
rect 2736 3667 2743 3773
rect 2756 3687 2763 3913
rect 2836 3907 2843 3991
rect 2776 3747 2783 3873
rect 2856 3847 2863 4296
rect 2896 4267 2903 4293
rect 2916 4287 2923 4303
rect 2896 4036 2903 4213
rect 2916 4167 2923 4273
rect 2976 4227 2983 4303
rect 3056 4247 3063 4293
rect 2916 4087 2923 4153
rect 2936 4047 2943 4133
rect 2956 4036 2963 4073
rect 2976 4067 2983 4213
rect 3076 4167 3083 4303
rect 3116 4267 3123 4303
rect 3076 4153 3093 4167
rect 3076 4068 3083 4153
rect 2876 3816 2883 3933
rect 2976 3907 2983 3993
rect 2996 3823 3003 4053
rect 3033 4040 3047 4053
rect 3116 4047 3123 4232
rect 3036 4036 3043 4040
rect 3136 4007 3143 4073
rect 3156 4047 3163 4513
rect 3176 4507 3183 4532
rect 3316 4527 3323 4593
rect 3336 4567 3343 4673
rect 3376 4663 3383 4776
rect 3416 4687 3423 4893
rect 3436 4867 3443 4913
rect 3516 4867 3523 4913
rect 3540 4883 3553 4887
rect 3536 4873 3553 4883
rect 3536 4856 3543 4873
rect 3456 4803 3463 4823
rect 3600 4823 3613 4827
rect 3456 4800 3483 4803
rect 3456 4796 3487 4800
rect 3436 4663 3443 4793
rect 3473 4787 3487 4796
rect 3376 4656 3403 4663
rect 3376 4556 3383 4633
rect 3396 4567 3403 4656
rect 3416 4656 3443 4663
rect 3216 4520 3223 4523
rect 3196 4336 3203 4513
rect 3213 4507 3227 4520
rect 3296 4487 3303 4513
rect 3356 4427 3363 4523
rect 3236 4336 3243 4373
rect 3320 4363 3333 4367
rect 3316 4353 3333 4363
rect 3316 4336 3323 4353
rect 3356 4336 3363 4373
rect 3396 4347 3403 4513
rect 3416 4307 3423 4656
rect 3436 4467 3443 4633
rect 3456 4567 3463 4773
rect 3476 4627 3483 4773
rect 3496 4587 3503 4813
rect 3556 4667 3563 4823
rect 3596 4816 3613 4823
rect 3600 4813 3613 4816
rect 3596 4727 3603 4773
rect 3596 4607 3603 4653
rect 3533 4560 3547 4573
rect 3587 4586 3600 4587
rect 3587 4573 3593 4586
rect 3553 4567 3567 4573
rect 3536 4556 3543 4560
rect 3616 4563 3623 4753
rect 3636 4647 3643 5033
rect 3676 5003 3683 5076
rect 3736 5007 3743 5043
rect 3656 4996 3683 5003
rect 3656 4867 3663 4996
rect 3676 4856 3683 4973
rect 3736 4967 3743 4993
rect 3756 4927 3763 4973
rect 3707 4876 3733 4883
rect 3747 4880 3763 4883
rect 3747 4876 3767 4880
rect 3753 4867 3767 4876
rect 3796 4863 3803 5033
rect 3816 5027 3823 5336
rect 3833 5327 3847 5340
rect 3836 5127 3843 5273
rect 3876 5247 3883 5343
rect 4016 5336 4043 5343
rect 3856 5087 3863 5113
rect 3896 5076 3903 5213
rect 3936 5147 3943 5253
rect 3956 5187 3963 5293
rect 4016 5267 4023 5313
rect 4036 5287 4043 5336
rect 4056 5267 4063 5393
rect 4076 5387 4083 5413
rect 4136 5407 4143 5473
rect 4176 5387 4183 5523
rect 4096 5287 4103 5343
rect 4136 5307 4143 5343
rect 3996 5107 4003 5153
rect 3927 5093 3933 5107
rect 4053 5080 4066 5093
rect 4076 5087 4083 5233
rect 4096 5127 4103 5273
rect 4096 5087 4103 5113
rect 4056 5076 4063 5080
rect 4136 5076 4143 5293
rect 4176 5227 4183 5333
rect 4196 5287 4203 5453
rect 4216 5447 4223 5473
rect 4576 5427 4583 5473
rect 4233 5380 4247 5393
rect 4273 5380 4287 5393
rect 4236 5376 4243 5380
rect 4276 5376 4283 5380
rect 4416 5376 4423 5413
rect 4556 5389 4563 5413
rect 4596 5376 4603 5453
rect 4256 5340 4263 5343
rect 4236 5303 4243 5333
rect 4253 5327 4267 5340
rect 4236 5296 4263 5303
rect 3836 4907 3843 5033
rect 3876 5007 3883 5043
rect 3916 5023 3923 5031
rect 3916 5016 3943 5023
rect 3893 4987 3907 4993
rect 3880 4986 3907 4987
rect 3887 4980 3907 4986
rect 3887 4976 3903 4980
rect 3887 4973 3900 4976
rect 3776 4856 3803 4863
rect 3696 4727 3703 4812
rect 3736 4767 3743 4823
rect 3753 4807 3767 4813
rect 3680 4706 3700 4707
rect 3680 4703 3693 4706
rect 3676 4693 3693 4703
rect 3656 4607 3663 4693
rect 3616 4556 3643 4563
rect 3676 4527 3683 4693
rect 3736 4556 3743 4593
rect 3756 4567 3763 4633
rect 3776 4587 3783 4856
rect 3876 4856 3883 4913
rect 3896 4867 3903 4953
rect 3916 4907 3923 4933
rect 3796 4563 3803 4813
rect 3856 4647 3863 4792
rect 3776 4556 3803 4563
rect 3813 4560 3827 4573
rect 3816 4556 3823 4560
rect 3456 4387 3463 4513
rect 3476 4336 3483 4490
rect 3516 4467 3523 4523
rect 3576 4487 3583 4513
rect 3776 4525 3783 4556
rect 3713 4507 3727 4512
rect 3847 4516 3863 4523
rect 3727 4493 3733 4507
rect 3656 4447 3663 4493
rect 3176 4127 3183 4253
rect 3216 4247 3223 4303
rect 3236 4247 3243 4293
rect 3176 4036 3183 4113
rect 3016 3887 3023 3993
rect 3096 3927 3103 4003
rect 3027 3876 3043 3883
rect 2996 3816 3023 3823
rect 2816 3707 2823 3783
rect 2747 3663 2760 3667
rect 2747 3653 2763 3663
rect 2356 3307 2363 3333
rect 2136 3227 2143 3253
rect 2156 3207 2163 3263
rect 2196 3243 2203 3263
rect 2233 3243 2247 3253
rect 2196 3240 2247 3243
rect 2196 3236 2243 3240
rect 2116 3167 2123 3192
rect 2036 3156 2083 3163
rect 1967 3060 1987 3067
rect 1967 3056 1983 3060
rect 1967 3053 1980 3056
rect 1876 2776 1883 2813
rect 1896 2807 1903 2953
rect 1916 2847 1923 2933
rect 1936 2823 1943 2963
rect 1996 2943 2003 3053
rect 2036 3008 2043 3156
rect 2076 3067 2083 3113
rect 2056 3007 2063 3053
rect 2136 3027 2143 3192
rect 2176 3087 2183 3233
rect 2193 3000 2207 3013
rect 2216 3007 2223 3213
rect 2256 3207 2263 3296
rect 2376 3267 2383 3433
rect 2436 3309 2443 3473
rect 2456 3347 2463 3373
rect 2276 3187 2283 3213
rect 2260 3186 2283 3187
rect 2267 3176 2283 3186
rect 2267 3173 2280 3176
rect 2396 3167 2403 3253
rect 2416 3227 2423 3263
rect 2576 3260 2583 3263
rect 2573 3247 2587 3260
rect 2196 2996 2203 3000
rect 2076 2956 2103 2963
rect 1976 2936 2003 2943
rect 1976 2887 1983 2936
rect 1936 2816 1963 2823
rect 1936 2747 1943 2793
rect 1956 2787 1963 2816
rect 1996 2776 2003 2913
rect 1747 2743 1760 2747
rect 1747 2736 1763 2743
rect 1747 2733 1760 2736
rect 1796 2627 1803 2743
rect 1836 2547 1843 2733
rect 2016 2740 2023 2743
rect 1936 2687 1943 2733
rect 876 2440 883 2443
rect 873 2427 887 2440
rect 956 2427 963 2473
rect 616 2256 623 2373
rect 676 2267 683 2313
rect 696 2256 703 2293
rect 733 2260 747 2273
rect 736 2256 743 2260
rect 856 2256 863 2293
rect 916 2227 923 2255
rect 516 1967 523 2013
rect 536 2003 543 2053
rect 536 1996 563 2003
rect 556 1968 563 1996
rect 436 1907 443 1954
rect 593 1747 607 1753
rect 496 1703 503 1734
rect 496 1696 543 1703
rect 456 1436 463 1493
rect 516 1407 523 1696
rect 576 1647 583 1703
rect 336 1400 343 1403
rect 333 1387 347 1400
rect 133 1220 147 1233
rect 136 1216 143 1220
rect 36 887 43 1173
rect 76 1087 83 1183
rect 196 1087 203 1273
rect 416 1216 423 1373
rect 436 1247 443 1403
rect 596 1287 603 1393
rect 616 1347 623 1893
rect 656 1867 663 1954
rect 676 1887 683 2213
rect 716 2187 723 2223
rect 756 2220 773 2223
rect 753 2216 773 2220
rect 753 2207 767 2216
rect 776 2147 783 2213
rect 876 2167 883 2223
rect 936 2187 943 2293
rect 956 2287 963 2373
rect 976 2327 983 2393
rect 996 2256 1003 2333
rect 1016 2287 1023 2313
rect 1016 2216 1043 2223
rect 976 2167 983 2212
rect 1016 2187 1023 2216
rect 736 1916 763 1923
rect 756 1827 763 1916
rect 776 1907 783 2133
rect 1016 2067 1023 2173
rect 1136 2047 1143 2513
rect 1296 2476 1303 2513
rect 1156 2347 1163 2433
rect 1196 2407 1203 2443
rect 1236 2263 1243 2433
rect 1336 2367 1343 2433
rect 1456 2387 1463 2513
rect 1327 2316 1353 2323
rect 1216 2256 1243 2263
rect 1156 2147 1163 2254
rect 1256 2227 1263 2293
rect 1336 2256 1343 2293
rect 733 1740 747 1753
rect 736 1736 743 1740
rect 636 1707 643 1734
rect 667 1703 680 1707
rect 776 1706 783 1872
rect 796 1747 803 2013
rect 996 1956 1003 2033
rect 1100 1963 1113 1967
rect 1096 1956 1113 1963
rect 1100 1953 1113 1956
rect 816 1767 823 1913
rect 916 1827 923 1953
rect 1136 1927 1143 1973
rect 1193 1960 1207 1973
rect 1196 1956 1203 1960
rect 976 1867 983 1923
rect 916 1787 923 1813
rect 916 1727 923 1773
rect 1016 1767 1023 1923
rect 667 1696 683 1703
rect 667 1693 680 1696
rect 816 1667 823 1703
rect 513 1220 527 1233
rect 516 1216 523 1220
rect 216 1187 223 1214
rect 316 1176 343 1183
rect 336 1107 343 1176
rect 93 920 107 933
rect 96 916 103 920
rect 116 827 123 883
rect 156 867 163 1073
rect 196 880 203 883
rect 193 867 207 880
rect 36 188 43 813
rect 113 740 127 753
rect 236 747 243 883
rect 276 807 283 933
rect 336 916 343 953
rect 396 943 403 1183
rect 436 1180 443 1183
rect 433 1167 447 1180
rect 576 1167 583 1233
rect 616 1216 623 1333
rect 636 1247 643 1633
rect 680 1463 693 1467
rect 676 1453 693 1463
rect 676 1436 683 1453
rect 716 1447 723 1533
rect 816 1527 823 1653
rect 956 1527 963 1703
rect 767 1463 780 1467
rect 767 1453 783 1463
rect 776 1436 783 1453
rect 816 1436 823 1473
rect 856 1443 863 1513
rect 856 1436 883 1443
rect 756 1347 763 1403
rect 736 1256 803 1263
rect 676 1147 683 1183
rect 716 1186 723 1233
rect 736 1227 743 1256
rect 753 1220 767 1233
rect 756 1216 763 1220
rect 796 1216 803 1256
rect 836 1227 843 1273
rect 856 1186 863 1293
rect 893 1220 907 1233
rect 896 1216 903 1220
rect 936 1216 943 1273
rect 696 967 703 1173
rect 376 940 403 943
rect 373 936 403 940
rect 373 927 387 936
rect 580 923 593 927
rect 576 916 593 923
rect 580 913 593 916
rect 356 876 373 883
rect 316 827 323 872
rect 116 736 123 740
rect 67 673 73 687
rect 76 396 83 453
rect 116 407 123 613
rect 296 507 303 733
rect 356 708 363 853
rect 376 807 383 872
rect 416 827 423 883
rect 476 807 483 913
rect 476 696 483 733
rect 516 696 523 753
rect 536 747 543 853
rect 556 847 563 883
rect 596 807 603 873
rect 616 767 623 953
rect 776 947 783 1033
rect 773 907 787 912
rect 316 666 323 693
rect 576 667 583 753
rect 676 696 683 753
rect 796 696 803 1133
rect 816 927 823 1151
rect 976 1147 983 1473
rect 996 1287 1003 1733
rect 1016 1667 1023 1753
rect 1076 1736 1083 1912
rect 1156 1907 1163 1954
rect 1176 1803 1183 1913
rect 1216 1867 1223 1923
rect 1176 1800 1223 1803
rect 1176 1796 1227 1800
rect 1213 1787 1227 1796
rect 1196 1736 1203 1773
rect 1236 1748 1243 1893
rect 1296 1867 1303 2033
rect 1336 1956 1343 2053
rect 1356 1967 1363 2223
rect 1396 2187 1403 2353
rect 1416 2268 1423 2373
rect 1476 2256 1483 2493
rect 1556 2488 1563 2513
rect 1576 2327 1583 2533
rect 1613 2480 1627 2493
rect 1616 2476 1623 2480
rect 1636 2343 1643 2432
rect 1656 2407 1663 2443
rect 1716 2446 1723 2473
rect 1696 2347 1703 2433
rect 1636 2336 1663 2343
rect 1593 2260 1607 2273
rect 1596 2256 1603 2260
rect 1416 2207 1423 2254
rect 1496 2220 1503 2223
rect 1456 2167 1463 2212
rect 1493 2207 1507 2220
rect 1616 2187 1623 2223
rect 1656 2063 1663 2336
rect 1716 2307 1723 2432
rect 1816 2427 1823 2513
rect 1873 2480 1887 2493
rect 1876 2476 1883 2480
rect 1916 2476 1923 2533
rect 1956 2487 1963 2733
rect 2013 2727 2027 2740
rect 2076 2727 2083 2933
rect 2096 2927 2103 2956
rect 2127 2843 2140 2847
rect 2127 2840 2143 2843
rect 2127 2833 2147 2840
rect 2133 2827 2147 2833
rect 2113 2780 2127 2793
rect 2156 2783 2163 2933
rect 2176 2867 2183 2963
rect 2213 2943 2227 2953
rect 2236 2947 2243 3013
rect 2276 2996 2283 3153
rect 2576 3127 2583 3193
rect 2596 3107 2603 3253
rect 2616 3223 2623 3373
rect 2636 3267 2643 3413
rect 2676 3407 2683 3473
rect 2696 3447 2703 3573
rect 2716 3567 2723 3612
rect 2720 3546 2740 3547
rect 2727 3533 2733 3546
rect 2756 3516 2763 3653
rect 2856 3607 2863 3783
rect 2896 3776 2923 3783
rect 2876 3727 2883 3753
rect 2896 3683 2903 3776
rect 2896 3676 2923 3683
rect 2876 3647 2883 3673
rect 2856 3567 2863 3593
rect 2873 3567 2887 3573
rect 2813 3547 2827 3553
rect 2916 3547 2923 3676
rect 2976 3667 2983 3733
rect 3016 3727 3023 3816
rect 3036 3747 3043 3876
rect 3116 3823 3123 3893
rect 3096 3816 3123 3823
rect 3116 3727 3123 3753
rect 3136 3723 3143 3953
rect 3156 3947 3163 3993
rect 3156 3743 3163 3912
rect 3256 3823 3263 4113
rect 3296 4047 3303 4273
rect 3336 4187 3343 4303
rect 3376 4267 3383 4303
rect 3436 4296 3463 4303
rect 3336 4067 3343 4173
rect 3396 4087 3403 4273
rect 3416 4167 3423 4272
rect 3436 4227 3443 4296
rect 3496 4267 3503 4303
rect 3513 4287 3527 4293
rect 3507 4256 3523 4263
rect 3276 3967 3283 3993
rect 3316 3967 3323 4003
rect 3356 3843 3363 3993
rect 3376 3867 3383 4053
rect 3416 4036 3423 4073
rect 3456 4036 3463 4193
rect 3496 4047 3503 4213
rect 3516 4147 3523 4256
rect 3536 4207 3543 4373
rect 3596 4347 3603 4433
rect 3616 4336 3623 4393
rect 3536 4067 3543 4172
rect 3556 4127 3563 4293
rect 3576 4283 3583 4293
rect 3576 4276 3613 4283
rect 3596 4127 3603 4253
rect 3616 4187 3623 4273
rect 3556 4087 3563 4113
rect 3576 4063 3583 4093
rect 3616 4067 3623 4152
rect 3636 4147 3643 4303
rect 3656 4247 3663 4293
rect 3636 4087 3643 4112
rect 3556 4056 3583 4063
rect 3556 4036 3563 4056
rect 3593 4040 3607 4053
rect 3596 4036 3603 4040
rect 3396 3927 3403 3993
rect 3476 3947 3483 4003
rect 3336 3836 3363 3843
rect 3256 3816 3283 3823
rect 3336 3816 3343 3836
rect 3156 3736 3183 3743
rect 3136 3716 3163 3723
rect 3036 3647 3043 3712
rect 2936 3527 2943 3633
rect 3056 3587 3063 3653
rect 3156 3627 3163 3716
rect 3176 3667 3183 3736
rect 2916 3516 2933 3523
rect 2973 3520 2987 3533
rect 2976 3516 2983 3520
rect 2836 3487 2843 3513
rect 2716 3363 2723 3473
rect 2736 3387 2743 3472
rect 2756 3367 2763 3433
rect 2776 3427 2783 3483
rect 2847 3476 2863 3483
rect 2696 3360 2723 3363
rect 2693 3356 2723 3360
rect 2693 3347 2707 3356
rect 2856 3347 2863 3476
rect 2936 3387 2943 3473
rect 2956 3427 2963 3453
rect 3076 3407 3083 3613
rect 3096 3547 3103 3593
rect 2700 3323 2713 3327
rect 2696 3313 2713 3323
rect 2696 3296 2703 3313
rect 2747 3296 2783 3303
rect 2840 3263 2853 3267
rect 2716 3260 2723 3263
rect 2713 3247 2727 3260
rect 2616 3216 2643 3223
rect 2636 3147 2643 3216
rect 2796 3207 2803 3263
rect 2836 3256 2853 3263
rect 2840 3253 2853 3256
rect 2316 2996 2323 3073
rect 2373 3000 2387 3013
rect 2376 2996 2383 3000
rect 2296 2960 2303 2963
rect 2293 2947 2307 2960
rect 2476 2963 2483 3013
rect 2616 3003 2623 3113
rect 2596 2996 2623 3003
rect 2456 2956 2483 2963
rect 2196 2940 2227 2943
rect 2196 2936 2223 2940
rect 2116 2776 2123 2780
rect 2156 2776 2183 2783
rect 2176 2743 2183 2776
rect 2196 2747 2203 2936
rect 2316 2827 2323 2893
rect 2356 2867 2363 2953
rect 2436 2747 2443 2774
rect 2156 2736 2183 2743
rect 2136 2607 2143 2732
rect 2156 2627 2163 2736
rect 2276 2727 2283 2743
rect 2316 2736 2343 2743
rect 1836 2407 1843 2433
rect 1796 2327 1803 2393
rect 1676 2267 1683 2293
rect 1816 2256 1823 2333
rect 1856 2267 1863 2443
rect 1896 2440 1903 2443
rect 1893 2427 1907 2440
rect 1716 2216 1733 2223
rect 1656 2056 1673 2063
rect 1476 1996 1523 2003
rect 1476 1963 1483 1996
rect 1456 1956 1483 1963
rect 1493 1960 1507 1973
rect 1516 1967 1523 1996
rect 1496 1956 1503 1960
rect 1416 1827 1423 1953
rect 1676 1947 1683 2053
rect 1716 2007 1723 2216
rect 1776 2187 1783 2253
rect 1840 2223 1853 2227
rect 1836 2213 1853 2223
rect 1667 1933 1683 1947
rect 1556 1827 1563 1932
rect 1616 1847 1623 1883
rect 1316 1736 1323 1773
rect 1356 1743 1363 1813
rect 1356 1736 1383 1743
rect 1236 1707 1243 1734
rect 1096 1547 1103 1693
rect 1096 1403 1103 1533
rect 1116 1527 1123 1673
rect 1336 1567 1343 1653
rect 1056 1396 1103 1403
rect 996 1187 1003 1233
rect 876 916 883 993
rect 827 883 840 887
rect 916 883 923 1133
rect 1036 1107 1043 1183
rect 933 928 947 933
rect 1016 916 1023 953
rect 1036 923 1043 1093
rect 1076 1047 1083 1273
rect 1116 1187 1123 1513
rect 1176 1436 1183 1533
rect 1273 1523 1287 1533
rect 1273 1520 1303 1523
rect 1276 1516 1303 1520
rect 1276 1448 1283 1493
rect 1296 1467 1303 1516
rect 1316 1436 1323 1533
rect 1156 1247 1163 1403
rect 1216 1187 1223 1313
rect 1236 1187 1243 1273
rect 1256 1247 1263 1403
rect 1296 1227 1303 1403
rect 1356 1247 1363 1633
rect 1436 1607 1443 1773
rect 1376 1287 1383 1593
rect 1413 1440 1427 1453
rect 1416 1436 1423 1440
rect 1456 1436 1463 1653
rect 1496 1627 1503 1703
rect 1556 1696 1583 1703
rect 1516 1567 1523 1593
rect 1436 1307 1443 1403
rect 1496 1400 1503 1403
rect 1493 1387 1507 1400
rect 1556 1307 1563 1473
rect 1576 1447 1583 1696
rect 1596 1627 1603 1753
rect 1636 1736 1643 1813
rect 1696 1703 1703 1953
rect 1716 1787 1723 1993
rect 1776 1956 1783 2033
rect 1816 1956 1823 2133
rect 1836 1967 1843 2213
rect 1876 2107 1883 2393
rect 1956 2147 1963 2213
rect 1756 1907 1763 1923
rect 1756 1896 1773 1907
rect 1760 1893 1773 1896
rect 1836 1887 1843 1911
rect 1856 1907 1863 2033
rect 1916 1956 1923 1993
rect 1976 1963 1983 2453
rect 1996 2347 2003 2493
rect 2196 2476 2203 2513
rect 2276 2507 2283 2713
rect 2316 2627 2323 2736
rect 2456 2627 2463 2956
rect 2556 2943 2563 2952
rect 2556 2936 2583 2943
rect 2576 2803 2583 2936
rect 2596 2907 2603 2996
rect 2716 2967 2723 3093
rect 2756 2996 2763 3133
rect 2836 3127 2843 3233
rect 2856 3147 2863 3232
rect 2876 3107 2883 3353
rect 2896 3307 2903 3373
rect 2933 3300 2947 3313
rect 2936 3296 2943 3300
rect 3016 3303 3023 3393
rect 3016 3296 3043 3303
rect 2896 3047 2903 3253
rect 2916 3167 2923 3263
rect 2956 3260 2963 3263
rect 2953 3247 2967 3260
rect 2936 3207 2943 3233
rect 2636 2927 2643 2963
rect 2636 2843 2643 2913
rect 2636 2836 2663 2843
rect 2596 2808 2603 2833
rect 2556 2796 2583 2803
rect 2536 2567 2543 2653
rect 2556 2647 2563 2796
rect 2627 2736 2643 2743
rect 2296 2476 2303 2513
rect 2473 2480 2487 2493
rect 2476 2476 2483 2480
rect 2236 2447 2243 2474
rect 2036 2407 2043 2443
rect 2016 2267 2023 2353
rect 2096 2267 2103 2333
rect 2136 2327 2143 2443
rect 2176 2367 2183 2443
rect 2236 2263 2243 2293
rect 2256 2287 2263 2474
rect 2516 2447 2523 2513
rect 2236 2256 2263 2263
rect 1996 2147 2003 2253
rect 2076 2107 2083 2223
rect 1956 1956 1983 1963
rect 2016 1956 2023 2033
rect 2116 1987 2123 2213
rect 2136 2187 2143 2223
rect 2176 2147 2183 2223
rect 2216 2167 2223 2253
rect 1896 1920 1903 1923
rect 1756 1767 1763 1813
rect 1776 1736 1783 1833
rect 1836 1707 1843 1873
rect 1656 1627 1663 1703
rect 1696 1696 1723 1703
rect 1616 1436 1623 1473
rect 1313 1220 1327 1233
rect 1393 1220 1407 1233
rect 1436 1227 1443 1293
rect 1316 1216 1323 1220
rect 1396 1216 1403 1220
rect 1036 916 1073 923
rect 1133 920 1147 933
rect 1136 916 1143 920
rect 827 876 843 883
rect 916 876 943 883
rect 827 873 840 876
rect 907 853 913 867
rect 936 843 943 876
rect 916 836 943 843
rect 856 667 863 813
rect 896 787 903 832
rect 916 696 923 836
rect 1056 767 1063 873
rect 1196 787 1203 1173
rect 1456 1167 1463 1233
rect 1576 1216 1583 1273
rect 1596 1227 1603 1253
rect 1696 1243 1703 1393
rect 1716 1387 1723 1696
rect 1747 1696 1763 1703
rect 1696 1236 1713 1243
rect 1476 1147 1483 1213
rect 1716 1207 1723 1233
rect 1556 1180 1563 1183
rect 1553 1167 1567 1180
rect 1676 1147 1683 1183
rect 1547 1136 1573 1143
rect 1396 927 1403 953
rect 1476 916 1483 953
rect 1496 947 1503 973
rect 1296 886 1303 913
rect 1296 807 1303 872
rect 1393 867 1407 873
rect 376 647 383 663
rect 376 636 393 647
rect 380 633 393 636
rect 196 146 203 493
rect 416 467 423 653
rect 453 647 467 653
rect 776 627 783 663
rect 313 400 327 413
rect 316 396 323 400
rect 416 396 423 453
rect 536 396 543 613
rect 816 567 823 663
rect 876 656 903 663
rect 876 627 883 656
rect 996 627 1003 663
rect 1096 627 1103 753
rect 1416 747 1423 913
rect 1456 847 1463 883
rect 1476 827 1483 853
rect 1556 847 1563 993
rect 1616 916 1623 973
rect 1656 916 1663 973
rect 1116 666 1123 733
rect 1256 696 1263 733
rect 1293 700 1307 713
rect 1296 696 1303 700
rect 1216 627 1223 694
rect 1476 703 1483 813
rect 1476 696 1503 703
rect 1356 666 1363 693
rect 1396 627 1403 663
rect 496 367 503 394
rect 396 360 403 363
rect 393 347 407 360
rect 356 147 363 213
rect 396 188 403 333
rect 436 176 443 213
rect 316 140 323 143
rect 196 87 203 132
rect 313 127 327 140
rect 496 146 503 173
rect 416 87 423 143
rect 696 127 703 413
rect 813 400 827 413
rect 816 396 823 400
rect 716 307 723 394
rect 853 347 867 352
rect 876 347 883 613
rect 996 367 1003 553
rect 1096 427 1103 613
rect 1116 403 1123 493
rect 1096 396 1123 403
rect 1133 400 1147 413
rect 1193 400 1207 413
rect 1136 396 1143 400
rect 1196 396 1203 400
rect 916 360 923 363
rect 913 347 927 360
rect 956 207 963 363
rect 1036 307 1043 363
rect 1076 327 1083 363
rect 953 180 967 193
rect 956 176 963 180
rect 1076 176 1083 233
rect 1236 207 1243 493
rect 1256 327 1263 533
rect 1556 507 1563 833
rect 1636 787 1643 883
rect 1676 827 1683 883
rect 1716 847 1723 933
rect 1736 927 1743 1633
rect 1756 1447 1763 1696
rect 1816 1527 1823 1693
rect 1856 1627 1863 1773
rect 1876 1747 1883 1913
rect 1893 1907 1907 1920
rect 1936 1887 1943 1923
rect 2036 1827 2043 1923
rect 1916 1736 1923 1813
rect 1953 1740 1967 1753
rect 1956 1736 1963 1740
rect 2016 1736 2023 1773
rect 2096 1747 2103 1953
rect 2116 1767 2123 1973
rect 2316 1967 2323 2443
rect 2296 1956 2313 1963
rect 2116 1707 2123 1753
rect 2176 1736 2183 1793
rect 2196 1767 2203 1923
rect 2236 1863 2243 1913
rect 2236 1856 2253 1863
rect 1876 1436 1883 1693
rect 1896 1683 1903 1703
rect 1896 1676 1923 1683
rect 1916 1403 1923 1676
rect 1936 1627 1943 1703
rect 1976 1607 1983 1693
rect 2036 1683 2043 1703
rect 2076 1700 2083 1703
rect 2016 1676 2043 1683
rect 2073 1687 2087 1700
rect 1956 1436 1963 1553
rect 2016 1527 2023 1676
rect 2196 1683 2203 1693
rect 2167 1676 2203 1683
rect 2216 1667 2223 1693
rect 2156 1567 2163 1613
rect 1996 1436 2003 1473
rect 1916 1396 1943 1403
rect 1816 1223 1823 1363
rect 1856 1227 1863 1273
rect 1816 1216 1843 1223
rect 1836 947 1843 1216
rect 1896 1216 1903 1253
rect 1936 1227 1943 1396
rect 1956 1187 1963 1373
rect 2036 1287 2043 1553
rect 2116 1436 2123 1493
rect 2156 1447 2163 1513
rect 2236 1507 2243 1793
rect 2256 1743 2263 1853
rect 2276 1767 2283 1923
rect 2256 1736 2283 1743
rect 2316 1736 2323 1913
rect 2336 1743 2343 2333
rect 2376 2256 2383 2293
rect 2416 2256 2423 2393
rect 2456 2307 2463 2443
rect 2556 2440 2563 2443
rect 2553 2427 2567 2440
rect 2467 2263 2480 2267
rect 2467 2256 2483 2263
rect 2516 2256 2523 2333
rect 2556 2267 2563 2353
rect 2467 2253 2480 2256
rect 2576 2247 2583 2293
rect 2616 2268 2623 2711
rect 2636 2367 2643 2736
rect 2656 2727 2663 2836
rect 2676 2787 2683 2813
rect 2756 2807 2763 2833
rect 2776 2827 2783 2963
rect 2836 2867 2843 2993
rect 2956 2967 2963 3013
rect 2856 2927 2863 2953
rect 2976 2966 2983 3033
rect 3013 3000 3027 3013
rect 3056 3008 3063 3153
rect 3016 2996 3023 3000
rect 3096 3003 3103 3533
rect 3176 3527 3183 3573
rect 3196 3387 3203 3783
rect 3216 3627 3223 3773
rect 3236 3747 3243 3783
rect 3236 3547 3243 3733
rect 3256 3523 3263 3653
rect 3276 3587 3283 3816
rect 3296 3587 3303 3753
rect 3356 3727 3363 3783
rect 3396 3687 3403 3773
rect 3416 3727 3423 3933
rect 3436 3827 3443 3933
rect 3476 3916 3483 3933
rect 3516 3887 3523 3933
rect 3536 3927 3543 4003
rect 3556 3907 3563 3973
rect 3576 3887 3583 4003
rect 3636 3967 3643 4052
rect 3656 4047 3663 4233
rect 3676 4167 3683 4473
rect 3696 4347 3703 4393
rect 3736 4336 3743 4453
rect 3756 4407 3763 4473
rect 3756 4363 3763 4393
rect 3756 4356 3783 4363
rect 3776 4336 3783 4356
rect 3816 4347 3823 4493
rect 3716 4300 3723 4303
rect 3713 4287 3727 4300
rect 3696 4036 3703 4233
rect 3736 4127 3743 4253
rect 3756 4127 3763 4303
rect 3776 4107 3783 4293
rect 3836 4247 3843 4413
rect 3856 4347 3863 4516
rect 3876 4487 3883 4753
rect 3896 4687 3903 4813
rect 3916 4747 3923 4893
rect 3936 4827 3943 5016
rect 3976 4887 3983 5073
rect 3996 4856 4003 5013
rect 4036 4987 4043 5043
rect 4076 5003 4083 5033
rect 4116 5007 4123 5043
rect 4056 4996 4083 5003
rect 4056 4927 4063 4996
rect 4156 4987 4163 5043
rect 4076 4856 4083 4893
rect 4156 4863 4163 4973
rect 4176 4967 4183 5033
rect 4196 4947 4203 5252
rect 4236 5087 4243 5273
rect 4256 5147 4263 5296
rect 4296 5076 4303 5193
rect 4316 5187 4323 5253
rect 4336 5167 4343 5373
rect 4387 5336 4403 5343
rect 4436 5340 4443 5343
rect 4316 5087 4323 5133
rect 4216 5043 4223 5073
rect 4336 5046 4343 5113
rect 4376 5088 4383 5333
rect 4433 5327 4447 5340
rect 4556 5343 4563 5375
rect 4516 5336 4563 5343
rect 4476 5227 4483 5333
rect 4416 5076 4423 5213
rect 4556 5087 4563 5193
rect 4656 5167 4663 5413
rect 5033 5380 5047 5393
rect 5036 5376 5043 5380
rect 4736 5307 4743 5333
rect 4716 5296 4733 5303
rect 4676 5207 4683 5233
rect 4216 5036 4243 5043
rect 4156 4856 4183 4863
rect 4216 4856 4223 5013
rect 4236 4927 4243 5036
rect 4256 4856 4263 5013
rect 4296 4867 4303 5013
rect 4396 4987 4403 5043
rect 4027 4816 4043 4823
rect 3936 4727 3943 4813
rect 3896 4347 3903 4673
rect 3936 4556 3943 4673
rect 3996 4607 4003 4673
rect 3916 4447 3923 4463
rect 3916 4336 3923 4433
rect 3956 4407 3963 4523
rect 3940 4303 3953 4307
rect 3936 4296 3953 4303
rect 3940 4293 3953 4296
rect 3760 4106 3783 4107
rect 3767 4096 3783 4106
rect 3767 4093 3780 4096
rect 3816 4083 3823 4193
rect 3876 4187 3883 4293
rect 3816 4076 3843 4083
rect 3713 4067 3727 4073
rect 3807 4053 3813 4067
rect 3836 4047 3843 4076
rect 3667 4003 3680 4007
rect 3667 3993 3683 4003
rect 3716 4000 3723 4003
rect 3456 3829 3463 3853
rect 3536 3828 3543 3853
rect 3596 3847 3603 3913
rect 3636 3786 3643 3833
rect 3656 3827 3663 3893
rect 3676 3867 3683 3993
rect 3713 3987 3727 4000
rect 3816 4000 3823 4003
rect 3680 3846 3700 3847
rect 3687 3843 3700 3846
rect 3687 3833 3703 3843
rect 3696 3816 3703 3833
rect 3736 3827 3743 3993
rect 3813 3987 3827 4000
rect 3816 3843 3823 3973
rect 3836 3887 3843 3993
rect 3856 3927 3863 4153
rect 3896 4127 3903 4273
rect 3916 4267 3923 4293
rect 3976 4287 3983 4433
rect 3996 4387 4003 4513
rect 4016 4507 4023 4773
rect 4036 4567 4043 4816
rect 4096 4803 4103 4823
rect 4076 4796 4103 4803
rect 4076 4647 4083 4796
rect 4136 4787 4143 4823
rect 4176 4807 4183 4856
rect 4056 4556 4063 4593
rect 4216 4576 4223 4693
rect 4236 4687 4243 4823
rect 4260 4805 4280 4807
rect 4267 4793 4273 4805
rect 4153 4560 4167 4573
rect 4156 4556 4163 4560
rect 4076 4520 4083 4523
rect 4036 4447 4043 4513
rect 4073 4507 4087 4520
rect 4196 4487 4203 4523
rect 4036 4407 4043 4433
rect 4196 4407 4203 4473
rect 4033 4340 4047 4353
rect 4036 4336 4043 4340
rect 4076 4336 4083 4393
rect 4107 4353 4113 4367
rect 4167 4363 4180 4367
rect 4167 4353 4183 4363
rect 4176 4336 4183 4353
rect 4216 4336 4223 4413
rect 3876 4047 3883 4073
rect 3896 4036 3903 4113
rect 3816 3836 3843 3843
rect 3836 3828 3843 3836
rect 3876 3807 3883 3973
rect 3916 3947 3923 4003
rect 3956 3947 3963 4213
rect 3976 4067 3983 4173
rect 3996 4047 4003 4153
rect 4016 4047 4023 4272
rect 4056 4107 4063 4303
rect 4087 4293 4093 4307
rect 4076 4067 4083 4113
rect 4053 4047 4067 4053
rect 4096 4043 4103 4153
rect 4116 4067 4123 4332
rect 4276 4307 4283 4473
rect 4296 4467 4303 4813
rect 4316 4767 4323 4933
rect 4416 4896 4423 4993
rect 4496 4987 4503 5043
rect 4536 5007 4543 5043
rect 4576 5007 4583 5093
rect 4596 4927 4603 5113
rect 4633 5080 4647 5093
rect 4636 5076 4643 5080
rect 4676 5076 4683 5193
rect 4696 5107 4703 5153
rect 4716 5087 4723 5296
rect 4736 5107 4743 5233
rect 4796 5167 4803 5373
rect 4856 5207 4863 5343
rect 4896 5287 4903 5343
rect 4756 5087 4763 5153
rect 4796 5076 4803 5113
rect 4876 5087 4883 5273
rect 4867 5076 4883 5087
rect 4916 5076 4923 5153
rect 4936 5087 4943 5375
rect 5336 5346 5343 5433
rect 5453 5380 5467 5393
rect 5513 5380 5527 5393
rect 5456 5376 5463 5380
rect 5516 5376 5523 5380
rect 4867 5073 4880 5076
rect 4616 4863 4623 5033
rect 4656 4987 4663 5043
rect 4656 4867 4663 4952
rect 4676 4907 4683 5013
rect 4736 4967 4743 5072
rect 4816 5040 4823 5043
rect 4813 5027 4827 5040
rect 4853 5027 4867 5033
rect 4616 4856 4643 4863
rect 4336 4827 4343 4854
rect 4336 4787 4343 4813
rect 4356 4767 4363 4793
rect 4396 4687 4403 4713
rect 4356 4568 4363 4673
rect 4416 4627 4423 4773
rect 4536 4767 4543 4812
rect 4596 4747 4603 4823
rect 4616 4787 4623 4813
rect 4636 4727 4643 4856
rect 4676 4856 4683 4893
rect 4316 4427 4323 4513
rect 4336 4367 4343 4523
rect 4376 4487 4383 4523
rect 4196 4296 4223 4303
rect 4196 4167 4203 4273
rect 4216 4267 4223 4296
rect 4136 4047 4143 4113
rect 4296 4083 4303 4353
rect 4333 4340 4347 4353
rect 4336 4336 4343 4340
rect 4376 4336 4383 4433
rect 4436 4367 4443 4713
rect 4696 4707 4703 4823
rect 4533 4627 4547 4633
rect 4476 4336 4483 4492
rect 4616 4427 4623 4553
rect 4636 4403 4643 4513
rect 4676 4487 4683 4523
rect 4716 4407 4723 4523
rect 4756 4507 4763 4733
rect 4776 4607 4783 4853
rect 4796 4826 4803 4973
rect 4896 4883 4903 5031
rect 4876 4876 4903 4883
rect 4876 4856 4883 4876
rect 4916 4867 4923 5013
rect 4936 4987 4943 5033
rect 4956 5027 4963 5313
rect 4976 5107 4983 5343
rect 5016 5340 5023 5343
rect 5013 5327 5027 5340
rect 5116 5247 5123 5343
rect 5156 5167 5163 5343
rect 5236 5340 5243 5343
rect 5233 5327 5247 5340
rect 5256 5336 5283 5343
rect 4973 5087 4987 5093
rect 5033 5080 5047 5093
rect 5036 5076 5043 5080
rect 5176 5076 5183 5253
rect 5016 5040 5023 5043
rect 5013 5027 5027 5040
rect 5096 5007 5103 5073
rect 4936 4867 4943 4913
rect 4956 4856 4963 4893
rect 4996 4868 5003 4993
rect 4816 4647 4823 4793
rect 4836 4647 4843 4813
rect 4856 4787 4863 4823
rect 4976 4787 4983 4812
rect 5016 4707 5023 4823
rect 5056 4747 5063 4893
rect 5116 4869 5123 5033
rect 5156 4856 5163 4893
rect 5216 4867 5223 5033
rect 5236 4887 5243 5113
rect 5256 5047 5263 5336
rect 5336 5127 5343 5332
rect 5356 5187 5363 5373
rect 5576 5267 5583 5343
rect 5296 5100 5353 5104
rect 5293 5093 5353 5100
rect 5293 5087 5307 5093
rect 5306 5080 5307 5087
rect 5353 5080 5367 5093
rect 5356 5076 5363 5080
rect 5416 5076 5423 5133
rect 5456 5076 5463 5113
rect 5473 5087 5487 5093
rect 5256 4856 5263 4993
rect 5296 4903 5303 5043
rect 5336 5007 5343 5043
rect 5436 4907 5443 5043
rect 5496 4963 5503 5133
rect 5516 5087 5523 5173
rect 5573 5080 5587 5093
rect 5616 5087 5623 5373
rect 5576 5076 5583 5080
rect 5516 5007 5523 5033
rect 5556 5007 5563 5043
rect 5496 4956 5523 4963
rect 5456 4936 5493 4943
rect 5296 4896 5323 4903
rect 5293 4860 5307 4873
rect 5316 4867 5323 4896
rect 5296 4856 5303 4860
rect 5193 4827 5207 4833
rect 5136 4820 5143 4823
rect 5133 4807 5147 4820
rect 5156 4707 5163 4813
rect 5336 4727 5343 4893
rect 5456 4856 5463 4936
rect 5476 4867 5483 4913
rect 4776 4567 4783 4593
rect 4793 4560 4807 4573
rect 4796 4556 4803 4560
rect 4836 4556 4843 4633
rect 4616 4396 4643 4403
rect 4616 4336 4623 4396
rect 4636 4343 4643 4396
rect 4636 4336 4663 4343
rect 4356 4247 4363 4303
rect 4296 4076 4323 4083
rect 4096 4036 4123 4043
rect 4153 4040 4167 4053
rect 4156 4036 4163 4040
rect 4316 4047 4323 4076
rect 3916 3867 3923 3933
rect 3976 3907 3983 4013
rect 4036 4000 4043 4003
rect 3940 3883 3953 3887
rect 3936 3873 3953 3883
rect 3936 3816 3943 3873
rect 3976 3823 3983 3853
rect 3996 3847 4003 3993
rect 4033 3987 4047 4000
rect 4016 3847 4023 3953
rect 4096 3927 4103 3993
rect 4136 3923 4143 4003
rect 4196 3967 4203 4034
rect 4136 3916 4163 3923
rect 4036 3828 4043 3893
rect 3976 3816 4003 3823
rect 3236 3516 3263 3523
rect 3216 3407 3223 3513
rect 3236 3303 3243 3516
rect 3396 3516 3403 3633
rect 3456 3527 3463 3613
rect 3256 3367 3263 3473
rect 3296 3447 3303 3483
rect 3367 3476 3383 3483
rect 3276 3307 3283 3393
rect 3356 3347 3363 3473
rect 3236 3296 3263 3303
rect 3116 3127 3123 3293
rect 3156 3227 3163 3263
rect 3216 3256 3243 3263
rect 3136 3107 3143 3193
rect 3096 2996 3113 3003
rect 3176 2996 3183 3033
rect 3236 3008 3243 3256
rect 3256 3187 3263 3296
rect 3336 3256 3363 3263
rect 3296 3107 3303 3253
rect 3356 3167 3363 3256
rect 3076 2867 3083 2963
rect 2656 2627 2663 2692
rect 2716 2607 2723 2743
rect 2816 2707 2823 2743
rect 2916 2667 2923 2853
rect 3096 2847 3103 2913
rect 3116 2776 3123 2873
rect 2936 2746 2943 2773
rect 3036 2727 3043 2753
rect 3056 2747 3063 2773
rect 3136 2740 3143 2743
rect 3133 2727 3147 2740
rect 2673 2480 2687 2493
rect 2676 2476 2683 2480
rect 2927 2483 2940 2487
rect 2927 2476 2943 2483
rect 2927 2473 2940 2476
rect 3036 2487 3043 2713
rect 3007 2474 3013 2487
rect 3000 2473 3013 2474
rect 3176 2487 3183 2933
rect 3236 2883 3243 2994
rect 3336 2887 3343 2993
rect 3356 2966 3363 3073
rect 3376 3027 3383 3353
rect 3416 3303 3423 3483
rect 3456 3447 3463 3473
rect 3396 3296 3423 3303
rect 3456 3296 3463 3393
rect 3476 3327 3483 3733
rect 3496 3647 3503 3753
rect 3516 3747 3523 3773
rect 3556 3747 3563 3783
rect 3556 3647 3563 3673
rect 3676 3667 3683 3773
rect 3716 3687 3723 3773
rect 3736 3727 3743 3773
rect 3996 3786 4003 3816
rect 4076 3816 4083 3873
rect 3516 3516 3523 3573
rect 3536 3527 3543 3613
rect 3556 3524 3563 3553
rect 3556 3517 3593 3524
rect 3656 3516 3663 3613
rect 3736 3523 3743 3593
rect 3736 3516 3763 3523
rect 3596 3487 3603 3514
rect 3496 3296 3503 3373
rect 3516 3307 3523 3453
rect 3396 3227 3403 3296
rect 3556 3296 3563 3333
rect 3596 3296 3603 3452
rect 3616 3407 3623 3493
rect 3636 3307 3643 3473
rect 3676 3407 3683 3483
rect 3716 3480 3743 3483
rect 3716 3476 3747 3480
rect 3456 3207 3463 3233
rect 3436 3008 3443 3173
rect 3476 3167 3483 3263
rect 3656 3266 3663 3313
rect 3696 3307 3703 3413
rect 3716 3347 3723 3476
rect 3733 3467 3747 3476
rect 3836 3403 3843 3473
rect 3856 3427 3863 3653
rect 3876 3627 3883 3772
rect 3916 3687 3923 3713
rect 3936 3707 3943 3773
rect 3956 3647 3963 3773
rect 3836 3396 3863 3403
rect 3516 3227 3523 3253
rect 3536 3167 3543 3253
rect 3616 3260 3623 3263
rect 3613 3247 3627 3260
rect 3676 3247 3683 3294
rect 3756 3307 3763 3393
rect 3796 3296 3803 3373
rect 3836 3347 3843 3373
rect 3856 3308 3863 3396
rect 3876 3387 3883 3573
rect 3956 3547 3963 3633
rect 3976 3467 3983 3773
rect 3380 3006 3400 3007
rect 3387 3003 3400 3006
rect 3387 2996 3403 3003
rect 3387 2993 3400 2996
rect 3556 2996 3563 3073
rect 3416 2927 3423 2963
rect 3496 2965 3503 2993
rect 3236 2876 3263 2883
rect 3216 2707 3223 2743
rect 3256 2707 3263 2876
rect 3456 2847 3463 2952
rect 3496 2867 3503 2951
rect 3596 2947 3603 3213
rect 3636 2996 3643 3153
rect 3696 3087 3703 3253
rect 3676 2996 3683 3053
rect 3716 3008 3723 3263
rect 3816 3260 3823 3263
rect 3813 3247 3827 3260
rect 3853 3187 3867 3193
rect 3876 3187 3883 3352
rect 3896 3347 3903 3393
rect 3976 3327 3983 3453
rect 3996 3367 4003 3733
rect 4036 3627 4043 3673
rect 4056 3667 4063 3772
rect 4136 3747 4143 3893
rect 4156 3827 4163 3916
rect 4196 3816 4203 3953
rect 4236 3907 4243 4003
rect 4276 4000 4283 4003
rect 4273 3987 4287 4000
rect 4236 3816 4243 3893
rect 4316 3848 4323 3993
rect 4336 3827 4343 4153
rect 4376 4047 4383 4273
rect 4416 4247 4423 4313
rect 4456 4300 4463 4303
rect 4453 4287 4467 4300
rect 4567 4293 4573 4307
rect 4456 4227 4463 4273
rect 4356 3887 4363 4034
rect 4436 4036 4443 4113
rect 4496 4087 4503 4293
rect 4596 4227 4603 4303
rect 4656 4127 4663 4336
rect 4756 4336 4763 4453
rect 4696 4227 4703 4303
rect 4736 4247 4743 4303
rect 4496 4047 4503 4073
rect 4536 4036 4543 4113
rect 4576 4036 4583 4073
rect 4373 3987 4387 3993
rect 4456 3967 4463 4003
rect 4396 3847 4403 3913
rect 4436 3843 4443 3873
rect 4436 3836 4463 3843
rect 4456 3816 4463 3836
rect 4496 3816 4503 3993
rect 4516 3967 4523 4003
rect 4516 3827 4523 3953
rect 4556 3847 4563 4003
rect 4616 3987 4623 4113
rect 4653 4040 4667 4053
rect 4656 4036 4663 4040
rect 4756 4005 4763 4113
rect 4796 4067 4803 4493
rect 4816 4487 4823 4523
rect 4856 4387 4863 4523
rect 4916 4447 4923 4573
rect 4956 4556 4963 4593
rect 5136 4556 5143 4633
rect 5296 4526 5303 4653
rect 5336 4556 5343 4692
rect 5356 4583 5363 4853
rect 5396 4707 5403 4823
rect 5436 4820 5443 4823
rect 5433 4807 5447 4820
rect 5356 4580 5383 4583
rect 5356 4576 5387 4580
rect 5373 4567 5387 4576
rect 5416 4556 5423 4653
rect 5476 4563 5483 4813
rect 5496 4807 5503 4873
rect 5516 4867 5523 4956
rect 5536 4856 5543 4933
rect 5596 4927 5603 5043
rect 5573 4860 5587 4873
rect 5616 4867 5623 5033
rect 5576 4856 5583 4860
rect 5656 4856 5663 5033
rect 5676 4887 5683 5043
rect 5556 4807 5563 4823
rect 5456 4556 5483 4563
rect 4976 4387 4983 4523
rect 5016 4467 5023 4523
rect 4956 4336 4963 4373
rect 5016 4347 5023 4373
rect 5056 4347 5063 4493
rect 5076 4467 5083 4523
rect 5116 4520 5123 4523
rect 5113 4507 5127 4520
rect 5096 4336 5103 4393
rect 5116 4367 5123 4453
rect 5216 4447 5223 4523
rect 5156 4347 5163 4393
rect 5236 4336 5243 4453
rect 4816 4267 4823 4313
rect 4856 4227 4863 4303
rect 4936 4267 4943 4303
rect 5013 4287 5027 4293
rect 5036 4247 5043 4333
rect 5176 4307 5183 4333
rect 5053 4287 5067 4293
rect 5076 4227 5083 4303
rect 5116 4300 5123 4303
rect 5016 4107 5023 4133
rect 5096 4107 5103 4293
rect 5113 4287 5127 4300
rect 5256 4267 5263 4293
rect 5296 4267 5303 4333
rect 5316 4247 5323 4413
rect 5396 4367 5403 4513
rect 5436 4487 5443 4523
rect 5476 4503 5483 4523
rect 5456 4496 5483 4503
rect 5456 4367 5463 4496
rect 5386 4353 5387 4360
rect 5373 4340 5387 4353
rect 5376 4336 5383 4340
rect 5476 4336 5483 4473
rect 5516 4407 5523 4713
rect 5556 4687 5563 4793
rect 5556 4556 5563 4673
rect 5576 4567 5583 4813
rect 5596 4556 5603 4813
rect 5633 4807 5647 4813
rect 5676 4747 5683 4823
rect 5716 4820 5723 4823
rect 5713 4807 5727 4820
rect 5513 4340 5527 4353
rect 5536 4347 5543 4513
rect 5616 4487 5623 4523
rect 5516 4336 5523 4340
rect 5333 4247 5347 4253
rect 5356 4247 5363 4303
rect 5240 4246 5260 4247
rect 5247 4233 5253 4246
rect 4796 4036 4803 4053
rect 4953 4040 4967 4053
rect 4956 4036 4963 4040
rect 5073 4040 5087 4053
rect 5076 4036 5083 4040
rect 4576 3823 4583 3973
rect 4596 3947 4603 3973
rect 4636 3947 4643 3973
rect 4716 3907 4723 4003
rect 4816 4000 4823 4003
rect 4813 3987 4827 4000
rect 4856 3907 4863 4003
rect 4616 3847 4623 3873
rect 4756 3847 4763 3893
rect 4556 3816 4583 3823
rect 4613 3820 4627 3833
rect 4616 3816 4623 3820
rect 4156 3627 4163 3792
rect 4176 3647 4183 3773
rect 4216 3727 4223 3783
rect 4256 3747 4263 3773
rect 4296 3747 4303 3783
rect 4356 3780 4363 3783
rect 4196 3627 4203 3713
rect 4033 3520 4047 3533
rect 4076 3527 4083 3613
rect 4216 3607 4223 3673
rect 4036 3516 4043 3520
rect 4176 3516 4223 3523
rect 4036 3387 4043 3453
rect 4056 3407 4063 3483
rect 4056 3328 4063 3393
rect 4216 3387 4223 3516
rect 3896 3227 3903 3253
rect 3896 3143 3903 3192
rect 3916 3187 3923 3263
rect 3896 3136 3923 3143
rect 3816 3008 3823 3093
rect 3916 3087 3923 3136
rect 3880 3063 3893 3067
rect 3876 3053 3893 3063
rect 3876 2966 3883 3053
rect 3913 3000 3927 3013
rect 3916 2996 3923 3000
rect 3556 2747 3563 2933
rect 3656 2789 3663 2963
rect 3776 2787 3783 2813
rect 3936 2776 3943 2813
rect 3976 2783 3983 3263
rect 4016 3207 4023 3313
rect 4096 3296 4103 3333
rect 4116 3207 4123 3263
rect 4156 3227 4163 3373
rect 4236 3363 4243 3693
rect 4336 3547 4343 3773
rect 4353 3767 4367 3780
rect 4376 3527 4383 3773
rect 4396 3747 4403 3812
rect 4436 3727 4443 3783
rect 4476 3780 4483 3783
rect 4473 3767 4487 3780
rect 4416 3516 4423 3613
rect 4436 3528 4443 3653
rect 4336 3483 4343 3512
rect 4296 3476 4343 3483
rect 4353 3467 4367 3473
rect 4456 3407 4463 3533
rect 4476 3527 4483 3732
rect 4516 3647 4523 3773
rect 4556 3528 4563 3816
rect 4756 3816 4763 3833
rect 4656 3747 4663 3813
rect 4796 3727 4803 3853
rect 4856 3816 4863 3893
rect 4896 3867 4903 4033
rect 4936 3847 4943 4003
rect 4896 3816 4943 3823
rect 4976 3816 4983 3893
rect 4996 3887 5003 4033
rect 5056 3927 5063 4003
rect 5007 3876 5023 3883
rect 5016 3827 5023 3876
rect 4856 3607 4863 3673
rect 4896 3647 4903 3816
rect 5096 3816 5103 4003
rect 5136 3987 5143 4193
rect 5156 3967 5163 4133
rect 5236 4047 5243 4133
rect 5000 3783 5013 3787
rect 4996 3776 5013 3783
rect 5000 3773 5013 3776
rect 5056 3747 5063 3783
rect 5116 3747 5123 3783
rect 4693 3520 4707 3533
rect 4793 3520 4807 3533
rect 4696 3516 4703 3520
rect 4796 3516 4803 3520
rect 4487 3483 4500 3487
rect 4487 3476 4503 3483
rect 4487 3473 4500 3476
rect 4476 3427 4483 3473
rect 4567 3453 4573 3467
rect 4216 3356 4243 3363
rect 4216 3307 4223 3356
rect 4516 3336 4523 3373
rect 4236 3296 4243 3333
rect 4196 3107 4203 3263
rect 4216 3127 4223 3193
rect 4036 2996 4043 3033
rect 4173 3000 4187 3013
rect 4176 2996 4183 3000
rect 4216 2996 4223 3113
rect 4236 3087 4243 3213
rect 4296 3187 4303 3293
rect 4567 3273 4573 3287
rect 4456 3260 4463 3263
rect 4356 3243 4363 3253
rect 4453 3247 4467 3260
rect 4356 3236 4393 3243
rect 4296 3067 4303 3113
rect 4016 2787 4023 2963
rect 4056 2823 4063 2963
rect 4116 2887 4123 2993
rect 4047 2816 4063 2823
rect 3976 2776 4003 2783
rect 3467 2736 3483 2743
rect 2716 2347 2723 2443
rect 2756 2427 2763 2473
rect 2976 2440 2983 2443
rect 2816 2387 2823 2431
rect 2373 1967 2387 1973
rect 2413 1960 2427 1973
rect 2456 1967 2463 2213
rect 2536 2220 2543 2223
rect 2533 2207 2547 2220
rect 2416 1956 2423 1960
rect 2356 1927 2363 1953
rect 2376 1747 2383 1913
rect 2436 1867 2443 1912
rect 2336 1736 2363 1743
rect 2256 1443 2263 1553
rect 2276 1467 2283 1573
rect 2296 1527 2303 1703
rect 2356 1567 2363 1736
rect 2387 1736 2403 1743
rect 2236 1436 2263 1443
rect 2056 1247 2063 1333
rect 2096 1223 2103 1403
rect 2276 1347 2283 1453
rect 2296 1307 2303 1473
rect 2376 1447 2383 1493
rect 2396 1443 2403 1573
rect 2416 1547 2423 1692
rect 2456 1547 2463 1753
rect 2476 1467 2483 1993
rect 2576 1967 2583 2193
rect 2596 2007 2603 2213
rect 2656 2147 2663 2223
rect 2676 1956 2683 2073
rect 2696 1967 2703 2212
rect 2536 1787 2543 1923
rect 2496 1747 2503 1773
rect 2553 1763 2567 1773
rect 2536 1760 2567 1763
rect 2536 1756 2563 1760
rect 2536 1736 2543 1756
rect 2596 1747 2603 1953
rect 2613 1903 2627 1913
rect 2613 1900 2643 1903
rect 2616 1896 2643 1900
rect 2636 1736 2643 1896
rect 2716 1743 2723 2333
rect 2776 2256 2783 2293
rect 2856 2227 2863 2293
rect 2876 2267 2883 2333
rect 2916 2287 2923 2433
rect 2973 2427 2987 2440
rect 2916 2256 2923 2273
rect 2953 2260 2967 2273
rect 2956 2256 2963 2260
rect 2796 2220 2803 2223
rect 2793 2207 2807 2220
rect 2896 2220 2903 2223
rect 2836 2087 2843 2213
rect 2893 2207 2907 2220
rect 3036 2147 3043 2433
rect 3076 2387 3083 2443
rect 3136 2427 3143 2473
rect 3156 2387 3163 2474
rect 3236 2476 3243 2573
rect 3296 2516 3393 2523
rect 3296 2487 3303 2516
rect 3327 2496 3373 2503
rect 3313 2480 3327 2493
rect 3316 2476 3323 2480
rect 3136 2216 3163 2223
rect 2793 1960 2807 1973
rect 2836 1967 2843 2073
rect 3156 2067 3163 2216
rect 2796 1956 2803 1960
rect 2696 1736 2723 1743
rect 2756 1736 2763 1893
rect 2776 1887 2783 1923
rect 2827 1916 2843 1923
rect 2796 1747 2803 1773
rect 2616 1547 2623 1703
rect 2480 1443 2493 1447
rect 2396 1436 2423 1443
rect 2476 1436 2493 1443
rect 2480 1433 2493 1436
rect 2096 1216 2123 1223
rect 2176 1216 2183 1293
rect 2216 1216 2223 1273
rect 2356 1228 2363 1293
rect 1876 1127 1883 1173
rect 1916 987 1923 1133
rect 1753 920 1767 933
rect 1793 920 1807 933
rect 1756 916 1763 920
rect 1796 916 1803 920
rect 1913 920 1927 933
rect 1936 927 1943 1173
rect 1976 1107 1983 1213
rect 2056 967 2063 1183
rect 2073 1147 2087 1153
rect 2096 1147 2103 1173
rect 2116 1167 2123 1216
rect 2133 1167 2147 1173
rect 2136 1087 2143 1132
rect 2156 1107 2163 1183
rect 2236 1176 2263 1183
rect 2316 1180 2323 1183
rect 2236 1107 2243 1176
rect 2313 1167 2327 1180
rect 1916 916 1923 920
rect 1776 880 1783 883
rect 1576 687 1583 733
rect 1596 707 1603 773
rect 1716 663 1723 812
rect 1736 703 1743 873
rect 1773 867 1787 880
rect 1816 787 1823 883
rect 1816 747 1823 773
rect 1736 696 1763 703
rect 1676 627 1683 663
rect 1696 656 1723 663
rect 1356 367 1363 413
rect 1476 396 1483 493
rect 1327 356 1343 363
rect 1336 327 1343 356
rect 716 146 723 173
rect 856 147 863 173
rect 996 147 1003 173
rect 816 140 823 143
rect 813 127 827 140
rect 936 127 943 143
rect 1013 127 1027 133
rect 936 116 953 127
rect 940 113 953 116
rect 1096 87 1103 143
rect 1136 140 1143 143
rect 1133 127 1147 140
rect 1236 87 1243 193
rect 1356 107 1363 174
rect 1376 127 1383 393
rect 1576 387 1583 513
rect 1696 507 1703 656
rect 1836 627 1843 873
rect 1936 787 1943 873
rect 1956 867 1963 933
rect 2236 916 2243 1072
rect 2276 916 2283 1033
rect 2316 927 2323 1013
rect 2356 987 2363 1214
rect 2336 927 2343 953
rect 2376 943 2383 1333
rect 2496 1327 2503 1393
rect 2516 1267 2523 1533
rect 2616 1507 2623 1533
rect 2536 1347 2543 1453
rect 2636 1403 2643 1693
rect 2656 1627 2663 1703
rect 2696 1647 2703 1736
rect 2716 1436 2723 1473
rect 2736 1467 2743 1703
rect 2816 1687 2823 1891
rect 2836 1767 2843 1916
rect 2856 1907 2863 1993
rect 2876 1967 2883 2013
rect 2893 1960 2907 1973
rect 2896 1956 2903 1960
rect 3076 1956 3083 2013
rect 3156 1983 3163 2053
rect 3136 1976 3163 1983
rect 3136 1956 3143 1976
rect 2876 1887 2883 1913
rect 2916 1847 2923 1923
rect 2956 1920 2963 1923
rect 2936 1867 2943 1913
rect 2953 1907 2967 1920
rect 3016 1847 3023 1893
rect 2856 1767 2863 1813
rect 2853 1740 2867 1753
rect 2856 1736 2863 1740
rect 2796 1447 2803 1493
rect 2836 1436 2843 1473
rect 2876 1467 2883 1673
rect 2896 1667 2903 1703
rect 2896 1627 2903 1653
rect 2936 1627 2943 1773
rect 3016 1736 3023 1773
rect 3076 1667 3083 1734
rect 2636 1396 2653 1403
rect 2416 987 2423 1073
rect 2356 936 2383 943
rect 2076 886 2083 913
rect 2076 847 2083 872
rect 2136 827 2143 883
rect 2067 816 2093 823
rect 1896 696 1903 773
rect 1956 727 1963 793
rect 2056 666 2063 773
rect 2196 747 2203 913
rect 2356 887 2363 936
rect 2396 923 2403 973
rect 2376 916 2403 923
rect 2416 916 2423 973
rect 2476 927 2483 1253
rect 2556 1216 2563 1313
rect 2576 1180 2583 1183
rect 2536 1163 2543 1172
rect 2573 1167 2587 1180
rect 2536 1156 2563 1163
rect 2256 727 2263 883
rect 2296 847 2303 883
rect 2196 696 2243 703
rect 2276 696 2283 773
rect 1416 176 1423 313
rect 1596 247 1603 473
rect 1636 396 1643 433
rect 1716 423 1723 613
rect 1756 547 1763 573
rect 1736 447 1743 493
rect 1696 416 1723 423
rect 1696 396 1703 416
rect 1736 366 1743 412
rect 1756 407 1763 533
rect 1776 456 1813 463
rect 1776 427 1783 456
rect 1796 396 1803 433
rect 1856 407 1863 493
rect 1816 327 1823 363
rect 1856 327 1863 353
rect 1876 347 1883 653
rect 1916 567 1923 653
rect 2156 627 2163 663
rect 2196 587 2203 696
rect 2300 663 2313 667
rect 2296 656 2313 663
rect 2300 653 2313 656
rect 2256 467 2263 613
rect 2336 607 2343 753
rect 2356 647 2363 852
rect 2376 827 2383 916
rect 2556 927 2563 1156
rect 2616 1147 2623 1214
rect 2636 1127 2643 1253
rect 2656 1227 2663 1392
rect 2696 1367 2703 1392
rect 2736 1228 2743 1392
rect 2816 1347 2823 1403
rect 2896 1396 2923 1403
rect 2896 1367 2903 1396
rect 2816 1307 2823 1333
rect 2596 923 2603 1053
rect 2676 987 2683 1093
rect 2676 928 2683 973
rect 2696 943 2703 1133
rect 2716 967 2723 1183
rect 2816 1167 2823 1183
rect 2853 1163 2867 1173
rect 2836 1160 2867 1163
rect 2836 1156 2863 1160
rect 2816 1027 2823 1153
rect 2836 967 2843 1156
rect 2876 1143 2883 1333
rect 2933 1220 2947 1233
rect 2936 1216 2943 1220
rect 2976 1216 2983 1533
rect 2996 1247 3003 1633
rect 3096 1543 3103 1773
rect 3176 1767 3183 2433
rect 3196 2007 3203 2393
rect 3256 2347 3263 2432
rect 3336 2387 3343 2443
rect 3476 2407 3483 2736
rect 3596 2583 3603 2743
rect 3756 2707 3763 2743
rect 3856 2740 3863 2743
rect 3596 2576 3613 2583
rect 3536 2476 3543 2513
rect 3616 2488 3623 2573
rect 3596 2476 3613 2483
rect 3756 2407 3763 2474
rect 3276 2268 3283 2293
rect 3336 2268 3343 2333
rect 3776 2327 3783 2733
rect 3853 2727 3867 2740
rect 3996 2707 4003 2776
rect 4036 2776 4043 2813
rect 4076 2776 4083 2873
rect 4136 2867 4143 2913
rect 3996 2527 4003 2693
rect 4016 2647 4023 2733
rect 4036 2487 4043 2713
rect 4056 2507 4063 2743
rect 4116 2547 4123 2813
rect 4156 2808 4163 2963
rect 4256 2947 4263 3013
rect 4396 3008 4403 3033
rect 4376 2927 4383 2963
rect 4416 2960 4423 2963
rect 4413 2947 4427 2960
rect 4476 2927 4483 3073
rect 4196 2776 4203 2813
rect 4336 2747 4343 2774
rect 4216 2740 4223 2743
rect 4213 2727 4227 2740
rect 4356 2743 4363 2813
rect 4356 2736 4403 2743
rect 4456 2736 4483 2743
rect 4076 2476 4083 2533
rect 3976 2445 3983 2473
rect 4136 2445 4143 2493
rect 4176 2476 4183 2513
rect 3956 2436 3973 2443
rect 3413 2267 3427 2273
rect 3796 2256 3843 2263
rect 3436 2226 3443 2253
rect 3236 2087 3243 2223
rect 3356 2167 3363 2223
rect 3456 2187 3463 2253
rect 3236 1967 3243 2073
rect 3396 1956 3403 1993
rect 3196 1925 3203 1953
rect 3236 1867 3243 1911
rect 3316 1827 3323 1953
rect 3136 1667 3143 1703
rect 3176 1700 3183 1703
rect 3173 1687 3187 1700
rect 3216 1667 3223 1703
rect 3276 1627 3283 1703
rect 3096 1536 3123 1543
rect 3116 1443 3123 1536
rect 3316 1527 3323 1753
rect 3336 1687 3343 1734
rect 3436 1707 3443 2113
rect 3496 1987 3503 2213
rect 3536 2027 3543 2213
rect 3556 2067 3563 2193
rect 3696 2187 3703 2223
rect 3753 2203 3767 2212
rect 3753 2196 3783 2203
rect 3556 2003 3563 2053
rect 3536 1996 3563 2003
rect 3536 1956 3543 1996
rect 3576 1749 3583 2013
rect 3633 1960 3647 1973
rect 3656 1967 3663 2033
rect 3776 1968 3783 2196
rect 3796 2087 3803 2256
rect 3896 2167 3903 2223
rect 3936 2187 3943 2254
rect 3636 1956 3643 1960
rect 3776 1847 3783 1954
rect 3796 1887 3803 1973
rect 3836 1956 3843 1993
rect 3936 1923 3943 2152
rect 3956 2107 3963 2436
rect 4056 2407 4063 2443
rect 4276 2347 4283 2573
rect 4013 2260 4027 2273
rect 4016 2256 4023 2260
rect 4056 2220 4063 2223
rect 4053 2207 4067 2220
rect 4116 2187 4123 2223
rect 3956 1927 3963 1993
rect 3996 1956 4003 2033
rect 4036 1956 4043 2053
rect 3916 1916 3943 1923
rect 3716 1787 3723 1833
rect 3716 1706 3723 1773
rect 3816 1743 3823 1913
rect 3816 1736 3843 1743
rect 3916 1736 3923 1916
rect 4056 1887 4063 1912
rect 3996 1748 4003 1853
rect 3336 1587 3343 1633
rect 3096 1436 3123 1443
rect 3136 1187 3143 1453
rect 2856 1136 2883 1143
rect 2696 936 2723 943
rect 2596 916 2623 923
rect 2476 807 2483 873
rect 2496 863 2503 913
rect 2496 856 2523 863
rect 2373 707 2387 713
rect 2496 667 2503 833
rect 2516 747 2523 856
rect 2556 787 2563 873
rect 2576 807 2583 883
rect 2596 847 2603 873
rect 2556 696 2563 773
rect 2636 696 2643 753
rect 2676 696 2683 813
rect 2696 727 2703 773
rect 2716 703 2723 936
rect 2736 827 2743 913
rect 2796 863 2803 883
rect 2796 856 2823 863
rect 2736 727 2743 813
rect 2816 767 2823 856
rect 2716 696 2743 703
rect 2396 567 2403 663
rect 2436 660 2443 663
rect 2433 647 2447 660
rect 2516 567 2523 593
rect 2376 467 2383 513
rect 1916 407 1923 453
rect 1956 396 1963 433
rect 1453 180 1467 193
rect 1456 176 1463 180
rect 1596 176 1603 233
rect 1496 146 1503 173
rect 1736 147 1743 213
rect 1876 207 1883 333
rect 1976 247 1983 353
rect 1816 196 1863 203
rect 1816 176 1823 196
rect 1856 183 1863 196
rect 1856 176 1883 183
rect 1436 140 1443 143
rect 1433 127 1447 140
rect 1576 140 1583 143
rect 1573 127 1587 140
rect 1876 146 1883 176
rect 1976 176 1983 233
rect 1996 227 2003 433
rect 2016 307 2023 453
rect 2207 416 2233 423
rect 2256 403 2263 453
rect 2256 396 2283 403
rect 2333 400 2347 413
rect 2336 396 2343 400
rect 2076 347 2083 363
rect 2136 347 2143 394
rect 2076 336 2093 347
rect 2080 333 2093 336
rect 1656 107 1663 133
rect 1693 127 1707 133
rect 1956 107 1963 143
rect 2136 146 2143 293
rect 2236 267 2243 363
rect 2376 287 2383 453
rect 2556 447 2563 573
rect 2656 527 2663 663
rect 2736 467 2743 696
rect 2756 667 2763 753
rect 2836 709 2843 953
rect 2856 807 2863 1136
rect 2916 1107 2923 1183
rect 2956 987 2963 1183
rect 2996 1180 3003 1183
rect 2993 1167 3007 1180
rect 3136 1127 3143 1173
rect 3156 1167 3163 1513
rect 3193 1440 3207 1453
rect 3336 1447 3343 1573
rect 3436 1507 3443 1693
rect 3516 1647 3523 1703
rect 3196 1436 3203 1440
rect 3176 1007 3183 1233
rect 3276 1186 3283 1433
rect 3336 1216 3343 1373
rect 3376 1347 3383 1433
rect 3536 1407 3543 1653
rect 3556 1527 3563 1703
rect 3676 1667 3683 1703
rect 3636 1447 3643 1593
rect 3716 1523 3723 1692
rect 3736 1607 3743 1734
rect 3836 1547 3843 1736
rect 3716 1516 3743 1523
rect 3716 1436 3723 1493
rect 3736 1448 3743 1516
rect 3876 1443 3883 1633
rect 3896 1607 3903 1703
rect 4016 1700 4023 1703
rect 4013 1687 4027 1700
rect 4056 1647 4063 1703
rect 3876 1436 3903 1443
rect 3436 1400 3443 1403
rect 3433 1387 3447 1400
rect 3576 1400 3583 1403
rect 3573 1387 3587 1400
rect 3636 1223 3643 1273
rect 3616 1216 3643 1223
rect 3196 1067 3203 1173
rect 3236 1107 3243 1183
rect 3196 947 3203 1053
rect 2973 920 2987 933
rect 2976 916 2983 920
rect 3236 923 3243 1093
rect 3216 916 3243 923
rect 3273 920 3287 933
rect 3316 927 3323 1183
rect 3356 1107 3363 1183
rect 3396 967 3403 1173
rect 3536 1183 3543 1213
rect 3496 1176 3543 1183
rect 3656 1167 3663 1393
rect 3696 1387 3703 1403
rect 3696 1347 3703 1373
rect 3696 1216 3703 1273
rect 3736 1228 3743 1333
rect 3796 1187 3803 1273
rect 3856 1228 3863 1273
rect 3276 916 3283 920
rect 2876 747 2883 873
rect 2916 747 2923 883
rect 2876 696 2883 733
rect 2920 723 2933 727
rect 2916 713 2933 723
rect 2916 696 2923 713
rect 2896 607 2903 663
rect 2976 647 2983 713
rect 2776 427 2783 593
rect 2396 327 2403 373
rect 2436 167 2443 253
rect 2456 147 2463 273
rect 2556 207 2563 363
rect 2516 176 2563 183
rect 2616 176 2623 353
rect 2636 287 2643 393
rect 2756 367 2763 393
rect 2916 396 2923 433
rect 2696 360 2703 363
rect 2693 347 2707 360
rect 2733 347 2747 353
rect 2776 327 2783 392
rect 2976 383 2983 612
rect 2996 407 3003 793
rect 3036 696 3043 813
rect 3076 767 3083 914
rect 3156 880 3163 883
rect 3096 847 3103 873
rect 3153 867 3167 880
rect 3076 696 3083 753
rect 3096 727 3103 833
rect 3196 707 3203 793
rect 3216 666 3223 916
rect 3373 920 3387 933
rect 3376 916 3383 920
rect 3416 916 3423 1033
rect 3456 927 3463 993
rect 3556 987 3563 1033
rect 3547 956 3573 963
rect 3476 916 3483 953
rect 3676 927 3683 953
rect 3116 660 3123 663
rect 3113 647 3127 660
rect 3047 636 3073 643
rect 3056 396 3063 433
rect 3096 396 3103 533
rect 3236 487 3243 873
rect 3256 847 3263 883
rect 3296 880 3303 883
rect 3293 867 3307 880
rect 3396 880 3403 883
rect 3393 867 3407 880
rect 3296 787 3303 853
rect 3293 700 3307 713
rect 3436 707 3443 853
rect 3296 696 3303 700
rect 3416 660 3423 663
rect 3413 647 3427 660
rect 3436 627 3443 653
rect 3196 408 3203 453
rect 2976 376 3003 383
rect 2896 360 2903 363
rect 2833 347 2847 352
rect 2893 347 2907 360
rect 1567 96 1593 103
rect 1996 87 2003 133
rect 2076 87 2083 143
rect 2296 107 2303 143
rect 2356 27 2363 133
rect 2396 67 2403 143
rect 2427 93 2433 107
rect 2487 93 2493 107
rect 2556 27 2563 176
rect 2696 146 2703 233
rect 2716 187 2723 273
rect 2756 176 2763 233
rect 2776 187 2783 313
rect 2936 287 2943 363
rect 2996 363 3003 376
rect 2996 356 3023 363
rect 2953 307 2967 313
rect 2976 283 2983 351
rect 2993 307 3007 313
rect 2976 276 3003 283
rect 2996 227 3003 276
rect 2856 176 2863 213
rect 3016 187 3023 356
rect 3076 287 3083 363
rect 2596 107 2603 143
rect 2727 143 2740 147
rect 2727 136 2743 143
rect 2836 140 2843 143
rect 2727 133 2740 136
rect 2833 127 2847 140
rect 3036 143 3043 273
rect 2996 136 3043 143
rect 2876 47 2883 132
rect 3056 47 3063 253
rect 3113 180 3127 193
rect 3116 176 3123 180
rect 3156 87 3163 313
rect 3176 207 3183 363
rect 3236 207 3243 473
rect 3256 267 3263 533
rect 3296 487 3303 533
rect 3296 396 3303 473
rect 3416 396 3423 553
rect 3456 407 3463 873
rect 3476 647 3483 773
rect 3576 708 3583 914
rect 3636 696 3643 753
rect 3656 727 3663 793
rect 3696 707 3703 1153
rect 3716 1107 3723 1183
rect 3836 1127 3843 1183
rect 3756 916 3763 993
rect 3896 967 3903 1436
rect 3916 1007 3923 1533
rect 3900 943 3913 947
rect 3896 933 3913 943
rect 3896 916 3903 933
rect 3936 927 3943 1313
rect 4016 1227 4023 1633
rect 4096 1527 4103 2093
rect 4176 1987 4183 2333
rect 4296 2287 4303 2513
rect 4316 2483 4323 2633
rect 4336 2507 4343 2733
rect 4476 2587 4483 2736
rect 4496 2667 4503 3173
rect 4596 3127 4603 3513
rect 4616 3487 4623 3514
rect 4620 3466 4633 3467
rect 4627 3453 4633 3466
rect 4676 3447 4683 3483
rect 4816 3407 4823 3483
rect 4636 3307 4643 3393
rect 4616 3247 4623 3294
rect 4656 3296 4663 3373
rect 4676 3107 4683 3263
rect 4536 3008 4543 3093
rect 4636 2967 4643 3033
rect 4736 3027 4743 3313
rect 4756 3307 4763 3353
rect 4776 3296 4783 3373
rect 4807 3315 4813 3327
rect 4876 3327 4883 3473
rect 4896 3308 4903 3633
rect 4996 3627 5003 3713
rect 4916 3527 4923 3573
rect 5056 3527 5063 3673
rect 5133 3520 5147 3533
rect 5156 3527 5163 3833
rect 5136 3516 5143 3520
rect 5047 3493 5053 3507
rect 5076 3467 5083 3513
rect 4936 3296 4943 3353
rect 4956 3307 4963 3393
rect 5076 3387 5083 3453
rect 4796 3127 4803 3263
rect 4916 3260 4923 3263
rect 4913 3247 4927 3260
rect 4936 3127 4943 3233
rect 4956 3227 4963 3253
rect 4696 3017 4733 3024
rect 4696 3000 4704 3017
rect 4796 3007 4803 3113
rect 4936 3027 4943 3113
rect 4976 3087 4983 3373
rect 4993 3327 5007 3333
rect 5176 3303 5183 3853
rect 5216 3847 5223 4003
rect 5276 3843 5283 4093
rect 5313 4040 5327 4053
rect 5316 4036 5323 4040
rect 5356 4036 5363 4173
rect 5376 4087 5383 4293
rect 5396 4267 5403 4303
rect 5416 4067 5423 4293
rect 5496 4247 5503 4303
rect 5556 4147 5563 4353
rect 5576 4347 5583 4393
rect 5616 4336 5623 4413
rect 5696 4363 5703 4553
rect 5716 4525 5723 4793
rect 5696 4356 5723 4363
rect 5596 4267 5603 4303
rect 5453 4040 5467 4053
rect 5456 4036 5463 4040
rect 5256 3836 5283 3843
rect 5256 3828 5263 3836
rect 5296 3827 5303 3993
rect 5416 3967 5423 4003
rect 5356 3816 5363 3853
rect 5216 3587 5223 3783
rect 5236 3523 5243 3773
rect 5276 3747 5283 3783
rect 5216 3516 5243 3523
rect 5256 3516 5263 3733
rect 5336 3727 5343 3783
rect 5376 3747 5383 3773
rect 5416 3523 5423 3833
rect 5456 3816 5463 3973
rect 5476 3827 5483 3993
rect 5496 3847 5503 4073
rect 5596 4047 5603 4173
rect 5536 3907 5543 4003
rect 5500 3783 5513 3787
rect 5496 3776 5513 3783
rect 5500 3773 5513 3776
rect 5476 3627 5483 3773
rect 5536 3587 5543 3853
rect 5556 3827 5563 3973
rect 5576 3967 5583 4003
rect 5596 3823 5603 3993
rect 5616 3867 5623 4293
rect 5696 4187 5703 4333
rect 5716 4067 5723 4356
rect 5736 4307 5743 4813
rect 5756 4283 5763 5113
rect 5736 4276 5763 4283
rect 5656 3947 5663 4003
rect 5596 3816 5613 3823
rect 5556 3527 5563 3773
rect 5576 3747 5583 3783
rect 5396 3516 5423 3523
rect 5236 3347 5243 3483
rect 5176 3296 5203 3303
rect 5296 3303 5303 3513
rect 5336 3480 5343 3483
rect 5333 3467 5347 3480
rect 5376 3367 5383 3473
rect 5396 3427 5403 3516
rect 5276 3296 5303 3303
rect 5156 3267 5163 3293
rect 4996 3256 5023 3263
rect 4996 3147 5003 3256
rect 5073 3167 5087 3173
rect 4776 2996 4793 3003
rect 4556 2887 4563 2963
rect 4576 2907 4583 2933
rect 4716 2927 4723 2963
rect 4776 2923 4783 2996
rect 4813 3000 4827 3013
rect 5060 3023 5073 3027
rect 4853 3000 4867 3013
rect 4816 2996 4823 3000
rect 4856 2996 4863 3000
rect 4973 3000 4987 3013
rect 5056 3013 5073 3023
rect 4976 2996 4983 3000
rect 5056 2996 5063 3013
rect 5096 2967 5103 3013
rect 4776 2916 4803 2923
rect 4696 2776 4703 2813
rect 4576 2587 4583 2733
rect 4616 2707 4623 2773
rect 4676 2667 4683 2743
rect 4716 2707 4723 2743
rect 4756 2667 4763 2773
rect 4776 2707 4783 2893
rect 4796 2787 4803 2916
rect 4876 2776 4883 2953
rect 4916 2907 4923 2953
rect 4956 2807 4963 2963
rect 5116 2927 5123 3073
rect 5153 3000 5167 3013
rect 5156 2996 5163 3000
rect 5196 2996 5203 3193
rect 5216 3027 5223 3263
rect 5276 3187 5283 3296
rect 5396 3267 5403 3413
rect 5416 3307 5423 3453
rect 5456 3296 5463 3413
rect 5496 3323 5503 3443
rect 5496 3320 5523 3323
rect 5496 3316 5527 3320
rect 5513 3307 5527 3316
rect 5316 3256 5343 3263
rect 5336 3207 5343 3256
rect 5276 2996 5283 3133
rect 5316 3007 5323 3173
rect 5073 2780 5087 2793
rect 5076 2776 5083 2780
rect 5116 2776 5123 2833
rect 4807 2746 4820 2747
rect 4807 2733 4813 2746
rect 4316 2476 4343 2483
rect 4376 2476 4383 2513
rect 4416 2476 4423 2553
rect 4436 2527 4443 2573
rect 4436 2483 4443 2513
rect 4436 2476 4463 2483
rect 4396 2407 4403 2443
rect 4556 2443 4563 2553
rect 4536 2436 4563 2443
rect 4436 2283 4443 2433
rect 4436 2276 4463 2283
rect 4233 2260 4247 2273
rect 4236 2256 4243 2260
rect 4276 2167 4283 2273
rect 4456 2268 4463 2276
rect 4296 2127 4303 2252
rect 4316 2027 4323 2213
rect 4376 2167 4383 2213
rect 4536 2187 4543 2436
rect 4576 2407 4583 2573
rect 4696 2476 4703 2513
rect 4636 2436 4663 2443
rect 4656 2287 4663 2436
rect 4733 2423 4747 2433
rect 4733 2420 4763 2423
rect 4736 2416 4763 2420
rect 4756 2256 4763 2416
rect 4796 2256 4803 2712
rect 4856 2707 4863 2743
rect 4916 2647 4923 2773
rect 4956 2687 4963 2743
rect 4996 2707 5003 2743
rect 5056 2740 5063 2743
rect 5036 2667 5043 2733
rect 5053 2727 5067 2740
rect 5133 2727 5147 2733
rect 5067 2716 5083 2723
rect 4816 2407 4823 2474
rect 5076 2476 5083 2716
rect 5156 2707 5163 2913
rect 5176 2787 5183 2963
rect 5296 2943 5303 2963
rect 5276 2940 5303 2943
rect 5273 2936 5303 2940
rect 5216 2776 5223 2873
rect 5236 2867 5243 2933
rect 5273 2927 5287 2936
rect 5286 2920 5287 2927
rect 5253 2780 5267 2793
rect 5276 2787 5283 2833
rect 5256 2776 5263 2780
rect 5176 2707 5183 2733
rect 5196 2667 5203 2743
rect 5236 2740 5243 2743
rect 5233 2727 5247 2740
rect 5256 2547 5263 2733
rect 5116 2476 5123 2533
rect 5173 2480 5187 2493
rect 5176 2476 5183 2480
rect 4936 2446 4943 2473
rect 4876 2440 4883 2443
rect 4873 2427 4887 2440
rect 4996 2440 5003 2443
rect 4993 2427 5007 2440
rect 4996 2327 5003 2413
rect 4893 2260 4907 2273
rect 4896 2256 4903 2260
rect 4993 2260 5007 2273
rect 4996 2256 5003 2260
rect 4213 1960 4227 1973
rect 4216 1956 4223 1960
rect 4276 1956 4283 2013
rect 4176 1827 4183 1923
rect 4116 1667 4123 1734
rect 4316 1706 4323 1973
rect 4396 1916 4423 1923
rect 4416 1887 4423 1916
rect 4276 1667 4283 1703
rect 4336 1567 4343 1813
rect 4416 1743 4423 1852
rect 4407 1736 4423 1743
rect 4436 1667 4443 2173
rect 4533 2047 4547 2053
rect 4473 1967 4487 1973
rect 4616 1963 4623 2013
rect 4636 1967 4643 2223
rect 4676 2127 4683 2233
rect 4836 2226 4843 2253
rect 4976 2220 4983 2223
rect 4656 1987 4663 2033
rect 4596 1956 4623 1963
rect 4696 1967 4703 2212
rect 4973 2207 4987 2220
rect 5036 2207 5043 2293
rect 5056 2287 5063 2432
rect 5096 2407 5103 2443
rect 5276 2347 5283 2474
rect 5073 2260 5087 2273
rect 5076 2256 5083 2260
rect 5116 2256 5123 2313
rect 5236 2256 5243 2293
rect 5296 2263 5303 2913
rect 5336 2907 5343 2963
rect 5316 2787 5323 2873
rect 5356 2776 5363 2833
rect 5376 2827 5383 3253
rect 5436 3147 5443 3263
rect 5476 3260 5483 3263
rect 5473 3247 5487 3260
rect 5516 3083 5523 3253
rect 5536 3207 5543 3313
rect 5576 3303 5583 3573
rect 5596 3527 5603 3653
rect 5616 3527 5623 3613
rect 5636 3523 5643 3783
rect 5676 3727 5683 3813
rect 5696 3567 5703 3953
rect 5736 3783 5743 4276
rect 5756 3967 5763 4053
rect 5716 3776 5743 3783
rect 5716 3547 5723 3776
rect 5636 3516 5653 3523
rect 5616 3327 5623 3453
rect 5636 3427 5643 3483
rect 5676 3476 5703 3483
rect 5556 3296 5583 3303
rect 5616 3296 5623 3313
rect 5507 3076 5523 3083
rect 5416 2960 5423 2963
rect 5413 2947 5427 2960
rect 5496 2803 5503 3073
rect 5556 3067 5563 3296
rect 5596 3260 5603 3263
rect 5593 3247 5607 3260
rect 5516 2927 5523 3053
rect 5676 3027 5683 3453
rect 5696 3407 5703 3476
rect 5716 3467 5723 3512
rect 5533 3007 5547 3013
rect 5696 3007 5703 3293
rect 5476 2796 5503 2803
rect 5400 2783 5413 2787
rect 5396 2776 5413 2783
rect 5400 2773 5413 2776
rect 5476 2776 5483 2796
rect 5516 2787 5523 2813
rect 5400 2768 5407 2773
rect 5336 2740 5343 2743
rect 5333 2727 5347 2740
rect 5376 2707 5383 2743
rect 5436 2727 5443 2774
rect 5367 2436 5383 2443
rect 5276 2256 5303 2263
rect 5156 2227 5163 2254
rect 4816 1956 4823 2113
rect 4716 1926 4723 1953
rect 4456 1687 4463 1873
rect 4496 1767 4503 1793
rect 4656 1787 4663 1912
rect 4496 1736 4503 1753
rect 4536 1736 4543 1773
rect 4716 1747 4723 1912
rect 4736 1747 4743 1913
rect 4773 1740 4787 1753
rect 4796 1747 4803 1923
rect 4776 1736 4783 1740
rect 4516 1683 4523 1703
rect 4516 1676 4543 1683
rect 4076 1436 4083 1493
rect 4153 1440 4167 1453
rect 4156 1436 4163 1440
rect 4056 1367 4063 1392
rect 3976 1107 3983 1183
rect 3956 1096 3973 1103
rect 3736 767 3743 883
rect 3816 807 3823 873
rect 3876 787 3883 883
rect 3576 667 3583 694
rect 3647 663 3660 667
rect 3647 656 3663 663
rect 3647 653 3660 656
rect 3593 627 3607 633
rect 3653 607 3667 613
rect 3516 408 3523 553
rect 3553 400 3567 413
rect 3556 396 3563 400
rect 3376 366 3383 393
rect 3436 287 3443 363
rect 3476 356 3503 363
rect 3476 327 3483 356
rect 3496 307 3503 333
rect 3536 307 3543 363
rect 3240 183 3253 187
rect 3236 176 3253 183
rect 3240 173 3253 176
rect 3276 67 3283 213
rect 3296 187 3303 273
rect 3316 140 3323 143
rect 2396 -24 2403 13
rect 2496 -24 2503 13
rect 3296 -24 3303 133
rect 3313 127 3327 140
rect 3336 -24 3343 133
rect 3356 87 3363 143
rect 3396 107 3403 233
rect 3456 176 3463 213
rect 3476 207 3483 253
rect 3496 176 3503 293
rect 3576 267 3583 353
rect 3596 327 3603 413
rect 3616 347 3623 553
rect 3676 403 3683 653
rect 3696 547 3703 653
rect 3667 396 3683 403
rect 3696 396 3703 433
rect 3716 407 3723 713
rect 3776 696 3783 753
rect 3816 667 3823 753
rect 3836 707 3843 773
rect 3956 727 3963 1096
rect 4036 1007 4043 1333
rect 4096 1287 4103 1403
rect 4196 1229 4203 1273
rect 4236 1216 4243 1393
rect 4256 1347 4263 1513
rect 4456 1436 4463 1493
rect 4336 1400 4343 1403
rect 4333 1387 4347 1400
rect 4376 1247 4383 1373
rect 4376 1216 4383 1233
rect 4396 1227 4403 1393
rect 4407 1216 4423 1223
rect 4116 1147 4123 1183
rect 4176 1176 4203 1183
rect 3973 927 3987 933
rect 4013 920 4027 933
rect 4016 916 4023 920
rect 4056 916 4063 953
rect 3976 696 3983 853
rect 4036 707 4043 883
rect 4096 747 4103 993
rect 4156 916 4163 1173
rect 4196 927 4203 1176
rect 4216 887 4223 933
rect 4276 916 4283 1033
rect 4316 916 4323 953
rect 4396 943 4403 1173
rect 4476 987 4483 1393
rect 4467 966 4480 967
rect 4467 953 4473 966
rect 4396 936 4423 943
rect 4416 916 4423 936
rect 4136 767 4143 883
rect 4176 876 4203 883
rect 3756 607 3763 653
rect 3896 607 3903 663
rect 3836 467 3843 593
rect 3936 567 3943 693
rect 3727 396 3743 403
rect 3676 327 3683 363
rect 3716 267 3723 353
rect 3836 307 3843 394
rect 3856 366 3863 433
rect 3467 96 3493 103
rect 3516 83 3523 133
rect 3596 107 3603 213
rect 3756 146 3763 253
rect 3956 247 3963 473
rect 3996 396 4003 473
rect 4036 396 4043 433
rect 4056 407 4063 733
rect 4076 627 4083 653
rect 4096 603 4103 633
rect 4076 596 4103 603
rect 4076 367 4083 596
rect 4136 427 4143 663
rect 4156 567 4163 613
rect 4176 587 4183 853
rect 4196 847 4203 876
rect 4236 867 4243 913
rect 4196 707 4203 733
rect 4193 647 4207 653
rect 4206 640 4207 647
rect 4196 563 4203 593
rect 4176 556 4203 563
rect 4176 543 4183 556
rect 4156 540 4183 543
rect 4153 536 4183 540
rect 4153 527 4167 536
rect 4096 347 4103 393
rect 4173 400 4187 413
rect 4196 407 4203 473
rect 4176 396 4183 400
rect 3873 187 3887 193
rect 3996 188 4003 233
rect 3776 147 3783 173
rect 3447 76 3523 83
rect 3656 67 3663 143
rect 3896 87 3903 174
rect 3927 143 3940 147
rect 3927 136 3943 143
rect 3927 133 3940 136
rect 4036 140 4043 143
rect 4033 127 4047 140
rect 4096 87 4103 143
rect 4116 -24 4123 353
rect 4156 287 4163 363
rect 4196 263 4203 353
rect 4216 267 4223 633
rect 4236 407 4243 513
rect 4256 487 4263 663
rect 4296 527 4303 883
rect 4336 847 4343 883
rect 4396 767 4403 883
rect 4336 707 4343 733
rect 4316 647 4323 694
rect 4416 696 4423 833
rect 4476 807 4483 873
rect 4496 867 4503 1673
rect 4516 1407 4523 1653
rect 4536 1447 4543 1676
rect 4596 1436 4603 1693
rect 4616 1647 4623 1703
rect 4716 1467 4723 1712
rect 4816 1707 4823 1893
rect 4856 1887 4863 1993
rect 4936 1956 4943 2013
rect 4976 1967 4983 2193
rect 5016 1987 5023 2033
rect 5013 1960 5027 1973
rect 5016 1956 5023 1960
rect 5056 1956 5063 2133
rect 5136 1926 5143 2133
rect 5216 2107 5223 2223
rect 5276 2187 5283 2256
rect 5376 2263 5383 2436
rect 5356 2256 5383 2263
rect 5296 2007 5303 2053
rect 5193 1960 5207 1973
rect 5273 1960 5287 1973
rect 5316 1967 5323 2093
rect 5336 1967 5343 2223
rect 5196 1956 5203 1960
rect 5276 1956 5283 1960
rect 4916 1807 4923 1923
rect 5036 1920 5043 1923
rect 5033 1907 5047 1920
rect 5013 1740 5027 1753
rect 5036 1747 5043 1853
rect 5076 1847 5083 1923
rect 5216 1920 5223 1923
rect 5213 1907 5227 1920
rect 5016 1736 5023 1740
rect 4736 1447 4743 1633
rect 4796 1503 4803 1693
rect 4876 1647 4883 1703
rect 4996 1696 5033 1703
rect 4916 1547 4923 1693
rect 4976 1647 4983 1693
rect 5056 1667 5063 1734
rect 5176 1707 5183 1793
rect 5196 1687 5203 1833
rect 5296 1736 5303 1923
rect 5336 1743 5343 1913
rect 5356 1767 5363 2013
rect 5376 1967 5383 2113
rect 5396 1987 5403 2473
rect 5416 2427 5423 2533
rect 5436 2487 5443 2513
rect 5456 2476 5463 2733
rect 5496 2476 5503 2553
rect 5516 2487 5523 2733
rect 5536 2647 5543 2833
rect 5596 2807 5603 2923
rect 5616 2707 5623 2743
rect 5556 2476 5563 2513
rect 5596 2487 5603 2593
rect 5436 2263 5443 2433
rect 5476 2347 5483 2443
rect 5576 2440 5583 2443
rect 5573 2427 5587 2440
rect 5416 2256 5443 2263
rect 5416 2027 5423 2256
rect 5436 2127 5443 2213
rect 5456 2147 5463 2223
rect 5436 2067 5443 2113
rect 5416 1956 5423 2013
rect 5376 1887 5383 1913
rect 5416 1747 5423 1893
rect 5436 1867 5443 1923
rect 5476 1827 5483 1913
rect 5496 1763 5503 2213
rect 5516 1787 5523 2293
rect 5536 2268 5543 2313
rect 5576 2256 5583 2293
rect 5636 2267 5643 2733
rect 5656 2287 5663 2773
rect 5676 2707 5683 2733
rect 5676 2256 5683 2313
rect 5696 2287 5703 2513
rect 5716 2487 5723 3432
rect 5736 2787 5743 3553
rect 5756 2503 5763 3893
rect 5736 2496 5763 2503
rect 5556 1956 5563 2173
rect 5596 2007 5603 2223
rect 5616 1983 5623 2213
rect 5656 2127 5663 2223
rect 5596 1976 5623 1983
rect 5596 1956 5603 1976
rect 5496 1760 5523 1763
rect 5496 1756 5527 1760
rect 5513 1747 5527 1756
rect 5336 1736 5363 1743
rect 5236 1700 5243 1703
rect 5233 1687 5247 1700
rect 5067 1656 5083 1663
rect 4776 1496 4803 1503
rect 4776 1443 4783 1496
rect 4916 1447 4923 1533
rect 4776 1436 4803 1443
rect 4533 1387 4547 1393
rect 4576 1307 4583 1403
rect 4616 1400 4623 1403
rect 4613 1387 4627 1400
rect 4516 1227 4523 1293
rect 4596 1176 4623 1183
rect 4616 1107 4623 1176
rect 4636 1147 4643 1393
rect 4656 1367 4663 1433
rect 4936 1406 4943 1553
rect 5016 1507 5023 1593
rect 5016 1436 5023 1493
rect 4656 1107 4663 1273
rect 4673 1227 4687 1233
rect 4716 1216 4723 1273
rect 4856 1247 4863 1363
rect 4876 1216 4883 1253
rect 4936 1223 4943 1392
rect 4916 1216 4943 1223
rect 4976 1216 4983 1253
rect 5016 1216 5023 1253
rect 5056 1227 5063 1553
rect 5076 1267 5083 1656
rect 5276 1567 5283 1692
rect 5116 1436 5123 1533
rect 5196 1367 5203 1403
rect 5096 1227 5103 1313
rect 4773 1207 4787 1213
rect 4736 1147 4743 1183
rect 4616 1067 4623 1093
rect 4736 1047 4743 1133
rect 4516 927 4523 973
rect 4547 953 4553 967
rect 4516 747 4523 873
rect 4536 807 4543 883
rect 4556 823 4563 853
rect 4576 847 4583 873
rect 4556 816 4583 823
rect 4576 787 4583 816
rect 4336 527 4343 653
rect 4356 607 4363 663
rect 4456 447 4463 733
rect 4556 696 4563 753
rect 4576 707 4583 773
rect 4596 727 4603 1033
rect 4616 927 4623 953
rect 4656 916 4663 973
rect 4616 703 4623 873
rect 4636 787 4643 883
rect 4707 883 4720 887
rect 4707 876 4723 883
rect 4707 873 4720 876
rect 4596 696 4623 703
rect 4656 696 4663 733
rect 4693 700 4707 713
rect 4696 696 4703 700
rect 4776 696 4783 1172
rect 4796 928 4803 1173
rect 4856 1147 4863 1183
rect 4916 1183 4923 1216
rect 5116 1216 5123 1253
rect 4916 1176 4943 1183
rect 4956 1180 4963 1183
rect 4896 1027 4903 1173
rect 4913 1147 4927 1153
rect 4916 923 4923 1053
rect 4896 916 4923 923
rect 4816 847 4823 873
rect 4936 867 4943 1176
rect 4953 1167 4967 1180
rect 5136 1147 5143 1183
rect 5176 1167 5183 1253
rect 5276 1247 5283 1493
rect 5296 1327 5303 1613
rect 5316 1507 5323 1693
rect 5376 1667 5383 1703
rect 5396 1367 5403 1693
rect 5496 1700 5503 1703
rect 5476 1667 5483 1693
rect 5493 1687 5507 1700
rect 5416 1447 5423 1653
rect 5516 1627 5523 1693
rect 5536 1607 5543 1912
rect 5576 1823 5583 1923
rect 5556 1816 5583 1823
rect 5556 1687 5563 1816
rect 5436 1436 5443 1493
rect 5476 1436 5483 1533
rect 5213 1227 5227 1233
rect 4960 1146 4980 1147
rect 4967 1133 4973 1146
rect 5156 1107 5163 1153
rect 5196 1127 5203 1214
rect 5296 1216 5303 1253
rect 5236 1180 5243 1183
rect 5013 920 5027 933
rect 5016 916 5023 920
rect 4976 880 4983 883
rect 4973 867 4987 880
rect 5056 867 5063 933
rect 5116 916 5123 1013
rect 5196 887 5203 914
rect 5096 880 5103 883
rect 5093 867 5107 880
rect 4916 696 4963 703
rect 4476 656 4503 663
rect 4476 627 4483 656
rect 4536 567 4543 663
rect 4576 443 4583 653
rect 4596 567 4603 696
rect 5016 667 5023 853
rect 5136 807 5143 883
rect 5056 707 5063 793
rect 5073 723 5087 733
rect 5216 728 5223 1173
rect 5233 1167 5247 1180
rect 5276 1163 5283 1183
rect 5276 1156 5303 1163
rect 5256 947 5263 1153
rect 5276 1067 5283 1133
rect 5296 1087 5303 1156
rect 5336 1147 5343 1183
rect 5396 1127 5403 1183
rect 5436 1167 5443 1313
rect 5516 1307 5523 1533
rect 5656 1467 5663 1773
rect 5676 1748 5683 2193
rect 5736 2023 5743 2496
rect 5716 2016 5743 2023
rect 5676 1507 5683 1734
rect 5716 1547 5723 2016
rect 5553 1440 5567 1453
rect 5556 1436 5563 1440
rect 5576 1223 5583 1403
rect 5596 1228 5603 1293
rect 5556 1216 5583 1223
rect 5276 987 5283 1053
rect 5456 1007 5463 1193
rect 5253 920 5267 933
rect 5300 923 5313 927
rect 5256 916 5263 920
rect 5296 916 5313 923
rect 5300 914 5313 916
rect 5413 920 5427 933
rect 5456 927 5463 993
rect 5416 916 5423 920
rect 5300 913 5320 914
rect 5267 856 5293 863
rect 5073 720 5103 723
rect 5076 716 5107 720
rect 5093 707 5107 716
rect 4636 527 4643 663
rect 4676 587 4683 663
rect 4556 436 4583 443
rect 4253 427 4267 433
rect 4276 420 4323 423
rect 4276 416 4327 420
rect 4276 396 4283 416
rect 4313 407 4327 416
rect 4396 396 4403 433
rect 4456 420 4513 423
rect 4453 416 4513 420
rect 4453 407 4467 416
rect 4536 407 4543 433
rect 4256 360 4263 363
rect 4236 327 4243 353
rect 4253 347 4267 360
rect 4156 256 4203 263
rect 4156 -24 4163 256
rect 4256 -24 4263 312
rect 4296 176 4303 313
rect 4356 267 4363 363
rect 4456 327 4463 353
rect 4476 146 4483 363
rect 4556 176 4563 436
rect 4573 407 4587 413
rect 4616 396 4623 453
rect 4656 403 4663 453
rect 4676 427 4683 573
rect 4756 567 4763 663
rect 4896 587 4903 663
rect 5080 663 5093 667
rect 5076 656 5093 663
rect 5080 653 5093 656
rect 5136 660 5143 663
rect 5016 507 5023 653
rect 5056 587 5063 653
rect 5133 647 5147 660
rect 4656 396 4683 403
rect 4596 147 4603 363
rect 4636 327 4643 363
rect 4676 267 4683 396
rect 4796 396 4803 453
rect 5076 447 5083 633
rect 5176 607 5183 713
rect 5256 696 5263 813
rect 5356 767 5363 883
rect 5396 880 5403 883
rect 5393 867 5407 880
rect 5336 756 5353 763
rect 5196 547 5203 653
rect 5236 643 5243 663
rect 5216 636 5243 643
rect 5116 408 5123 533
rect 4696 327 4703 393
rect 4736 188 4743 363
rect 4756 176 4763 213
rect 4796 176 4803 213
rect 4876 176 4883 253
rect 4916 187 4923 393
rect 4996 287 5003 363
rect 5056 243 5063 393
rect 5096 287 5103 352
rect 5056 236 5083 243
rect 5007 213 5013 227
rect 5013 180 5027 192
rect 5016 176 5023 180
rect 4936 147 4943 174
rect 5056 147 5063 213
rect 5076 207 5083 236
rect 5116 227 5123 333
rect 5156 227 5163 493
rect 5216 408 5223 636
rect 5276 607 5283 663
rect 5316 507 5323 713
rect 5336 707 5343 756
rect 5376 696 5383 813
rect 5436 703 5443 873
rect 5536 827 5543 933
rect 5556 928 5563 1216
rect 5616 1087 5623 1183
rect 5656 928 5663 953
rect 5436 696 5463 703
rect 5396 567 5403 663
rect 5676 663 5683 873
rect 5636 656 5683 663
rect 5436 587 5443 652
rect 5276 396 5283 433
rect 5176 223 5183 393
rect 5236 360 5243 363
rect 5233 347 5247 360
rect 5376 267 5383 394
rect 5396 347 5403 493
rect 5496 408 5503 553
rect 5656 396 5663 633
rect 5676 447 5683 656
rect 5696 647 5703 1392
rect 5716 847 5723 1434
rect 5736 1007 5743 1993
rect 5756 1927 5763 2473
rect 5496 363 5503 394
rect 5476 356 5503 363
rect 5176 216 5203 223
rect 5087 196 5183 203
rect 5176 176 5183 196
rect 5196 187 5203 216
rect 5436 176 5443 213
rect 5456 187 5463 253
rect 4336 -24 4343 143
rect 4956 107 4963 133
rect 5076 67 5083 172
rect 5116 107 5123 143
rect 5236 67 5243 143
rect 5296 107 5303 143
rect 5336 127 5343 175
rect 5476 147 5483 356
rect 5636 287 5643 363
rect 5676 327 5683 363
rect 5527 216 5563 223
rect 5556 203 5563 216
rect 5556 196 5583 203
rect 5533 180 5547 193
rect 5536 176 5543 180
rect 5576 176 5583 196
rect 5420 143 5433 147
rect 5376 67 5383 143
rect 5416 136 5433 143
rect 5420 133 5433 136
rect 5556 140 5563 143
rect 5493 127 5507 133
rect 5553 127 5567 140
rect 5596 107 5603 143
rect 5407 96 5433 103
<< m3contact >>
rect 313 5473 327 5487
rect 593 5473 607 5487
rect 1553 5473 1567 5487
rect 2033 5473 2047 5487
rect 2893 5473 2907 5487
rect 2933 5473 2947 5487
rect 213 5413 227 5427
rect 33 5373 47 5387
rect 73 5375 87 5389
rect 113 5375 127 5389
rect 213 5375 227 5389
rect 253 5375 267 5389
rect 293 5375 307 5389
rect 93 5313 107 5327
rect 113 5333 127 5347
rect 133 5333 147 5347
rect 233 5333 247 5347
rect 193 5313 207 5327
rect 273 5333 287 5347
rect 193 5213 207 5227
rect 333 5453 347 5467
rect 333 5413 347 5427
rect 393 5413 407 5427
rect 573 5413 587 5427
rect 493 5375 507 5389
rect 553 5373 567 5387
rect 313 5333 327 5347
rect 373 5333 387 5347
rect 413 5333 427 5347
rect 473 5333 487 5347
rect 413 5253 427 5267
rect 293 5153 307 5167
rect 113 5113 127 5127
rect 213 5113 227 5127
rect 313 5113 327 5127
rect 73 5074 87 5088
rect 253 5074 267 5088
rect 293 5073 307 5087
rect 33 5013 47 5027
rect 13 4933 27 4947
rect 73 4933 87 4947
rect 33 4873 47 4887
rect 133 5013 147 5027
rect 193 5013 207 5027
rect 273 5033 287 5047
rect 273 4993 287 5007
rect 233 4953 247 4967
rect 113 4933 127 4947
rect 213 4933 227 4947
rect 93 4873 107 4887
rect 253 4855 267 4869
rect 33 4813 47 4827
rect 93 4813 107 4827
rect 193 4813 207 4827
rect 213 4793 227 4807
rect 133 4713 147 4727
rect 33 4613 47 4627
rect 193 4613 207 4627
rect 73 4554 87 4568
rect 133 4553 147 4567
rect 273 4813 287 4827
rect 233 4713 247 4727
rect 253 4693 267 4707
rect 233 4653 247 4667
rect 213 4553 227 4567
rect 253 4613 267 4627
rect 353 5074 367 5088
rect 313 5033 327 5047
rect 373 4993 387 5007
rect 333 4953 347 4967
rect 313 4893 327 4907
rect 353 4933 367 4947
rect 333 4853 347 4867
rect 393 4893 407 4907
rect 373 4873 387 4887
rect 553 5333 567 5347
rect 513 5293 527 5307
rect 613 5453 627 5467
rect 753 5453 767 5467
rect 893 5453 907 5467
rect 1473 5453 1487 5467
rect 593 5373 607 5387
rect 653 5393 667 5407
rect 813 5393 827 5407
rect 753 5375 767 5389
rect 633 5333 647 5347
rect 573 5313 587 5327
rect 753 5313 767 5327
rect 553 5253 567 5267
rect 733 5253 747 5267
rect 553 5213 567 5227
rect 473 5173 487 5187
rect 533 5153 547 5167
rect 473 5113 487 5127
rect 513 5073 527 5087
rect 653 5113 667 5127
rect 613 5073 627 5087
rect 693 5093 707 5107
rect 733 5074 747 5088
rect 793 5313 807 5327
rect 773 5293 787 5307
rect 853 5374 867 5388
rect 1153 5413 1167 5427
rect 1233 5413 1247 5427
rect 1393 5413 1407 5427
rect 973 5373 987 5387
rect 1053 5374 1067 5388
rect 1233 5375 1247 5389
rect 1293 5375 1307 5389
rect 1333 5375 1347 5389
rect 813 5293 827 5307
rect 793 5253 807 5267
rect 1013 5332 1027 5346
rect 1113 5313 1127 5327
rect 1113 5253 1127 5267
rect 1233 5313 1247 5327
rect 1273 5253 1287 5267
rect 973 5213 987 5227
rect 1053 5213 1067 5227
rect 1133 5213 1147 5227
rect 1173 5213 1187 5227
rect 453 5031 467 5045
rect 553 5033 567 5047
rect 493 4973 507 4987
rect 693 5033 707 5047
rect 633 4973 647 4987
rect 813 5073 827 5087
rect 973 5173 987 5187
rect 1053 5153 1067 5167
rect 973 5113 987 5127
rect 912 5093 926 5107
rect 933 5093 947 5107
rect 1013 5073 1027 5087
rect 713 5013 727 5027
rect 773 5013 787 5027
rect 693 4953 707 4967
rect 593 4913 607 4927
rect 473 4893 487 4907
rect 533 4893 547 4907
rect 413 4873 427 4887
rect 453 4873 467 4887
rect 353 4813 367 4827
rect 313 4773 327 4787
rect 293 4753 307 4767
rect 273 4593 287 4607
rect 373 4753 387 4767
rect 493 4855 507 4869
rect 533 4855 547 4869
rect 633 4855 647 4869
rect 493 4813 507 4827
rect 473 4773 487 4787
rect 593 4812 607 4826
rect 553 4793 567 4807
rect 513 4773 527 4787
rect 493 4753 507 4767
rect 613 4773 627 4787
rect 653 4772 667 4786
rect 393 4653 407 4667
rect 453 4653 467 4667
rect 593 4653 607 4667
rect 353 4573 367 4587
rect 333 4554 347 4568
rect 33 4512 47 4526
rect 93 4512 107 4526
rect 133 4453 147 4467
rect 93 4373 107 4387
rect 213 4511 227 4525
rect 253 4511 267 4525
rect 313 4512 327 4526
rect 373 4513 387 4527
rect 313 4433 327 4447
rect 233 4373 247 4387
rect 293 4373 307 4387
rect 93 4334 107 4348
rect 133 4333 147 4347
rect 193 4334 207 4348
rect 453 4613 467 4627
rect 573 4613 587 4627
rect 493 4553 507 4567
rect 533 4553 547 4567
rect 613 4593 627 4607
rect 413 4513 427 4527
rect 393 4453 407 4467
rect 373 4353 387 4367
rect 333 4334 347 4348
rect 73 4253 87 4267
rect 13 4113 27 4127
rect 213 4292 227 4306
rect 313 4292 327 4306
rect 373 4293 387 4307
rect 353 4273 367 4287
rect 173 4253 187 4267
rect 353 4233 367 4247
rect 173 4133 187 4147
rect 133 4053 147 4067
rect 193 4053 207 4067
rect 133 4032 147 4046
rect 373 4053 387 4067
rect 233 4033 247 4047
rect 293 4033 307 4047
rect 353 4033 367 4047
rect 553 4511 567 4525
rect 593 4511 607 4525
rect 633 4511 647 4525
rect 453 4493 467 4507
rect 493 4493 507 4507
rect 433 4373 447 4387
rect 533 4433 547 4447
rect 513 4373 527 4387
rect 413 4333 427 4347
rect 453 4335 467 4349
rect 493 4335 507 4349
rect 413 4233 427 4247
rect 393 4033 407 4047
rect 473 4273 487 4287
rect 433 4213 447 4227
rect 513 4213 527 4227
rect 473 4133 487 4147
rect 513 4073 527 4087
rect 913 5033 927 5047
rect 1033 5033 1047 5047
rect 993 5013 1007 5027
rect 833 4973 847 4987
rect 1033 4973 1047 4987
rect 793 4953 807 4967
rect 1093 5073 1107 5087
rect 1193 5193 1207 5207
rect 1173 5133 1187 5147
rect 1073 5033 1087 5047
rect 1053 4953 1067 4967
rect 833 4933 847 4947
rect 933 4933 947 4947
rect 793 4893 807 4907
rect 733 4853 747 4867
rect 793 4854 807 4868
rect 833 4854 847 4868
rect 873 4853 887 4867
rect 1053 4893 1067 4907
rect 973 4854 987 4868
rect 1113 4993 1127 5007
rect 1153 4953 1167 4967
rect 1113 4853 1127 4867
rect 1273 5173 1287 5187
rect 1333 5333 1347 5347
rect 1333 5253 1347 5267
rect 1353 5133 1367 5147
rect 1233 5113 1247 5127
rect 1313 5113 1327 5127
rect 1193 5093 1207 5107
rect 1753 5433 1767 5447
rect 2013 5433 2027 5447
rect 1553 5413 1567 5427
rect 1473 5374 1487 5388
rect 1593 5375 1607 5389
rect 1652 5375 1666 5389
rect 1433 5313 1447 5327
rect 1413 5233 1427 5247
rect 1333 5093 1347 5107
rect 1393 5093 1407 5107
rect 1273 5074 1287 5088
rect 1313 5073 1327 5087
rect 1253 5032 1267 5046
rect 1313 4993 1327 5007
rect 1213 4893 1227 4907
rect 1373 5074 1387 5088
rect 1513 5193 1527 5207
rect 1592 5333 1606 5347
rect 1613 5333 1627 5347
rect 1573 5233 1587 5247
rect 1533 5133 1547 5147
rect 1513 5074 1527 5088
rect 1673 5373 1687 5387
rect 1713 5375 1727 5389
rect 1853 5413 1867 5427
rect 2393 5453 2407 5467
rect 2853 5453 2867 5467
rect 2633 5433 2647 5447
rect 2033 5393 2047 5407
rect 2073 5393 2087 5407
rect 2313 5393 2327 5407
rect 2393 5393 2407 5407
rect 1853 5375 1867 5389
rect 1973 5375 1987 5389
rect 2013 5375 2027 5389
rect 1653 5273 1667 5287
rect 1913 5353 1927 5367
rect 1733 5333 1747 5347
rect 1773 5273 1787 5287
rect 1873 5333 1887 5347
rect 1873 5312 1887 5326
rect 1833 5233 1847 5247
rect 1673 5093 1687 5107
rect 1813 5093 1827 5107
rect 1233 4873 1247 4887
rect 1333 4873 1347 4887
rect 1173 4853 1187 4867
rect 773 4773 787 4787
rect 753 4753 767 4767
rect 813 4753 827 4767
rect 913 4812 927 4826
rect 973 4793 987 4807
rect 953 4773 967 4787
rect 993 4773 1007 4787
rect 973 4733 987 4747
rect 873 4713 887 4727
rect 933 4713 947 4727
rect 753 4693 767 4707
rect 733 4653 747 4667
rect 793 4673 807 4687
rect 753 4633 767 4647
rect 673 4593 687 4607
rect 712 4593 726 4607
rect 733 4593 747 4607
rect 672 4553 686 4567
rect 693 4552 707 4566
rect 733 4553 747 4567
rect 833 4633 847 4647
rect 873 4573 887 4587
rect 913 4573 927 4587
rect 853 4553 867 4567
rect 593 4373 607 4387
rect 653 4373 667 4387
rect 773 4513 787 4527
rect 813 4511 827 4525
rect 813 4473 827 4487
rect 773 4453 787 4467
rect 853 4453 867 4467
rect 713 4433 727 4447
rect 972 4554 986 4568
rect 1033 4713 1047 4727
rect 993 4553 1007 4567
rect 993 4513 1007 4527
rect 1033 4513 1047 4527
rect 973 4473 987 4487
rect 933 4393 947 4407
rect 673 4332 687 4346
rect 713 4333 727 4347
rect 753 4335 767 4349
rect 873 4335 887 4349
rect 913 4335 927 4349
rect 613 4293 627 4307
rect 573 4273 587 4287
rect 613 4113 627 4127
rect 553 4073 567 4087
rect 573 4052 587 4066
rect 613 4053 627 4067
rect 533 4033 547 4047
rect 113 3991 127 4005
rect 213 3991 227 4005
rect 213 3913 227 3927
rect 73 3893 87 3907
rect 133 3893 147 3907
rect 13 3853 27 3867
rect 93 3853 107 3867
rect 33 3833 47 3847
rect 173 3833 187 3847
rect 133 3813 147 3827
rect 333 3993 347 4007
rect 33 3773 47 3787
rect 73 3772 87 3786
rect 13 3733 27 3747
rect 13 3593 27 3607
rect 53 3553 67 3567
rect 33 3513 47 3527
rect 153 3773 167 3787
rect 193 3773 207 3787
rect 253 3773 267 3787
rect 213 3673 227 3687
rect 133 3533 147 3547
rect 393 3991 407 4005
rect 433 3993 447 4007
rect 353 3973 367 3987
rect 373 3893 387 3907
rect 333 3853 347 3867
rect 333 3814 347 3828
rect 413 3853 427 3867
rect 353 3772 367 3786
rect 373 3753 387 3767
rect 313 3733 327 3747
rect 273 3653 287 3667
rect 233 3533 247 3547
rect 213 3513 227 3527
rect 493 3973 507 3987
rect 453 3893 467 3907
rect 433 3813 447 3827
rect 553 3913 567 3927
rect 633 4033 647 4047
rect 713 4293 727 4307
rect 693 4133 707 4147
rect 733 4273 747 4287
rect 853 4293 867 4307
rect 793 4193 807 4207
rect 853 4133 867 4147
rect 713 4113 727 4127
rect 813 4113 827 4127
rect 733 4073 747 4087
rect 673 4033 687 4047
rect 713 4033 727 4047
rect 633 3973 647 3987
rect 953 4333 967 4347
rect 1033 4473 1047 4487
rect 993 4393 1007 4407
rect 953 4293 967 4307
rect 933 4273 947 4287
rect 893 4193 907 4207
rect 913 4113 927 4127
rect 873 4093 887 4107
rect 853 4033 867 4047
rect 993 4273 1007 4287
rect 1073 4813 1087 4827
rect 1073 4773 1087 4787
rect 1293 4855 1307 4869
rect 1113 4673 1127 4687
rect 1113 4593 1127 4607
rect 1073 4553 1087 4567
rect 1232 4813 1246 4827
rect 1253 4813 1267 4827
rect 1193 4613 1207 4627
rect 1273 4693 1287 4707
rect 1213 4573 1227 4587
rect 1253 4573 1267 4587
rect 1133 4553 1147 4567
rect 1233 4553 1247 4567
rect 1313 4653 1327 4667
rect 1313 4613 1327 4627
rect 1133 4511 1147 4525
rect 1113 4493 1127 4507
rect 1093 4413 1107 4427
rect 1053 4373 1067 4387
rect 1093 4335 1107 4349
rect 1273 4511 1287 4525
rect 1293 4473 1307 4487
rect 1233 4453 1247 4467
rect 1173 4413 1187 4427
rect 1153 4373 1167 4387
rect 1133 4333 1147 4347
rect 1093 4293 1107 4307
rect 1093 4233 1107 4247
rect 1073 4153 1087 4167
rect 1273 4373 1287 4387
rect 1233 4334 1247 4348
rect 1193 4293 1207 4307
rect 1173 4213 1187 4227
rect 1053 4133 1067 4147
rect 1112 4133 1126 4147
rect 1133 4133 1147 4147
rect 1033 4113 1047 4127
rect 993 4053 1007 4067
rect 953 4033 967 4047
rect 733 4013 747 4027
rect 713 3973 727 3987
rect 673 3953 687 3967
rect 773 3973 787 3987
rect 833 3992 847 4006
rect 893 3992 907 4006
rect 733 3913 747 3927
rect 573 3853 587 3867
rect 653 3853 667 3867
rect 493 3815 507 3829
rect 533 3815 547 3829
rect 593 3815 607 3829
rect 633 3815 647 3829
rect 813 3893 827 3907
rect 773 3833 787 3847
rect 673 3814 687 3828
rect 713 3814 727 3828
rect 753 3814 767 3828
rect 453 3773 467 3787
rect 413 3713 427 3727
rect 433 3653 447 3667
rect 53 3433 67 3447
rect 33 3353 47 3367
rect 113 3471 127 3485
rect 213 3471 227 3485
rect 253 3471 267 3485
rect 293 3473 307 3487
rect 133 3433 147 3447
rect 93 3333 107 3347
rect 33 3313 47 3327
rect 73 3313 87 3327
rect 13 3253 27 3267
rect 13 3093 27 3107
rect 13 3033 27 3047
rect 13 2993 27 3007
rect 293 3452 307 3466
rect 353 3453 367 3467
rect 253 3333 267 3347
rect 233 3294 247 3308
rect 373 3353 387 3367
rect 333 3294 347 3308
rect 173 3252 187 3266
rect 133 3053 147 3067
rect 73 3033 87 3047
rect 113 3033 127 3047
rect 313 3252 327 3266
rect 273 3213 287 3227
rect 313 3213 327 3227
rect 233 3153 247 3167
rect 273 3153 287 3167
rect 73 2994 87 3008
rect 173 3013 187 3027
rect 233 3013 247 3027
rect 153 2993 167 3007
rect 53 2953 67 2967
rect 33 2933 47 2947
rect 33 2793 47 2807
rect 153 2953 167 2967
rect 293 3133 307 3147
rect 293 3093 307 3107
rect 133 2933 147 2947
rect 93 2813 107 2827
rect 73 2793 87 2807
rect 113 2775 127 2789
rect 193 2893 207 2907
rect 253 2913 267 2927
rect 173 2813 187 2827
rect 213 2813 227 2827
rect 273 2813 287 2827
rect 153 2773 167 2787
rect 33 2733 47 2747
rect 92 2733 106 2747
rect 112 2733 126 2747
rect 133 2733 147 2747
rect 13 2633 27 2647
rect 193 2773 207 2787
rect 233 2793 247 2807
rect 213 2732 227 2746
rect 253 2733 267 2747
rect 193 2613 207 2627
rect 33 2553 47 2567
rect 173 2553 187 2567
rect 433 3473 447 3487
rect 473 3753 487 3767
rect 573 3753 587 3767
rect 513 3713 527 3727
rect 653 3773 667 3787
rect 613 3713 627 3727
rect 953 3973 967 3987
rect 893 3933 907 3947
rect 933 3933 947 3947
rect 933 3893 947 3907
rect 913 3873 927 3887
rect 873 3833 887 3847
rect 973 3953 987 3967
rect 993 3933 1007 3947
rect 1153 4113 1167 4127
rect 1133 4093 1147 4107
rect 1093 4073 1107 4087
rect 1073 4053 1087 4067
rect 1053 4033 1067 4047
rect 1113 4053 1127 4067
rect 1093 4033 1107 4047
rect 1033 3993 1047 4007
rect 1053 3913 1067 3927
rect 1113 3913 1127 3927
rect 973 3873 987 3887
rect 1033 3873 1047 3887
rect 973 3852 987 3866
rect 1013 3853 1027 3867
rect 1093 3893 1107 3907
rect 1093 3872 1107 3886
rect 1012 3832 1026 3846
rect 1053 3833 1067 3847
rect 973 3813 987 3827
rect 953 3793 967 3807
rect 733 3772 747 3786
rect 693 3753 707 3767
rect 673 3733 687 3747
rect 693 3713 707 3727
rect 813 3772 827 3786
rect 813 3713 827 3727
rect 653 3673 667 3687
rect 773 3673 787 3687
rect 793 3653 807 3667
rect 573 3633 587 3647
rect 773 3633 787 3647
rect 893 3773 907 3787
rect 853 3753 867 3767
rect 973 3773 987 3787
rect 1033 3773 1047 3787
rect 1073 3773 1087 3787
rect 953 3753 967 3767
rect 833 3673 847 3687
rect 933 3633 947 3647
rect 813 3613 827 3627
rect 793 3593 807 3607
rect 833 3593 847 3607
rect 513 3553 527 3567
rect 733 3553 747 3567
rect 773 3553 787 3567
rect 593 3513 607 3527
rect 653 3513 667 3527
rect 693 3513 707 3527
rect 493 3471 507 3485
rect 613 3453 627 3467
rect 593 3433 607 3447
rect 573 3413 587 3427
rect 473 3393 487 3407
rect 553 3393 567 3407
rect 453 3373 467 3387
rect 393 3333 407 3347
rect 533 3353 547 3367
rect 513 3333 527 3347
rect 413 3295 427 3309
rect 453 3295 467 3309
rect 373 3113 387 3127
rect 473 3213 487 3227
rect 413 3093 427 3107
rect 433 3093 447 3107
rect 373 3053 387 3067
rect 373 3012 387 3026
rect 453 3073 467 3087
rect 433 3053 447 3067
rect 553 3333 567 3347
rect 533 3293 547 3307
rect 573 3294 587 3308
rect 673 3471 687 3485
rect 673 3433 687 3447
rect 873 3553 887 3567
rect 913 3533 927 3547
rect 793 3513 807 3527
rect 833 3512 847 3526
rect 873 3513 887 3527
rect 953 3533 967 3547
rect 813 3471 827 3485
rect 853 3473 867 3487
rect 793 3433 807 3447
rect 733 3393 747 3407
rect 773 3393 787 3407
rect 693 3373 707 3387
rect 653 3333 667 3347
rect 653 3293 667 3307
rect 733 3333 747 3347
rect 532 3253 546 3267
rect 513 3173 527 3187
rect 553 3252 567 3266
rect 593 3252 607 3266
rect 613 3133 627 3147
rect 593 3073 607 3087
rect 533 3053 547 3067
rect 433 2993 447 3007
rect 473 3013 487 3027
rect 513 3013 527 3027
rect 893 3453 907 3467
rect 853 3433 867 3447
rect 1093 3733 1107 3747
rect 1072 3633 1086 3647
rect 1093 3633 1107 3647
rect 1093 3612 1107 3626
rect 1053 3593 1067 3607
rect 1013 3553 1027 3567
rect 973 3513 987 3527
rect 1093 3573 1107 3587
rect 1213 4233 1227 4247
rect 1253 4193 1267 4207
rect 1433 4933 1447 4947
rect 1593 5033 1607 5047
rect 1593 4993 1607 5007
rect 1673 5072 1687 5086
rect 1713 5073 1727 5087
rect 1773 5073 1787 5087
rect 1613 4953 1627 4967
rect 1573 4933 1587 4947
rect 1693 5031 1707 5045
rect 1793 4993 1807 5007
rect 1813 4953 1827 4967
rect 1573 4912 1587 4926
rect 1653 4913 1667 4927
rect 1533 4893 1547 4907
rect 1673 4893 1687 4907
rect 1753 4893 1767 4907
rect 1433 4855 1447 4869
rect 1473 4855 1487 4869
rect 1513 4855 1527 4869
rect 1613 4855 1627 4869
rect 1653 4853 1667 4867
rect 1393 4813 1407 4827
rect 1453 4813 1467 4827
rect 1553 4772 1567 4786
rect 1493 4753 1507 4767
rect 1713 4855 1727 4869
rect 1713 4813 1727 4827
rect 1673 4793 1687 4807
rect 1613 4773 1627 4787
rect 1593 4753 1607 4767
rect 1573 4733 1587 4747
rect 1553 4673 1567 4687
rect 1453 4653 1467 4667
rect 1513 4653 1527 4667
rect 1573 4653 1587 4667
rect 1413 4554 1427 4568
rect 1353 4413 1367 4427
rect 1313 4373 1327 4387
rect 1313 4335 1327 4349
rect 1433 4513 1447 4527
rect 1413 4493 1427 4507
rect 1393 4393 1407 4407
rect 1373 4353 1387 4367
rect 1553 4554 1567 4568
rect 1533 4512 1547 4526
rect 1573 4493 1587 4507
rect 1473 4473 1487 4487
rect 1453 4453 1467 4467
rect 1433 4413 1447 4427
rect 1593 4453 1607 4467
rect 1493 4433 1507 4447
rect 1473 4373 1487 4387
rect 1413 4334 1427 4348
rect 1533 4413 1547 4427
rect 1293 4293 1307 4307
rect 1273 4173 1287 4187
rect 1373 4293 1387 4307
rect 1353 4273 1367 4287
rect 1413 4253 1427 4267
rect 1373 4233 1387 4247
rect 1473 4233 1487 4247
rect 1333 4213 1347 4227
rect 1393 4213 1407 4227
rect 1333 4192 1347 4206
rect 1293 4113 1307 4127
rect 1253 4093 1267 4107
rect 1313 4053 1327 4067
rect 1353 4173 1367 4187
rect 1333 4033 1347 4047
rect 1213 3991 1227 4005
rect 1273 3993 1287 4007
rect 1193 3953 1207 3967
rect 1193 3913 1207 3927
rect 1153 3833 1167 3847
rect 1133 3813 1147 3827
rect 1273 3873 1287 3887
rect 1233 3853 1247 3867
rect 1233 3813 1247 3827
rect 1292 3833 1306 3847
rect 1313 3833 1327 3847
rect 1673 4713 1687 4727
rect 1673 4613 1687 4627
rect 1653 4593 1667 4607
rect 1772 4813 1786 4827
rect 1793 4813 1807 4827
rect 1733 4713 1747 4727
rect 1713 4693 1727 4707
rect 1713 4653 1727 4667
rect 1713 4593 1727 4607
rect 1853 5013 1867 5027
rect 1913 5293 1927 5307
rect 1993 5313 2007 5327
rect 2033 5273 2047 5287
rect 1953 5233 1967 5247
rect 1913 5093 1927 5107
rect 1933 5031 1947 5045
rect 1873 4993 1887 5007
rect 2093 5373 2107 5387
rect 2153 5374 2167 5388
rect 2233 5375 2247 5389
rect 2293 5375 2307 5389
rect 2093 5332 2107 5346
rect 2133 5332 2147 5346
rect 2193 5233 2207 5247
rect 2073 5193 2087 5207
rect 2133 5173 2147 5187
rect 2433 5375 2447 5389
rect 2493 5375 2507 5389
rect 2593 5374 2607 5388
rect 2693 5413 2707 5427
rect 2353 5332 2367 5346
rect 2433 5333 2447 5347
rect 2333 5313 2347 5327
rect 2333 5273 2347 5287
rect 2473 5293 2487 5307
rect 2453 5273 2467 5287
rect 2493 5253 2507 5267
rect 2313 5233 2327 5247
rect 2353 5233 2367 5247
rect 2473 5233 2487 5247
rect 2293 5213 2307 5227
rect 2253 5193 2267 5207
rect 2213 5173 2227 5187
rect 2193 5153 2207 5167
rect 2213 5133 2227 5147
rect 2453 5173 2467 5187
rect 2413 5133 2427 5147
rect 2233 5113 2247 5127
rect 2293 5113 2307 5127
rect 2133 5093 2147 5107
rect 2133 5072 2147 5086
rect 2393 5093 2407 5107
rect 2233 5073 2247 5087
rect 2273 5073 2287 5087
rect 2313 5073 2327 5087
rect 2053 5033 2067 5047
rect 2173 5033 2187 5047
rect 2113 5013 2127 5027
rect 2033 4953 2047 4967
rect 2193 4953 2207 4967
rect 1933 4913 1947 4927
rect 1973 4913 1987 4927
rect 1833 4893 1847 4907
rect 1893 4893 1907 4907
rect 1832 4853 1846 4867
rect 1853 4855 1867 4869
rect 2253 5031 2267 5045
rect 2313 5031 2327 5045
rect 2353 5031 2367 5045
rect 2433 5031 2447 5045
rect 2393 4993 2407 5007
rect 2253 4973 2267 4987
rect 2433 4973 2447 4987
rect 2573 5333 2587 5347
rect 2753 5375 2767 5389
rect 2653 5332 2667 5346
rect 2693 5332 2707 5346
rect 2753 5333 2767 5347
rect 2673 5273 2687 5287
rect 2733 5273 2747 5287
rect 2573 5213 2587 5227
rect 2613 5213 2627 5227
rect 2533 5133 2547 5147
rect 2493 5073 2507 5087
rect 2593 5073 2607 5087
rect 2733 5252 2747 5266
rect 2753 5233 2767 5247
rect 2793 5333 2807 5347
rect 2773 5213 2787 5227
rect 2733 5133 2747 5147
rect 2713 5093 2727 5107
rect 2673 5073 2687 5087
rect 2813 5253 2827 5267
rect 2932 5433 2946 5447
rect 3013 5413 3027 5427
rect 2893 5393 2907 5407
rect 2953 5393 2967 5407
rect 3013 5374 3027 5388
rect 3072 5473 3086 5487
rect 3093 5473 3107 5487
rect 3053 5373 3067 5387
rect 2873 5333 2887 5347
rect 2913 5332 2927 5346
rect 2993 5333 3007 5347
rect 2893 5293 2907 5307
rect 2853 5233 2867 5247
rect 2953 5313 2967 5327
rect 2933 5293 2947 5307
rect 2913 5273 2927 5287
rect 2933 5253 2947 5267
rect 2893 5193 2907 5207
rect 2853 5153 2867 5167
rect 2813 5133 2827 5147
rect 2813 5093 2827 5107
rect 2213 4933 2227 4947
rect 2313 4933 2327 4947
rect 2453 4933 2467 4947
rect 2113 4893 2127 4907
rect 2193 4893 2207 4907
rect 2013 4873 2027 4887
rect 2073 4873 2087 4887
rect 1932 4853 1946 4867
rect 1973 4854 1987 4868
rect 1913 4793 1927 4807
rect 1933 4813 1947 4827
rect 1953 4813 1967 4827
rect 1893 4773 1907 4787
rect 1873 4713 1887 4727
rect 2033 4812 2047 4826
rect 2113 4854 2127 4868
rect 2173 4855 2187 4869
rect 2233 4855 2247 4869
rect 2273 4855 2287 4869
rect 2133 4812 2147 4826
rect 2173 4793 2187 4807
rect 1893 4693 1907 4707
rect 1813 4673 1827 4687
rect 1853 4673 1867 4687
rect 1813 4633 1827 4647
rect 1873 4633 1887 4647
rect 1853 4613 1867 4627
rect 1793 4573 1807 4587
rect 1693 4554 1707 4568
rect 1813 4554 1827 4568
rect 1853 4553 1867 4567
rect 1613 4413 1627 4427
rect 1593 4393 1607 4407
rect 1713 4512 1727 4526
rect 1773 4493 1787 4507
rect 1733 4393 1747 4407
rect 1573 4334 1587 4348
rect 1633 4333 1647 4347
rect 1693 4335 1707 4349
rect 1913 4613 1927 4627
rect 1953 4753 1967 4767
rect 2073 4753 2087 4767
rect 1953 4732 1967 4746
rect 2253 4813 2267 4827
rect 2033 4713 2047 4727
rect 2213 4713 2227 4727
rect 1953 4593 1967 4607
rect 1932 4553 1946 4567
rect 1953 4553 1967 4567
rect 1993 4553 2007 4567
rect 2073 4653 2087 4667
rect 2493 4993 2507 5007
rect 2333 4913 2347 4927
rect 2473 4913 2487 4927
rect 2393 4893 2407 4907
rect 2513 4913 2527 4927
rect 2613 5031 2627 5045
rect 2653 5031 2667 5045
rect 2693 5033 2707 5047
rect 2693 4993 2707 5007
rect 2633 4973 2647 4987
rect 2593 4893 2607 4907
rect 2893 5073 2907 5087
rect 2833 4993 2847 5007
rect 2753 4953 2767 4967
rect 2813 4953 2827 4967
rect 2713 4893 2727 4907
rect 2673 4873 2687 4887
rect 2333 4812 2347 4826
rect 2373 4812 2387 4826
rect 2493 4853 2507 4867
rect 2533 4854 2547 4868
rect 2573 4854 2587 4868
rect 2633 4854 2647 4868
rect 2733 4873 2747 4887
rect 2372 4753 2386 4767
rect 2393 4753 2407 4767
rect 2253 4633 2267 4647
rect 2313 4633 2327 4647
rect 2093 4613 2107 4627
rect 2073 4553 2087 4567
rect 2133 4593 2147 4607
rect 2193 4573 2207 4587
rect 2132 4553 2146 4567
rect 2153 4553 2167 4567
rect 1933 4511 1947 4525
rect 1873 4493 1887 4507
rect 1973 4493 1987 4507
rect 2073 4513 2087 4527
rect 2113 4513 2127 4527
rect 1993 4473 2007 4487
rect 2053 4473 2067 4487
rect 1973 4453 1987 4467
rect 1933 4433 1947 4447
rect 1773 4373 1787 4387
rect 1853 4373 1867 4387
rect 1533 4173 1547 4187
rect 1393 4133 1407 4147
rect 1613 4133 1627 4147
rect 1593 4113 1607 4127
rect 1493 4093 1507 4107
rect 1393 4053 1407 4067
rect 1433 4033 1447 4047
rect 1453 3991 1467 4005
rect 1553 4034 1567 4048
rect 1473 3913 1487 3927
rect 1413 3873 1427 3887
rect 1393 3833 1407 3847
rect 1153 3773 1167 3787
rect 1133 3693 1147 3707
rect 1133 3553 1147 3567
rect 1213 3773 1227 3787
rect 1353 3813 1367 3827
rect 1433 3833 1447 3847
rect 1493 3833 1507 3847
rect 1473 3813 1487 3827
rect 1253 3732 1267 3746
rect 1233 3713 1247 3727
rect 1173 3673 1187 3687
rect 1173 3633 1187 3647
rect 1153 3533 1167 3547
rect 1193 3553 1207 3567
rect 1332 3773 1346 3787
rect 1353 3773 1367 3787
rect 1333 3713 1347 3727
rect 1333 3673 1347 3687
rect 1273 3653 1287 3667
rect 1293 3633 1307 3647
rect 1273 3613 1287 3627
rect 1393 3733 1407 3747
rect 1353 3613 1367 3627
rect 1293 3573 1307 3587
rect 1353 3553 1367 3567
rect 1273 3533 1287 3547
rect 1093 3492 1107 3506
rect 873 3413 887 3427
rect 953 3413 967 3427
rect 833 3353 847 3367
rect 793 3293 807 3307
rect 1033 3472 1047 3486
rect 1253 3513 1267 3527
rect 1293 3513 1307 3527
rect 1173 3471 1187 3485
rect 1213 3471 1227 3485
rect 1113 3453 1127 3467
rect 1173 3433 1187 3447
rect 1033 3373 1047 3387
rect 1072 3373 1086 3387
rect 1093 3373 1107 3387
rect 993 3353 1007 3367
rect 973 3333 987 3347
rect 873 3295 887 3309
rect 933 3295 947 3309
rect 1133 3333 1147 3347
rect 713 3252 727 3266
rect 773 3253 787 3267
rect 813 3252 827 3266
rect 653 3213 667 3227
rect 693 3213 707 3227
rect 713 3193 727 3207
rect 653 3133 667 3147
rect 633 3053 647 3067
rect 593 3033 607 3047
rect 1033 3293 1047 3307
rect 1073 3295 1087 3309
rect 1333 3433 1347 3447
rect 1273 3413 1287 3427
rect 1253 3373 1267 3387
rect 1213 3313 1227 3327
rect 1193 3295 1207 3309
rect 1453 3772 1467 3786
rect 1413 3693 1427 3707
rect 1413 3672 1427 3686
rect 1453 3593 1467 3607
rect 1533 3913 1547 3927
rect 1653 4293 1667 4307
rect 1673 4253 1687 4267
rect 1713 4252 1727 4266
rect 1653 4233 1667 4247
rect 1633 4053 1647 4067
rect 1673 4093 1687 4107
rect 1753 4173 1767 4187
rect 1673 4053 1687 4067
rect 1713 4053 1727 4067
rect 1653 4033 1667 4047
rect 1633 3993 1647 4007
rect 1633 3933 1647 3947
rect 1613 3913 1627 3927
rect 1593 3853 1607 3867
rect 1633 3853 1647 3867
rect 1553 3815 1567 3829
rect 1693 3991 1707 4005
rect 1733 3993 1747 4007
rect 1853 4335 1867 4349
rect 1913 4335 1927 4349
rect 1793 4293 1807 4307
rect 1833 4273 1847 4287
rect 1792 4233 1806 4247
rect 1813 4233 1827 4247
rect 1793 4173 1807 4187
rect 1853 4253 1867 4267
rect 1913 4293 1927 4307
rect 1852 4213 1866 4227
rect 1873 4213 1887 4227
rect 1833 4153 1847 4167
rect 1993 4335 2007 4349
rect 2052 4333 2066 4347
rect 2073 4333 2087 4347
rect 2213 4511 2227 4525
rect 2213 4473 2227 4487
rect 2173 4433 2187 4447
rect 2213 4433 2227 4447
rect 2153 4393 2167 4407
rect 2173 4373 2187 4387
rect 2193 4353 2207 4367
rect 2173 4333 2187 4347
rect 1973 4293 1987 4307
rect 1953 4193 1967 4207
rect 1833 4132 1847 4146
rect 1932 4133 1946 4147
rect 1953 4133 1967 4147
rect 1773 4113 1787 4127
rect 1793 4034 1807 4048
rect 1913 4093 1927 4107
rect 1853 4073 1867 4087
rect 2053 4292 2067 4306
rect 2093 4292 2107 4306
rect 2013 4273 2027 4287
rect 2073 4253 2087 4267
rect 2053 4213 2067 4227
rect 2033 4173 2047 4187
rect 2013 4093 2027 4107
rect 1973 4053 1987 4067
rect 1953 4033 1967 4047
rect 1732 3933 1746 3947
rect 1753 3933 1767 3947
rect 1793 3933 1807 3947
rect 1632 3813 1646 3827
rect 1653 3813 1667 3827
rect 1693 3815 1707 3829
rect 1753 3912 1767 3926
rect 1733 3813 1747 3827
rect 1773 3893 1787 3907
rect 1513 3772 1527 3786
rect 1553 3773 1567 3787
rect 1493 3733 1507 3747
rect 1513 3593 1527 3607
rect 1513 3572 1527 3586
rect 1473 3553 1487 3567
rect 1413 3513 1427 3527
rect 1453 3513 1467 3527
rect 1413 3473 1427 3487
rect 1393 3413 1407 3427
rect 1353 3393 1367 3407
rect 1333 3353 1347 3367
rect 1293 3313 1307 3327
rect 1373 3333 1387 3347
rect 1353 3313 1367 3327
rect 1453 3471 1467 3485
rect 1493 3473 1507 3487
rect 1493 3373 1507 3387
rect 1673 3773 1687 3787
rect 1733 3773 1747 3787
rect 1593 3753 1607 3767
rect 1573 3733 1587 3747
rect 1613 3733 1627 3747
rect 1593 3573 1607 3587
rect 1733 3673 1747 3687
rect 1753 3653 1767 3667
rect 1673 3593 1687 3607
rect 1592 3513 1606 3527
rect 1613 3513 1627 3527
rect 1653 3513 1667 3527
rect 1593 3453 1607 3467
rect 1273 3273 1287 3287
rect 873 3173 887 3187
rect 733 3133 747 3147
rect 713 3113 727 3127
rect 673 3093 687 3107
rect 733 3093 747 3107
rect 713 3053 727 3067
rect 573 2993 587 3007
rect 633 2994 647 3008
rect 673 2994 687 3008
rect 393 2951 407 2965
rect 453 2951 467 2965
rect 533 2951 547 2965
rect 573 2953 587 2967
rect 553 2933 567 2947
rect 492 2913 506 2927
rect 513 2913 527 2927
rect 433 2893 447 2907
rect 413 2873 427 2887
rect 313 2793 327 2807
rect 353 2793 367 2807
rect 333 2733 347 2747
rect 273 2513 287 2527
rect 93 2473 107 2487
rect 133 2473 147 2487
rect 193 2473 207 2487
rect 373 2713 387 2727
rect 433 2853 447 2867
rect 473 2774 487 2788
rect 533 2893 547 2907
rect 453 2732 467 2746
rect 413 2693 427 2707
rect 493 2693 507 2707
rect 413 2513 427 2527
rect 292 2473 306 2487
rect 313 2474 327 2488
rect 373 2474 387 2488
rect 53 2433 67 2447
rect 33 2353 47 2367
rect 113 2431 127 2445
rect 213 2431 227 2445
rect 73 2393 87 2407
rect 113 2353 127 2367
rect 213 2353 227 2367
rect 133 2293 147 2307
rect 93 2254 107 2268
rect 293 2433 307 2447
rect 253 2313 267 2327
rect 373 2413 387 2427
rect 293 2293 307 2307
rect 173 2255 187 2269
rect 213 2255 227 2269
rect 353 2255 367 2269
rect 433 2473 447 2487
rect 413 2353 427 2367
rect 613 2933 627 2947
rect 693 2953 707 2967
rect 873 3013 887 3027
rect 733 2994 747 3008
rect 773 2994 787 3008
rect 813 2994 827 3008
rect 1053 3253 1067 3267
rect 1153 3253 1167 3267
rect 953 3233 967 3247
rect 1013 3233 1027 3247
rect 1113 3233 1127 3247
rect 973 3193 987 3207
rect 993 3173 1007 3187
rect 973 3113 987 3127
rect 1013 3133 1027 3147
rect 993 3053 1007 3067
rect 953 3013 967 3027
rect 873 2992 887 3006
rect 733 2953 747 2967
rect 793 2952 807 2966
rect 713 2933 727 2947
rect 693 2873 707 2887
rect 653 2853 667 2867
rect 1013 2973 1027 2987
rect 893 2953 907 2967
rect 873 2933 887 2947
rect 933 2951 947 2965
rect 913 2933 927 2947
rect 853 2893 867 2907
rect 893 2893 907 2907
rect 853 2813 867 2827
rect 593 2775 607 2789
rect 633 2775 647 2789
rect 693 2773 707 2787
rect 733 2775 747 2789
rect 773 2775 787 2789
rect 1053 2893 1067 2907
rect 1033 2813 1047 2827
rect 913 2774 927 2788
rect 953 2774 967 2788
rect 993 2774 1007 2788
rect 633 2733 647 2747
rect 653 2733 667 2747
rect 613 2713 627 2727
rect 633 2693 647 2707
rect 553 2613 567 2627
rect 653 2513 667 2527
rect 613 2473 627 2487
rect 793 2693 807 2707
rect 753 2573 767 2587
rect 753 2513 767 2527
rect 793 2473 807 2487
rect 553 2413 567 2427
rect 513 2353 527 2367
rect 513 2313 527 2327
rect 433 2273 447 2287
rect 33 2213 47 2227
rect 73 2212 87 2226
rect 112 2213 126 2227
rect 133 2213 147 2227
rect 193 2213 207 2227
rect 273 2213 287 2227
rect 353 2213 367 2227
rect 333 2193 347 2207
rect 253 2073 267 2087
rect 353 2073 367 2087
rect 193 2053 207 2067
rect 73 2033 87 2047
rect 113 2033 127 2047
rect 33 2013 47 2027
rect 13 1993 27 2007
rect 13 1953 27 1967
rect 233 2013 247 2027
rect 113 1953 127 1967
rect 193 1953 207 1967
rect 373 1993 387 2007
rect 253 1953 267 1967
rect 313 1954 327 1968
rect 413 2253 427 2267
rect 473 2254 487 2268
rect 393 1953 407 1967
rect 33 1913 47 1927
rect 93 1911 107 1925
rect 253 1911 267 1925
rect 93 1873 107 1887
rect 173 1873 187 1887
rect 33 1734 47 1748
rect 53 1313 67 1327
rect 113 1734 127 1748
rect 393 1893 407 1907
rect 373 1813 387 1827
rect 233 1733 247 1747
rect 153 1692 167 1706
rect 333 1692 347 1706
rect 213 1653 227 1667
rect 153 1434 167 1448
rect 273 1653 287 1667
rect 313 1433 327 1447
rect 493 2212 507 2226
rect 453 2193 467 2207
rect 633 2431 647 2445
rect 693 2431 707 2445
rect 773 2431 787 2445
rect 872 2732 886 2746
rect 893 2733 907 2747
rect 893 2513 907 2527
rect 1033 2773 1047 2787
rect 1013 2732 1027 2746
rect 973 2693 987 2707
rect 973 2653 987 2667
rect 933 2633 947 2647
rect 953 2613 967 2627
rect 913 2493 927 2507
rect 893 2474 907 2488
rect 973 2573 987 2587
rect 1073 2833 1087 2847
rect 1093 2774 1107 2788
rect 1173 3013 1187 3027
rect 1213 3253 1227 3267
rect 1253 3253 1267 3267
rect 1313 3253 1327 3267
rect 1213 3073 1227 3087
rect 1253 3073 1267 3087
rect 1293 3213 1307 3227
rect 1273 3053 1287 3067
rect 1353 3193 1367 3207
rect 1373 3093 1387 3107
rect 1373 3053 1387 3067
rect 1293 3033 1307 3047
rect 1253 3013 1267 3027
rect 1313 2993 1327 3007
rect 1473 3312 1487 3326
rect 1533 3353 1547 3367
rect 1573 3353 1587 3367
rect 1553 3333 1567 3347
rect 1573 3293 1587 3307
rect 1613 3433 1627 3447
rect 1713 3573 1727 3587
rect 1933 3991 1947 4005
rect 1853 3933 1867 3947
rect 1973 3933 1987 3947
rect 1833 3893 1847 3907
rect 1813 3853 1827 3867
rect 1873 3853 1887 3867
rect 1933 3853 1947 3867
rect 1993 3853 2007 3867
rect 1833 3773 1847 3787
rect 1793 3673 1807 3687
rect 1793 3633 1807 3647
rect 1773 3533 1787 3547
rect 1893 3833 1907 3847
rect 1933 3815 1947 3829
rect 2053 4133 2067 4147
rect 2113 4233 2127 4247
rect 2173 4293 2187 4307
rect 2153 4253 2167 4267
rect 2133 4193 2147 4207
rect 2113 4153 2127 4167
rect 2153 4113 2167 4127
rect 2132 4053 2146 4067
rect 2153 4053 2167 4067
rect 2033 3991 2047 4005
rect 2093 3992 2107 4006
rect 2153 3993 2167 4007
rect 2053 3913 2067 3927
rect 2013 3813 2027 3827
rect 2073 3815 2087 3829
rect 2133 3953 2147 3967
rect 2133 3893 2147 3907
rect 2133 3853 2147 3867
rect 1913 3753 1927 3767
rect 1913 3673 1927 3687
rect 1893 3593 1907 3607
rect 1813 3553 1827 3567
rect 1873 3553 1887 3567
rect 1793 3513 1807 3527
rect 1733 3472 1747 3486
rect 1773 3472 1787 3486
rect 1673 3413 1687 3427
rect 1633 3294 1647 3308
rect 1793 3393 1807 3407
rect 1733 3373 1747 3387
rect 1713 3353 1727 3367
rect 2033 3773 2047 3787
rect 2073 3773 2087 3787
rect 2053 3733 2067 3747
rect 1973 3653 1987 3667
rect 1993 3633 2007 3647
rect 1973 3613 1987 3627
rect 1953 3513 1967 3527
rect 1993 3513 2007 3527
rect 1873 3433 1887 3447
rect 1932 3473 1946 3487
rect 1953 3473 1967 3487
rect 1933 3433 1947 3447
rect 1892 3413 1906 3427
rect 1913 3413 1927 3427
rect 1833 3373 1847 3387
rect 1813 3353 1827 3367
rect 1753 3333 1767 3347
rect 1793 3333 1807 3347
rect 1733 3313 1747 3327
rect 1413 3273 1427 3287
rect 1893 3353 1907 3367
rect 1893 3332 1907 3346
rect 1933 3333 1947 3347
rect 1853 3313 1867 3327
rect 1793 3295 1807 3309
rect 1833 3292 1847 3306
rect 1553 3252 1567 3266
rect 1533 3233 1547 3247
rect 1433 3193 1447 3207
rect 1413 3013 1427 3027
rect 1393 2993 1407 3007
rect 1453 3173 1467 3187
rect 1473 3053 1487 3067
rect 1433 2993 1447 3007
rect 1173 2951 1187 2965
rect 1213 2873 1227 2887
rect 1173 2833 1187 2847
rect 1073 2733 1087 2747
rect 1053 2653 1067 2667
rect 1093 2713 1107 2727
rect 1073 2613 1087 2627
rect 993 2553 1007 2567
rect 1113 2693 1127 2707
rect 1113 2633 1127 2647
rect 1133 2593 1147 2607
rect 1113 2553 1127 2567
rect 1353 2951 1367 2965
rect 1413 2953 1427 2967
rect 1233 2813 1247 2827
rect 1373 2933 1387 2947
rect 1393 2893 1407 2907
rect 1373 2793 1387 2807
rect 1173 2573 1187 2587
rect 1253 2775 1267 2789
rect 1353 2775 1367 2789
rect 1433 2853 1447 2867
rect 1453 2833 1467 2847
rect 1613 3233 1627 3247
rect 1672 3253 1686 3267
rect 1693 3253 1707 3267
rect 1733 3253 1747 3267
rect 1653 3173 1667 3187
rect 1793 3233 1807 3247
rect 1693 3193 1707 3207
rect 1833 3173 1847 3187
rect 1793 3133 1807 3147
rect 1833 3133 1847 3147
rect 1693 3113 1707 3127
rect 1653 2993 1667 3007
rect 1833 2972 1847 2986
rect 1993 3471 2007 3485
rect 2093 3693 2107 3707
rect 2273 4613 2287 4627
rect 2293 4573 2307 4587
rect 2353 4573 2367 4587
rect 2313 4553 2327 4567
rect 2513 4812 2527 4826
rect 2493 4773 2507 4787
rect 2473 4753 2487 4767
rect 2453 4713 2467 4727
rect 2413 4693 2427 4707
rect 2433 4673 2447 4687
rect 2473 4673 2487 4687
rect 2393 4653 2407 4667
rect 2413 4593 2427 4607
rect 2373 4553 2387 4567
rect 2453 4593 2467 4607
rect 2433 4573 2447 4587
rect 2513 4733 2527 4747
rect 2593 4813 2607 4827
rect 2553 4753 2567 4767
rect 2533 4693 2547 4707
rect 2513 4653 2527 4667
rect 2513 4593 2527 4607
rect 2493 4553 2507 4567
rect 2273 4513 2287 4527
rect 2252 4353 2266 4367
rect 2273 4353 2287 4367
rect 2333 4511 2347 4525
rect 2433 4493 2447 4507
rect 2473 4453 2487 4467
rect 2693 4773 2707 4787
rect 2653 4753 2667 4767
rect 2673 4733 2687 4747
rect 2653 4713 2667 4727
rect 2633 4613 2647 4627
rect 2533 4573 2547 4587
rect 2753 4853 2767 4867
rect 2793 4855 2807 4869
rect 2933 4993 2947 5007
rect 2913 4973 2927 4987
rect 2873 4933 2887 4947
rect 2873 4853 2887 4867
rect 3093 5373 3107 5387
rect 3133 5375 3147 5389
rect 3193 5373 3207 5387
rect 3093 5333 3107 5347
rect 3073 5253 3087 5267
rect 3093 5173 3107 5187
rect 3173 5333 3187 5347
rect 3433 5473 3447 5487
rect 3413 5453 3427 5467
rect 3772 5473 3786 5487
rect 3453 5453 3467 5467
rect 3733 5453 3747 5467
rect 3293 5433 3307 5447
rect 3433 5433 3447 5447
rect 3273 5412 3287 5426
rect 3233 5373 3247 5387
rect 3553 5413 3567 5427
rect 3633 5413 3647 5427
rect 3293 5393 3307 5407
rect 3313 5375 3327 5389
rect 3413 5375 3427 5389
rect 3453 5375 3467 5389
rect 3493 5373 3507 5387
rect 3373 5333 3387 5347
rect 3233 5313 3247 5327
rect 3333 5313 3347 5327
rect 3213 5293 3227 5307
rect 3193 5233 3207 5247
rect 3193 5193 3207 5207
rect 3193 5153 3207 5167
rect 3413 5333 3427 5347
rect 3393 5293 3407 5307
rect 3233 5273 3247 5287
rect 3292 5253 3306 5267
rect 3313 5253 3327 5267
rect 3393 5233 3407 5247
rect 3313 5213 3327 5227
rect 3233 5173 3247 5187
rect 3373 5173 3387 5187
rect 3213 5112 3227 5126
rect 2993 5073 3007 5087
rect 3073 5093 3087 5107
rect 3173 5093 3187 5107
rect 3053 5038 3067 5052
rect 3013 5013 3027 5027
rect 3073 5013 3087 5027
rect 3052 4993 3066 5007
rect 3073 4992 3087 5006
rect 2993 4973 3007 4987
rect 2973 4893 2987 4907
rect 2953 4873 2967 4887
rect 3053 4953 3067 4967
rect 2673 4693 2687 4707
rect 2733 4693 2747 4707
rect 2733 4613 2747 4627
rect 2653 4553 2667 4567
rect 2813 4813 2827 4827
rect 2753 4573 2767 4587
rect 2933 4813 2947 4827
rect 2913 4793 2927 4807
rect 2853 4773 2867 4787
rect 2893 4693 2907 4707
rect 2793 4613 2807 4627
rect 2873 4593 2887 4607
rect 2793 4573 2807 4587
rect 2733 4553 2747 4567
rect 2533 4453 2547 4467
rect 2433 4413 2447 4427
rect 2473 4413 2487 4427
rect 2513 4413 2527 4427
rect 2373 4393 2387 4407
rect 2293 4335 2307 4349
rect 2333 4335 2347 4349
rect 2373 4333 2387 4347
rect 2313 4292 2327 4306
rect 2213 4153 2227 4167
rect 2193 4073 2207 4087
rect 2333 4153 2347 4167
rect 2313 4133 2327 4147
rect 2373 4133 2387 4147
rect 2333 4093 2347 4107
rect 2433 4373 2447 4387
rect 2413 4353 2427 4367
rect 2433 4334 2447 4348
rect 2493 4292 2507 4306
rect 2473 4233 2487 4247
rect 2533 4233 2547 4247
rect 2453 4193 2467 4207
rect 2393 4093 2407 4107
rect 2313 4073 2327 4087
rect 2373 4073 2387 4087
rect 2233 4033 2247 4047
rect 2273 4033 2287 4047
rect 2213 3973 2227 3987
rect 2253 3973 2267 3987
rect 2173 3853 2187 3867
rect 2173 3833 2187 3847
rect 2152 3813 2166 3827
rect 2173 3813 2187 3827
rect 2353 4053 2367 4067
rect 2393 4034 2407 4048
rect 2453 4034 2467 4048
rect 2573 4493 2587 4507
rect 2613 4473 2627 4487
rect 2713 4473 2727 4487
rect 2653 4433 2667 4447
rect 2593 4373 2607 4387
rect 2593 4335 2607 4349
rect 2593 4293 2607 4307
rect 2573 4213 2587 4227
rect 2553 4173 2567 4187
rect 2533 4153 2547 4167
rect 2513 4133 2527 4147
rect 2513 4093 2527 4107
rect 2553 4113 2567 4127
rect 2633 4293 2647 4307
rect 2613 4153 2627 4167
rect 2613 4093 2627 4107
rect 2573 4073 2587 4087
rect 2713 4334 2727 4348
rect 2813 4553 2827 4567
rect 2913 4573 2927 4587
rect 2893 4553 2907 4567
rect 2953 4773 2967 4787
rect 3033 4873 3047 4887
rect 3213 5073 3227 5087
rect 3113 4953 3127 4967
rect 3233 5033 3247 5047
rect 3193 4953 3207 4967
rect 3233 4953 3247 4967
rect 3153 4933 3167 4947
rect 3173 4893 3187 4907
rect 3073 4873 3087 4887
rect 3053 4853 3067 4867
rect 3093 4855 3107 4869
rect 3073 4813 3087 4827
rect 3053 4793 3067 4807
rect 2973 4593 2987 4607
rect 2933 4553 2947 4567
rect 3033 4753 3047 4767
rect 3013 4733 3027 4747
rect 3073 4713 3087 4727
rect 3093 4673 3107 4687
rect 3073 4653 3087 4667
rect 3053 4633 3067 4647
rect 2993 4573 3007 4587
rect 3033 4573 3047 4587
rect 2793 4473 2807 4487
rect 3113 4653 3127 4667
rect 3093 4633 3107 4647
rect 3133 4593 3147 4607
rect 3113 4573 3127 4587
rect 3133 4554 3147 4568
rect 3353 5093 3367 5107
rect 3313 5073 3327 5087
rect 3453 5333 3467 5347
rect 3493 5333 3507 5347
rect 3433 5233 3447 5247
rect 3413 5193 3427 5207
rect 3493 5253 3507 5267
rect 3573 5313 3587 5327
rect 3533 5233 3547 5247
rect 3493 5213 3507 5227
rect 3473 5173 3487 5187
rect 3453 5093 3467 5107
rect 3333 5038 3347 5052
rect 3313 5013 3327 5027
rect 3353 5013 3367 5027
rect 3273 4993 3287 5007
rect 3353 4953 3367 4967
rect 3253 4893 3267 4907
rect 3433 5073 3447 5087
rect 3793 5413 3807 5427
rect 3873 5413 3887 5427
rect 3733 5393 3747 5407
rect 3653 5373 3667 5387
rect 3713 5374 3727 5388
rect 3753 5374 3767 5388
rect 3633 5293 3647 5307
rect 3573 5153 3587 5167
rect 3613 5153 3627 5167
rect 3493 5073 3507 5087
rect 3613 5113 3627 5127
rect 3693 5313 3707 5327
rect 3773 5333 3787 5347
rect 4033 5473 4047 5487
rect 4133 5473 4147 5487
rect 3993 5453 4007 5467
rect 3933 5433 3947 5447
rect 3833 5393 3847 5407
rect 3853 5393 3867 5407
rect 3913 5393 3927 5407
rect 3893 5374 3907 5388
rect 4053 5433 4067 5447
rect 4093 5433 4107 5447
rect 4073 5413 4087 5427
rect 4053 5393 4067 5407
rect 4033 5374 4047 5388
rect 3933 5353 3947 5367
rect 3753 5273 3767 5287
rect 3673 5233 3687 5247
rect 3733 5233 3747 5247
rect 3693 5213 3707 5227
rect 3652 5173 3666 5187
rect 3673 5173 3687 5187
rect 3653 5133 3667 5147
rect 3633 5093 3647 5107
rect 3673 5113 3687 5127
rect 3753 5153 3767 5167
rect 3473 5031 3487 5045
rect 3513 5033 3527 5047
rect 3453 5013 3467 5027
rect 3413 4992 3427 5006
rect 3393 4953 3407 4967
rect 3533 4993 3547 5007
rect 3453 4973 3467 4987
rect 3513 4973 3527 4987
rect 3413 4933 3427 4947
rect 3593 5032 3607 5046
rect 3653 5033 3667 5047
rect 3613 5013 3627 5027
rect 3553 4973 3567 4987
rect 3433 4913 3447 4927
rect 3492 4913 3506 4927
rect 3513 4913 3527 4927
rect 3613 4913 3627 4927
rect 3413 4893 3427 4907
rect 3313 4873 3327 4887
rect 3373 4873 3387 4887
rect 3253 4813 3267 4827
rect 3353 4812 3367 4826
rect 3253 4773 3267 4787
rect 3353 4733 3367 4747
rect 3333 4673 3347 4687
rect 3273 4613 3287 4627
rect 3173 4553 3187 4567
rect 3233 4554 3247 4568
rect 3313 4593 3327 4607
rect 3173 4532 3187 4546
rect 2833 4513 2847 4527
rect 2813 4453 2827 4467
rect 2773 4433 2787 4447
rect 2833 4373 2847 4387
rect 2893 4511 2907 4525
rect 2993 4511 3007 4525
rect 2873 4493 2887 4507
rect 2853 4333 2867 4347
rect 2733 4292 2747 4306
rect 2813 4293 2827 4307
rect 3013 4473 3027 4487
rect 2993 4433 3007 4447
rect 2973 4393 2987 4407
rect 2953 4373 2967 4387
rect 2893 4353 2907 4367
rect 2993 4353 3007 4367
rect 2953 4335 2967 4349
rect 3073 4513 3087 4527
rect 3153 4513 3167 4527
rect 3113 4453 3127 4467
rect 3033 4413 3047 4427
rect 3093 4413 3107 4427
rect 3093 4335 3107 4349
rect 3013 4313 3027 4327
rect 2693 4273 2707 4287
rect 2833 4233 2847 4247
rect 2673 4173 2687 4187
rect 2653 4133 2667 4147
rect 2593 4053 2607 4067
rect 2633 4053 2647 4067
rect 2553 4033 2567 4047
rect 2373 3973 2387 3987
rect 2373 3933 2387 3947
rect 2373 3912 2387 3926
rect 2433 3913 2447 3927
rect 2313 3873 2327 3887
rect 2413 3893 2427 3907
rect 2293 3813 2307 3827
rect 2353 3815 2367 3829
rect 2153 3773 2167 3787
rect 2153 3733 2167 3747
rect 2133 3633 2147 3647
rect 2113 3573 2127 3587
rect 2073 3533 2087 3547
rect 2233 3772 2247 3786
rect 2333 3773 2347 3787
rect 2373 3773 2387 3787
rect 2293 3753 2307 3767
rect 2233 3693 2247 3707
rect 2213 3673 2227 3687
rect 2333 3673 2347 3687
rect 2453 3853 2467 3867
rect 2573 3993 2587 4007
rect 2533 3933 2547 3947
rect 2493 3873 2507 3887
rect 2753 4053 2767 4067
rect 2673 4034 2687 4048
rect 2813 4053 2827 4067
rect 2833 3991 2847 4005
rect 2693 3973 2707 3987
rect 2732 3973 2746 3987
rect 2753 3973 2767 3987
rect 2793 3973 2807 3987
rect 2653 3953 2667 3967
rect 2633 3933 2647 3947
rect 2613 3873 2627 3887
rect 2573 3853 2587 3867
rect 2473 3833 2487 3847
rect 2493 3815 2507 3829
rect 2633 3815 2647 3829
rect 2732 3913 2746 3927
rect 2753 3913 2767 3927
rect 2793 3913 2807 3927
rect 2693 3833 2707 3847
rect 2733 3813 2747 3827
rect 2433 3773 2447 3787
rect 2193 3533 2207 3547
rect 2053 3453 2067 3467
rect 2053 3373 2067 3387
rect 2033 3353 2047 3367
rect 2053 3333 2067 3347
rect 1953 3313 1967 3327
rect 2033 3313 2047 3327
rect 1893 3294 1907 3308
rect 1933 3294 1947 3308
rect 2013 3295 2027 3309
rect 2093 3472 2107 3486
rect 2073 3293 2087 3307
rect 1893 3113 1907 3127
rect 1853 2953 1867 2967
rect 1633 2933 1647 2947
rect 1553 2913 1567 2927
rect 1453 2793 1467 2807
rect 1493 2793 1507 2807
rect 1253 2733 1267 2747
rect 1273 2673 1287 2687
rect 1213 2633 1227 2647
rect 1253 2633 1267 2647
rect 1413 2733 1427 2747
rect 1413 2693 1427 2707
rect 1513 2775 1527 2789
rect 1613 2913 1627 2927
rect 1773 2873 1787 2887
rect 1813 2873 1827 2887
rect 1713 2853 1727 2867
rect 1793 2853 1807 2867
rect 1633 2833 1647 2847
rect 1713 2813 1727 2827
rect 1653 2793 1667 2807
rect 1593 2773 1607 2787
rect 1693 2793 1707 2807
rect 1453 2653 1467 2667
rect 1533 2733 1547 2747
rect 1573 2733 1587 2747
rect 1373 2633 1387 2647
rect 1493 2633 1507 2647
rect 1633 2733 1647 2747
rect 1693 2733 1707 2747
rect 1673 2693 1687 2707
rect 1593 2613 1607 2627
rect 1253 2593 1267 2607
rect 1333 2593 1347 2607
rect 1493 2593 1507 2607
rect 1213 2553 1227 2567
rect 1793 2793 1807 2807
rect 1953 3253 1967 3267
rect 1993 3253 2007 3267
rect 2053 3253 2067 3267
rect 1953 3193 1967 3207
rect 1993 3173 2007 3187
rect 1973 3073 1987 3087
rect 2053 3173 2067 3187
rect 2133 3433 2147 3447
rect 2113 3413 2127 3427
rect 2133 3393 2147 3407
rect 2113 3373 2127 3387
rect 2293 3653 2307 3667
rect 2253 3513 2267 3527
rect 2313 3633 2327 3647
rect 2333 3613 2347 3627
rect 2373 3593 2387 3607
rect 2313 3573 2327 3587
rect 2333 3553 2347 3567
rect 2273 3471 2287 3485
rect 2233 3453 2247 3467
rect 2213 3433 2227 3447
rect 2193 3393 2207 3407
rect 2233 3392 2247 3406
rect 2212 3294 2226 3308
rect 2253 3373 2267 3387
rect 2253 3352 2267 3366
rect 2233 3293 2247 3307
rect 2313 3413 2327 3427
rect 2413 3653 2427 3667
rect 2413 3573 2427 3587
rect 2393 3513 2407 3527
rect 2473 3753 2487 3767
rect 2493 3673 2507 3687
rect 2453 3633 2467 3647
rect 2493 3633 2507 3647
rect 2533 3773 2547 3787
rect 2593 3772 2607 3786
rect 2633 3773 2647 3787
rect 2553 3733 2567 3747
rect 2533 3713 2547 3727
rect 2513 3533 2527 3547
rect 2553 3693 2567 3707
rect 2573 3653 2587 3667
rect 2733 3773 2747 3787
rect 2713 3753 2727 3767
rect 2713 3713 2727 3727
rect 2673 3693 2687 3707
rect 2653 3633 2667 3647
rect 2633 3613 2647 3627
rect 2653 3593 2667 3607
rect 2612 3553 2626 3567
rect 2633 3553 2647 3567
rect 2613 3532 2627 3546
rect 2573 3513 2587 3527
rect 2693 3673 2707 3687
rect 2833 3893 2847 3907
rect 2773 3873 2787 3887
rect 2913 4273 2927 4287
rect 2893 4253 2907 4267
rect 2893 4213 2907 4227
rect 3053 4293 3067 4307
rect 3053 4233 3067 4247
rect 2973 4213 2987 4227
rect 2913 4153 2927 4167
rect 2933 4133 2947 4147
rect 2913 4073 2927 4087
rect 2953 4073 2967 4087
rect 2933 4033 2947 4047
rect 3113 4253 3127 4267
rect 3113 4232 3127 4246
rect 3093 4153 3107 4167
rect 2993 4053 3007 4067
rect 3073 4054 3087 4068
rect 2913 3991 2927 4005
rect 2973 3993 2987 4007
rect 2873 3933 2887 3947
rect 2853 3833 2867 3847
rect 2833 3814 2847 3828
rect 2973 3893 2987 3907
rect 3133 4073 3147 4087
rect 3073 4033 3087 4047
rect 3113 4033 3127 4047
rect 3473 4854 3487 4868
rect 3553 4873 3567 4887
rect 3513 4853 3527 4867
rect 3573 4854 3587 4868
rect 3433 4793 3447 4807
rect 3493 4813 3507 4827
rect 3413 4673 3427 4687
rect 3452 4773 3466 4787
rect 3473 4773 3487 4787
rect 3373 4633 3387 4647
rect 3173 4493 3187 4507
rect 3253 4512 3267 4526
rect 3313 4513 3327 4527
rect 3213 4493 3227 4507
rect 3293 4473 3307 4487
rect 3393 4513 3407 4527
rect 3353 4413 3367 4427
rect 3233 4373 3247 4387
rect 3353 4373 3367 4387
rect 3333 4353 3347 4367
rect 3433 4633 3447 4647
rect 3473 4613 3487 4627
rect 3613 4813 3627 4827
rect 3593 4773 3607 4787
rect 3613 4753 3627 4767
rect 3593 4713 3607 4727
rect 3553 4653 3567 4667
rect 3593 4653 3607 4667
rect 3593 4593 3607 4607
rect 3493 4573 3507 4587
rect 3453 4553 3467 4567
rect 3493 4552 3507 4566
rect 3553 4573 3567 4587
rect 3593 4572 3607 4586
rect 3713 5073 3727 5087
rect 3773 5073 3787 5087
rect 3733 4993 3747 5007
rect 3673 4973 3687 4987
rect 3653 4853 3667 4867
rect 3753 4973 3767 4987
rect 3733 4953 3747 4967
rect 3753 4913 3767 4927
rect 3693 4873 3707 4887
rect 3733 4873 3747 4887
rect 3713 4854 3727 4868
rect 3833 5273 3847 5287
rect 4013 5313 4027 5327
rect 3953 5293 3967 5307
rect 3933 5253 3947 5267
rect 3873 5233 3887 5247
rect 3893 5213 3907 5227
rect 3832 5113 3846 5127
rect 3853 5113 3867 5127
rect 3853 5073 3867 5087
rect 4033 5273 4047 5287
rect 4133 5393 4147 5407
rect 4073 5373 4087 5387
rect 4113 5374 4127 5388
rect 4152 5374 4166 5388
rect 4213 5473 4227 5487
rect 4573 5473 4587 5487
rect 4193 5453 4207 5467
rect 4173 5373 4187 5387
rect 4173 5333 4187 5347
rect 4133 5293 4147 5307
rect 4093 5273 4107 5287
rect 4013 5253 4027 5267
rect 4053 5253 4067 5267
rect 4073 5233 4087 5247
rect 3953 5173 3967 5187
rect 3993 5153 4007 5167
rect 3933 5133 3947 5147
rect 3913 5093 3927 5107
rect 4053 5093 4067 5107
rect 4013 5073 4027 5087
rect 4093 5113 4107 5127
rect 4072 5073 4086 5087
rect 4093 5073 4107 5087
rect 4213 5433 4227 5447
rect 4593 5453 4607 5467
rect 4413 5413 4427 5427
rect 4552 5413 4566 5427
rect 4573 5413 4587 5427
rect 4233 5393 4247 5407
rect 4273 5393 4287 5407
rect 4333 5373 4347 5387
rect 4373 5375 4387 5389
rect 4493 5374 4507 5388
rect 4553 5375 4567 5389
rect 5333 5433 5347 5447
rect 4653 5413 4667 5427
rect 4233 5333 4247 5347
rect 4293 5333 4307 5347
rect 4253 5313 4267 5327
rect 4193 5273 4207 5287
rect 4233 5273 4247 5287
rect 4193 5252 4207 5266
rect 4173 5213 4187 5227
rect 3833 5033 3847 5047
rect 3813 5013 3827 5027
rect 3913 5031 3927 5045
rect 3872 4993 3886 5007
rect 3893 4993 3907 5007
rect 3873 4972 3887 4986
rect 3893 4953 3907 4967
rect 3873 4913 3887 4927
rect 3833 4893 3847 4907
rect 3693 4812 3707 4826
rect 3753 4813 3767 4827
rect 3733 4753 3747 4767
rect 3693 4713 3707 4727
rect 3653 4693 3667 4707
rect 3633 4633 3647 4647
rect 3653 4593 3667 4607
rect 3693 4692 3707 4706
rect 3753 4633 3767 4647
rect 3733 4593 3747 4607
rect 3833 4855 3847 4869
rect 3913 4933 3927 4947
rect 3913 4893 3927 4907
rect 3893 4853 3907 4867
rect 3813 4813 3827 4827
rect 3853 4813 3867 4827
rect 3893 4813 3907 4827
rect 3773 4573 3787 4587
rect 3753 4553 3767 4567
rect 3873 4753 3887 4767
rect 3853 4633 3867 4647
rect 3813 4573 3827 4587
rect 3433 4453 3447 4467
rect 3473 4511 3487 4525
rect 3473 4490 3487 4504
rect 3453 4373 3467 4387
rect 3573 4513 3587 4527
rect 3613 4511 3627 4525
rect 3673 4513 3687 4527
rect 3713 4512 3727 4526
rect 3773 4511 3787 4525
rect 3833 4511 3847 4525
rect 3733 4493 3747 4507
rect 3813 4493 3827 4507
rect 3573 4473 3587 4487
rect 3513 4453 3527 4467
rect 3673 4473 3687 4487
rect 3753 4473 3767 4487
rect 3593 4433 3607 4447
rect 3653 4433 3667 4447
rect 3533 4373 3547 4387
rect 3173 4253 3187 4267
rect 3232 4293 3246 4307
rect 3253 4293 3267 4307
rect 3293 4273 3307 4287
rect 3212 4233 3226 4247
rect 3233 4233 3247 4247
rect 3173 4113 3187 4127
rect 3253 4113 3267 4127
rect 3213 4033 3227 4047
rect 3013 3993 3027 4007
rect 3053 3992 3067 4006
rect 3133 3993 3147 4007
rect 3133 3953 3147 3967
rect 3093 3913 3107 3927
rect 3113 3893 3127 3907
rect 3013 3873 3027 3887
rect 2773 3733 2787 3747
rect 2813 3693 2827 3707
rect 2753 3673 2767 3687
rect 2733 3653 2747 3667
rect 2713 3633 2727 3647
rect 2713 3612 2727 3626
rect 2693 3573 2707 3587
rect 2673 3513 2687 3527
rect 2393 3471 2407 3485
rect 2453 3473 2467 3487
rect 2373 3433 2387 3447
rect 2333 3353 2347 3367
rect 2353 3333 2367 3347
rect 2133 3253 2147 3267
rect 2133 3213 2147 3227
rect 2173 3233 2187 3247
rect 2153 3193 2167 3207
rect 2013 3113 2027 3127
rect 1953 3053 1967 3067
rect 1993 3053 2007 3067
rect 1893 2993 1907 3007
rect 1953 2993 1967 3007
rect 1893 2953 1907 2967
rect 1873 2853 1887 2867
rect 1873 2813 1887 2827
rect 1773 2774 1787 2788
rect 1813 2774 1827 2788
rect 1913 2933 1927 2947
rect 1913 2833 1927 2847
rect 2092 3153 2106 3167
rect 2113 3153 2127 3167
rect 2073 3113 2087 3127
rect 2052 3053 2066 3067
rect 2073 3053 2087 3067
rect 2032 2994 2046 3008
rect 2213 3213 2227 3227
rect 2173 3073 2187 3087
rect 2133 3013 2147 3027
rect 2053 2993 2067 3007
rect 2153 2994 2167 3008
rect 2513 3472 2527 3486
rect 2553 3472 2567 3486
rect 2633 3471 2647 3485
rect 2673 3473 2687 3487
rect 2633 3413 2647 3427
rect 2453 3373 2467 3387
rect 2613 3373 2627 3387
rect 2453 3333 2467 3347
rect 2433 3295 2447 3309
rect 2553 3295 2567 3309
rect 2293 3253 2307 3267
rect 2333 3253 2347 3267
rect 2373 3253 2387 3267
rect 2273 3213 2287 3227
rect 2253 3193 2267 3207
rect 2253 3172 2267 3186
rect 2473 3253 2487 3267
rect 2533 3253 2547 3267
rect 2593 3253 2607 3267
rect 2573 3233 2587 3247
rect 2413 3213 2427 3227
rect 2573 3193 2587 3207
rect 2273 3153 2287 3167
rect 2393 3153 2407 3167
rect 2213 2993 2227 3007
rect 2073 2933 2087 2947
rect 1993 2913 2007 2927
rect 1973 2873 1987 2887
rect 1893 2793 1907 2807
rect 1933 2793 1947 2807
rect 2033 2775 2047 2789
rect 1713 2633 1727 2647
rect 1833 2733 1847 2747
rect 1793 2613 1807 2627
rect 1893 2732 1907 2746
rect 1933 2733 1947 2747
rect 1973 2733 1987 2747
rect 1933 2673 1947 2687
rect 1573 2533 1587 2547
rect 1693 2533 1707 2547
rect 1833 2533 1847 2547
rect 1913 2533 1927 2547
rect 1133 2513 1147 2527
rect 1193 2513 1207 2527
rect 1293 2513 1307 2527
rect 1453 2513 1467 2527
rect 1553 2513 1567 2527
rect 1113 2493 1127 2507
rect 913 2432 927 2446
rect 1053 2432 1067 2446
rect 873 2413 887 2427
rect 953 2413 967 2427
rect 973 2393 987 2407
rect 613 2373 627 2387
rect 733 2373 747 2387
rect 833 2373 847 2387
rect 953 2373 967 2387
rect 593 2313 607 2327
rect 673 2313 687 2327
rect 693 2293 707 2307
rect 853 2293 867 2307
rect 933 2293 947 2307
rect 673 2253 687 2267
rect 733 2273 747 2287
rect 773 2255 787 2269
rect 913 2255 927 2269
rect 593 2212 607 2226
rect 673 2213 687 2227
rect 553 2153 567 2167
rect 453 2053 467 2067
rect 533 2053 547 2067
rect 513 2013 527 2027
rect 433 1954 447 1968
rect 513 1953 527 1967
rect 553 1954 567 1968
rect 613 1954 627 1968
rect 653 1954 667 1968
rect 493 1912 507 1926
rect 433 1893 447 1907
rect 613 1893 627 1907
rect 413 1813 427 1827
rect 593 1753 607 1767
rect 453 1734 467 1748
rect 493 1734 507 1748
rect 553 1735 567 1749
rect 393 1653 407 1667
rect 453 1493 467 1507
rect 573 1633 587 1647
rect 573 1434 587 1448
rect 333 1373 347 1387
rect 413 1373 427 1387
rect 113 1313 127 1327
rect 93 1273 107 1287
rect 193 1273 207 1287
rect 133 1233 147 1247
rect 53 1214 67 1228
rect 33 1173 47 1187
rect 213 1214 227 1228
rect 473 1392 487 1406
rect 513 1393 527 1407
rect 553 1392 567 1406
rect 593 1393 607 1407
rect 773 2213 787 2227
rect 833 2213 847 2227
rect 753 2193 767 2207
rect 713 2173 727 2187
rect 913 2213 927 2227
rect 1033 2392 1047 2406
rect 993 2333 1007 2347
rect 973 2313 987 2327
rect 953 2273 967 2287
rect 1013 2313 1027 2327
rect 1013 2273 1027 2287
rect 973 2212 987 2226
rect 933 2173 947 2187
rect 1093 2212 1107 2226
rect 1013 2173 1027 2187
rect 873 2153 887 2167
rect 973 2153 987 2167
rect 773 2133 787 2147
rect 673 1873 687 1887
rect 653 1853 667 1867
rect 1013 2053 1027 2067
rect 1173 2473 1187 2487
rect 1213 2473 1227 2487
rect 1353 2474 1367 2488
rect 1413 2474 1427 2488
rect 1153 2433 1167 2447
rect 1233 2433 1247 2447
rect 1193 2393 1207 2407
rect 1153 2333 1167 2347
rect 1153 2254 1167 2268
rect 1273 2432 1287 2446
rect 1333 2433 1347 2447
rect 1473 2493 1487 2507
rect 1413 2373 1427 2387
rect 1453 2373 1467 2387
rect 1333 2353 1347 2367
rect 1393 2353 1407 2367
rect 1313 2313 1327 2327
rect 1353 2313 1367 2327
rect 1253 2293 1267 2307
rect 1333 2293 1347 2307
rect 1293 2254 1307 2268
rect 1253 2213 1267 2227
rect 1313 2212 1327 2226
rect 1153 2133 1167 2147
rect 1333 2053 1347 2067
rect 993 2033 1007 2047
rect 1133 2033 1147 2047
rect 1293 2033 1307 2047
rect 793 2013 807 2027
rect 773 1893 787 1907
rect 773 1872 787 1886
rect 753 1813 767 1827
rect 733 1753 747 1767
rect 633 1734 647 1748
rect 693 1734 707 1748
rect 633 1693 647 1707
rect 833 1953 847 1967
rect 873 1953 887 1967
rect 913 1953 927 1967
rect 953 1954 967 1968
rect 813 1913 827 1927
rect 853 1911 867 1925
rect 1153 1954 1167 1968
rect 1233 1954 1247 1968
rect 973 1853 987 1867
rect 913 1813 927 1827
rect 913 1773 927 1787
rect 813 1753 827 1767
rect 793 1733 807 1747
rect 1073 1912 1087 1926
rect 1133 1913 1147 1927
rect 1013 1753 1027 1767
rect 993 1733 1007 1747
rect 913 1713 927 1727
rect 713 1692 727 1706
rect 773 1692 787 1706
rect 813 1653 827 1667
rect 633 1633 647 1647
rect 613 1333 627 1347
rect 593 1273 607 1287
rect 433 1233 447 1247
rect 513 1233 527 1247
rect 573 1233 587 1247
rect 213 1173 227 1187
rect 253 1172 267 1186
rect 333 1093 347 1107
rect 73 1073 87 1087
rect 153 1073 167 1087
rect 193 1073 207 1087
rect 93 933 107 947
rect 33 873 47 887
rect 73 872 87 886
rect 333 953 347 967
rect 273 933 287 947
rect 213 914 227 928
rect 153 853 167 867
rect 193 853 207 867
rect 33 813 47 827
rect 113 813 127 827
rect 113 753 127 767
rect 533 1172 547 1186
rect 713 1533 727 1547
rect 813 1513 827 1527
rect 853 1513 867 1527
rect 953 1513 967 1527
rect 813 1473 827 1487
rect 713 1433 727 1447
rect 973 1473 987 1487
rect 933 1434 947 1448
rect 693 1392 707 1406
rect 793 1392 807 1406
rect 753 1333 767 1347
rect 853 1293 867 1307
rect 833 1273 847 1287
rect 633 1233 647 1247
rect 713 1233 727 1247
rect 653 1214 667 1228
rect 633 1172 647 1186
rect 433 1153 447 1167
rect 573 1153 587 1167
rect 753 1233 767 1247
rect 833 1213 847 1227
rect 933 1273 947 1287
rect 893 1233 907 1247
rect 673 1133 687 1147
rect 713 1172 727 1186
rect 773 1172 787 1186
rect 813 1172 827 1186
rect 853 1172 867 1186
rect 913 1172 927 1186
rect 813 1151 827 1165
rect 793 1133 807 1147
rect 773 1033 787 1047
rect 613 953 627 967
rect 693 953 707 967
rect 373 913 387 927
rect 433 914 447 928
rect 473 913 487 927
rect 533 914 547 928
rect 313 872 327 886
rect 373 872 387 886
rect 353 853 367 867
rect 313 813 327 827
rect 273 793 287 807
rect 233 733 247 747
rect 293 733 307 747
rect 233 694 247 708
rect 53 673 67 687
rect 173 652 187 666
rect 253 652 267 666
rect 113 613 127 627
rect 73 453 87 467
rect 413 813 427 827
rect 513 872 527 886
rect 533 853 547 867
rect 373 793 387 807
rect 473 793 487 807
rect 513 753 527 767
rect 473 733 487 747
rect 313 693 327 707
rect 353 694 367 708
rect 393 694 407 708
rect 553 833 567 847
rect 593 793 607 807
rect 653 914 667 928
rect 653 893 667 907
rect 773 893 787 907
rect 713 853 727 867
rect 573 753 587 767
rect 613 753 627 767
rect 673 753 687 767
rect 533 733 547 747
rect 653 712 667 726
rect 1153 1893 1167 1907
rect 1253 1912 1267 1926
rect 1233 1893 1247 1907
rect 1213 1853 1227 1867
rect 1192 1773 1206 1787
rect 1213 1773 1227 1787
rect 1153 1734 1167 1748
rect 1413 2254 1427 2268
rect 1553 2474 1567 2488
rect 1533 2432 1547 2446
rect 1813 2513 1827 2527
rect 1613 2493 1627 2507
rect 1673 2473 1687 2487
rect 1713 2473 1727 2487
rect 1773 2474 1787 2488
rect 1633 2432 1647 2446
rect 1692 2433 1706 2447
rect 1653 2393 1667 2407
rect 1713 2432 1727 2446
rect 1753 2432 1767 2446
rect 1573 2313 1587 2327
rect 1593 2273 1607 2287
rect 1553 2254 1567 2268
rect 1453 2212 1467 2226
rect 1413 2193 1427 2207
rect 1393 2173 1407 2187
rect 1573 2212 1587 2226
rect 1493 2193 1507 2207
rect 1613 2173 1627 2187
rect 1453 2153 1467 2167
rect 1693 2333 1707 2347
rect 1873 2493 1887 2507
rect 2133 2952 2147 2966
rect 2153 2933 2167 2947
rect 2093 2913 2107 2927
rect 2113 2833 2127 2847
rect 2133 2813 2147 2827
rect 2113 2793 2127 2807
rect 2213 2953 2227 2967
rect 2573 3113 2587 3127
rect 2713 3553 2727 3567
rect 2733 3532 2747 3546
rect 2873 3753 2887 3767
rect 2873 3713 2887 3727
rect 2873 3673 2887 3687
rect 2973 3772 2987 3786
rect 2973 3733 2987 3747
rect 2873 3633 2887 3647
rect 2853 3593 2867 3607
rect 2873 3573 2887 3587
rect 2853 3553 2867 3567
rect 3113 3753 3127 3767
rect 3033 3733 3047 3747
rect 3012 3713 3026 3727
rect 3033 3712 3047 3726
rect 3113 3713 3127 3727
rect 3193 3991 3207 4005
rect 3153 3933 3167 3947
rect 3153 3912 3167 3926
rect 3213 3815 3227 3829
rect 3413 4293 3427 4307
rect 3393 4273 3407 4287
rect 3373 4253 3387 4267
rect 3333 4173 3347 4187
rect 3513 4293 3527 4307
rect 3493 4253 3507 4267
rect 3433 4213 3447 4227
rect 3493 4213 3507 4227
rect 3453 4193 3467 4207
rect 3413 4153 3427 4167
rect 3413 4073 3427 4087
rect 3333 4032 3347 4046
rect 3273 3953 3287 3967
rect 3313 3953 3327 3967
rect 3613 4393 3627 4407
rect 3593 4333 3607 4347
rect 3553 4293 3567 4307
rect 3533 4193 3547 4207
rect 3533 4172 3547 4186
rect 3513 4133 3527 4147
rect 3613 4273 3627 4287
rect 3593 4253 3607 4267
rect 3613 4173 3627 4187
rect 3613 4152 3627 4166
rect 3553 4113 3567 4127
rect 3593 4113 3607 4127
rect 3573 4093 3587 4107
rect 3553 4073 3567 4087
rect 3533 4053 3547 4067
rect 3653 4293 3667 4307
rect 3653 4233 3667 4247
rect 3633 4133 3647 4147
rect 3633 4112 3647 4126
rect 3633 4073 3647 4087
rect 3493 4033 3507 4047
rect 3613 4053 3627 4067
rect 3393 3993 3407 4007
rect 3433 3992 3447 4006
rect 3412 3933 3426 3947
rect 3433 3933 3447 3947
rect 3473 3933 3487 3947
rect 3513 3933 3527 3947
rect 3393 3913 3407 3927
rect 3373 3853 3387 3867
rect 2973 3653 2987 3667
rect 3053 3653 3067 3667
rect 2933 3633 2947 3647
rect 3033 3633 3047 3647
rect 2813 3533 2827 3547
rect 2913 3533 2927 3547
rect 2793 3514 2807 3528
rect 3173 3653 3187 3667
rect 3073 3613 3087 3627
rect 3153 3613 3167 3627
rect 3053 3573 3067 3587
rect 2973 3533 2987 3547
rect 2933 3513 2947 3527
rect 3033 3514 3047 3528
rect 2693 3433 2707 3447
rect 2673 3393 2687 3407
rect 2733 3472 2747 3486
rect 2753 3433 2767 3447
rect 2733 3373 2747 3387
rect 2833 3473 2847 3487
rect 2773 3413 2787 3427
rect 2753 3353 2767 3367
rect 2893 3471 2907 3485
rect 2933 3473 2947 3487
rect 2953 3453 2967 3467
rect 2953 3413 2967 3427
rect 3093 3593 3107 3607
rect 3173 3573 3187 3587
rect 3093 3533 3107 3547
rect 3013 3393 3027 3407
rect 3073 3393 3087 3407
rect 2893 3373 2907 3387
rect 2933 3373 2947 3387
rect 2873 3353 2887 3367
rect 2693 3333 2707 3347
rect 2853 3333 2867 3347
rect 2713 3313 2727 3327
rect 2733 3293 2747 3307
rect 2813 3294 2827 3308
rect 2633 3253 2647 3267
rect 2673 3253 2687 3267
rect 2713 3233 2727 3247
rect 2853 3253 2867 3267
rect 2793 3193 2807 3207
rect 2633 3133 2647 3147
rect 2753 3133 2767 3147
rect 2613 3113 2627 3127
rect 2593 3093 2607 3107
rect 2313 3073 2327 3087
rect 2373 3013 2387 3027
rect 2473 3013 2487 3027
rect 2433 2994 2447 3008
rect 2353 2953 2367 2967
rect 2713 3093 2727 3107
rect 2173 2853 2187 2867
rect 2133 2732 2147 2746
rect 2233 2933 2247 2947
rect 2293 2933 2307 2947
rect 2313 2893 2327 2907
rect 2353 2853 2367 2867
rect 2313 2813 2327 2827
rect 2253 2774 2267 2788
rect 2293 2774 2307 2788
rect 2433 2774 2447 2788
rect 2013 2713 2027 2727
rect 2073 2713 2087 2727
rect 2193 2733 2207 2747
rect 2233 2732 2247 2746
rect 2273 2713 2287 2727
rect 2153 2613 2167 2627
rect 2133 2593 2147 2607
rect 2193 2513 2207 2527
rect 1993 2493 2007 2507
rect 1953 2473 1967 2487
rect 1973 2453 1987 2467
rect 1833 2433 1847 2447
rect 1813 2413 1827 2427
rect 1793 2393 1807 2407
rect 1833 2393 1847 2407
rect 1813 2333 1827 2347
rect 1793 2313 1807 2327
rect 1673 2293 1687 2307
rect 1713 2293 1727 2307
rect 1673 2253 1687 2267
rect 1713 2255 1727 2269
rect 1773 2253 1787 2267
rect 1933 2431 1947 2445
rect 1893 2413 1907 2427
rect 1873 2393 1887 2407
rect 1693 2213 1707 2227
rect 1673 2053 1687 2067
rect 1353 1953 1367 1967
rect 1493 1973 1507 1987
rect 1513 1953 1527 1967
rect 1353 1911 1367 1925
rect 1293 1853 1307 1867
rect 1733 2213 1747 2227
rect 1773 2173 1787 2187
rect 1813 2133 1827 2147
rect 1773 2033 1787 2047
rect 1713 1993 1727 2007
rect 1693 1953 1707 1967
rect 1473 1911 1487 1925
rect 1613 1833 1627 1847
rect 1353 1813 1367 1827
rect 1413 1813 1427 1827
rect 1553 1813 1567 1827
rect 1633 1813 1647 1827
rect 1313 1773 1327 1787
rect 1233 1734 1247 1748
rect 1273 1734 1287 1748
rect 1433 1773 1447 1787
rect 1053 1693 1067 1707
rect 1093 1693 1107 1707
rect 1013 1653 1027 1667
rect 1173 1692 1187 1706
rect 1233 1693 1247 1707
rect 1293 1692 1307 1706
rect 1113 1673 1127 1687
rect 1093 1533 1107 1547
rect 1333 1653 1347 1667
rect 1353 1633 1367 1647
rect 1333 1553 1347 1567
rect 1173 1533 1187 1547
rect 1273 1533 1287 1547
rect 1313 1533 1327 1547
rect 1113 1513 1127 1527
rect 993 1273 1007 1287
rect 1073 1273 1087 1287
rect 993 1233 1007 1247
rect 993 1173 1007 1187
rect 913 1133 927 1147
rect 973 1133 987 1147
rect 873 993 887 1007
rect 813 913 827 927
rect 1033 1093 1047 1107
rect 1013 953 1027 967
rect 933 914 947 928
rect 973 914 987 928
rect 1273 1493 1287 1507
rect 1293 1453 1307 1467
rect 1273 1434 1287 1448
rect 1193 1392 1207 1406
rect 1213 1313 1227 1327
rect 1153 1233 1167 1247
rect 1233 1273 1247 1287
rect 1253 1233 1267 1247
rect 1593 1753 1607 1767
rect 1453 1653 1467 1667
rect 1373 1593 1387 1607
rect 1433 1593 1447 1607
rect 1413 1453 1427 1467
rect 1493 1613 1507 1627
rect 1513 1593 1527 1607
rect 1513 1553 1527 1567
rect 1553 1473 1567 1487
rect 1493 1373 1507 1387
rect 1913 2254 1927 2268
rect 1933 2212 1947 2226
rect 1953 2133 1967 2147
rect 1873 2093 1887 2107
rect 1853 2033 1867 2047
rect 1833 1953 1847 1967
rect 1793 1911 1807 1925
rect 1833 1911 1847 1925
rect 1913 1993 1927 2007
rect 2053 2474 2067 2488
rect 2153 2474 2167 2488
rect 2393 2732 2407 2746
rect 2433 2733 2447 2747
rect 2553 2952 2567 2966
rect 2673 2994 2687 3008
rect 2853 3232 2867 3246
rect 2853 3133 2867 3147
rect 2833 3113 2847 3127
rect 2933 3313 2947 3327
rect 2893 3293 2907 3307
rect 2973 3295 2987 3309
rect 2893 3253 2907 3267
rect 2873 3093 2887 3107
rect 2953 3233 2967 3247
rect 2933 3193 2947 3207
rect 2913 3153 2927 3167
rect 3053 3153 3067 3167
rect 2893 3033 2907 3047
rect 2973 3033 2987 3047
rect 2793 2993 2807 3007
rect 2833 2993 2847 3007
rect 2873 2993 2887 3007
rect 2913 2993 2927 3007
rect 2713 2953 2727 2967
rect 2633 2913 2647 2927
rect 2593 2893 2607 2907
rect 2593 2833 2607 2847
rect 2513 2774 2527 2788
rect 2533 2653 2547 2667
rect 2313 2613 2327 2627
rect 2453 2613 2467 2627
rect 2593 2794 2607 2808
rect 2593 2773 2607 2787
rect 2613 2732 2627 2746
rect 2613 2711 2627 2725
rect 2553 2633 2567 2647
rect 2533 2553 2547 2567
rect 2293 2513 2307 2527
rect 2513 2513 2527 2527
rect 2273 2493 2287 2507
rect 2232 2474 2246 2488
rect 2253 2474 2267 2488
rect 2473 2493 2487 2507
rect 2333 2474 2347 2488
rect 2433 2474 2447 2488
rect 2073 2432 2087 2446
rect 2033 2393 2047 2407
rect 2013 2353 2027 2367
rect 1993 2333 2007 2347
rect 2093 2333 2107 2347
rect 1993 2253 2007 2267
rect 2053 2255 2067 2269
rect 2233 2433 2247 2447
rect 2173 2353 2187 2367
rect 2133 2313 2147 2327
rect 2233 2293 2247 2307
rect 2093 2253 2107 2267
rect 2153 2255 2167 2269
rect 2213 2253 2227 2267
rect 2573 2474 2587 2488
rect 2253 2273 2267 2287
rect 2033 2213 2047 2227
rect 1993 2133 2007 2147
rect 2113 2213 2127 2227
rect 2073 2093 2087 2107
rect 2013 2033 2027 2047
rect 2133 2173 2147 2187
rect 2273 2212 2287 2226
rect 2213 2153 2227 2167
rect 2173 2133 2187 2147
rect 2113 1973 2127 1987
rect 2053 1953 2067 1967
rect 2093 1953 2107 1967
rect 1873 1913 1887 1927
rect 1833 1873 1847 1887
rect 1773 1833 1787 1847
rect 1753 1813 1767 1827
rect 1713 1773 1727 1787
rect 1753 1753 1767 1767
rect 1853 1773 1867 1787
rect 1593 1613 1607 1627
rect 1653 1613 1667 1627
rect 1613 1473 1627 1487
rect 1573 1433 1587 1447
rect 1673 1434 1687 1448
rect 1693 1393 1707 1407
rect 1433 1293 1447 1307
rect 1553 1293 1567 1307
rect 1373 1273 1387 1287
rect 1313 1233 1327 1247
rect 1353 1233 1367 1247
rect 1393 1233 1407 1247
rect 1293 1213 1307 1227
rect 1573 1273 1587 1287
rect 1453 1233 1467 1247
rect 1433 1213 1447 1227
rect 1113 1173 1127 1187
rect 1173 1173 1187 1187
rect 1213 1173 1227 1187
rect 1073 1033 1087 1047
rect 1133 933 1147 947
rect 1073 914 1087 928
rect 893 853 907 867
rect 893 832 907 846
rect 953 872 967 886
rect 993 872 1007 886
rect 1053 873 1067 887
rect 853 813 867 827
rect 893 773 907 787
rect 1273 1172 1287 1186
rect 1373 1173 1387 1187
rect 1413 1173 1427 1187
rect 1473 1213 1487 1227
rect 1533 1214 1547 1228
rect 1593 1253 1607 1267
rect 1733 1693 1747 1707
rect 1733 1633 1747 1647
rect 1713 1373 1727 1387
rect 1713 1233 1727 1247
rect 1593 1213 1607 1227
rect 1453 1153 1467 1167
rect 1713 1193 1727 1207
rect 1513 1172 1527 1186
rect 1613 1172 1627 1186
rect 1553 1153 1567 1167
rect 1473 1133 1487 1147
rect 1533 1133 1547 1147
rect 1573 1133 1587 1147
rect 1673 1133 1687 1147
rect 1553 993 1567 1007
rect 1493 973 1507 987
rect 1393 953 1407 967
rect 1473 953 1487 967
rect 1293 913 1307 927
rect 1333 913 1347 927
rect 1373 913 1387 927
rect 1413 913 1427 927
rect 1493 933 1507 947
rect 1513 914 1527 928
rect 1253 872 1267 886
rect 1293 872 1307 886
rect 1353 871 1367 885
rect 1393 853 1407 867
rect 1293 793 1307 807
rect 1193 773 1207 787
rect 1053 753 1067 767
rect 1093 753 1107 767
rect 313 652 327 666
rect 413 653 427 667
rect 453 653 467 667
rect 493 653 507 667
rect 533 653 547 667
rect 193 493 207 507
rect 293 493 307 507
rect 113 393 127 407
rect 93 352 107 366
rect 133 352 147 366
rect 33 174 47 188
rect 93 174 107 188
rect 133 174 147 188
rect 713 652 727 666
rect 533 613 547 627
rect 773 613 787 627
rect 413 453 427 467
rect 313 413 327 427
rect 253 394 267 408
rect 453 394 467 408
rect 493 394 507 408
rect 853 653 867 667
rect 933 653 947 667
rect 1053 652 1067 666
rect 1493 872 1507 886
rect 1473 853 1487 867
rect 1453 833 1467 847
rect 1613 973 1627 987
rect 1653 973 1667 987
rect 1713 933 1727 947
rect 1553 833 1567 847
rect 1473 813 1487 827
rect 1113 733 1127 747
rect 1253 733 1267 747
rect 1413 733 1427 747
rect 1173 694 1187 708
rect 1213 694 1227 708
rect 1293 713 1307 727
rect 1113 652 1127 666
rect 1353 693 1367 707
rect 1413 695 1427 709
rect 1273 652 1287 666
rect 1313 652 1327 666
rect 1353 652 1367 666
rect 1433 653 1447 667
rect 873 613 887 627
rect 993 613 1007 627
rect 1093 613 1107 627
rect 1213 613 1227 627
rect 1393 613 1407 627
rect 813 553 827 567
rect 693 413 707 427
rect 813 413 827 427
rect 573 393 587 407
rect 433 352 447 366
rect 493 353 507 367
rect 553 351 567 365
rect 633 352 647 366
rect 393 333 407 347
rect 353 213 367 227
rect 433 213 447 227
rect 393 174 407 188
rect 493 173 507 187
rect 553 175 567 189
rect 633 174 647 188
rect 73 132 87 146
rect 193 132 207 146
rect 253 132 267 146
rect 353 133 367 147
rect 313 113 327 127
rect 453 132 467 146
rect 493 132 507 146
rect 533 133 547 147
rect 573 133 587 147
rect 713 394 727 408
rect 753 394 767 408
rect 853 352 867 366
rect 993 553 1007 567
rect 933 394 947 408
rect 1253 533 1267 547
rect 1113 493 1127 507
rect 1233 493 1247 507
rect 1093 413 1107 427
rect 1053 393 1067 407
rect 1133 413 1147 427
rect 1193 413 1207 427
rect 873 333 887 347
rect 713 293 727 307
rect 993 353 1007 367
rect 1073 313 1087 327
rect 1033 293 1047 307
rect 1073 233 1087 247
rect 953 193 967 207
rect 713 173 727 187
rect 853 173 867 187
rect 913 174 927 188
rect 993 173 1007 187
rect 1033 175 1047 189
rect 1793 1693 1807 1707
rect 1833 1693 1847 1707
rect 1893 1893 1907 1907
rect 1933 1873 1947 1887
rect 1913 1813 1927 1827
rect 2033 1813 2047 1827
rect 2013 1773 2027 1787
rect 1953 1753 1967 1767
rect 2053 1734 2067 1748
rect 2153 1954 2167 1968
rect 2353 2432 2367 2446
rect 2413 2432 2427 2446
rect 2413 2393 2427 2407
rect 2333 2333 2347 2347
rect 2253 1953 2267 1967
rect 2313 1953 2327 1967
rect 2173 1793 2187 1807
rect 2113 1753 2127 1767
rect 2093 1733 2107 1747
rect 2233 1913 2247 1927
rect 2253 1853 2267 1867
rect 2233 1793 2247 1807
rect 2193 1753 2207 1767
rect 1873 1693 1887 1707
rect 1853 1613 1867 1627
rect 1813 1513 1827 1527
rect 1973 1693 1987 1707
rect 1933 1613 1947 1627
rect 2113 1693 2127 1707
rect 2153 1693 2167 1707
rect 2213 1693 2227 1707
rect 1973 1593 1987 1607
rect 1953 1553 1967 1567
rect 2213 1653 2227 1667
rect 2153 1613 2167 1627
rect 2033 1553 2047 1567
rect 2153 1553 2167 1567
rect 2013 1513 2027 1527
rect 1993 1473 2007 1487
rect 1793 1214 1807 1228
rect 1853 1273 1867 1287
rect 1893 1253 1907 1267
rect 1853 1213 1867 1227
rect 1973 1391 1987 1405
rect 1953 1373 1967 1387
rect 2153 1513 2167 1527
rect 2113 1493 2127 1507
rect 2073 1434 2087 1448
rect 2313 1913 2327 1927
rect 2373 2293 2387 2307
rect 2513 2433 2527 2447
rect 2553 2413 2567 2427
rect 2553 2353 2567 2367
rect 2513 2333 2527 2347
rect 2453 2293 2467 2307
rect 2453 2253 2467 2267
rect 2573 2293 2587 2307
rect 2553 2253 2567 2267
rect 2753 2833 2767 2847
rect 2673 2813 2687 2827
rect 2853 2953 2867 2967
rect 2893 2951 2907 2965
rect 2952 2953 2966 2967
rect 3053 2994 3067 3008
rect 3173 3513 3187 3527
rect 3153 3472 3167 3486
rect 3213 3773 3227 3787
rect 3233 3733 3247 3747
rect 3213 3613 3227 3627
rect 3253 3653 3267 3667
rect 3213 3513 3227 3527
rect 3373 3814 3387 3828
rect 3313 3772 3327 3786
rect 3293 3753 3307 3767
rect 3393 3773 3407 3787
rect 3353 3713 3367 3727
rect 3553 3973 3567 3987
rect 3533 3913 3547 3927
rect 3553 3893 3567 3907
rect 3733 4453 3747 4467
rect 3693 4393 3707 4407
rect 3693 4333 3707 4347
rect 3753 4393 3767 4407
rect 3833 4413 3847 4427
rect 3713 4273 3727 4287
rect 3733 4253 3747 4267
rect 3693 4233 3707 4247
rect 3673 4153 3687 4167
rect 3653 4033 3667 4047
rect 3773 4293 3787 4307
rect 3732 4113 3746 4127
rect 3753 4113 3767 4127
rect 3993 5013 4007 5027
rect 3973 4873 3987 4887
rect 4072 5033 4086 5047
rect 4033 4973 4047 4987
rect 4113 4993 4127 5007
rect 4173 5033 4187 5047
rect 4153 4973 4167 4987
rect 4053 4913 4067 4927
rect 4073 4893 4087 4907
rect 4113 4854 4127 4868
rect 4173 4953 4187 4967
rect 4313 5253 4327 5267
rect 4293 5193 4307 5207
rect 4253 5133 4267 5147
rect 4233 5073 4247 5087
rect 4313 5173 4327 5187
rect 4373 5333 4387 5347
rect 4333 5153 4347 5167
rect 4313 5133 4327 5147
rect 4333 5113 4347 5127
rect 4473 5333 4487 5347
rect 4433 5313 4447 5327
rect 4613 5332 4627 5346
rect 4413 5213 4427 5227
rect 4473 5213 4487 5227
rect 4373 5074 4387 5088
rect 4553 5193 4567 5207
rect 4513 5074 4527 5088
rect 5033 5393 5047 5407
rect 4713 5375 4727 5389
rect 4753 5375 4767 5389
rect 4793 5373 4807 5387
rect 4833 5374 4847 5388
rect 4873 5374 4887 5388
rect 4933 5375 4947 5389
rect 4993 5375 5007 5389
rect 5133 5375 5147 5389
rect 5253 5375 5267 5389
rect 5293 5375 5307 5389
rect 4693 5333 4707 5347
rect 4733 5333 4747 5347
rect 4673 5233 4687 5247
rect 4673 5193 4687 5207
rect 4653 5153 4667 5167
rect 4593 5113 4607 5127
rect 4573 5093 4587 5107
rect 4213 5013 4227 5027
rect 4193 4933 4207 4947
rect 4273 5031 4287 5045
rect 4333 5032 4347 5046
rect 4253 5013 4267 5027
rect 4233 4913 4247 4927
rect 4433 5032 4447 5046
rect 4413 4993 4427 5007
rect 4393 4973 4407 4987
rect 4313 4933 4327 4947
rect 4013 4813 4027 4827
rect 3913 4733 3927 4747
rect 4013 4773 4027 4787
rect 3933 4713 3947 4727
rect 3893 4673 3907 4687
rect 3933 4673 3947 4687
rect 3993 4673 4007 4687
rect 3873 4473 3887 4487
rect 3993 4593 4007 4607
rect 3973 4553 3987 4567
rect 3913 4433 3927 4447
rect 3853 4333 3867 4347
rect 3893 4333 3907 4347
rect 3993 4513 4007 4527
rect 3973 4433 3987 4447
rect 3953 4393 3967 4407
rect 3913 4293 3927 4307
rect 3833 4233 3847 4247
rect 3813 4193 3827 4207
rect 3753 4092 3767 4106
rect 3713 4073 3727 4087
rect 3893 4273 3907 4287
rect 3873 4173 3887 4187
rect 3853 4153 3867 4167
rect 3813 4053 3827 4067
rect 3793 4032 3807 4046
rect 3833 4033 3847 4047
rect 3653 3993 3667 4007
rect 3633 3953 3647 3967
rect 3593 3913 3607 3927
rect 3513 3873 3527 3887
rect 3573 3873 3587 3887
rect 3453 3853 3467 3867
rect 3533 3853 3547 3867
rect 3432 3813 3446 3827
rect 3453 3815 3467 3829
rect 3653 3893 3667 3907
rect 3593 3833 3607 3847
rect 3533 3814 3547 3828
rect 3573 3814 3587 3828
rect 3473 3773 3487 3787
rect 3513 3773 3527 3787
rect 3733 3993 3747 4007
rect 3713 3973 3727 3987
rect 3673 3853 3687 3867
rect 3653 3813 3667 3827
rect 3813 3973 3827 3987
rect 4293 4853 4307 4867
rect 4173 4793 4187 4807
rect 4133 4773 4147 4787
rect 4213 4693 4227 4707
rect 4073 4633 4087 4647
rect 4053 4593 4067 4607
rect 4033 4553 4047 4567
rect 4153 4573 4167 4587
rect 4272 4813 4286 4827
rect 4293 4813 4307 4827
rect 4253 4791 4267 4805
rect 4233 4673 4247 4687
rect 4093 4553 4107 4567
rect 4033 4513 4047 4527
rect 4013 4493 4027 4507
rect 4073 4493 4087 4507
rect 4193 4473 4207 4487
rect 4273 4473 4287 4487
rect 4033 4433 4047 4447
rect 4213 4413 4227 4427
rect 4033 4393 4047 4407
rect 4073 4393 4087 4407
rect 4193 4393 4207 4407
rect 3993 4373 4007 4387
rect 4033 4353 4047 4367
rect 4093 4353 4107 4367
rect 4113 4332 4127 4346
rect 4013 4293 4027 4307
rect 3973 4273 3987 4287
rect 4013 4272 4027 4286
rect 3913 4253 3927 4267
rect 3953 4213 3967 4227
rect 3893 4113 3907 4127
rect 3873 4073 3887 4087
rect 3873 3973 3887 3987
rect 3853 3913 3867 3927
rect 3833 3873 3847 3887
rect 3793 3814 3807 3828
rect 3833 3814 3847 3828
rect 3973 4173 3987 4187
rect 3993 4153 4007 4167
rect 3973 4053 3987 4067
rect 4073 4293 4087 4307
rect 4093 4153 4107 4167
rect 4073 4113 4087 4127
rect 4053 4093 4067 4107
rect 4073 4053 4087 4067
rect 3993 4033 4007 4047
rect 4053 4033 4067 4047
rect 4533 4993 4547 5007
rect 4573 4993 4587 5007
rect 4493 4973 4507 4987
rect 4633 5093 4647 5107
rect 4693 5153 4707 5167
rect 4733 5293 4747 5307
rect 4733 5233 4747 5247
rect 4873 5273 4887 5287
rect 4893 5273 4907 5287
rect 4853 5193 4867 5207
rect 4753 5153 4767 5167
rect 4793 5153 4807 5167
rect 4733 5093 4747 5107
rect 4793 5113 4807 5127
rect 4713 5073 4727 5087
rect 4753 5073 4767 5087
rect 4913 5153 4927 5167
rect 4853 5073 4867 5087
rect 5453 5393 5467 5407
rect 5353 5373 5367 5387
rect 5413 5374 5427 5388
rect 5513 5393 5527 5407
rect 5553 5374 5567 5388
rect 5613 5373 5627 5387
rect 4933 5073 4947 5087
rect 4593 4913 4607 4927
rect 4333 4854 4347 4868
rect 4553 4854 4567 4868
rect 4693 5032 4707 5046
rect 4673 5013 4687 5027
rect 4653 4973 4667 4987
rect 4653 4952 4667 4966
rect 4773 5032 4787 5046
rect 4853 5033 4867 5047
rect 4893 5031 4907 5045
rect 4793 4973 4807 4987
rect 4733 4953 4747 4967
rect 4673 4893 4687 4907
rect 4473 4812 4487 4826
rect 4533 4812 4547 4826
rect 4333 4773 4347 4787
rect 4413 4773 4427 4787
rect 4313 4753 4327 4767
rect 4353 4753 4367 4767
rect 4393 4713 4407 4727
rect 4353 4673 4367 4687
rect 4393 4673 4407 4687
rect 4533 4753 4547 4767
rect 4613 4773 4627 4787
rect 4593 4733 4607 4747
rect 4713 4854 4727 4868
rect 4773 4853 4787 4867
rect 4433 4713 4447 4727
rect 4633 4713 4647 4727
rect 4413 4613 4427 4627
rect 4353 4554 4367 4568
rect 4393 4554 4407 4568
rect 4293 4453 4307 4467
rect 4313 4413 4327 4427
rect 4373 4473 4387 4487
rect 4373 4433 4387 4447
rect 4293 4353 4307 4367
rect 4333 4353 4347 4367
rect 4193 4273 4207 4287
rect 4213 4253 4227 4267
rect 4193 4153 4207 4167
rect 4133 4113 4147 4127
rect 4733 4812 4747 4826
rect 4753 4733 4767 4747
rect 4693 4693 4707 4707
rect 4533 4613 4547 4627
rect 4473 4553 4487 4567
rect 4653 4553 4667 4567
rect 4693 4553 4707 4567
rect 4473 4492 4487 4506
rect 4433 4353 4447 4367
rect 4633 4513 4647 4527
rect 4613 4413 4627 4427
rect 4673 4473 4687 4487
rect 4913 5013 4927 5027
rect 4833 4855 4847 4869
rect 5113 5233 5127 5247
rect 5233 5313 5247 5327
rect 5173 5253 5187 5267
rect 5153 5153 5167 5167
rect 4973 5093 4987 5107
rect 5033 5093 5047 5107
rect 4993 5073 5007 5087
rect 5093 5073 5107 5087
rect 5133 5073 5147 5087
rect 5233 5113 5247 5127
rect 5053 5031 5067 5045
rect 4953 5013 4967 5027
rect 5013 5013 5027 5027
rect 5113 5033 5127 5047
rect 4993 4993 5007 5007
rect 5093 4993 5107 5007
rect 4933 4973 4947 4987
rect 4933 4913 4947 4927
rect 4953 4893 4967 4907
rect 4912 4853 4926 4867
rect 4933 4853 4947 4867
rect 5053 4893 5067 4907
rect 4993 4854 5007 4868
rect 4793 4812 4807 4826
rect 4833 4813 4847 4827
rect 4813 4793 4827 4807
rect 4893 4813 4907 4827
rect 4973 4812 4987 4826
rect 4853 4773 4867 4787
rect 4973 4773 4987 4787
rect 5153 5031 5167 5045
rect 5193 5031 5207 5045
rect 5153 4893 5167 4907
rect 5113 4855 5127 4869
rect 5333 5332 5347 5346
rect 5393 5332 5407 5346
rect 5433 5332 5447 5346
rect 5533 5332 5547 5346
rect 5573 5253 5587 5267
rect 5353 5173 5367 5187
rect 5513 5173 5527 5187
rect 5413 5133 5427 5147
rect 5493 5133 5507 5147
rect 5333 5113 5347 5127
rect 5353 5093 5367 5107
rect 5292 5073 5306 5087
rect 5313 5072 5327 5086
rect 5453 5113 5467 5127
rect 5473 5073 5487 5087
rect 5253 4993 5267 5007
rect 5233 4873 5247 4887
rect 5213 4853 5227 4867
rect 5333 4993 5347 5007
rect 5533 5073 5547 5087
rect 5753 5113 5767 5127
rect 5613 5073 5627 5087
rect 5693 5074 5707 5088
rect 5513 4993 5527 5007
rect 5553 4993 5567 5007
rect 5293 4873 5307 4887
rect 5333 4893 5347 4907
rect 5433 4893 5447 4907
rect 5313 4853 5327 4867
rect 5193 4833 5207 4847
rect 5093 4813 5107 4827
rect 5153 4813 5167 4827
rect 5273 4813 5287 4827
rect 5133 4793 5147 4807
rect 5053 4733 5067 4747
rect 5353 4853 5367 4867
rect 5413 4854 5427 4868
rect 5493 4933 5507 4947
rect 5473 4913 5487 4927
rect 5493 4873 5507 4887
rect 5473 4853 5487 4867
rect 5333 4713 5347 4727
rect 5013 4693 5027 4707
rect 5153 4693 5167 4707
rect 5333 4692 5347 4706
rect 5293 4653 5307 4667
rect 4812 4633 4826 4647
rect 4833 4633 4847 4647
rect 5133 4633 5147 4647
rect 4773 4593 4787 4607
rect 4793 4573 4807 4587
rect 4773 4553 4787 4567
rect 4953 4593 4967 4607
rect 4913 4573 4927 4587
rect 4753 4493 4767 4507
rect 4793 4493 4807 4507
rect 4753 4453 4767 4467
rect 4573 4335 4587 4349
rect 4713 4393 4727 4407
rect 4413 4313 4427 4327
rect 4373 4273 4387 4287
rect 4353 4233 4367 4247
rect 4333 4153 4347 4167
rect 4153 4053 4167 4067
rect 4133 4033 4147 4047
rect 4193 4034 4207 4048
rect 4253 4034 4267 4048
rect 4293 4034 4307 4048
rect 3973 4013 3987 4027
rect 3913 3933 3927 3947
rect 3953 3933 3967 3947
rect 3973 3893 3987 3907
rect 3953 3873 3967 3887
rect 3913 3853 3927 3867
rect 3973 3853 3987 3867
rect 4093 3993 4107 4007
rect 4033 3973 4047 3987
rect 4013 3953 4027 3967
rect 4093 3913 4107 3927
rect 4193 3953 4207 3967
rect 4033 3893 4047 3907
rect 4133 3893 4147 3907
rect 4013 3833 4027 3847
rect 4073 3873 4087 3887
rect 3493 3753 3507 3767
rect 3473 3733 3487 3747
rect 3413 3713 3427 3727
rect 3393 3673 3407 3687
rect 3393 3633 3407 3647
rect 3272 3573 3286 3587
rect 3293 3573 3307 3587
rect 3213 3393 3227 3407
rect 3193 3373 3207 3387
rect 3113 3293 3127 3307
rect 3273 3513 3287 3527
rect 3313 3513 3327 3527
rect 3453 3613 3467 3627
rect 3433 3514 3447 3528
rect 3353 3473 3367 3487
rect 3293 3433 3307 3447
rect 3273 3393 3287 3407
rect 3253 3353 3267 3367
rect 3373 3353 3387 3367
rect 3353 3333 3367 3347
rect 3153 3213 3167 3227
rect 3133 3193 3147 3207
rect 3113 3113 3127 3127
rect 3133 3093 3147 3107
rect 3173 3033 3187 3047
rect 3113 2994 3127 3008
rect 3273 3293 3287 3307
rect 3313 3295 3327 3309
rect 3293 3253 3307 3267
rect 3253 3173 3267 3187
rect 3353 3153 3367 3167
rect 3293 3093 3307 3107
rect 3353 3073 3367 3087
rect 3233 2994 3247 3008
rect 2973 2952 2987 2966
rect 3033 2952 3047 2966
rect 2853 2913 2867 2927
rect 3173 2933 3187 2947
rect 3093 2913 3107 2927
rect 2833 2853 2847 2867
rect 2913 2853 2927 2867
rect 3073 2853 3087 2867
rect 2773 2813 2787 2827
rect 2753 2793 2767 2807
rect 2672 2773 2686 2787
rect 2693 2774 2707 2788
rect 2733 2774 2747 2788
rect 2653 2713 2667 2727
rect 2653 2692 2667 2706
rect 2653 2613 2667 2627
rect 2753 2732 2767 2746
rect 2873 2732 2887 2746
rect 2813 2693 2827 2707
rect 3113 2873 3127 2887
rect 3093 2833 3107 2847
rect 2933 2773 2947 2787
rect 2993 2774 3007 2788
rect 3053 2773 3067 2787
rect 3033 2753 3047 2767
rect 2933 2732 2947 2746
rect 3053 2733 3067 2747
rect 3093 2733 3107 2747
rect 3033 2713 3047 2727
rect 3133 2713 3147 2727
rect 2913 2653 2927 2667
rect 2713 2593 2727 2607
rect 2673 2493 2687 2507
rect 2753 2473 2767 2487
rect 2793 2473 2807 2487
rect 2993 2474 3007 2488
rect 3033 2473 3047 2487
rect 3093 2473 3107 2487
rect 3132 2473 3146 2487
rect 3153 2474 3167 2488
rect 3293 2952 3307 2966
rect 3453 3473 3467 3487
rect 3453 3433 3467 3447
rect 3453 3393 3467 3407
rect 3593 3772 3607 3786
rect 3633 3772 3647 3786
rect 3673 3773 3687 3787
rect 3733 3773 3747 3787
rect 3513 3733 3527 3747
rect 3553 3733 3567 3747
rect 3553 3673 3567 3687
rect 3813 3772 3827 3786
rect 3873 3772 3887 3786
rect 3933 3773 3947 3787
rect 3973 3773 3987 3787
rect 4033 3814 4047 3828
rect 3733 3713 3747 3727
rect 3713 3673 3727 3687
rect 3673 3653 3687 3667
rect 3853 3653 3867 3667
rect 3493 3633 3507 3647
rect 3553 3633 3567 3647
rect 3533 3613 3547 3627
rect 3653 3613 3667 3627
rect 3513 3573 3527 3587
rect 3553 3553 3567 3567
rect 3533 3513 3547 3527
rect 3593 3514 3607 3528
rect 3733 3593 3747 3607
rect 3693 3514 3707 3528
rect 3813 3514 3827 3528
rect 3613 3493 3627 3507
rect 3533 3471 3547 3485
rect 3493 3373 3507 3387
rect 3473 3313 3487 3327
rect 3593 3452 3607 3466
rect 3553 3333 3567 3347
rect 3513 3293 3527 3307
rect 3613 3393 3627 3407
rect 3693 3413 3707 3427
rect 3673 3393 3687 3407
rect 3653 3313 3667 3327
rect 3633 3293 3647 3307
rect 3433 3252 3447 3266
rect 3453 3233 3467 3247
rect 3393 3213 3407 3227
rect 3453 3193 3467 3207
rect 3433 3173 3447 3187
rect 3373 3013 3387 3027
rect 3512 3253 3526 3267
rect 3533 3253 3547 3267
rect 3673 3294 3687 3308
rect 3833 3473 3847 3487
rect 3733 3453 3747 3467
rect 3753 3393 3767 3407
rect 3913 3713 3927 3727
rect 3933 3693 3947 3707
rect 3913 3673 3927 3687
rect 3953 3633 3967 3647
rect 3873 3613 3887 3627
rect 3873 3573 3887 3587
rect 3853 3413 3867 3427
rect 3713 3333 3727 3347
rect 3513 3213 3527 3227
rect 3573 3252 3587 3266
rect 3653 3252 3667 3266
rect 3732 3294 3746 3308
rect 3793 3373 3807 3387
rect 3833 3373 3847 3387
rect 3753 3293 3767 3307
rect 3953 3533 3967 3547
rect 3933 3472 3947 3486
rect 3993 3772 4007 3786
rect 4053 3772 4067 3786
rect 4093 3772 4107 3786
rect 3993 3733 4007 3747
rect 3973 3453 3987 3467
rect 3893 3393 3907 3407
rect 3873 3373 3887 3387
rect 3873 3352 3887 3366
rect 3832 3294 3846 3308
rect 3853 3294 3867 3308
rect 3613 3233 3627 3247
rect 3673 3233 3687 3247
rect 3593 3213 3607 3227
rect 3473 3153 3487 3167
rect 3533 3153 3547 3167
rect 3553 3073 3567 3087
rect 3433 2994 3447 3008
rect 3493 2993 3507 3007
rect 3353 2952 3367 2966
rect 3453 2952 3467 2966
rect 3413 2913 3427 2927
rect 3333 2873 3347 2887
rect 3493 2951 3507 2965
rect 3533 2951 3547 2965
rect 3633 3153 3647 3167
rect 3693 3073 3707 3087
rect 3673 3053 3687 3067
rect 3813 3233 3827 3247
rect 3853 3193 3867 3207
rect 4033 3673 4047 3687
rect 4273 3973 4287 3987
rect 4233 3893 4247 3907
rect 4313 3834 4327 3848
rect 4353 4034 4367 4048
rect 4573 4293 4587 4307
rect 4453 4273 4467 4287
rect 4413 4233 4427 4247
rect 4453 4213 4467 4227
rect 4433 4113 4447 4127
rect 4393 4034 4407 4048
rect 4593 4213 4607 4227
rect 4713 4335 4727 4349
rect 4733 4233 4747 4247
rect 4693 4213 4707 4227
rect 4533 4113 4547 4127
rect 4613 4113 4627 4127
rect 4653 4113 4667 4127
rect 4753 4113 4767 4127
rect 4493 4073 4507 4087
rect 4493 4033 4507 4047
rect 4573 4073 4587 4087
rect 4413 3992 4427 4006
rect 4373 3973 4387 3987
rect 4493 3993 4507 4007
rect 4453 3953 4467 3967
rect 4393 3913 4407 3927
rect 4353 3873 4367 3887
rect 4433 3873 4447 3887
rect 4312 3813 4326 3827
rect 4333 3813 4347 3827
rect 4393 3812 4407 3826
rect 4513 3953 4527 3967
rect 4653 4053 4667 4067
rect 4693 4033 4707 4047
rect 4813 4473 4827 4487
rect 4993 4554 5007 4568
rect 5093 4554 5107 4568
rect 5233 4554 5247 4568
rect 5473 4813 5487 4827
rect 5433 4793 5447 4807
rect 5393 4693 5407 4707
rect 5413 4653 5427 4667
rect 5373 4553 5387 4567
rect 5533 4933 5547 4947
rect 5513 4853 5527 4867
rect 5613 5033 5627 5047
rect 5653 5033 5667 5047
rect 5593 4913 5607 4927
rect 5573 4873 5587 4887
rect 5613 4853 5627 4867
rect 5673 4873 5687 4887
rect 5693 4854 5707 4868
rect 5572 4813 5586 4827
rect 5593 4813 5607 4827
rect 5633 4813 5647 4827
rect 5493 4793 5507 4807
rect 5513 4713 5527 4727
rect 4913 4433 4927 4447
rect 5053 4493 5067 4507
rect 5013 4453 5027 4467
rect 4853 4373 4867 4387
rect 4952 4373 4966 4387
rect 4973 4373 4987 4387
rect 5013 4373 5027 4387
rect 4873 4334 4887 4348
rect 4993 4335 5007 4349
rect 5113 4493 5127 4507
rect 5073 4453 5087 4467
rect 5113 4453 5127 4467
rect 5093 4393 5107 4407
rect 5033 4333 5047 4347
rect 5053 4333 5067 4347
rect 5293 4512 5307 4526
rect 5353 4512 5367 4526
rect 5393 4513 5407 4527
rect 5233 4453 5247 4467
rect 5213 4433 5227 4447
rect 5153 4393 5167 4407
rect 5113 4353 5127 4367
rect 5133 4335 5147 4349
rect 5173 4333 5187 4347
rect 5313 4413 5327 4427
rect 5293 4333 5307 4347
rect 4813 4313 4827 4327
rect 4813 4253 4827 4267
rect 4973 4293 4987 4307
rect 5013 4293 5027 4307
rect 4933 4253 4947 4267
rect 5053 4293 5067 4307
rect 5033 4233 5047 4247
rect 5093 4293 5107 4307
rect 4853 4213 4867 4227
rect 5073 4213 5087 4227
rect 5013 4133 5027 4147
rect 5173 4293 5187 4307
rect 5253 4293 5267 4307
rect 5253 4253 5267 4267
rect 5433 4473 5447 4487
rect 5473 4473 5487 4487
rect 5372 4353 5386 4367
rect 5393 4353 5407 4367
rect 5453 4353 5467 4367
rect 5553 4673 5567 4687
rect 5573 4553 5587 4567
rect 5733 4813 5747 4827
rect 5713 4793 5727 4807
rect 5673 4733 5687 4747
rect 5693 4553 5707 4567
rect 5533 4513 5547 4527
rect 5513 4393 5527 4407
rect 5513 4353 5527 4367
rect 5573 4511 5587 4525
rect 5613 4473 5627 4487
rect 5613 4413 5627 4427
rect 5573 4393 5587 4407
rect 5553 4353 5567 4367
rect 5533 4333 5547 4347
rect 5373 4293 5387 4307
rect 5233 4232 5247 4246
rect 5333 4233 5347 4247
rect 5133 4193 5147 4207
rect 5013 4093 5027 4107
rect 5093 4093 5107 4107
rect 4793 4053 4807 4067
rect 4953 4053 4967 4067
rect 4833 4033 4847 4047
rect 4893 4033 4907 4047
rect 5073 4053 5087 4067
rect 4673 3991 4687 4005
rect 4573 3973 4587 3987
rect 4613 3973 4627 3987
rect 4553 3833 4567 3847
rect 4513 3813 4527 3827
rect 4593 3933 4607 3947
rect 4633 3933 4647 3947
rect 4753 3991 4767 4005
rect 4813 3973 4827 3987
rect 4713 3893 4727 3907
rect 4753 3893 4767 3907
rect 4853 3893 4867 3907
rect 4613 3873 4627 3887
rect 4793 3853 4807 3867
rect 4613 3833 4627 3847
rect 4753 3833 4767 3847
rect 4153 3792 4167 3806
rect 4133 3733 4147 3747
rect 4053 3653 4067 3667
rect 4253 3773 4267 3787
rect 4333 3773 4347 3787
rect 4253 3733 4267 3747
rect 4293 3733 4307 3747
rect 4192 3713 4206 3727
rect 4213 3713 4227 3727
rect 4173 3633 4187 3647
rect 4233 3693 4247 3707
rect 4213 3673 4227 3687
rect 4033 3613 4047 3627
rect 4073 3613 4087 3627
rect 4153 3613 4167 3627
rect 4193 3613 4207 3627
rect 4033 3533 4047 3547
rect 4213 3593 4227 3607
rect 4073 3513 4087 3527
rect 4113 3514 4127 3528
rect 4033 3453 4047 3467
rect 4053 3393 4067 3407
rect 4033 3373 4047 3387
rect 3993 3353 4007 3367
rect 4153 3373 4167 3387
rect 4213 3373 4227 3387
rect 4093 3333 4107 3347
rect 3973 3313 3987 3327
rect 4013 3313 4027 3327
rect 4053 3314 4067 3328
rect 3933 3294 3947 3308
rect 3893 3253 3907 3267
rect 3893 3213 3907 3227
rect 3873 3173 3887 3187
rect 3913 3173 3927 3187
rect 3813 3093 3827 3107
rect 3913 3073 3927 3087
rect 3893 3053 3907 3067
rect 3713 2994 3727 3008
rect 3753 2994 3767 3008
rect 3813 2994 3827 3008
rect 3913 3013 3927 3027
rect 3553 2933 3567 2947
rect 3593 2933 3607 2947
rect 3493 2853 3507 2867
rect 3453 2833 3467 2847
rect 3693 2952 3707 2966
rect 3773 2952 3787 2966
rect 3873 2952 3887 2966
rect 3933 2952 3947 2966
rect 3773 2813 3787 2827
rect 3933 2813 3947 2827
rect 3653 2775 3667 2789
rect 3713 2775 3727 2789
rect 3773 2773 3787 2787
rect 3813 2774 3827 2788
rect 4053 3293 4067 3307
rect 4073 3252 4087 3266
rect 4353 3753 4367 3767
rect 4513 3773 4527 3787
rect 4473 3753 4487 3767
rect 4433 3713 4447 3727
rect 4433 3653 4447 3667
rect 4413 3613 4427 3627
rect 4333 3512 4347 3526
rect 4373 3513 4387 3527
rect 4453 3533 4467 3547
rect 4433 3514 4447 3528
rect 4393 3471 4407 3485
rect 4353 3453 4367 3467
rect 4513 3633 4527 3647
rect 4653 3813 4667 3827
rect 4713 3814 4727 3828
rect 4593 3772 4607 3786
rect 4693 3772 4707 3786
rect 4733 3772 4747 3786
rect 4653 3733 4667 3747
rect 4893 3853 4907 3867
rect 4973 3893 4987 3907
rect 4933 3833 4947 3847
rect 5053 3913 5067 3927
rect 4993 3873 5007 3887
rect 4833 3772 4847 3786
rect 4793 3713 4807 3727
rect 4853 3673 4867 3687
rect 5013 3813 5027 3827
rect 5353 4173 5367 4187
rect 5153 4133 5167 4147
rect 5233 4133 5247 4147
rect 5133 3973 5147 3987
rect 5273 4093 5287 4107
rect 5193 4033 5207 4047
rect 5153 3953 5167 3967
rect 5173 3853 5187 3867
rect 5153 3833 5167 3847
rect 4953 3773 4967 3787
rect 5013 3773 5027 3787
rect 5053 3733 5067 3747
rect 5113 3733 5127 3747
rect 4993 3713 5007 3727
rect 4893 3633 4907 3647
rect 4853 3593 4867 3607
rect 4693 3533 4707 3547
rect 4513 3514 4527 3528
rect 4553 3514 4567 3528
rect 4592 3513 4606 3527
rect 4613 3514 4627 3528
rect 4653 3514 4667 3528
rect 4793 3533 4807 3547
rect 4533 3472 4547 3486
rect 4553 3453 4567 3467
rect 4473 3413 4487 3427
rect 4453 3393 4467 3407
rect 4513 3373 4527 3387
rect 4233 3333 4247 3347
rect 4213 3293 4227 3307
rect 4293 3293 4307 3307
rect 4373 3295 4387 3309
rect 4153 3213 4167 3227
rect 4013 3193 4027 3207
rect 4113 3193 4127 3207
rect 4253 3253 4267 3267
rect 4233 3213 4247 3227
rect 4213 3193 4227 3207
rect 4213 3113 4227 3127
rect 4193 3093 4207 3107
rect 4033 3033 4047 3047
rect 4573 3273 4587 3287
rect 4353 3253 4367 3267
rect 4393 3253 4407 3267
rect 4293 3173 4307 3187
rect 4493 3173 4507 3187
rect 4293 3113 4307 3127
rect 4233 3073 4247 3087
rect 4473 3073 4487 3087
rect 4293 3053 4307 3067
rect 4393 3033 4407 3047
rect 4033 2813 4047 2827
rect 4133 2913 4147 2927
rect 4073 2873 4087 2887
rect 4113 2873 4127 2887
rect 3353 2733 3367 2747
rect 3453 2733 3467 2747
rect 3213 2693 3227 2707
rect 3253 2693 3267 2707
rect 3233 2573 3247 2587
rect 2633 2353 2647 2367
rect 2813 2431 2827 2445
rect 2913 2433 2927 2447
rect 2753 2413 2767 2427
rect 2813 2373 2827 2387
rect 2713 2333 2727 2347
rect 2873 2333 2887 2347
rect 2613 2254 2627 2268
rect 2573 2233 2587 2247
rect 2393 2212 2407 2226
rect 2453 2213 2467 2227
rect 2373 1973 2387 1987
rect 2353 1953 2367 1967
rect 2413 1973 2427 1987
rect 2493 2212 2507 2226
rect 2593 2213 2607 2227
rect 2533 2193 2547 2207
rect 2573 2193 2587 2207
rect 2473 1993 2487 2007
rect 2453 1953 2467 1967
rect 2353 1913 2367 1927
rect 2393 1912 2407 1926
rect 2433 1912 2447 1926
rect 2433 1853 2447 1867
rect 2453 1753 2467 1767
rect 2273 1573 2287 1587
rect 2253 1553 2267 1567
rect 2233 1493 2247 1507
rect 2152 1433 2166 1447
rect 2173 1434 2187 1448
rect 2373 1733 2387 1747
rect 2413 1692 2427 1706
rect 2393 1573 2407 1587
rect 2353 1553 2367 1567
rect 2293 1513 2307 1527
rect 2373 1493 2387 1507
rect 2293 1473 2307 1487
rect 2273 1453 2287 1467
rect 2053 1333 2067 1347
rect 2033 1273 2047 1287
rect 2053 1233 2067 1247
rect 1973 1213 1987 1227
rect 2033 1214 2047 1228
rect 2073 1214 2087 1228
rect 2133 1392 2147 1406
rect 2273 1333 2287 1347
rect 2373 1433 2387 1447
rect 2413 1533 2427 1547
rect 2453 1533 2467 1547
rect 2693 2212 2707 2226
rect 2653 2133 2667 2147
rect 2673 2073 2687 2087
rect 2593 1993 2607 2007
rect 2513 1953 2527 1967
rect 2553 1953 2567 1967
rect 2593 1953 2607 1967
rect 2633 1953 2647 1967
rect 2693 1953 2707 1967
rect 2493 1773 2507 1787
rect 2532 1773 2546 1787
rect 2553 1773 2567 1787
rect 2493 1733 2507 1747
rect 2653 1911 2667 1925
rect 2593 1733 2607 1747
rect 2773 2293 2787 2307
rect 2853 2293 2867 2307
rect 2813 2254 2827 2268
rect 3033 2433 3047 2447
rect 2973 2413 2987 2427
rect 2913 2273 2927 2287
rect 2953 2273 2967 2287
rect 2873 2253 2887 2267
rect 2753 2212 2767 2226
rect 2832 2213 2846 2227
rect 2853 2213 2867 2227
rect 2793 2193 2807 2207
rect 2893 2193 2907 2207
rect 3133 2413 3147 2427
rect 3193 2474 3207 2488
rect 3393 2513 3407 2527
rect 3313 2493 3327 2507
rect 3373 2493 3387 2507
rect 3293 2473 3307 2487
rect 3353 2473 3367 2487
rect 3073 2373 3087 2387
rect 3153 2373 3167 2387
rect 3073 2212 3087 2226
rect 3033 2133 3047 2147
rect 2833 2073 2847 2087
rect 2793 1973 2807 1987
rect 2753 1954 2767 1968
rect 3153 2053 3167 2067
rect 2873 2013 2887 2027
rect 3073 2013 3087 2027
rect 2853 1993 2867 2007
rect 2833 1953 2847 1967
rect 2753 1893 2767 1907
rect 2813 1912 2827 1926
rect 2813 1891 2827 1905
rect 2773 1873 2787 1887
rect 2793 1773 2807 1787
rect 2513 1693 2527 1707
rect 2553 1693 2567 1707
rect 2633 1693 2647 1707
rect 2513 1533 2527 1547
rect 2613 1533 2627 1547
rect 2473 1453 2487 1467
rect 2493 1433 2507 1447
rect 2353 1392 2367 1406
rect 2493 1393 2507 1407
rect 2373 1333 2387 1347
rect 2173 1293 2187 1307
rect 2293 1293 2307 1307
rect 2353 1293 2367 1307
rect 2213 1273 2227 1287
rect 1873 1173 1887 1187
rect 1913 1173 1927 1187
rect 1953 1173 1967 1187
rect 1913 1133 1927 1147
rect 1873 1113 1887 1127
rect 1913 973 1927 987
rect 1753 933 1767 947
rect 1733 913 1747 927
rect 1793 933 1807 947
rect 1833 933 1847 947
rect 1913 933 1927 947
rect 1853 914 1867 928
rect 2013 1172 2027 1186
rect 1973 1093 1987 1107
rect 2093 1173 2107 1187
rect 2353 1214 2367 1228
rect 2133 1173 2147 1187
rect 2113 1153 2127 1167
rect 2073 1133 2087 1147
rect 2193 1172 2207 1186
rect 2313 1153 2327 1167
rect 2153 1093 2167 1107
rect 2233 1093 2247 1107
rect 2133 1073 2147 1087
rect 2233 1072 2247 1086
rect 2053 953 2067 967
rect 1953 933 1967 947
rect 1933 913 1947 927
rect 1733 873 1747 887
rect 1713 833 1727 847
rect 1673 813 1687 827
rect 1713 812 1727 826
rect 1593 773 1607 787
rect 1633 773 1647 787
rect 1573 733 1587 747
rect 1593 693 1607 707
rect 1573 673 1587 687
rect 1613 652 1627 666
rect 1773 853 1787 867
rect 1833 873 1847 887
rect 1933 873 1947 887
rect 1813 773 1827 787
rect 1813 733 1827 747
rect 1673 613 1687 627
rect 1573 513 1587 527
rect 1473 493 1487 507
rect 1553 493 1567 507
rect 1353 413 1367 427
rect 1373 393 1387 407
rect 1433 393 1447 407
rect 1313 352 1327 366
rect 1353 353 1367 367
rect 1253 313 1267 327
rect 1333 313 1347 327
rect 1233 193 1247 207
rect 713 132 727 146
rect 753 132 767 146
rect 853 133 867 147
rect 693 113 707 127
rect 813 113 827 127
rect 992 133 1006 147
rect 1013 133 1027 147
rect 1053 133 1067 147
rect 1193 132 1207 146
rect 1133 113 1147 127
rect 1313 174 1327 188
rect 1353 174 1367 188
rect 1793 652 1807 666
rect 2273 1033 2287 1047
rect 2313 1013 2327 1027
rect 2353 973 2367 987
rect 2333 953 2347 967
rect 2493 1313 2507 1327
rect 2613 1493 2627 1507
rect 2533 1453 2547 1467
rect 2593 1392 2607 1406
rect 2793 1733 2807 1747
rect 2693 1633 2707 1647
rect 2653 1613 2667 1627
rect 2713 1473 2727 1487
rect 2893 1973 2907 1987
rect 2873 1953 2887 1967
rect 2873 1913 2887 1927
rect 2853 1893 2867 1907
rect 2873 1873 2887 1887
rect 2933 1913 2947 1927
rect 2953 1893 2967 1907
rect 3013 1893 3027 1907
rect 2933 1853 2947 1867
rect 2913 1833 2927 1847
rect 3013 1833 3027 1847
rect 2853 1813 2867 1827
rect 2933 1773 2947 1787
rect 3013 1773 3027 1787
rect 3093 1773 3107 1787
rect 2853 1753 2867 1767
rect 2813 1673 2827 1687
rect 2873 1673 2887 1687
rect 2793 1493 2807 1507
rect 2733 1453 2747 1467
rect 2833 1473 2847 1487
rect 2793 1433 2807 1447
rect 2893 1653 2907 1667
rect 2973 1734 2987 1748
rect 3073 1734 3087 1748
rect 2993 1692 3007 1706
rect 3033 1692 3047 1706
rect 3073 1653 3087 1667
rect 2993 1633 3007 1647
rect 2893 1613 2907 1627
rect 2933 1613 2947 1627
rect 2973 1533 2987 1547
rect 2873 1453 2887 1467
rect 2653 1392 2667 1406
rect 2693 1392 2707 1406
rect 2733 1392 2747 1406
rect 2533 1333 2547 1347
rect 2553 1313 2567 1327
rect 2473 1253 2487 1267
rect 2513 1253 2527 1267
rect 2433 1214 2447 1228
rect 2413 1073 2427 1087
rect 2392 973 2406 987
rect 2413 973 2427 987
rect 2313 913 2327 927
rect 2033 872 2047 886
rect 2073 872 2087 886
rect 1953 853 1967 867
rect 2073 833 2087 847
rect 2053 813 2067 827
rect 2093 813 2107 827
rect 2133 813 2147 827
rect 1953 793 1967 807
rect 1893 773 1907 787
rect 1933 773 1947 787
rect 2053 773 2067 787
rect 1953 713 1967 727
rect 1973 694 1987 708
rect 1873 653 1887 667
rect 1913 653 1927 667
rect 2513 1214 2527 1228
rect 2633 1253 2647 1267
rect 2613 1214 2627 1228
rect 2533 1172 2547 1186
rect 2193 733 2207 747
rect 2353 873 2367 887
rect 2293 833 2307 847
rect 2273 773 2287 787
rect 2253 713 2267 727
rect 2333 753 2347 767
rect 1713 613 1727 627
rect 1833 613 1847 627
rect 1693 493 1707 507
rect 1593 473 1607 487
rect 1573 373 1587 387
rect 1413 351 1427 365
rect 1453 351 1467 365
rect 1513 352 1527 366
rect 1413 313 1427 327
rect 1633 433 1647 447
rect 1753 573 1767 587
rect 1753 533 1767 547
rect 1733 493 1747 507
rect 1733 433 1747 447
rect 1853 493 1867 507
rect 1813 453 1827 467
rect 1793 433 1807 447
rect 1753 393 1767 407
rect 1833 394 1847 408
rect 1733 352 1747 366
rect 1773 352 1787 366
rect 2053 652 2067 666
rect 2093 652 2107 666
rect 2153 613 2167 627
rect 2253 652 2267 666
rect 2253 613 2267 627
rect 2193 573 2207 587
rect 1913 553 1927 567
rect 2493 913 2507 927
rect 2532 914 2546 928
rect 2573 1153 2587 1167
rect 2613 1133 2627 1147
rect 2693 1353 2707 1367
rect 2853 1391 2867 1405
rect 2893 1353 2907 1367
rect 2813 1333 2827 1347
rect 2873 1333 2887 1347
rect 2813 1293 2827 1307
rect 2653 1213 2667 1227
rect 2693 1214 2707 1228
rect 2733 1214 2747 1228
rect 2793 1214 2807 1228
rect 2833 1214 2847 1228
rect 2673 1172 2687 1186
rect 2693 1133 2707 1147
rect 2633 1113 2647 1127
rect 2673 1093 2687 1107
rect 2593 1053 2607 1067
rect 2553 913 2567 927
rect 2673 973 2687 987
rect 2853 1173 2867 1187
rect 2813 1153 2827 1167
rect 2813 1013 2827 1027
rect 2933 1233 2947 1247
rect 3213 2432 3227 2446
rect 3253 2432 3267 2446
rect 3193 2393 3207 2407
rect 3413 2432 3427 2446
rect 3553 2733 3567 2747
rect 3693 2733 3707 2747
rect 3773 2733 3787 2747
rect 3753 2693 3767 2707
rect 3613 2573 3627 2587
rect 3533 2513 3547 2527
rect 3613 2474 3627 2488
rect 3653 2474 3667 2488
rect 3713 2474 3727 2488
rect 3753 2474 3767 2488
rect 3473 2393 3487 2407
rect 3753 2393 3767 2407
rect 3333 2373 3347 2387
rect 3253 2333 3267 2347
rect 3333 2333 3347 2347
rect 3273 2293 3287 2307
rect 3953 2732 3967 2746
rect 3853 2713 3867 2727
rect 4133 2853 4147 2867
rect 4113 2813 4127 2827
rect 3993 2693 4007 2707
rect 4033 2713 4047 2727
rect 4013 2633 4027 2647
rect 3993 2513 4007 2527
rect 3933 2474 3947 2488
rect 4193 2951 4207 2965
rect 4293 2994 4307 3008
rect 4393 2994 4407 3008
rect 4433 2994 4447 3008
rect 4313 2952 4327 2966
rect 4253 2933 4267 2947
rect 4413 2933 4427 2947
rect 4373 2913 4387 2927
rect 4473 2913 4487 2927
rect 4193 2813 4207 2827
rect 4353 2813 4367 2827
rect 4153 2794 4167 2808
rect 4153 2773 4167 2787
rect 4273 2774 4287 2788
rect 4333 2774 4347 2788
rect 4173 2732 4187 2746
rect 4333 2733 4347 2747
rect 4213 2713 4227 2727
rect 4313 2633 4327 2647
rect 4273 2573 4287 2587
rect 4073 2533 4087 2547
rect 4113 2533 4127 2547
rect 4053 2493 4067 2507
rect 3973 2473 3987 2487
rect 4033 2473 4047 2487
rect 4173 2513 4187 2527
rect 4133 2493 4147 2507
rect 3833 2432 3847 2446
rect 3913 2432 3927 2446
rect 4233 2473 4247 2487
rect 3773 2313 3787 2327
rect 3413 2273 3427 2287
rect 3273 2254 3287 2268
rect 3333 2254 3347 2268
rect 3373 2254 3387 2268
rect 3433 2253 3447 2267
rect 3513 2255 3527 2269
rect 3573 2254 3587 2268
rect 3393 2212 3407 2226
rect 3433 2212 3447 2226
rect 3493 2213 3507 2227
rect 3533 2213 3547 2227
rect 3453 2173 3467 2187
rect 3353 2153 3367 2167
rect 3433 2113 3447 2127
rect 3233 2073 3247 2087
rect 3193 1993 3207 2007
rect 3393 1993 3407 2007
rect 3193 1953 3207 1967
rect 3233 1953 3247 1967
rect 3273 1953 3287 1967
rect 3313 1953 3327 1967
rect 3193 1911 3207 1925
rect 3233 1911 3247 1925
rect 3233 1853 3247 1867
rect 3313 1813 3327 1827
rect 3173 1753 3187 1767
rect 3313 1753 3327 1767
rect 3153 1735 3167 1749
rect 3173 1673 3187 1687
rect 3133 1653 3147 1667
rect 3213 1653 3227 1667
rect 3273 1613 3287 1627
rect 3033 1434 3047 1448
rect 3333 1734 3347 1748
rect 3393 1734 3407 1748
rect 3553 2193 3567 2207
rect 3753 2212 3767 2226
rect 3693 2173 3707 2187
rect 3553 2053 3567 2067
rect 3533 2013 3547 2027
rect 3653 2033 3667 2047
rect 3573 2013 3587 2027
rect 3493 1973 3507 1987
rect 3633 1973 3647 1987
rect 3873 2254 3887 2268
rect 3933 2254 3947 2268
rect 3853 2212 3867 2226
rect 3933 2173 3947 2187
rect 3793 2073 3807 2087
rect 3833 1993 3847 2007
rect 3793 1973 3807 1987
rect 3653 1953 3667 1967
rect 3673 1953 3687 1967
rect 3773 1954 3787 1968
rect 3652 1911 3666 1925
rect 3713 1912 3727 1926
rect 3893 1954 3907 1968
rect 3813 1913 3827 1927
rect 3973 2431 3987 2445
rect 4013 2431 4027 2445
rect 4093 2431 4107 2445
rect 4133 2431 4147 2445
rect 4213 2431 4227 2445
rect 4053 2393 4067 2407
rect 4293 2513 4307 2527
rect 4173 2333 4187 2347
rect 4273 2333 4287 2347
rect 4013 2273 4027 2287
rect 3993 2212 4007 2226
rect 4053 2193 4067 2207
rect 4113 2173 4127 2187
rect 3953 2093 3967 2107
rect 4093 2093 4107 2107
rect 4033 2053 4047 2067
rect 3993 2033 4007 2047
rect 3953 1993 3967 2007
rect 3793 1873 3807 1887
rect 3713 1833 3727 1847
rect 3773 1833 3787 1847
rect 3713 1773 3727 1787
rect 3493 1735 3507 1749
rect 3533 1735 3547 1749
rect 3573 1735 3587 1749
rect 3733 1734 3747 1748
rect 3793 1734 3807 1748
rect 3953 1913 3967 1927
rect 4013 1912 4027 1926
rect 4053 1912 4067 1926
rect 4053 1873 4067 1887
rect 3993 1853 4007 1867
rect 3333 1673 3347 1687
rect 3333 1633 3347 1647
rect 3333 1573 3347 1587
rect 3153 1513 3167 1527
rect 3313 1513 3327 1527
rect 3133 1453 3147 1467
rect 2993 1233 3007 1247
rect 2713 953 2727 967
rect 2833 953 2847 967
rect 2673 914 2687 928
rect 2453 872 2467 886
rect 2373 813 2387 827
rect 2553 873 2567 887
rect 2493 833 2507 847
rect 2473 793 2487 807
rect 2373 713 2387 727
rect 2413 694 2427 708
rect 2453 694 2467 708
rect 2593 873 2607 887
rect 2593 833 2607 847
rect 2673 813 2687 827
rect 2573 793 2587 807
rect 2553 773 2567 787
rect 2513 733 2527 747
rect 2633 753 2647 767
rect 2693 773 2707 787
rect 2733 913 2747 927
rect 2733 813 2747 827
rect 2753 753 2767 767
rect 2813 753 2827 767
rect 2733 713 2747 727
rect 2353 633 2367 647
rect 2333 593 2347 607
rect 2493 653 2507 667
rect 2533 652 2547 666
rect 2613 653 2627 667
rect 2433 633 2447 647
rect 2513 593 2527 607
rect 2553 573 2567 587
rect 2393 553 2407 567
rect 2513 553 2527 567
rect 2373 513 2387 527
rect 1913 453 1927 467
rect 2013 453 2027 467
rect 2253 453 2267 467
rect 2373 453 2387 467
rect 1953 433 1967 447
rect 1993 433 2007 447
rect 1913 393 1927 407
rect 1933 351 1947 365
rect 1973 353 1987 367
rect 1873 333 1887 347
rect 1813 313 1827 327
rect 1853 313 1867 327
rect 1593 233 1607 247
rect 1453 193 1467 207
rect 1493 173 1507 187
rect 1553 174 1567 188
rect 1733 213 1747 227
rect 1673 175 1687 189
rect 1973 233 1987 247
rect 1873 193 1887 207
rect 1493 132 1507 146
rect 1533 132 1547 146
rect 1373 113 1387 127
rect 1433 113 1447 127
rect 1653 133 1667 147
rect 1793 133 1807 147
rect 1833 133 1847 147
rect 1933 174 1947 188
rect 2193 413 2207 427
rect 2233 413 2247 427
rect 2053 393 2067 407
rect 2093 393 2107 407
rect 2133 394 2147 408
rect 2173 394 2187 408
rect 2213 394 2227 408
rect 2333 413 2347 427
rect 2193 352 2207 366
rect 2013 293 2027 307
rect 2133 293 2147 307
rect 1993 213 2007 227
rect 1573 113 1587 127
rect 1873 132 1887 146
rect 1913 132 1927 146
rect 1693 113 1707 127
rect 1992 133 2006 147
rect 2653 513 2667 527
rect 2913 1093 2927 1107
rect 3093 1173 3107 1187
rect 3133 1173 3147 1187
rect 2993 1153 3007 1167
rect 3193 1453 3207 1467
rect 3533 1653 3547 1667
rect 3513 1633 3527 1647
rect 3433 1493 3447 1507
rect 3273 1433 3287 1447
rect 3333 1433 3347 1447
rect 3373 1433 3387 1447
rect 3413 1433 3427 1447
rect 3453 1433 3467 1447
rect 3173 1233 3187 1247
rect 3153 1153 3167 1167
rect 3133 1113 3147 1127
rect 3193 1173 3207 1187
rect 3333 1373 3347 1387
rect 3613 1692 3627 1706
rect 3713 1692 3727 1706
rect 3673 1653 3687 1667
rect 3633 1593 3647 1607
rect 3553 1513 3567 1527
rect 3593 1434 3607 1448
rect 3733 1593 3747 1607
rect 3993 1734 4007 1748
rect 4033 1734 4047 1748
rect 3873 1633 3887 1647
rect 3833 1533 3847 1547
rect 3713 1493 3727 1507
rect 3633 1433 3647 1447
rect 3673 1433 3687 1447
rect 3733 1434 3747 1448
rect 3793 1434 3807 1448
rect 3853 1434 3867 1448
rect 3933 1693 3947 1707
rect 4013 1673 4027 1687
rect 4013 1633 4027 1647
rect 4053 1633 4067 1647
rect 3893 1593 3907 1607
rect 3913 1533 3927 1547
rect 3473 1391 3487 1405
rect 3533 1393 3547 1407
rect 3433 1373 3447 1387
rect 3613 1392 3627 1406
rect 3653 1393 3667 1407
rect 3573 1373 3587 1387
rect 3373 1333 3387 1347
rect 3633 1273 3647 1287
rect 3373 1215 3387 1229
rect 3533 1213 3547 1227
rect 3273 1172 3287 1186
rect 3233 1093 3247 1107
rect 3193 1053 3207 1067
rect 3173 993 3187 1007
rect 2953 973 2967 987
rect 2973 933 2987 947
rect 3193 933 3207 947
rect 2893 913 2907 927
rect 2933 913 2947 927
rect 3033 914 3047 928
rect 3073 914 3087 928
rect 3273 933 3287 947
rect 3393 1173 3407 1187
rect 3353 1093 3367 1107
rect 3433 1172 3447 1186
rect 3733 1391 3747 1405
rect 3693 1373 3707 1387
rect 3693 1333 3707 1347
rect 3733 1333 3747 1347
rect 3693 1273 3707 1287
rect 3793 1273 3807 1287
rect 3853 1273 3867 1287
rect 3733 1214 3747 1228
rect 3853 1214 3867 1228
rect 3653 1153 3667 1167
rect 3693 1153 3707 1167
rect 3413 1033 3427 1047
rect 3553 1033 3567 1047
rect 3393 953 3407 967
rect 3373 933 3387 947
rect 2873 873 2887 887
rect 2853 793 2867 807
rect 3033 813 3047 827
rect 2993 793 3007 807
rect 2873 733 2887 747
rect 2913 733 2927 747
rect 2793 695 2807 709
rect 2833 695 2847 709
rect 2933 713 2947 727
rect 2973 713 2987 727
rect 2753 653 2767 667
rect 2813 653 2827 667
rect 2933 652 2947 666
rect 2973 633 2987 647
rect 2973 612 2987 626
rect 2773 593 2787 607
rect 2893 593 2907 607
rect 2733 453 2747 467
rect 2553 433 2567 447
rect 2913 433 2927 447
rect 2533 393 2547 407
rect 2573 393 2587 407
rect 2633 393 2647 407
rect 2393 373 2407 387
rect 2453 352 2467 366
rect 2393 313 2407 327
rect 2373 273 2387 287
rect 2453 273 2467 287
rect 2233 253 2247 267
rect 2433 253 2447 267
rect 2193 174 2207 188
rect 2273 174 2287 188
rect 2373 174 2387 188
rect 2433 153 2447 167
rect 2593 351 2607 365
rect 2553 193 2567 207
rect 2773 392 2787 406
rect 2813 394 2827 408
rect 2693 333 2707 347
rect 2753 353 2767 367
rect 2733 333 2747 347
rect 3093 873 3107 887
rect 3153 853 3167 867
rect 3093 833 3107 847
rect 3073 753 3087 767
rect 3193 793 3207 807
rect 3093 713 3107 727
rect 3193 693 3207 707
rect 3313 913 3327 927
rect 3453 993 3467 1007
rect 3553 973 3567 987
rect 3473 953 3487 967
rect 3533 953 3547 967
rect 3573 953 3587 967
rect 3673 953 3687 967
rect 3453 913 3467 927
rect 3533 914 3547 928
rect 3573 914 3587 928
rect 3233 873 3247 887
rect 3053 652 3067 666
rect 3173 652 3187 666
rect 3213 652 3227 666
rect 3033 633 3047 647
rect 3073 633 3087 647
rect 3113 633 3127 647
rect 3093 533 3107 547
rect 3053 433 3067 447
rect 2993 393 3007 407
rect 3353 872 3367 886
rect 3293 853 3307 867
rect 3453 873 3467 887
rect 3393 853 3407 867
rect 3433 853 3447 867
rect 3253 833 3267 847
rect 3293 773 3307 787
rect 3293 713 3307 727
rect 3433 693 3447 707
rect 3353 652 3367 666
rect 3433 653 3447 667
rect 3413 633 3427 647
rect 3433 613 3447 627
rect 3413 553 3427 567
rect 3253 533 3267 547
rect 3293 533 3307 547
rect 3233 473 3247 487
rect 3193 453 3207 467
rect 3193 394 3207 408
rect 2833 352 2847 366
rect 2773 313 2787 327
rect 2633 273 2647 287
rect 2713 273 2727 287
rect 2693 233 2707 247
rect 1353 93 1367 107
rect 1553 93 1567 107
rect 1593 93 1607 107
rect 1653 93 1667 107
rect 1953 93 1967 107
rect 2013 132 2027 146
rect 2133 132 2147 146
rect 2353 133 2367 147
rect 2293 93 2307 107
rect 193 73 207 87
rect 413 73 427 87
rect 1093 73 1107 87
rect 1233 73 1247 87
rect 1993 73 2007 87
rect 2073 73 2087 87
rect 2453 133 2467 147
rect 2493 132 2507 146
rect 2413 93 2427 107
rect 2493 93 2507 107
rect 2393 53 2407 67
rect 2653 174 2667 188
rect 2753 233 2767 247
rect 2973 351 2987 365
rect 2953 293 2967 307
rect 2933 273 2947 287
rect 2993 293 3007 307
rect 2853 213 2867 227
rect 2993 213 3007 227
rect 2773 173 2787 187
rect 2813 174 2827 188
rect 3033 351 3047 365
rect 3113 351 3127 365
rect 3153 313 3167 327
rect 3033 273 3047 287
rect 3073 273 3087 287
rect 3013 173 3027 187
rect 2633 132 2647 146
rect 2693 132 2707 146
rect 2873 132 2887 146
rect 2933 132 2947 146
rect 3053 253 3067 267
rect 2833 113 2847 127
rect 2593 93 2607 107
rect 3113 193 3127 207
rect 3293 473 3307 487
rect 3373 393 3387 407
rect 3473 773 3487 787
rect 3673 913 3687 927
rect 3653 872 3667 886
rect 3653 793 3667 807
rect 3633 753 3647 767
rect 3533 694 3547 708
rect 3573 694 3587 708
rect 3653 713 3667 727
rect 3673 695 3687 709
rect 3793 1173 3807 1187
rect 3833 1113 3847 1127
rect 3713 1093 3727 1107
rect 3753 993 3767 1007
rect 3973 1392 3987 1406
rect 3933 1313 3947 1327
rect 3913 993 3927 1007
rect 3893 953 3907 967
rect 3793 914 3807 928
rect 4833 3513 4847 3527
rect 4613 3473 4627 3487
rect 4633 3453 4647 3467
rect 4713 3472 4727 3486
rect 4773 3471 4787 3485
rect 4673 3433 4687 3447
rect 4853 3471 4867 3485
rect 4633 3393 4647 3407
rect 4813 3393 4827 3407
rect 4613 3294 4627 3308
rect 4653 3373 4667 3387
rect 4773 3373 4787 3387
rect 4753 3353 4767 3367
rect 4733 3313 4747 3327
rect 4693 3294 4707 3308
rect 4613 3233 4627 3247
rect 4593 3113 4607 3127
rect 4533 3093 4547 3107
rect 4673 3093 4687 3107
rect 4633 3033 4647 3047
rect 4533 2994 4547 3008
rect 4573 2994 4587 3008
rect 4753 3293 4767 3307
rect 4793 3313 4807 3327
rect 5053 3673 5067 3687
rect 4913 3573 4927 3587
rect 5133 3533 5147 3547
rect 5073 3513 5087 3527
rect 5153 3513 5167 3527
rect 4933 3493 4947 3507
rect 5053 3493 5067 3507
rect 5113 3472 5127 3486
rect 5073 3453 5087 3467
rect 4953 3393 4967 3407
rect 4933 3353 4947 3367
rect 4813 3294 4827 3308
rect 4893 3294 4907 3308
rect 4973 3373 4987 3387
rect 5073 3373 5087 3387
rect 4953 3293 4967 3307
rect 4833 3253 4847 3267
rect 4953 3253 4967 3267
rect 4913 3233 4927 3247
rect 4953 3213 4967 3227
rect 4793 3113 4807 3127
rect 4933 3113 4947 3127
rect 4733 3013 4747 3027
rect 4993 3333 5007 3347
rect 5153 3293 5167 3307
rect 5213 3833 5227 3847
rect 5313 4053 5327 4067
rect 5413 4293 5427 4307
rect 5453 4293 5467 4307
rect 5393 4253 5407 4267
rect 5373 4073 5387 4087
rect 5493 4233 5507 4247
rect 5573 4333 5587 4347
rect 5713 4511 5727 4525
rect 5653 4335 5667 4349
rect 5693 4333 5707 4347
rect 5612 4293 5626 4307
rect 5633 4293 5647 4307
rect 5593 4253 5607 4267
rect 5593 4173 5607 4187
rect 5553 4133 5567 4147
rect 5493 4073 5507 4087
rect 5413 4053 5427 4067
rect 5453 4053 5467 4067
rect 5253 3814 5267 3828
rect 5333 3991 5347 4005
rect 5473 3993 5487 4007
rect 5453 3973 5467 3987
rect 5413 3953 5427 3967
rect 5353 3853 5367 3867
rect 5293 3813 5307 3827
rect 5413 3833 5427 3847
rect 5233 3773 5247 3787
rect 5213 3573 5227 3587
rect 5253 3733 5267 3747
rect 5273 3733 5287 3747
rect 5373 3773 5387 3787
rect 5373 3733 5387 3747
rect 5333 3713 5347 3727
rect 5293 3513 5307 3527
rect 5353 3514 5367 3528
rect 5553 4034 5567 4048
rect 5593 4033 5607 4047
rect 5553 3973 5567 3987
rect 5533 3893 5547 3907
rect 5533 3853 5547 3867
rect 5493 3833 5507 3847
rect 5473 3813 5487 3827
rect 5473 3773 5487 3787
rect 5513 3773 5527 3787
rect 5473 3613 5487 3627
rect 5593 3993 5607 4007
rect 5573 3953 5587 3967
rect 5693 4173 5707 4187
rect 5733 4293 5747 4307
rect 5713 4053 5727 4067
rect 5693 4034 5707 4048
rect 5693 3953 5707 3967
rect 5653 3933 5667 3947
rect 5613 3853 5627 3867
rect 5613 3815 5627 3829
rect 5673 3813 5687 3827
rect 5533 3573 5547 3587
rect 5573 3733 5587 3747
rect 5593 3653 5607 3667
rect 5573 3573 5587 3587
rect 5233 3333 5247 3347
rect 5233 3294 5247 3308
rect 5373 3473 5387 3487
rect 5333 3453 5347 3467
rect 5553 3513 5567 3527
rect 5433 3493 5447 3507
rect 5413 3453 5427 3467
rect 5393 3413 5407 3427
rect 5373 3353 5387 3367
rect 5193 3193 5207 3207
rect 5073 3153 5087 3167
rect 4993 3133 5007 3147
rect 4973 3073 4987 3087
rect 5113 3073 5127 3087
rect 4593 2952 4607 2966
rect 4633 2953 4647 2967
rect 4673 2951 4687 2965
rect 4573 2933 4587 2947
rect 4713 2913 4727 2927
rect 4973 3013 4987 3027
rect 5093 3013 5107 3027
rect 4833 2951 4847 2965
rect 4873 2953 4887 2967
rect 4573 2893 4587 2907
rect 4773 2893 4787 2907
rect 4553 2873 4567 2887
rect 4693 2813 4707 2827
rect 4553 2775 4567 2789
rect 4613 2773 4627 2787
rect 4653 2774 4667 2788
rect 4753 2773 4767 2787
rect 4533 2733 4547 2747
rect 4573 2733 4587 2747
rect 4493 2653 4507 2667
rect 4613 2693 4627 2707
rect 4713 2693 4727 2707
rect 4833 2774 4847 2788
rect 4913 2893 4927 2907
rect 5033 2952 5047 2966
rect 5093 2953 5107 2967
rect 5333 3295 5347 3309
rect 5453 3413 5467 3427
rect 5493 3295 5507 3309
rect 5533 3313 5547 3327
rect 5353 3253 5367 3267
rect 5393 3253 5407 3267
rect 5333 3193 5347 3207
rect 5273 3173 5287 3187
rect 5313 3173 5327 3187
rect 5273 3133 5287 3147
rect 5213 3013 5227 3027
rect 5313 2993 5327 3007
rect 5113 2913 5127 2927
rect 5153 2913 5167 2927
rect 5113 2833 5127 2847
rect 4953 2793 4967 2807
rect 5073 2793 5087 2807
rect 4913 2773 4927 2787
rect 4973 2775 4987 2789
rect 4813 2732 4827 2746
rect 4793 2712 4807 2726
rect 4773 2693 4787 2707
rect 4673 2653 4687 2667
rect 4753 2653 4767 2667
rect 4433 2573 4447 2587
rect 4473 2573 4487 2587
rect 4573 2573 4587 2587
rect 4413 2553 4427 2567
rect 4373 2513 4387 2527
rect 4333 2493 4347 2507
rect 4553 2553 4567 2567
rect 4433 2513 4447 2527
rect 4513 2474 4527 2488
rect 4353 2431 4367 2445
rect 4433 2433 4447 2447
rect 4393 2393 4407 2407
rect 4233 2273 4247 2287
rect 4273 2273 4287 2287
rect 4293 2252 4307 2266
rect 4353 2255 4367 2269
rect 4453 2254 4467 2268
rect 4273 2153 4287 2167
rect 4333 2213 4347 2227
rect 4373 2213 4387 2227
rect 4293 2113 4307 2127
rect 4433 2212 4447 2226
rect 4493 2212 4507 2226
rect 4693 2513 4707 2527
rect 4753 2474 4767 2488
rect 4573 2393 4587 2407
rect 4733 2433 4747 2447
rect 4653 2273 4667 2287
rect 4613 2255 4627 2269
rect 4853 2693 4867 2707
rect 5033 2733 5047 2747
rect 4993 2693 5007 2707
rect 4953 2673 4967 2687
rect 5093 2733 5107 2747
rect 5133 2733 5147 2747
rect 5053 2713 5067 2727
rect 5033 2653 5047 2667
rect 4913 2633 4927 2647
rect 4813 2474 4827 2488
rect 4933 2473 4947 2487
rect 4973 2474 4987 2488
rect 5213 2952 5227 2966
rect 5233 2933 5247 2947
rect 5213 2873 5227 2887
rect 5272 2913 5286 2927
rect 5293 2913 5307 2927
rect 5233 2853 5247 2867
rect 5273 2833 5287 2847
rect 5253 2793 5267 2807
rect 5273 2773 5287 2787
rect 5173 2733 5187 2747
rect 5152 2693 5166 2707
rect 5173 2693 5187 2707
rect 5253 2733 5267 2747
rect 5193 2653 5207 2667
rect 5113 2533 5127 2547
rect 5253 2533 5267 2547
rect 5173 2493 5187 2507
rect 5233 2474 5247 2488
rect 5273 2474 5287 2488
rect 4933 2432 4947 2446
rect 4873 2413 4887 2427
rect 5053 2432 5067 2446
rect 4993 2413 5007 2427
rect 4813 2393 4827 2407
rect 4993 2313 5007 2327
rect 5033 2293 5047 2307
rect 4893 2273 4907 2287
rect 4833 2253 4847 2267
rect 4953 2254 4967 2268
rect 4673 2233 4687 2247
rect 4573 2213 4587 2227
rect 4433 2173 4447 2187
rect 4533 2173 4547 2187
rect 4373 2153 4387 2167
rect 4273 2013 4287 2027
rect 4313 2013 4327 2027
rect 4173 1973 4187 1987
rect 4213 1973 4227 1987
rect 4133 1954 4147 1968
rect 4313 1973 4327 1987
rect 4173 1813 4187 1827
rect 4113 1734 4127 1748
rect 4173 1734 4187 1748
rect 4413 1873 4427 1887
rect 4413 1852 4427 1866
rect 4333 1813 4347 1827
rect 4153 1692 4167 1706
rect 4213 1692 4227 1706
rect 4313 1692 4327 1706
rect 4113 1653 4127 1667
rect 4273 1653 4287 1667
rect 4393 1734 4407 1748
rect 4533 2033 4547 2047
rect 4613 2013 4627 2027
rect 4473 1973 4487 1987
rect 4693 2212 4707 2226
rect 4733 2212 4747 2226
rect 4773 2212 4787 2226
rect 4833 2212 4847 2226
rect 4873 2212 4887 2226
rect 4673 2113 4687 2127
rect 4653 2033 4667 2047
rect 4653 1973 4667 1987
rect 4633 1953 4647 1967
rect 4673 1954 4687 1968
rect 5093 2393 5107 2407
rect 5273 2333 5287 2347
rect 5113 2313 5127 2327
rect 5073 2273 5087 2287
rect 5233 2293 5247 2307
rect 5153 2254 5167 2268
rect 5193 2254 5207 2268
rect 5333 2893 5347 2907
rect 5313 2873 5327 2887
rect 5353 2833 5367 2847
rect 5313 2773 5327 2787
rect 5473 3233 5487 3247
rect 5433 3133 5447 3147
rect 5493 3073 5507 3087
rect 5613 3613 5627 3627
rect 5613 3513 5627 3527
rect 5673 3713 5687 3727
rect 5753 4053 5767 4067
rect 5753 3953 5767 3967
rect 5753 3893 5767 3907
rect 5693 3553 5707 3567
rect 5733 3553 5747 3567
rect 5653 3513 5667 3527
rect 5713 3512 5727 3526
rect 5613 3453 5627 3467
rect 5673 3453 5687 3467
rect 5633 3413 5647 3427
rect 5613 3313 5627 3327
rect 5533 3193 5547 3207
rect 5453 2994 5467 3008
rect 5413 2933 5427 2947
rect 5373 2813 5387 2827
rect 5593 3233 5607 3247
rect 5513 3053 5527 3067
rect 5553 3053 5567 3067
rect 5713 3453 5727 3467
rect 5693 3393 5707 3407
rect 5693 3293 5707 3307
rect 5533 3013 5547 3027
rect 5673 3013 5687 3027
rect 5513 2913 5527 2927
rect 5533 2833 5547 2847
rect 5513 2813 5527 2827
rect 5433 2774 5447 2788
rect 5333 2713 5347 2727
rect 5433 2713 5447 2727
rect 5373 2693 5387 2707
rect 5413 2533 5427 2547
rect 5393 2473 5407 2487
rect 5353 2432 5367 2446
rect 5093 2212 5107 2226
rect 5153 2213 5167 2227
rect 4973 2193 4987 2207
rect 5033 2193 5047 2207
rect 4813 2113 4827 2127
rect 4713 1953 4727 1967
rect 4773 1954 4787 1968
rect 4933 2013 4947 2027
rect 4853 1993 4867 2007
rect 4653 1912 4667 1926
rect 4713 1912 4727 1926
rect 4453 1873 4467 1887
rect 4493 1793 4507 1807
rect 4533 1773 4547 1787
rect 4653 1773 4667 1787
rect 4493 1753 4507 1767
rect 4633 1734 4647 1748
rect 4673 1734 4687 1748
rect 4753 1912 4767 1926
rect 4773 1753 4787 1767
rect 4713 1733 4727 1747
rect 4813 1893 4827 1907
rect 4593 1693 4607 1707
rect 4433 1653 4447 1667
rect 4333 1553 4347 1567
rect 4093 1513 4107 1527
rect 4253 1513 4267 1527
rect 4073 1493 4087 1507
rect 4153 1453 4167 1467
rect 4213 1434 4227 1448
rect 4053 1392 4067 1406
rect 4053 1353 4067 1367
rect 4033 1333 4047 1347
rect 4013 1213 4027 1227
rect 3933 913 3947 927
rect 3773 872 3787 886
rect 3813 873 3827 887
rect 3813 793 3827 807
rect 3913 872 3927 886
rect 3833 773 3847 787
rect 3873 773 3887 787
rect 3733 753 3747 767
rect 3773 753 3787 767
rect 3813 753 3827 767
rect 3713 713 3727 727
rect 3633 653 3647 667
rect 3673 653 3687 667
rect 3473 633 3487 647
rect 3593 633 3607 647
rect 3653 593 3667 607
rect 3513 553 3527 567
rect 3613 553 3627 567
rect 3453 393 3467 407
rect 3513 394 3527 408
rect 3333 352 3347 366
rect 3373 352 3387 366
rect 3493 333 3507 347
rect 3473 313 3487 327
rect 3573 353 3587 367
rect 3493 293 3507 307
rect 3533 293 3547 307
rect 3293 273 3307 287
rect 3433 273 3447 287
rect 3253 253 3267 267
rect 3273 213 3287 227
rect 3173 193 3187 207
rect 3233 193 3247 207
rect 3213 132 3227 146
rect 3153 73 3167 87
rect 3473 253 3487 267
rect 3393 233 3407 247
rect 3293 173 3307 187
rect 3333 175 3347 189
rect 3273 53 3287 67
rect 2873 33 2887 47
rect 3053 33 3067 47
rect 2353 13 2367 27
rect 2393 13 2407 27
rect 2493 13 2507 27
rect 2553 13 2567 27
rect 3333 133 3347 147
rect 3313 113 3327 127
rect 3453 213 3467 227
rect 3473 193 3487 207
rect 3653 394 3667 408
rect 3693 533 3707 547
rect 3693 433 3707 447
rect 3973 1093 3987 1107
rect 4233 1393 4247 1407
rect 4093 1273 4107 1287
rect 4193 1273 4207 1287
rect 4093 1215 4107 1229
rect 4193 1215 4207 1229
rect 4453 1493 4467 1507
rect 4413 1433 4427 1447
rect 4393 1393 4407 1407
rect 4333 1373 4347 1387
rect 4373 1373 4387 1387
rect 4253 1333 4267 1347
rect 4373 1233 4387 1247
rect 4333 1214 4347 1228
rect 4433 1391 4447 1405
rect 4473 1393 4487 1407
rect 4393 1213 4407 1227
rect 4073 1173 4087 1187
rect 4153 1173 4167 1187
rect 4113 1133 4127 1147
rect 4033 993 4047 1007
rect 4093 993 4107 1007
rect 4053 953 4067 967
rect 3973 913 3987 927
rect 4013 933 4027 947
rect 3993 872 4007 886
rect 3973 853 3987 867
rect 3953 713 3967 727
rect 3833 693 3847 707
rect 3873 695 3887 709
rect 3933 693 3947 707
rect 4213 1173 4227 1187
rect 4353 1172 4367 1186
rect 4393 1173 4407 1187
rect 4273 1033 4287 1047
rect 4213 933 4227 947
rect 4313 953 4327 967
rect 4473 973 4487 987
rect 4453 953 4467 967
rect 4453 914 4467 928
rect 4173 853 4187 867
rect 4133 753 4147 767
rect 4053 733 4067 747
rect 4093 733 4107 747
rect 4033 693 4047 707
rect 3753 653 3767 667
rect 3813 653 3827 667
rect 3853 653 3867 667
rect 3753 593 3767 607
rect 3833 593 3847 607
rect 3893 593 3907 607
rect 4013 652 4027 666
rect 3933 553 3947 567
rect 3953 473 3967 487
rect 3993 473 4007 487
rect 3833 453 3847 467
rect 3853 433 3867 447
rect 3713 393 3727 407
rect 3793 394 3807 408
rect 3833 394 3847 408
rect 3613 333 3627 347
rect 3713 353 3727 367
rect 3593 313 3607 327
rect 3673 313 3687 327
rect 3853 352 3867 366
rect 3913 352 3927 366
rect 3833 293 3847 307
rect 3573 253 3587 267
rect 3713 253 3727 267
rect 3753 253 3767 267
rect 3593 213 3607 227
rect 3533 174 3547 188
rect 3433 132 3447 146
rect 3473 132 3487 146
rect 3513 133 3527 147
rect 3393 93 3407 107
rect 3453 93 3467 107
rect 3493 93 3507 107
rect 4033 433 4047 447
rect 4093 694 4107 708
rect 4073 653 4087 667
rect 4093 633 4107 647
rect 4073 613 4087 627
rect 4053 393 4067 407
rect 4153 613 4167 627
rect 4213 873 4227 887
rect 4233 853 4247 867
rect 4193 833 4207 847
rect 4193 733 4207 747
rect 4213 694 4227 708
rect 4192 633 4206 647
rect 4213 633 4227 647
rect 4193 593 4207 607
rect 4173 573 4187 587
rect 4153 553 4167 567
rect 4153 513 4167 527
rect 4193 473 4207 487
rect 4173 413 4187 427
rect 4093 393 4107 407
rect 4013 351 4027 365
rect 4073 353 4087 367
rect 4133 392 4147 406
rect 4193 393 4207 407
rect 4093 333 4107 347
rect 3953 233 3967 247
rect 3993 233 4007 247
rect 3873 193 3887 207
rect 3773 173 3787 187
rect 3833 175 3847 189
rect 3893 174 3907 188
rect 3953 174 3967 188
rect 3993 174 4007 188
rect 3593 93 3607 107
rect 3713 132 3727 146
rect 3753 132 3767 146
rect 3853 133 3867 147
rect 3973 132 3987 146
rect 4033 113 4047 127
rect 3893 73 3907 87
rect 4093 73 4107 87
rect 3653 53 3667 67
rect 4193 353 4207 367
rect 4153 273 4167 287
rect 4233 513 4247 527
rect 4333 833 4347 847
rect 4433 872 4447 886
rect 4473 873 4487 887
rect 4413 833 4427 847
rect 4393 753 4407 767
rect 4333 733 4347 747
rect 4313 694 4327 708
rect 4373 694 4387 708
rect 4513 1653 4527 1667
rect 4553 1434 4567 1448
rect 4653 1692 4667 1706
rect 4613 1633 4627 1647
rect 5053 2133 5067 2147
rect 5133 2133 5147 2147
rect 5013 2033 5027 2047
rect 5013 1973 5027 1987
rect 4973 1953 4987 1967
rect 5313 2254 5327 2268
rect 5273 2173 5287 2187
rect 5213 2093 5227 2107
rect 5313 2093 5327 2107
rect 5293 2053 5307 2067
rect 5293 1993 5307 2007
rect 5193 1973 5207 1987
rect 5273 1973 5287 1987
rect 5373 2113 5387 2127
rect 5353 2013 5367 2027
rect 5313 1953 5327 1967
rect 4853 1873 4867 1887
rect 4953 1912 4967 1926
rect 5033 1893 5047 1907
rect 5033 1853 5047 1867
rect 4913 1793 4927 1807
rect 5013 1753 5027 1767
rect 4853 1734 4867 1748
rect 4893 1734 4907 1748
rect 4973 1735 4987 1749
rect 5133 1912 5147 1926
rect 5173 1912 5187 1926
rect 5213 1893 5227 1907
rect 5073 1833 5087 1847
rect 5193 1833 5207 1847
rect 5173 1793 5187 1807
rect 5053 1734 5067 1748
rect 5093 1734 5107 1748
rect 5133 1734 5147 1748
rect 4753 1692 4767 1706
rect 4813 1693 4827 1707
rect 4733 1633 4747 1647
rect 4713 1453 4727 1467
rect 4913 1693 4927 1707
rect 4952 1693 4966 1707
rect 4973 1693 4987 1707
rect 4873 1633 4887 1647
rect 5113 1692 5127 1706
rect 5173 1693 5187 1707
rect 5253 1734 5267 1748
rect 5333 1913 5347 1927
rect 5433 2513 5447 2527
rect 5433 2473 5447 2487
rect 5493 2732 5507 2746
rect 5493 2553 5507 2567
rect 5593 2793 5607 2807
rect 5573 2774 5587 2788
rect 5653 2773 5667 2787
rect 5633 2733 5647 2747
rect 5613 2693 5627 2707
rect 5533 2633 5547 2647
rect 5593 2593 5607 2607
rect 5553 2513 5567 2527
rect 5513 2473 5527 2487
rect 5593 2473 5607 2487
rect 5433 2433 5447 2447
rect 5413 2413 5427 2427
rect 5573 2413 5587 2427
rect 5473 2333 5487 2347
rect 5533 2313 5547 2327
rect 5513 2293 5527 2307
rect 5473 2254 5487 2268
rect 5433 2213 5447 2227
rect 5453 2133 5467 2147
rect 5433 2113 5447 2127
rect 5433 2053 5447 2067
rect 5413 2013 5427 2027
rect 5393 1973 5407 1987
rect 5373 1953 5387 1967
rect 5453 1954 5467 1968
rect 5393 1912 5407 1926
rect 5413 1893 5427 1907
rect 5373 1873 5387 1887
rect 5353 1753 5367 1767
rect 5473 1913 5487 1927
rect 5433 1853 5447 1867
rect 5473 1813 5487 1827
rect 5573 2293 5587 2307
rect 5533 2254 5547 2268
rect 5673 2733 5687 2747
rect 5673 2693 5687 2707
rect 5693 2513 5707 2527
rect 5673 2313 5687 2327
rect 5653 2273 5667 2287
rect 5633 2253 5647 2267
rect 5733 2773 5747 2787
rect 5713 2473 5727 2487
rect 5693 2273 5707 2287
rect 5553 2173 5567 2187
rect 5613 2213 5627 2227
rect 5593 1993 5607 2007
rect 5693 2213 5707 2227
rect 5673 2193 5687 2207
rect 5653 2113 5667 2127
rect 5533 1912 5547 1926
rect 5513 1773 5527 1787
rect 5413 1733 5427 1747
rect 5513 1733 5527 1747
rect 5273 1692 5287 1706
rect 5313 1693 5327 1707
rect 5193 1673 5207 1687
rect 5233 1673 5247 1687
rect 5053 1653 5067 1667
rect 4973 1633 4987 1647
rect 5013 1593 5027 1607
rect 4933 1553 4947 1567
rect 4913 1533 4927 1547
rect 4653 1433 4667 1447
rect 4693 1433 4707 1447
rect 4733 1433 4747 1447
rect 4513 1393 4527 1407
rect 4533 1373 4547 1387
rect 4633 1393 4647 1407
rect 4613 1373 4627 1387
rect 4513 1293 4527 1307
rect 4573 1293 4587 1307
rect 4513 1213 4527 1227
rect 4533 1172 4547 1186
rect 5053 1553 5067 1567
rect 5013 1493 5027 1507
rect 4713 1391 4727 1405
rect 4933 1392 4947 1406
rect 4973 1392 4987 1406
rect 4653 1353 4667 1367
rect 4653 1273 4667 1287
rect 4713 1273 4727 1287
rect 4633 1133 4647 1147
rect 4673 1233 4687 1247
rect 4873 1253 4887 1267
rect 4853 1233 4867 1247
rect 4773 1213 4787 1227
rect 4833 1214 4847 1228
rect 4973 1253 4987 1267
rect 5013 1253 5027 1267
rect 5293 1613 5307 1627
rect 5273 1553 5287 1567
rect 5113 1533 5127 1547
rect 5273 1493 5287 1507
rect 5213 1434 5227 1448
rect 5133 1392 5147 1406
rect 5233 1392 5247 1406
rect 5193 1353 5207 1367
rect 5093 1313 5107 1327
rect 5073 1253 5087 1267
rect 5113 1253 5127 1267
rect 5173 1253 5187 1267
rect 4773 1172 4787 1186
rect 4733 1133 4747 1147
rect 4613 1093 4627 1107
rect 4653 1093 4667 1107
rect 4613 1053 4627 1067
rect 4593 1033 4607 1047
rect 4733 1033 4747 1047
rect 4513 973 4527 987
rect 4553 953 4567 967
rect 4513 913 4527 927
rect 4553 914 4567 928
rect 4513 873 4527 887
rect 4493 853 4507 867
rect 4473 793 4487 807
rect 4573 873 4587 887
rect 4553 853 4567 867
rect 4573 833 4587 847
rect 4533 793 4547 807
rect 4573 773 4587 787
rect 4553 753 4567 767
rect 4453 733 4467 747
rect 4513 733 4527 747
rect 4313 633 4327 647
rect 4393 652 4407 666
rect 4353 593 4367 607
rect 4293 513 4307 527
rect 4333 513 4347 527
rect 4253 473 4267 487
rect 4513 694 4527 708
rect 4653 973 4667 987
rect 4613 953 4627 967
rect 4613 913 4627 927
rect 4613 873 4627 887
rect 4593 713 4607 727
rect 4573 693 4587 707
rect 4693 873 4707 887
rect 4633 773 4647 787
rect 4653 733 4667 747
rect 4693 713 4707 727
rect 4813 1172 4827 1186
rect 4893 1173 4907 1187
rect 5053 1213 5067 1227
rect 5093 1213 5107 1227
rect 4853 1133 4867 1147
rect 4913 1133 4927 1147
rect 4913 1053 4927 1067
rect 4893 1013 4907 1027
rect 4793 914 4807 928
rect 4833 914 4847 928
rect 4813 873 4827 887
rect 4993 1172 5007 1186
rect 5073 1173 5087 1187
rect 4953 1153 4967 1167
rect 5393 1693 5407 1707
rect 5373 1653 5387 1667
rect 5313 1493 5327 1507
rect 5333 1434 5347 1448
rect 5353 1392 5367 1406
rect 5433 1692 5447 1706
rect 5473 1693 5487 1707
rect 5513 1693 5527 1707
rect 5493 1673 5507 1687
rect 5413 1653 5427 1667
rect 5473 1653 5487 1667
rect 5513 1613 5527 1627
rect 5613 1912 5627 1926
rect 5653 1773 5667 1787
rect 5613 1734 5627 1748
rect 5553 1673 5567 1687
rect 5533 1593 5547 1607
rect 5473 1533 5487 1547
rect 5513 1533 5527 1547
rect 5433 1493 5447 1507
rect 5413 1433 5427 1447
rect 5453 1391 5467 1405
rect 5393 1353 5407 1367
rect 5293 1313 5307 1327
rect 5433 1313 5447 1327
rect 5293 1253 5307 1267
rect 5213 1233 5227 1247
rect 5273 1233 5287 1247
rect 5193 1214 5207 1228
rect 5173 1153 5187 1167
rect 4973 1132 4987 1146
rect 5133 1133 5147 1147
rect 5253 1214 5267 1228
rect 5193 1113 5207 1127
rect 5153 1093 5167 1107
rect 5113 1013 5127 1027
rect 5013 933 5027 947
rect 5053 933 5067 947
rect 5153 914 5167 928
rect 5193 914 5207 928
rect 4933 853 4947 867
rect 4973 853 4987 867
rect 5013 853 5027 867
rect 5053 853 5067 867
rect 5093 853 5107 867
rect 4813 833 4827 847
rect 4473 613 4487 627
rect 4573 653 4587 667
rect 4533 553 4547 567
rect 4253 433 4267 447
rect 4393 433 4407 447
rect 4453 433 4467 447
rect 4533 433 4547 447
rect 5193 873 5207 887
rect 5053 793 5067 807
rect 5133 793 5147 807
rect 5073 733 5087 747
rect 5253 1153 5267 1167
rect 5273 1133 5287 1147
rect 5333 1133 5347 1147
rect 5753 2473 5767 2487
rect 5673 1734 5687 1748
rect 5733 1993 5747 2007
rect 5713 1533 5727 1547
rect 5673 1493 5687 1507
rect 5553 1453 5567 1467
rect 5653 1453 5667 1467
rect 5593 1434 5607 1448
rect 5713 1434 5727 1448
rect 5513 1293 5527 1307
rect 5513 1214 5527 1228
rect 5613 1392 5627 1406
rect 5693 1392 5707 1406
rect 5593 1293 5607 1307
rect 5453 1193 5467 1207
rect 5433 1153 5447 1167
rect 5393 1113 5407 1127
rect 5293 1073 5307 1087
rect 5273 1053 5287 1067
rect 5453 993 5467 1007
rect 5273 973 5287 987
rect 5253 933 5267 947
rect 5413 933 5427 947
rect 5313 914 5327 928
rect 5373 914 5387 928
rect 5533 933 5547 947
rect 5453 913 5467 927
rect 5273 871 5287 885
rect 5253 853 5267 867
rect 5293 853 5307 867
rect 5253 813 5267 827
rect 5173 713 5187 727
rect 5213 714 5227 728
rect 5053 693 5067 707
rect 5093 693 5107 707
rect 4593 553 4607 567
rect 4673 573 4687 587
rect 4633 513 4647 527
rect 4613 453 4627 467
rect 4653 453 4667 467
rect 4233 393 4247 407
rect 4313 393 4327 407
rect 4453 393 4467 407
rect 4493 394 4507 408
rect 4533 393 4547 407
rect 4233 353 4247 367
rect 4293 352 4307 366
rect 4253 333 4267 347
rect 4233 313 4247 327
rect 4293 313 4307 327
rect 4213 253 4227 267
rect 4213 174 4227 188
rect 4453 353 4467 367
rect 4453 313 4467 327
rect 4353 253 4367 267
rect 4413 174 4427 188
rect 4513 352 4527 366
rect 4513 174 4527 188
rect 4573 393 4587 407
rect 4793 653 4807 667
rect 5013 653 5027 667
rect 5053 653 5067 667
rect 5093 653 5107 667
rect 4893 573 4907 587
rect 4753 553 4767 567
rect 5073 633 5087 647
rect 5133 633 5147 647
rect 5053 573 5067 587
rect 5013 493 5027 507
rect 4793 453 4807 467
rect 4673 413 4687 427
rect 4633 313 4647 327
rect 4693 393 4707 407
rect 4753 393 4767 407
rect 5213 693 5227 707
rect 5433 873 5447 887
rect 5393 853 5407 867
rect 5373 813 5387 827
rect 5313 713 5327 727
rect 5193 653 5207 667
rect 5173 593 5187 607
rect 5113 533 5127 547
rect 5193 533 5207 547
rect 5073 433 5087 447
rect 5153 493 5167 507
rect 4873 394 4887 408
rect 4913 393 4927 407
rect 4953 393 4967 407
rect 5013 393 5027 407
rect 5053 393 5067 407
rect 5113 394 5127 408
rect 4693 313 4707 327
rect 4673 253 4687 267
rect 4773 351 4787 365
rect 4853 352 4867 366
rect 4873 253 4887 267
rect 4753 213 4767 227
rect 4793 213 4807 227
rect 4673 174 4687 188
rect 4733 174 4747 188
rect 4993 273 5007 287
rect 5093 352 5107 366
rect 5113 333 5127 347
rect 5093 273 5107 287
rect 4993 213 5007 227
rect 4933 174 4947 188
rect 4973 174 4987 188
rect 5273 593 5287 607
rect 5353 753 5367 767
rect 5333 693 5347 707
rect 5473 872 5487 886
rect 5593 1214 5607 1228
rect 5613 1073 5627 1087
rect 5653 953 5667 967
rect 5553 914 5567 928
rect 5593 914 5607 928
rect 5653 914 5667 928
rect 5673 873 5687 887
rect 5533 813 5547 827
rect 5353 653 5367 667
rect 5433 652 5447 666
rect 5573 652 5587 666
rect 5653 633 5667 647
rect 5433 573 5447 587
rect 5393 553 5407 567
rect 5493 553 5507 567
rect 5313 493 5327 507
rect 5393 493 5407 507
rect 5273 433 5287 447
rect 5173 393 5187 407
rect 5213 394 5227 408
rect 5333 394 5347 408
rect 5373 394 5387 408
rect 5113 213 5127 227
rect 5153 213 5167 227
rect 5233 333 5247 347
rect 5493 394 5507 408
rect 5553 394 5567 408
rect 5753 1913 5767 1927
rect 5733 993 5747 1007
rect 5713 833 5727 847
rect 5693 633 5707 647
rect 5673 433 5687 447
rect 5453 352 5467 366
rect 5393 333 5407 347
rect 5373 253 5387 267
rect 5453 253 5467 267
rect 5073 172 5087 186
rect 5133 174 5147 188
rect 5433 213 5447 227
rect 5193 173 5207 187
rect 5253 174 5267 188
rect 5333 175 5347 189
rect 5393 175 5407 189
rect 4433 132 4447 146
rect 4473 132 4487 146
rect 4533 132 4547 146
rect 4593 133 4607 147
rect 4653 132 4667 146
rect 4773 133 4787 147
rect 4813 133 4827 147
rect 4893 132 4907 146
rect 4933 133 4947 147
rect 4993 132 5007 146
rect 5053 133 5067 147
rect 4953 93 4967 107
rect 5153 132 5167 146
rect 5113 93 5127 107
rect 5533 352 5547 366
rect 5673 313 5687 327
rect 5633 273 5647 287
rect 5513 213 5527 227
rect 5533 193 5547 207
rect 5333 113 5347 127
rect 5293 93 5307 107
rect 5433 133 5447 147
rect 5473 133 5487 147
rect 5513 133 5527 147
rect 5493 113 5507 127
rect 5553 113 5567 127
rect 5393 93 5407 107
rect 5433 93 5447 107
rect 5593 93 5607 107
rect 5073 53 5087 67
rect 5233 53 5247 67
rect 5373 53 5387 67
<< metal3 >>
rect 327 5476 593 5484
rect 1567 5476 2033 5484
rect 2096 5476 2893 5484
rect 347 5456 613 5464
rect 767 5456 893 5464
rect 2096 5464 2104 5476
rect 2947 5476 3072 5484
rect 3107 5476 3185 5484
rect 1487 5456 2104 5464
rect 2407 5456 2853 5464
rect 3177 5464 3185 5476
rect 3447 5476 3772 5484
rect 4047 5476 4133 5484
rect 4227 5476 4573 5484
rect 3177 5456 3413 5464
rect 3467 5456 3733 5464
rect 4007 5456 4193 5464
rect 4207 5456 4593 5464
rect 1767 5436 2013 5444
rect 2647 5436 2932 5444
rect 3307 5436 3433 5444
rect 3947 5436 4053 5444
rect 4107 5436 4213 5444
rect 4396 5436 5333 5444
rect 227 5416 333 5424
rect 407 5416 573 5424
rect 1167 5416 1233 5424
rect 1407 5416 1553 5424
rect 1867 5416 2693 5424
rect 3027 5416 3273 5424
rect 3567 5416 3633 5424
rect 3807 5416 3873 5424
rect 4396 5424 4404 5436
rect 4087 5416 4404 5424
rect 4427 5416 4552 5424
rect 4587 5416 4653 5424
rect 667 5396 813 5404
rect 2047 5396 2073 5404
rect 2327 5396 2393 5404
rect 2907 5396 2953 5404
rect 3133 5396 3293 5404
rect 3133 5389 3147 5396
rect 3847 5393 3853 5407
rect 3927 5396 4053 5404
rect 4147 5396 4233 5404
rect 4416 5404 4424 5413
rect 4287 5396 4424 5404
rect 5047 5396 5453 5404
rect 5467 5396 5513 5404
rect 47 5376 73 5384
rect 136 5376 213 5384
rect 116 5347 124 5375
rect 136 5347 144 5376
rect 267 5378 293 5386
rect 507 5376 553 5384
rect 607 5376 753 5384
rect 856 5364 864 5374
rect 987 5376 1053 5384
rect 1247 5378 1293 5386
rect 656 5356 864 5364
rect 247 5336 273 5344
rect 327 5336 373 5344
rect 427 5336 473 5344
rect 567 5336 633 5344
rect 656 5344 664 5356
rect 1336 5347 1344 5375
rect 1487 5376 1584 5384
rect 1576 5364 1584 5376
rect 1607 5378 1652 5386
rect 1687 5376 1713 5384
rect 1936 5376 1973 5384
rect 1576 5360 1603 5364
rect 1576 5356 1607 5360
rect 1593 5347 1607 5356
rect 647 5336 664 5344
rect 756 5336 1013 5344
rect 756 5327 764 5336
rect 1606 5340 1607 5347
rect 1627 5336 1733 5344
rect 1856 5344 1864 5375
rect 1876 5360 1913 5364
rect 1747 5336 1864 5344
rect 1873 5356 1913 5360
rect 1873 5347 1887 5356
rect 1936 5364 1944 5376
rect 2027 5376 2093 5384
rect 2167 5376 2233 5384
rect 2247 5378 2293 5386
rect 2447 5378 2493 5386
rect 2996 5376 3013 5384
rect 1927 5356 1944 5364
rect 2596 5347 2604 5374
rect 2756 5347 2764 5375
rect 2996 5347 3004 5376
rect 3147 5376 3184 5384
rect 2107 5335 2133 5343
rect 2367 5336 2433 5344
rect 2587 5336 2604 5347
rect 2587 5333 2600 5336
rect 2667 5335 2693 5343
rect 2807 5336 2873 5344
rect 2887 5336 2913 5344
rect 107 5316 193 5324
rect 587 5316 753 5324
rect 807 5316 1113 5324
rect 1247 5316 1433 5324
rect 1447 5316 1873 5324
rect 576 5304 584 5313
rect 527 5296 584 5304
rect 787 5296 813 5304
rect 1236 5304 1244 5313
rect 2007 5316 2333 5324
rect 3056 5324 3064 5373
rect 3096 5347 3104 5373
rect 3176 5347 3184 5376
rect 3207 5376 3233 5384
rect 3467 5376 3493 5384
rect 3316 5344 3324 5375
rect 3416 5364 3424 5375
rect 3667 5376 3713 5384
rect 3736 5364 3744 5393
rect 3767 5376 3893 5384
rect 3907 5377 4033 5385
rect 3416 5356 3724 5364
rect 3736 5356 3933 5364
rect 3416 5347 3424 5356
rect 3316 5336 3373 5344
rect 3467 5336 3493 5344
rect 3716 5344 3724 5356
rect 3716 5336 3773 5344
rect 2967 5316 3064 5324
rect 3247 5316 3324 5324
rect 827 5296 1244 5304
rect 1927 5296 2473 5304
rect 2487 5296 2893 5304
rect 2947 5296 3213 5304
rect 3316 5304 3324 5316
rect 3347 5316 3573 5324
rect 3587 5316 3693 5324
rect 4076 5324 4084 5373
rect 4116 5364 4124 5374
rect 4027 5316 4084 5324
rect 4096 5356 4124 5364
rect 3316 5296 3364 5304
rect 1667 5276 1773 5284
rect 1787 5276 2033 5284
rect 2347 5276 2453 5284
rect 2687 5276 2733 5284
rect 2927 5276 3233 5284
rect 3356 5284 3364 5296
rect 3407 5296 3633 5304
rect 4096 5304 4104 5356
rect 4156 5347 4164 5374
rect 4187 5384 4200 5387
rect 4187 5373 4204 5384
rect 4347 5376 4373 5384
rect 4567 5378 4713 5386
rect 4767 5376 4793 5384
rect 4196 5364 4204 5373
rect 4196 5356 4224 5364
rect 4216 5347 4224 5356
rect 4496 5347 4504 5374
rect 4887 5376 4924 5384
rect 4156 5336 4173 5347
rect 4160 5333 4173 5336
rect 4216 5336 4233 5347
rect 4220 5333 4233 5336
rect 4307 5336 4373 5344
rect 4487 5336 4504 5347
rect 4487 5333 4500 5336
rect 4627 5336 4693 5344
rect 4836 5344 4844 5374
rect 4916 5364 4924 5376
rect 4947 5378 4993 5386
rect 5147 5376 5253 5384
rect 5307 5376 5344 5384
rect 5336 5364 5344 5376
rect 5367 5376 5413 5384
rect 5567 5376 5613 5384
rect 4916 5356 4984 5364
rect 5336 5356 5444 5364
rect 4747 5336 4844 5344
rect 4976 5344 4984 5356
rect 5436 5346 5444 5356
rect 4976 5336 5004 5344
rect 4267 5316 4433 5324
rect 4613 5324 4627 5332
rect 4447 5316 4627 5324
rect 4996 5324 5004 5336
rect 5347 5335 5393 5343
rect 5447 5336 5533 5344
rect 4996 5316 5233 5324
rect 3967 5296 4104 5304
rect 4147 5296 4733 5304
rect 3356 5276 3753 5284
rect 3847 5276 4033 5284
rect 4107 5276 4193 5284
rect 4247 5276 4873 5284
rect 4887 5276 4893 5284
rect 427 5256 553 5264
rect 747 5256 793 5264
rect 1127 5256 1273 5264
rect 1347 5256 2364 5264
rect 2356 5247 2364 5256
rect 2507 5256 2733 5264
rect 2827 5256 2933 5264
rect 3087 5256 3292 5264
rect 3327 5256 3493 5264
rect 3947 5256 4013 5264
rect 4067 5256 4193 5264
rect 4327 5256 5173 5264
rect 5187 5256 5573 5264
rect 1427 5236 1573 5244
rect 1847 5236 1953 5244
rect 2207 5236 2313 5244
rect 2367 5236 2473 5244
rect 2487 5236 2753 5244
rect 2867 5236 3193 5244
rect 3207 5236 3393 5244
rect 3447 5236 3533 5244
rect 3547 5236 3673 5244
rect 3747 5236 3873 5244
rect 3887 5236 4073 5244
rect 4087 5236 4673 5244
rect 4747 5236 5113 5244
rect 207 5216 553 5224
rect 987 5216 1053 5224
rect 1147 5216 1173 5224
rect 1836 5224 1844 5233
rect 1187 5216 1844 5224
rect 2307 5216 2573 5224
rect 2627 5216 2773 5224
rect 3056 5216 3313 5224
rect 1207 5196 1513 5204
rect 2087 5196 2253 5204
rect 2267 5196 2724 5204
rect 487 5176 973 5184
rect 1287 5176 2133 5184
rect 2227 5176 2453 5184
rect 2716 5184 2724 5196
rect 3056 5204 3064 5216
rect 3507 5216 3693 5224
rect 3707 5216 3884 5224
rect 2907 5196 3064 5204
rect 3207 5196 3413 5204
rect 3876 5204 3884 5216
rect 3907 5216 4173 5224
rect 4187 5216 4413 5224
rect 4427 5216 4473 5224
rect 3876 5196 4293 5204
rect 4307 5196 4553 5204
rect 4687 5196 4853 5204
rect 2716 5176 3093 5184
rect 3247 5176 3373 5184
rect 3487 5176 3652 5184
rect 3687 5176 3953 5184
rect 3976 5176 4313 5184
rect 307 5156 533 5164
rect 1067 5156 2193 5164
rect 2867 5156 3193 5164
rect 3587 5156 3613 5164
rect 3976 5164 3984 5176
rect 5367 5176 5513 5184
rect 3767 5156 3984 5164
rect 4007 5156 4333 5164
rect 4667 5156 4693 5164
rect 4767 5156 4793 5164
rect 4807 5156 4913 5164
rect 4927 5156 5153 5164
rect 1076 5136 1173 5144
rect 127 5116 213 5124
rect 227 5116 313 5124
rect 487 5116 653 5124
rect 1076 5124 1084 5136
rect 1187 5136 1353 5144
rect 1367 5136 1533 5144
rect 1547 5136 2213 5144
rect 2427 5136 2533 5144
rect 2547 5136 2733 5144
rect 2747 5136 2813 5144
rect 3667 5136 3933 5144
rect 4267 5136 4313 5144
rect 5427 5136 5493 5144
rect 987 5116 1084 5124
rect 1247 5116 1313 5124
rect 2247 5116 2293 5124
rect 3227 5116 3613 5124
rect 3687 5116 3832 5124
rect 3867 5116 3944 5124
rect 707 5096 912 5104
rect 947 5096 1193 5104
rect 1347 5096 1393 5104
rect 1687 5096 1813 5104
rect 267 5076 293 5084
rect 76 5064 84 5074
rect 307 5076 353 5084
rect 527 5076 613 5084
rect 747 5076 813 5084
rect 1027 5076 1093 5084
rect 76 5056 104 5064
rect 96 5044 104 5056
rect 1076 5047 1084 5076
rect 1287 5076 1313 5084
rect 1527 5077 1673 5085
rect 96 5036 273 5044
rect 327 5036 453 5044
rect 567 5036 693 5044
rect 927 5036 1033 5044
rect 1376 5044 1384 5074
rect 1267 5036 1593 5044
rect 1696 5045 1704 5096
rect 1827 5096 1913 5104
rect 2147 5096 2393 5104
rect 2727 5096 2813 5104
rect 3087 5096 3173 5104
rect 3367 5096 3453 5104
rect 3647 5096 3913 5104
rect 3936 5104 3944 5116
rect 4107 5116 4333 5124
rect 4607 5116 4793 5124
rect 5247 5116 5333 5124
rect 5467 5116 5753 5124
rect 3936 5096 4053 5104
rect 4587 5096 4633 5104
rect 4647 5096 4733 5104
rect 4987 5096 5033 5104
rect 5367 5100 5484 5104
rect 5367 5096 5487 5100
rect 1727 5076 1773 5084
rect 1787 5076 1804 5084
rect 1796 5064 1804 5076
rect 2147 5076 2233 5084
rect 2287 5076 2313 5084
rect 2507 5076 2584 5084
rect 2576 5064 2584 5076
rect 2607 5076 2673 5084
rect 3007 5076 3064 5084
rect 2893 5064 2907 5073
rect 1796 5056 1924 5064
rect 2576 5056 2664 5064
rect 2696 5060 2907 5064
rect 3056 5064 3064 5076
rect 3447 5076 3484 5084
rect 3213 5064 3227 5073
rect 1916 5044 1924 5056
rect 1916 5036 1933 5044
rect 1947 5036 2053 5044
rect 2656 5045 2664 5056
rect 2693 5056 2904 5060
rect 3056 5056 3124 5064
rect 2693 5047 2707 5056
rect 3056 5052 3067 5056
rect 2187 5036 2253 5044
rect 2327 5034 2353 5042
rect 2447 5034 2613 5042
rect 3116 5044 3124 5056
rect 3196 5060 3227 5064
rect 3196 5056 3224 5060
rect 3196 5044 3204 5056
rect 3116 5036 3204 5044
rect 3316 5044 3324 5073
rect 3247 5036 3324 5044
rect 3476 5045 3484 5076
rect 3727 5076 3764 5084
rect 3496 5047 3504 5073
rect 3756 5064 3764 5076
rect 3787 5076 3853 5084
rect 4000 5084 4013 5087
rect 3996 5073 4013 5084
rect 4107 5076 4184 5084
rect 3756 5060 3844 5064
rect 3756 5056 3847 5060
rect 3833 5047 3847 5056
rect 3347 5038 3473 5044
rect 3333 5036 3473 5038
rect 3496 5036 3513 5047
rect 3500 5033 3513 5036
rect 3607 5036 3653 5044
rect 3996 5044 4004 5073
rect 4075 5047 4083 5073
rect 4176 5047 4184 5076
rect 4356 5076 4373 5084
rect 3927 5036 4004 5044
rect 47 5016 133 5024
rect 147 5016 193 5024
rect 727 5016 773 5024
rect 787 5016 993 5024
rect 1796 5016 1853 5024
rect 1796 5007 1804 5016
rect 2316 5024 2324 5031
rect 4236 5027 4244 5073
rect 4356 5064 4364 5076
rect 5473 5087 5487 5096
rect 4700 5084 4713 5087
rect 4527 5076 4564 5084
rect 4316 5056 4364 5064
rect 4556 5064 4564 5076
rect 4696 5073 4713 5084
rect 4767 5084 4780 5087
rect 4767 5073 4784 5084
rect 4916 5076 4933 5084
rect 4556 5056 4644 5064
rect 4316 5044 4324 5056
rect 4287 5036 4324 5044
rect 4347 5035 4433 5043
rect 4636 5044 4644 5056
rect 4696 5046 4704 5073
rect 4776 5046 4784 5073
rect 4856 5047 4864 5073
rect 4636 5040 4684 5044
rect 4636 5036 4687 5040
rect 4673 5027 4687 5036
rect 4916 5044 4924 5076
rect 4947 5076 4993 5084
rect 5107 5076 5133 5084
rect 5256 5076 5292 5084
rect 4907 5036 4924 5044
rect 5067 5036 5113 5044
rect 5127 5036 5153 5044
rect 5256 5044 5264 5076
rect 5656 5076 5693 5084
rect 5313 5064 5327 5072
rect 5533 5064 5547 5073
rect 5313 5060 5564 5064
rect 5316 5056 5564 5060
rect 5207 5036 5264 5044
rect 2127 5016 2324 5024
rect 2776 5016 3013 5024
rect 287 4996 373 5004
rect 1127 4996 1313 5004
rect 1607 4996 1793 5004
rect 1887 4996 2393 5004
rect 2507 4996 2693 5004
rect 2776 5004 2784 5016
rect 3087 5016 3313 5024
rect 3367 5016 3453 5024
rect 3627 5016 3813 5024
rect 4007 5016 4213 5024
rect 4236 5016 4253 5027
rect 4240 5013 4253 5016
rect 4927 5016 4953 5024
rect 4967 5016 5013 5024
rect 5556 5024 5564 5056
rect 5616 5047 5624 5073
rect 5656 5047 5664 5076
rect 5656 5024 5664 5033
rect 5556 5016 5664 5024
rect 2716 4996 2784 5004
rect 507 4976 633 4984
rect 647 4976 833 4984
rect 1116 4984 1124 4993
rect 1047 4976 1124 4984
rect 2267 4976 2433 4984
rect 2716 4984 2724 4996
rect 2847 4996 2933 5004
rect 2947 4996 3052 5004
rect 3087 4996 3273 5004
rect 3296 4996 3413 5004
rect 2647 4976 2724 4984
rect 2927 4976 2993 4984
rect 3296 4984 3304 4996
rect 3547 4996 3584 5004
rect 3016 4976 3304 4984
rect 247 4956 333 4964
rect 707 4956 793 4964
rect 1067 4956 1153 4964
rect 1627 4956 1813 4964
rect 2047 4956 2193 4964
rect 2767 4956 2813 4964
rect 3016 4964 3024 4976
rect 3467 4976 3513 4984
rect 3527 4976 3553 4984
rect 3576 4984 3584 4996
rect 3747 4996 3872 5004
rect 3907 4996 4113 5004
rect 4427 4996 4533 5004
rect 4547 4996 4573 5004
rect 5007 4996 5093 5004
rect 5107 4996 5253 5004
rect 5347 4996 5513 5004
rect 5527 4996 5553 5004
rect 3576 4976 3673 4984
rect 3767 4976 3873 4984
rect 4047 4976 4153 4984
rect 4407 4976 4493 4984
rect 4667 4976 4793 4984
rect 4807 4976 4933 4984
rect 2827 4956 3024 4964
rect 3067 4956 3113 4964
rect 3127 4956 3193 4964
rect 3247 4956 3353 4964
rect 3407 4956 3733 4964
rect 3907 4956 4173 4964
rect 4667 4956 4733 4964
rect 27 4936 73 4944
rect 127 4936 213 4944
rect 227 4936 353 4944
rect 847 4936 933 4944
rect 1447 4936 1573 4944
rect 1587 4936 2213 4944
rect 2327 4936 2453 4944
rect 2887 4936 3153 4944
rect 3427 4936 3664 4944
rect 396 4916 593 4924
rect 396 4907 404 4916
rect 1587 4916 1653 4924
rect 1947 4916 1973 4924
rect 2347 4916 2473 4924
rect 2487 4916 2513 4924
rect 3447 4916 3492 4924
rect 3527 4916 3613 4924
rect 3656 4924 3664 4936
rect 3927 4936 4164 4944
rect 3656 4916 3753 4924
rect 3887 4916 4053 4924
rect 4156 4924 4164 4936
rect 4207 4936 4313 4944
rect 5507 4936 5533 4944
rect 4156 4916 4233 4924
rect 4607 4916 4933 4924
rect 5487 4916 5593 4924
rect 327 4896 393 4904
rect 487 4896 533 4904
rect 807 4896 1053 4904
rect 1067 4896 1213 4904
rect 1547 4896 1673 4904
rect 1687 4896 1753 4904
rect 1847 4896 1893 4904
rect 1907 4896 2113 4904
rect 2207 4896 2393 4904
rect 2607 4896 2713 4904
rect 2987 4896 3173 4904
rect 3267 4896 3413 4904
rect 3847 4896 3913 4904
rect 3956 4896 4073 4904
rect 47 4876 93 4884
rect 427 4876 453 4884
rect 1247 4876 1333 4884
rect 2027 4876 2073 4884
rect 2687 4876 2733 4884
rect 3047 4876 3073 4884
rect 3327 4876 3373 4884
rect 3567 4876 3693 4884
rect 3956 4884 3964 4896
rect 4687 4896 4953 4904
rect 5067 4896 5153 4904
rect 5347 4896 5433 4904
rect 3747 4876 3964 4884
rect 3987 4876 4024 4884
rect 267 4856 284 4864
rect 276 4827 284 4856
rect 347 4864 360 4867
rect 347 4853 364 4864
rect 356 4827 364 4853
rect 47 4816 93 4824
rect 107 4816 193 4824
rect 376 4804 384 4873
rect 547 4856 633 4864
rect 496 4827 504 4855
rect 747 4856 793 4864
rect 847 4856 873 4864
rect 607 4815 913 4823
rect 976 4807 984 4854
rect 1127 4856 1173 4864
rect 1256 4856 1293 4864
rect 1256 4827 1264 4856
rect 1307 4856 1433 4864
rect 1487 4858 1513 4866
rect 1627 4856 1653 4864
rect 1775 4856 1832 4864
rect 1716 4827 1724 4855
rect 1775 4827 1783 4856
rect 1856 4844 1864 4855
rect 2036 4856 2113 4864
rect 1796 4840 1864 4844
rect 1793 4836 1864 4840
rect 1793 4827 1807 4836
rect 1935 4827 1943 4853
rect 1976 4827 1984 4854
rect 1087 4816 1232 4824
rect 1407 4816 1453 4824
rect 1967 4816 1984 4827
rect 2036 4826 2044 4856
rect 2187 4858 2233 4866
rect 2287 4856 2493 4864
rect 2507 4856 2524 4864
rect 1967 4813 1980 4816
rect 2147 4816 2253 4824
rect 2516 4826 2524 4856
rect 2547 4856 2564 4864
rect 2556 4844 2564 4856
rect 2587 4856 2633 4864
rect 2767 4856 2793 4864
rect 2816 4856 2873 4864
rect 2556 4840 2604 4844
rect 2556 4836 2607 4840
rect 2593 4827 2607 4836
rect 2816 4827 2824 4856
rect 2956 4844 2964 4873
rect 3356 4856 3473 4864
rect 2936 4840 2964 4844
rect 2933 4836 2964 4840
rect 2933 4827 2947 4836
rect 2347 4815 2373 4823
rect 3056 4827 3064 4853
rect 3056 4816 3073 4827
rect 3060 4813 3073 4816
rect 3096 4824 3104 4855
rect 3096 4816 3253 4824
rect 3356 4826 3364 4856
rect 3587 4856 3604 4864
rect 3516 4827 3524 4853
rect 227 4796 553 4804
rect 1016 4796 1584 4804
rect 327 4776 473 4784
rect 527 4776 613 4784
rect 667 4776 773 4784
rect 967 4776 993 4784
rect 1016 4784 1024 4796
rect 1007 4776 1024 4784
rect 1087 4776 1553 4784
rect 1576 4784 1584 4796
rect 1687 4796 1913 4804
rect 1927 4796 2173 4804
rect 2816 4804 2824 4813
rect 3507 4816 3524 4827
rect 3507 4813 3520 4816
rect 2816 4796 2913 4804
rect 3067 4796 3433 4804
rect 3596 4804 3604 4856
rect 3616 4856 3653 4864
rect 3616 4827 3624 4856
rect 3856 4856 3893 4864
rect 3716 4844 3724 4854
rect 3716 4840 3824 4844
rect 3716 4836 3827 4840
rect 3813 4827 3827 4836
rect 3707 4816 3753 4824
rect 3836 4804 3844 4855
rect 3856 4827 3864 4856
rect 4016 4827 4024 4876
rect 5247 4876 5284 4884
rect 4127 4856 4144 4864
rect 3907 4816 4013 4824
rect 4136 4824 4144 4856
rect 4347 4857 4553 4865
rect 4727 4856 4773 4864
rect 4296 4827 4304 4853
rect 4836 4827 4844 4855
rect 4947 4856 4984 4864
rect 4915 4827 4923 4853
rect 4136 4816 4272 4824
rect 4487 4816 4533 4824
rect 4747 4815 4793 4823
rect 4907 4816 4923 4827
rect 4976 4826 4984 4856
rect 5007 4856 5044 4864
rect 4907 4813 4920 4816
rect 3596 4796 3844 4804
rect 4187 4796 4253 4804
rect 4896 4804 4904 4813
rect 5036 4824 5044 4856
rect 5127 4856 5184 4864
rect 5176 4847 5184 4856
rect 5176 4836 5193 4847
rect 5180 4833 5193 4836
rect 5036 4816 5093 4824
rect 5216 4824 5224 4853
rect 5276 4827 5284 4876
rect 5307 4876 5493 4884
rect 5507 4876 5573 4884
rect 5327 4864 5340 4867
rect 5327 4853 5344 4864
rect 5367 4856 5413 4864
rect 5600 4864 5613 4867
rect 5527 4856 5583 4864
rect 5167 4816 5224 4824
rect 4827 4796 4904 4804
rect 5276 4804 5284 4813
rect 5147 4796 5284 4804
rect 5336 4804 5344 4853
rect 5476 4827 5484 4853
rect 5575 4827 5583 4856
rect 5596 4853 5613 4864
rect 5596 4827 5604 4853
rect 5676 4844 5684 4873
rect 5707 4856 5744 4864
rect 5656 4836 5684 4844
rect 5656 4827 5664 4836
rect 5736 4827 5744 4856
rect 5647 4816 5664 4827
rect 5647 4813 5660 4816
rect 5336 4796 5433 4804
rect 5507 4796 5713 4804
rect 1576 4776 1613 4784
rect 1627 4776 1893 4784
rect 2507 4776 2693 4784
rect 2707 4776 2853 4784
rect 2867 4776 2953 4784
rect 3267 4776 3452 4784
rect 3487 4776 3593 4784
rect 4027 4776 4133 4784
rect 4147 4776 4333 4784
rect 4427 4776 4613 4784
rect 4867 4776 4973 4784
rect 307 4756 373 4764
rect 656 4764 664 4772
rect 507 4756 664 4764
rect 767 4756 813 4764
rect 1507 4756 1593 4764
rect 1607 4756 1953 4764
rect 2087 4756 2372 4764
rect 2407 4756 2473 4764
rect 2567 4756 2653 4764
rect 2667 4756 3033 4764
rect 3456 4764 3464 4773
rect 3456 4756 3613 4764
rect 3747 4756 3784 4764
rect 987 4736 1573 4744
rect 1967 4736 2513 4744
rect 2687 4736 3013 4744
rect 3776 4744 3784 4756
rect 3887 4756 4313 4764
rect 4367 4756 4533 4764
rect 3367 4736 3764 4744
rect 3776 4736 3913 4744
rect 147 4716 233 4724
rect 247 4716 873 4724
rect 947 4716 1033 4724
rect 1047 4716 1673 4724
rect 1747 4716 1873 4724
rect 1887 4716 2033 4724
rect 2047 4716 2213 4724
rect 2467 4716 2653 4724
rect 3087 4716 3584 4724
rect 267 4696 753 4704
rect 1287 4696 1713 4704
rect 1907 4696 2413 4704
rect 2547 4696 2673 4704
rect 2747 4696 2893 4704
rect 3576 4704 3584 4716
rect 3607 4716 3693 4724
rect 3756 4724 3764 4736
rect 4607 4736 4753 4744
rect 5067 4736 5673 4744
rect 3756 4716 3933 4724
rect 4196 4716 4393 4724
rect 3576 4696 3653 4704
rect 4196 4704 4204 4716
rect 4447 4716 4633 4724
rect 5347 4716 5513 4724
rect 3707 4696 4204 4704
rect 4227 4696 4693 4704
rect 4707 4696 5013 4704
rect 5027 4696 5153 4704
rect 5347 4696 5393 4704
rect 807 4676 1113 4684
rect 1567 4676 1813 4684
rect 1867 4676 2433 4684
rect 2487 4676 3093 4684
rect 3347 4676 3413 4684
rect 3427 4676 3893 4684
rect 3947 4676 3993 4684
rect 4247 4676 4353 4684
rect 4407 4676 5553 4684
rect 247 4656 393 4664
rect 407 4656 453 4664
rect 467 4656 593 4664
rect 747 4656 1313 4664
rect 1327 4656 1453 4664
rect 1467 4656 1513 4664
rect 1587 4656 1713 4664
rect 2087 4656 2393 4664
rect 2527 4656 3073 4664
rect 3127 4656 3553 4664
rect 3607 4656 5293 4664
rect 5307 4656 5413 4664
rect 767 4636 833 4644
rect 1827 4636 1873 4644
rect 2096 4636 2253 4644
rect 2096 4627 2104 4636
rect 2327 4636 3053 4644
rect 3107 4636 3304 4644
rect 47 4616 193 4624
rect 207 4616 253 4624
rect 467 4616 573 4624
rect 1207 4616 1313 4624
rect 1687 4616 1853 4624
rect 1927 4616 2093 4624
rect 2287 4616 2633 4624
rect 2647 4616 2733 4624
rect 2807 4616 3273 4624
rect 3296 4624 3304 4636
rect 3387 4636 3433 4644
rect 3647 4636 3753 4644
rect 3867 4636 4073 4644
rect 4536 4640 4812 4644
rect 4533 4636 4812 4640
rect 4533 4627 4547 4636
rect 4847 4636 5133 4644
rect 3296 4616 3473 4624
rect 4400 4624 4413 4627
rect 4396 4613 4413 4624
rect 287 4596 613 4604
rect 687 4596 712 4604
rect 747 4596 1113 4604
rect 1127 4596 1653 4604
rect 1727 4596 1953 4604
rect 2147 4596 2413 4604
rect 2467 4596 2513 4604
rect 2887 4596 2973 4604
rect 2987 4596 3133 4604
rect 3327 4596 3593 4604
rect 3667 4596 3733 4604
rect 4007 4596 4053 4604
rect 4396 4604 4404 4613
rect 4067 4596 4404 4604
rect 4787 4596 4953 4604
rect 367 4576 424 4584
rect 87 4556 133 4564
rect 47 4515 93 4523
rect 216 4525 224 4553
rect 336 4544 344 4554
rect 336 4540 384 4544
rect 336 4536 387 4540
rect 373 4527 387 4536
rect 416 4527 424 4576
rect 887 4576 913 4584
rect 1227 4576 1253 4584
rect 1716 4576 1793 4584
rect 507 4556 533 4564
rect 267 4516 313 4524
rect 427 4516 553 4524
rect 607 4514 633 4522
rect 676 4524 684 4553
rect 747 4556 853 4564
rect 876 4556 972 4564
rect 693 4544 707 4552
rect 876 4544 884 4556
rect 1036 4556 1073 4564
rect 693 4540 884 4544
rect 696 4536 884 4540
rect 676 4516 773 4524
rect 816 4525 824 4536
rect 996 4527 1004 4553
rect 1036 4527 1044 4556
rect 1120 4564 1133 4567
rect 1116 4553 1133 4564
rect 1567 4556 1693 4564
rect 1116 4544 1124 4553
rect 1233 4544 1247 4553
rect 1096 4536 1124 4544
rect 1136 4540 1247 4544
rect 1136 4536 1244 4540
rect 1096 4507 1104 4536
rect 1136 4525 1144 4536
rect 1416 4524 1424 4554
rect 1287 4520 1424 4524
rect 1287 4516 1427 4520
rect 1413 4507 1427 4516
rect 1716 4526 1724 4576
rect 2207 4576 2293 4584
rect 2307 4576 2353 4584
rect 2447 4576 2533 4584
rect 2767 4576 2793 4584
rect 2927 4576 2993 4584
rect 3047 4576 3113 4584
rect 3396 4576 3493 4584
rect 1827 4556 1853 4564
rect 1967 4556 1993 4564
rect 2146 4553 2147 4560
rect 2387 4556 2493 4564
rect 2667 4564 2680 4567
rect 2667 4553 2684 4564
rect 2747 4556 2813 4564
rect 3147 4556 3164 4564
rect 1447 4516 1533 4524
rect 1936 4525 1944 4553
rect 2076 4527 2084 4553
rect 2133 4544 2147 4553
rect 2096 4540 2147 4544
rect 2096 4536 2143 4540
rect 467 4496 493 4504
rect 1096 4496 1113 4507
rect 1100 4493 1113 4496
rect 1713 4504 1727 4512
rect 1587 4496 1727 4504
rect 1787 4496 1873 4504
rect 2096 4504 2104 4536
rect 2156 4524 2164 4553
rect 2313 4544 2327 4553
rect 2256 4540 2327 4544
rect 2676 4544 2684 4553
rect 2256 4536 2324 4540
rect 2676 4536 2724 4544
rect 2127 4516 2164 4524
rect 2256 4524 2264 4536
rect 2227 4516 2264 4524
rect 2287 4516 2333 4524
rect 2716 4524 2724 4536
rect 2716 4516 2833 4524
rect 2896 4525 2904 4553
rect 2933 4544 2947 4553
rect 3156 4547 3164 4556
rect 3187 4557 3233 4565
rect 3156 4546 3180 4547
rect 2933 4540 3024 4544
rect 2936 4536 3024 4540
rect 3156 4536 3173 4546
rect 2907 4516 2993 4524
rect 1987 4496 2104 4504
rect 2447 4496 2573 4504
rect 3016 4504 3024 4536
rect 3160 4533 3173 4536
rect 3396 4527 3404 4576
rect 3580 4586 3600 4587
rect 3580 4584 3593 4586
rect 3087 4516 3153 4524
rect 3267 4516 3313 4524
rect 3456 4524 3464 4553
rect 3553 4564 3567 4573
rect 3507 4560 3567 4564
rect 3576 4573 3593 4584
rect 3507 4556 3563 4560
rect 3456 4516 3473 4524
rect 2887 4496 3024 4504
rect 3187 4496 3213 4504
rect 3496 4504 3504 4552
rect 3576 4527 3584 4573
rect 3787 4576 3813 4584
rect 3827 4576 3984 4584
rect 3976 4567 3984 4576
rect 4167 4576 4464 4584
rect 3987 4564 4000 4567
rect 3987 4553 4004 4564
rect 4047 4556 4093 4564
rect 4216 4556 4353 4564
rect 3753 4544 3767 4553
rect 3716 4540 3767 4544
rect 3716 4536 3764 4540
rect 3627 4516 3673 4524
rect 3716 4526 3724 4536
rect 3996 4527 4004 4553
rect 3787 4514 3833 4522
rect 4216 4524 4224 4556
rect 4456 4567 4464 4576
rect 4656 4576 4793 4584
rect 4656 4567 4664 4576
rect 4807 4576 4913 4584
rect 4456 4556 4473 4567
rect 4047 4516 4224 4524
rect 3487 4490 3504 4504
rect 3747 4496 3813 4504
rect 4027 4496 4073 4504
rect 4396 4504 4404 4554
rect 4460 4553 4473 4556
rect 4707 4556 4773 4564
rect 5007 4556 5093 4564
rect 5107 4556 5233 4564
rect 5387 4564 5400 4567
rect 5387 4553 5404 4564
rect 5587 4556 5693 4564
rect 4656 4527 4664 4553
rect 5396 4527 5404 4553
rect 4647 4516 4664 4527
rect 4647 4513 4660 4516
rect 5307 4515 5353 4523
rect 5547 4516 5573 4524
rect 5587 4514 5713 4522
rect 4396 4496 4473 4504
rect 4767 4496 4793 4504
rect 5067 4496 5113 4504
rect 827 4476 973 4484
rect 987 4476 1033 4484
rect 1307 4476 1473 4484
rect 2007 4476 2053 4484
rect 2067 4476 2213 4484
rect 2627 4476 2713 4484
rect 2727 4476 2793 4484
rect 3027 4476 3293 4484
rect 3587 4476 3673 4484
rect 3767 4476 3873 4484
rect 4207 4476 4273 4484
rect 4387 4476 4673 4484
rect 4687 4476 4813 4484
rect 5447 4476 5473 4484
rect 5487 4476 5613 4484
rect 147 4456 393 4464
rect 787 4456 853 4464
rect 1247 4456 1453 4464
rect 1607 4456 1973 4464
rect 2487 4456 2533 4464
rect 2827 4456 3113 4464
rect 3447 4456 3513 4464
rect 3747 4456 4293 4464
rect 3916 4447 3924 4456
rect 4767 4456 5013 4464
rect 5027 4456 5073 4464
rect 5127 4456 5233 4464
rect 327 4436 533 4444
rect 547 4436 713 4444
rect 1507 4436 1933 4444
rect 2187 4436 2213 4444
rect 2667 4436 2773 4444
rect 2787 4436 2993 4444
rect 3607 4436 3653 4444
rect 3927 4436 3973 4444
rect 4047 4436 4373 4444
rect 4927 4436 5213 4444
rect 1107 4416 1173 4424
rect 1367 4416 1433 4424
rect 1547 4416 1613 4424
rect 2447 4416 2473 4424
rect 2527 4416 3033 4424
rect 3107 4416 3353 4424
rect 3847 4416 4213 4424
rect 4227 4416 4313 4424
rect 4327 4416 4613 4424
rect 5327 4416 5613 4424
rect 947 4396 993 4404
rect 1407 4396 1593 4404
rect 1747 4396 1904 4404
rect 107 4376 233 4384
rect 247 4376 293 4384
rect 447 4376 513 4384
rect 527 4376 593 4384
rect 607 4376 653 4384
rect 1067 4376 1153 4384
rect 1287 4376 1313 4384
rect 1487 4376 1724 4384
rect 316 4356 373 4364
rect 96 4284 104 4334
rect 147 4336 193 4344
rect 316 4306 324 4356
rect 347 4336 384 4344
rect 376 4307 384 4336
rect 507 4336 673 4344
rect 413 4324 427 4333
rect 413 4320 444 4324
rect 416 4316 444 4320
rect 227 4296 313 4304
rect 96 4276 353 4284
rect 436 4284 444 4316
rect 456 4304 464 4335
rect 887 4338 913 4346
rect 716 4307 724 4333
rect 456 4296 613 4304
rect 756 4304 764 4335
rect 956 4307 964 4333
rect 1096 4307 1104 4335
rect 1147 4344 1160 4347
rect 1147 4333 1164 4344
rect 1296 4336 1313 4344
rect 1156 4324 1164 4333
rect 1156 4320 1204 4324
rect 1156 4316 1207 4320
rect 1193 4307 1207 4316
rect 756 4296 853 4304
rect 436 4276 473 4284
rect 487 4276 573 4284
rect 616 4284 624 4293
rect 616 4276 733 4284
rect 947 4276 993 4284
rect 1236 4284 1244 4334
rect 1296 4307 1304 4336
rect 1376 4307 1384 4353
rect 1427 4337 1573 4345
rect 1576 4324 1584 4334
rect 1647 4336 1693 4344
rect 1716 4324 1724 4376
rect 1787 4376 1853 4384
rect 1896 4384 1904 4396
rect 2167 4396 2373 4404
rect 2987 4396 3464 4404
rect 3456 4387 3464 4396
rect 3627 4396 3693 4404
rect 3707 4396 3753 4404
rect 3967 4396 4033 4404
rect 4087 4396 4193 4404
rect 4727 4396 5093 4404
rect 5107 4396 5153 4404
rect 5527 4396 5573 4404
rect 1896 4376 2173 4384
rect 2447 4376 2593 4384
rect 2847 4376 2953 4384
rect 3247 4376 3353 4384
rect 3467 4376 3533 4384
rect 4007 4376 4204 4384
rect 2207 4356 2252 4364
rect 2287 4356 2413 4364
rect 3007 4356 3304 4364
rect 1867 4338 1913 4346
rect 2007 4336 2052 4344
rect 2087 4336 2164 4344
rect 1576 4320 1664 4324
rect 1576 4316 1667 4320
rect 1716 4316 1764 4324
rect 1653 4307 1667 4316
rect 1756 4304 1764 4316
rect 2156 4307 2164 4336
rect 2187 4336 2284 4344
rect 2276 4324 2284 4336
rect 2307 4338 2333 4346
rect 2387 4336 2433 4344
rect 2636 4336 2713 4344
rect 2276 4316 2584 4324
rect 1756 4296 1793 4304
rect 1927 4296 1973 4304
rect 2067 4295 2093 4303
rect 2156 4296 2173 4307
rect 2160 4293 2173 4296
rect 2327 4295 2493 4303
rect 1236 4276 1353 4284
rect 1847 4276 2013 4284
rect 2576 4284 2584 4316
rect 2596 4307 2604 4335
rect 2636 4307 2644 4336
rect 2736 4336 2853 4344
rect 2736 4306 2744 4336
rect 2893 4344 2907 4353
rect 2893 4340 2953 4344
rect 2896 4336 2953 4340
rect 3296 4344 3304 4356
rect 3347 4356 3644 4364
rect 3107 4336 3244 4344
rect 3296 4336 3593 4344
rect 2816 4320 3013 4324
rect 2813 4316 3013 4320
rect 2813 4307 2827 4316
rect 3236 4324 3244 4336
rect 3636 4324 3644 4356
rect 4047 4356 4093 4364
rect 4196 4364 4204 4376
rect 4867 4376 4952 4384
rect 4987 4376 5013 4384
rect 4196 4356 4293 4364
rect 4347 4356 4433 4364
rect 5100 4364 5113 4367
rect 5096 4353 5113 4364
rect 5316 4356 5372 4364
rect 3707 4344 3720 4347
rect 3707 4333 3724 4344
rect 3236 4320 3264 4324
rect 3556 4320 3644 4324
rect 3236 4316 3267 4320
rect 3253 4307 3267 4316
rect 3553 4316 3644 4320
rect 3553 4307 3567 4316
rect 3067 4296 3232 4304
rect 3427 4296 3513 4304
rect 3716 4304 3724 4333
rect 3816 4336 3853 4344
rect 3816 4324 3824 4336
rect 3907 4336 4113 4344
rect 4456 4336 4573 4344
rect 3776 4320 4144 4324
rect 3773 4316 4144 4320
rect 3773 4307 3787 4316
rect 3667 4296 3744 4304
rect 2576 4276 2693 4284
rect 2927 4276 3293 4284
rect 3407 4276 3524 4284
rect 87 4256 173 4264
rect 1427 4256 1673 4264
rect 1687 4256 1713 4264
rect 1867 4256 2073 4264
rect 2167 4256 2644 4264
rect 367 4236 413 4244
rect 427 4236 1093 4244
rect 1227 4236 1373 4244
rect 1387 4236 1473 4244
rect 1667 4236 1792 4244
rect 1827 4236 2113 4244
rect 2487 4236 2533 4244
rect 2636 4244 2644 4256
rect 2716 4256 2893 4264
rect 2716 4244 2724 4256
rect 3127 4256 3173 4264
rect 3387 4256 3493 4264
rect 3516 4264 3524 4276
rect 3627 4276 3713 4284
rect 3736 4284 3744 4296
rect 3927 4296 4013 4304
rect 4027 4296 4073 4304
rect 3736 4276 3893 4284
rect 3987 4276 4013 4284
rect 4136 4284 4144 4316
rect 4456 4324 4464 4336
rect 4427 4316 4464 4324
rect 4716 4304 4724 4335
rect 5007 4336 5033 4344
rect 4876 4324 4884 4334
rect 4827 4316 4884 4324
rect 5056 4307 5064 4333
rect 5096 4307 5104 4353
rect 5316 4347 5324 4356
rect 5147 4336 5173 4344
rect 5307 4336 5324 4347
rect 5393 4344 5407 4353
rect 5376 4340 5407 4344
rect 5416 4356 5453 4364
rect 5376 4336 5404 4340
rect 5307 4333 5320 4336
rect 5376 4307 5384 4336
rect 5416 4307 5424 4356
rect 5527 4356 5553 4364
rect 5456 4336 5533 4344
rect 5456 4307 5464 4336
rect 5587 4336 5623 4344
rect 5615 4307 5623 4336
rect 5667 4336 5693 4344
rect 4587 4296 4724 4304
rect 4987 4296 5013 4304
rect 5187 4296 5253 4304
rect 5647 4296 5733 4304
rect 4136 4276 4193 4284
rect 4387 4276 4453 4284
rect 3516 4256 3593 4264
rect 3747 4256 3913 4264
rect 4227 4256 4813 4264
rect 4827 4256 4933 4264
rect 5267 4256 5393 4264
rect 5407 4256 5593 4264
rect 2636 4236 2724 4244
rect 2847 4236 3053 4244
rect 3127 4236 3212 4244
rect 3247 4236 3653 4244
rect 3707 4236 3833 4244
rect 4367 4236 4413 4244
rect 4427 4236 4733 4244
rect 5047 4236 5233 4244
rect 5347 4236 5493 4244
rect 447 4216 513 4224
rect 1187 4216 1333 4224
rect 1407 4216 1852 4224
rect 1887 4216 2053 4224
rect 2587 4216 2893 4224
rect 2987 4216 3433 4224
rect 3507 4216 3953 4224
rect 4467 4216 4593 4224
rect 4607 4216 4693 4224
rect 4867 4216 5073 4224
rect 807 4196 893 4204
rect 907 4196 1253 4204
rect 1347 4196 1953 4204
rect 2147 4196 2453 4204
rect 3467 4196 3533 4204
rect 3547 4196 3813 4204
rect 4136 4196 5133 4204
rect 1287 4176 1353 4184
rect 1547 4176 1753 4184
rect 1807 4176 2033 4184
rect 2567 4176 2624 4184
rect 2616 4167 2624 4176
rect 2687 4176 3333 4184
rect 3547 4176 3613 4184
rect 3887 4176 3964 4184
rect 1087 4156 1833 4164
rect 2127 4156 2213 4164
rect 2347 4156 2533 4164
rect 2627 4156 2913 4164
rect 3107 4156 3413 4164
rect 3427 4156 3613 4164
rect 3687 4156 3853 4164
rect 3956 4164 3964 4176
rect 4136 4184 4144 4196
rect 3987 4176 4144 4184
rect 5367 4176 5593 4184
rect 5607 4176 5693 4184
rect 3956 4156 3993 4164
rect 4007 4156 4093 4164
rect 4207 4156 4333 4164
rect 187 4136 473 4144
rect 707 4136 853 4144
rect 1067 4136 1112 4144
rect 1147 4136 1393 4144
rect 1456 4136 1613 4144
rect 27 4116 613 4124
rect 727 4116 813 4124
rect 827 4116 913 4124
rect 1047 4116 1153 4124
rect 1456 4124 1464 4136
rect 1847 4136 1932 4144
rect 1967 4136 2044 4144
rect 1307 4116 1464 4124
rect 1607 4116 1773 4124
rect 2036 4124 2044 4136
rect 2067 4136 2313 4144
rect 2387 4136 2513 4144
rect 2667 4136 2933 4144
rect 3527 4136 3633 4144
rect 3647 4136 3664 4144
rect 2036 4116 2153 4124
rect 2567 4116 3173 4124
rect 3187 4116 3253 4124
rect 3276 4116 3444 4124
rect 887 4096 1133 4104
rect 1267 4096 1493 4104
rect 1687 4096 1913 4104
rect 2027 4096 2333 4104
rect 2407 4096 2513 4104
rect 3276 4104 3284 4116
rect 2627 4096 3284 4104
rect 3436 4104 3444 4116
rect 3476 4116 3553 4124
rect 3476 4104 3484 4116
rect 3607 4116 3633 4124
rect 3656 4124 3664 4136
rect 5027 4136 5153 4144
rect 5247 4136 5553 4144
rect 3656 4116 3732 4124
rect 3767 4116 3884 4124
rect 3436 4096 3484 4104
rect 3587 4096 3753 4104
rect 3876 4104 3884 4116
rect 3907 4116 4073 4124
rect 4147 4116 4433 4124
rect 4447 4116 4533 4124
rect 4547 4116 4613 4124
rect 4667 4116 4753 4124
rect 3876 4096 4053 4104
rect 4096 4096 5013 4104
rect 527 4076 553 4084
rect 747 4076 1093 4084
rect 2207 4076 2313 4084
rect 2387 4076 2573 4084
rect 2927 4076 2953 4084
rect 3147 4076 3413 4084
rect 3647 4076 3713 4084
rect 4096 4084 4104 4096
rect 5107 4096 5273 4104
rect 3887 4076 4104 4084
rect 4507 4076 4573 4084
rect 5387 4076 5493 4084
rect 5536 4076 5804 4084
rect 116 4056 133 4064
rect 116 4005 124 4056
rect 147 4056 193 4064
rect 516 4064 524 4073
rect 387 4056 524 4064
rect 587 4056 613 4064
rect 1007 4056 1073 4064
rect 1127 4056 1313 4064
rect 1327 4056 1393 4064
rect 1647 4056 1673 4064
rect 1853 4064 1867 4073
rect 1727 4060 1867 4064
rect 1727 4056 1864 4060
rect 1987 4056 2132 4064
rect 2167 4056 2353 4064
rect 247 4036 293 4044
rect 340 4044 353 4047
rect 336 4033 353 4044
rect 436 4036 533 4044
rect 136 4004 144 4032
rect 336 4007 344 4033
rect 136 3996 213 4004
rect 396 4005 404 4033
rect 436 4007 444 4036
rect 687 4036 713 4044
rect 840 4044 853 4047
rect 836 4033 853 4044
rect 1276 4036 1333 4044
rect 633 4024 647 4033
rect 633 4020 733 4024
rect 636 4016 733 4020
rect 213 3984 227 3991
rect 836 4006 844 4033
rect 847 3996 893 4004
rect 213 3976 353 3984
rect 393 3984 407 3991
rect 956 3987 964 4033
rect 1053 4024 1067 4033
rect 1036 4020 1067 4024
rect 1033 4016 1064 4020
rect 1033 4007 1047 4016
rect 1096 4004 1104 4033
rect 1276 4007 1284 4036
rect 1447 4036 1553 4044
rect 1653 4024 1667 4033
rect 1653 4020 1704 4024
rect 1656 4016 1704 4020
rect 1096 3996 1213 4004
rect 1467 3996 1633 4004
rect 1696 4005 1704 4016
rect 1796 4004 1804 4034
rect 1967 4036 2104 4044
rect 2096 4006 2104 4036
rect 1747 3996 1804 4004
rect 1947 3994 2033 4002
rect 2216 4004 2224 4056
rect 2607 4056 2633 4064
rect 2767 4056 2804 4064
rect 2407 4037 2453 4045
rect 2167 3996 2224 4004
rect 2236 4004 2244 4033
rect 2273 4024 2287 4033
rect 2687 4036 2784 4044
rect 2553 4024 2567 4033
rect 2273 4020 2304 4024
rect 2553 4020 2604 4024
rect 2276 4016 2304 4020
rect 2556 4016 2604 4020
rect 2296 4004 2304 4016
rect 2236 3996 2284 4004
rect 2296 3996 2573 4004
rect 393 3976 493 3984
rect 647 3976 713 3984
rect 727 3976 773 3984
rect 2227 3976 2253 3984
rect 2276 3984 2284 3996
rect 2596 4004 2604 4016
rect 2596 4000 2764 4004
rect 2596 3996 2767 4000
rect 2753 3987 2767 3996
rect 2276 3976 2373 3984
rect 2707 3976 2732 3984
rect 687 3956 764 3964
rect 756 3944 764 3956
rect 987 3956 1193 3964
rect 2147 3956 2184 3964
rect 756 3936 893 3944
rect 947 3936 993 3944
rect 1647 3936 1732 3944
rect 1767 3936 1793 3944
rect 1867 3936 1973 3944
rect 2176 3944 2184 3956
rect 2776 3964 2784 4036
rect 2796 3987 2804 4056
rect 2827 4056 2993 4064
rect 3007 4056 3073 4064
rect 3553 4064 3567 4073
rect 3553 4060 3584 4064
rect 3556 4056 3584 4060
rect 2947 4036 2984 4044
rect 2976 4007 2984 4036
rect 3016 4036 3073 4044
rect 3016 4007 3024 4036
rect 3227 4036 3333 4044
rect 2847 3994 2913 4002
rect 3116 4004 3124 4033
rect 3333 4024 3347 4032
rect 3436 4036 3493 4044
rect 3333 4020 3404 4024
rect 3336 4016 3407 4020
rect 3393 4007 3407 4016
rect 3067 3996 3124 4004
rect 3147 3996 3193 4004
rect 3436 4006 3444 4036
rect 3536 4004 3544 4053
rect 3576 4044 3584 4056
rect 3627 4056 3764 4064
rect 3576 4036 3604 4044
rect 3596 4004 3604 4036
rect 3756 4044 3764 4056
rect 3827 4056 3973 4064
rect 4087 4056 4153 4064
rect 4667 4056 4793 4064
rect 4967 4056 5073 4064
rect 5327 4056 5413 4064
rect 5427 4056 5444 4064
rect 3667 4036 3744 4044
rect 3756 4036 3793 4044
rect 3736 4007 3744 4036
rect 3847 4036 3964 4044
rect 3956 4027 3964 4036
rect 4067 4036 4104 4044
rect 3956 4016 3973 4027
rect 3960 4013 3973 4016
rect 3536 4000 3564 4004
rect 3536 3996 3567 4000
rect 3596 3996 3653 4004
rect 3553 3987 3567 3996
rect 3996 4004 4004 4033
rect 4096 4007 4104 4036
rect 4207 4037 4253 4045
rect 4367 4037 4393 4045
rect 3916 3996 4004 4004
rect 3727 3976 3813 3984
rect 3916 3984 3924 3996
rect 3887 3976 3924 3984
rect 4136 3984 4144 4033
rect 4296 4004 4304 4034
rect 4707 4036 4833 4044
rect 4847 4036 4893 4044
rect 4496 4007 4504 4033
rect 4296 3996 4413 4004
rect 4687 3994 4753 4002
rect 5196 4004 5204 4033
rect 5436 4024 5444 4056
rect 5536 4064 5544 4076
rect 5467 4056 5544 4064
rect 5727 4056 5753 4064
rect 5436 4020 5484 4024
rect 5436 4016 5487 4020
rect 5473 4007 5487 4016
rect 5196 3996 5333 4004
rect 4047 3976 4144 3984
rect 4287 3976 4373 3984
rect 4587 3976 4613 3984
rect 4756 3984 4764 3991
rect 5556 3987 5564 4034
rect 5707 4036 5804 4044
rect 5596 4007 5604 4033
rect 4756 3976 4813 3984
rect 5147 3976 5453 3984
rect 2667 3956 2784 3964
rect 3147 3956 3273 3964
rect 3327 3956 3633 3964
rect 4027 3956 4193 3964
rect 4467 3956 4513 3964
rect 5167 3956 5413 3964
rect 5587 3956 5693 3964
rect 5707 3956 5753 3964
rect 2176 3936 2373 3944
rect 2547 3936 2633 3944
rect 2887 3936 3153 3944
rect 3167 3936 3412 3944
rect 3447 3936 3473 3944
rect 3527 3936 3913 3944
rect 3967 3936 4593 3944
rect 4647 3936 5653 3944
rect 227 3916 553 3924
rect 567 3916 733 3924
rect 1067 3916 1113 3924
rect 1207 3916 1473 3924
rect 1487 3916 1533 3924
rect 1627 3916 1753 3924
rect 2067 3916 2373 3924
rect 2447 3916 2732 3924
rect 2767 3916 2793 3924
rect 3107 3916 3153 3924
rect 3476 3924 3484 3933
rect 3407 3916 3533 3924
rect 3607 3916 3853 3924
rect 4107 3916 4393 3924
rect 4976 3916 5053 3924
rect 4976 3907 4984 3916
rect 87 3896 133 3904
rect 387 3896 453 3904
rect 467 3896 813 3904
rect 947 3896 1093 3904
rect 1787 3896 1833 3904
rect 1847 3896 2133 3904
rect 2427 3896 2833 3904
rect 2987 3896 3113 3904
rect 3567 3896 3653 3904
rect 3987 3896 4033 3904
rect 4147 3896 4233 3904
rect 4727 3896 4753 3904
rect 4867 3896 4973 3904
rect 5547 3896 5753 3904
rect 927 3876 973 3884
rect 1047 3876 1093 3884
rect 1287 3876 1413 3884
rect 2327 3876 2493 3884
rect 2627 3876 2773 3884
rect 3027 3876 3513 3884
rect 3587 3876 3833 3884
rect 3967 3876 4044 3884
rect 27 3856 93 3864
rect 347 3856 413 3864
rect 587 3856 653 3864
rect 987 3856 1013 3864
rect 1247 3856 1324 3864
rect 1316 3847 1324 3856
rect 1607 3856 1633 3864
rect 1827 3856 1873 3864
rect 1947 3856 1993 3864
rect 2147 3856 2173 3864
rect 2440 3864 2453 3867
rect 2436 3853 2453 3864
rect 2587 3856 2664 3864
rect 47 3836 173 3844
rect 787 3836 873 3844
rect 887 3836 1012 3844
rect 1040 3844 1053 3847
rect 1036 3833 1053 3844
rect 1306 3833 1307 3840
rect 1327 3836 1393 3844
rect 1447 3836 1493 3844
rect 2187 3836 2384 3844
rect 147 3824 160 3827
rect 147 3813 164 3824
rect 347 3816 384 3824
rect 156 3787 164 3813
rect 47 3776 73 3784
rect 207 3776 253 3784
rect 267 3776 353 3784
rect 376 3767 384 3816
rect 447 3824 460 3827
rect 447 3813 464 3824
rect 507 3818 533 3826
rect 547 3816 593 3824
rect 456 3787 464 3813
rect 636 3804 644 3815
rect 687 3817 713 3825
rect 756 3804 764 3814
rect 636 3800 664 3804
rect 636 3796 667 3800
rect 756 3796 953 3804
rect 653 3787 667 3796
rect 893 3787 907 3796
rect 976 3787 984 3813
rect 1036 3787 1044 3833
rect 1076 3816 1133 3824
rect 1076 3787 1084 3816
rect 1156 3787 1164 3833
rect 1220 3824 1233 3827
rect 1216 3813 1233 3824
rect 1293 3824 1307 3833
rect 1293 3820 1343 3824
rect 1296 3816 1343 3820
rect 1216 3787 1224 3813
rect 1335 3787 1343 3816
rect 1460 3824 1473 3827
rect 1456 3813 1473 3824
rect 1516 3816 1553 3824
rect 1356 3787 1364 3813
rect 747 3775 813 3783
rect 1456 3786 1464 3813
rect 1516 3786 1524 3816
rect 1576 3816 1632 3824
rect 1576 3804 1584 3816
rect 1667 3824 1680 3827
rect 1667 3813 1684 3824
rect 1720 3824 1733 3827
rect 1556 3800 1584 3804
rect 1553 3796 1584 3800
rect 1553 3787 1567 3796
rect 1676 3787 1684 3813
rect 487 3756 573 3764
rect 707 3756 853 3764
rect 867 3756 953 3764
rect 1696 3764 1704 3815
rect 1607 3756 1704 3764
rect 1716 3813 1733 3824
rect 1893 3824 1907 3833
rect 1893 3820 1933 3824
rect 1896 3816 1933 3820
rect 2027 3824 2040 3827
rect 2027 3813 2044 3824
rect 27 3736 313 3744
rect 327 3736 673 3744
rect 1107 3736 1253 3744
rect 1407 3736 1493 3744
rect 1507 3736 1573 3744
rect 1716 3744 1724 3813
rect 2036 3804 2044 3813
rect 1836 3800 2044 3804
rect 1833 3796 2044 3800
rect 1833 3787 1847 3796
rect 2036 3787 2044 3796
rect 2076 3787 2084 3815
rect 2166 3813 2167 3820
rect 2307 3816 2353 3824
rect 2153 3804 2167 3813
rect 2136 3800 2167 3804
rect 2136 3796 2163 3800
rect 1747 3776 1833 3784
rect 2136 3764 2144 3796
rect 2176 3787 2184 3813
rect 2376 3787 2384 3836
rect 2436 3787 2444 3853
rect 2656 3844 2664 3856
rect 3387 3856 3453 3864
rect 3547 3856 3673 3864
rect 3927 3856 3973 3864
rect 4036 3864 4044 3876
rect 4087 3876 4353 3884
rect 4367 3876 4433 3884
rect 4627 3876 4993 3884
rect 4036 3856 4104 3864
rect 2656 3836 2693 3844
rect 2867 3844 2880 3847
rect 2867 3833 2884 3844
rect 3607 3844 3620 3847
rect 3607 3833 3624 3844
rect 2167 3776 2184 3787
rect 2167 3773 2180 3776
rect 2247 3776 2333 3784
rect 2476 3784 2484 3833
rect 2507 3818 2633 3826
rect 2736 3787 2744 3813
rect 2836 3804 2844 3814
rect 2876 3804 2884 3833
rect 3227 3816 3324 3824
rect 2836 3796 2864 3804
rect 2876 3796 3144 3804
rect 2476 3776 2533 3784
rect 2607 3776 2633 3784
rect 2856 3784 2864 3796
rect 2856 3776 2973 3784
rect 3136 3784 3144 3796
rect 3136 3776 3213 3784
rect 3316 3786 3324 3816
rect 3387 3816 3432 3824
rect 3376 3784 3384 3814
rect 3467 3816 3524 3824
rect 3516 3787 3524 3816
rect 3336 3776 3384 3784
rect 1927 3756 2144 3764
rect 2307 3756 2473 3764
rect 2727 3756 2873 3764
rect 3127 3756 3293 3764
rect 1627 3736 1724 3744
rect 2067 3736 2153 3744
rect 2567 3736 2773 3744
rect 2987 3736 3033 3744
rect 3336 3744 3344 3776
rect 3407 3776 3473 3784
rect 3536 3764 3544 3814
rect 3576 3804 3584 3814
rect 3616 3804 3624 3833
rect 3956 3836 4013 3844
rect 3667 3824 3680 3827
rect 3667 3813 3684 3824
rect 3576 3796 3624 3804
rect 3676 3787 3684 3813
rect 3756 3816 3793 3824
rect 3756 3787 3764 3816
rect 3956 3824 3964 3836
rect 3847 3816 3964 3824
rect 3975 3816 4033 3824
rect 3936 3787 3944 3816
rect 3975 3787 3983 3816
rect 3607 3775 3633 3783
rect 3747 3776 3764 3787
rect 3747 3773 3760 3776
rect 3827 3776 3873 3784
rect 4096 3786 4104 3856
rect 4807 3856 4893 3864
rect 5187 3856 5353 3864
rect 5547 3856 5613 3864
rect 4236 3836 4313 3844
rect 4236 3804 4244 3836
rect 4567 3836 4613 3844
rect 4767 3836 4933 3844
rect 4947 3836 4964 3844
rect 4347 3816 4393 3824
rect 4167 3796 4244 3804
rect 4316 3804 4324 3813
rect 4667 3816 4713 3824
rect 4316 3800 4344 3804
rect 4316 3796 4347 3800
rect 4333 3787 4347 3796
rect 4516 3787 4524 3813
rect 4956 3787 4964 3836
rect 5167 3836 5213 3844
rect 5427 3836 5493 3844
rect 5236 3816 5253 3824
rect 5016 3787 5024 3813
rect 5236 3787 5244 3816
rect 5307 3816 5384 3824
rect 5376 3787 5384 3816
rect 5627 3816 5673 3824
rect 5476 3787 5484 3813
rect 4007 3775 4053 3783
rect 4107 3776 4253 3784
rect 4607 3776 4693 3784
rect 4747 3776 4833 3784
rect 5527 3776 5804 3784
rect 3507 3756 3544 3764
rect 4367 3756 4473 3764
rect 3247 3736 3344 3744
rect 3487 3736 3513 3744
rect 3527 3736 3553 3744
rect 4007 3736 4133 3744
rect 4267 3736 4293 3744
rect 4667 3736 5053 3744
rect 5127 3736 5253 3744
rect 5267 3736 5273 3744
rect 5387 3736 5573 3744
rect 427 3716 513 3724
rect 527 3716 613 3724
rect 707 3716 813 3724
rect 1247 3716 1333 3724
rect 2547 3716 2713 3724
rect 2887 3716 3012 3724
rect 3047 3716 3113 3724
rect 3367 3716 3413 3724
rect 3427 3716 3733 3724
rect 3927 3716 4192 3724
rect 4227 3716 4433 3724
rect 4807 3716 4993 3724
rect 5347 3716 5673 3724
rect 1147 3696 1413 3704
rect 2107 3696 2233 3704
rect 2256 3696 2553 3704
rect 227 3676 653 3684
rect 667 3676 773 3684
rect 847 3676 1173 3684
rect 1347 3676 1413 3684
rect 1427 3676 1733 3684
rect 1807 3676 1913 3684
rect 2256 3684 2264 3696
rect 2687 3696 2813 3704
rect 3947 3696 4233 3704
rect 2227 3676 2264 3684
rect 2347 3676 2493 3684
rect 2707 3676 2753 3684
rect 2887 3676 3393 3684
rect 3407 3676 3553 3684
rect 3727 3676 3913 3684
rect 4047 3676 4213 3684
rect 4867 3676 5053 3684
rect 287 3656 433 3664
rect 807 3656 1273 3664
rect 1767 3656 1824 3664
rect 587 3636 773 3644
rect 947 3636 1072 3644
rect 1107 3636 1173 3644
rect 1307 3636 1793 3644
rect 1816 3644 1824 3656
rect 1987 3656 2293 3664
rect 2307 3656 2413 3664
rect 2587 3656 2733 3664
rect 2776 3656 2973 3664
rect 1816 3636 1993 3644
rect 2007 3636 2133 3644
rect 2327 3636 2453 3644
rect 2507 3636 2653 3644
rect 2776 3644 2784 3656
rect 3067 3656 3104 3664
rect 2727 3636 2784 3644
rect 2836 3636 2873 3644
rect 827 3616 1093 3624
rect 1287 3616 1353 3624
rect 1987 3616 2333 3624
rect 2620 3624 2633 3627
rect 2376 3616 2444 3624
rect 2376 3607 2384 3616
rect 27 3596 793 3604
rect 847 3596 1053 3604
rect 1067 3596 1453 3604
rect 1527 3596 1673 3604
rect 1907 3596 2373 3604
rect 2436 3604 2444 3616
rect 2616 3613 2633 3624
rect 2616 3604 2624 3613
rect 2836 3624 2844 3636
rect 2947 3636 3033 3644
rect 3096 3644 3104 3656
rect 3187 3656 3253 3664
rect 3687 3656 3853 3664
rect 4067 3656 4433 3664
rect 5236 3656 5593 3664
rect 3096 3636 3393 3644
rect 3407 3636 3493 3644
rect 3567 3636 3953 3644
rect 4187 3636 4513 3644
rect 5236 3644 5244 3656
rect 4907 3636 5244 3644
rect 2727 3616 2844 3624
rect 3087 3616 3153 3624
rect 3227 3616 3453 3624
rect 3547 3616 3653 3624
rect 3887 3616 4033 3624
rect 4087 3616 4153 3624
rect 4207 3616 4413 3624
rect 5487 3616 5613 3624
rect 2436 3596 2624 3604
rect 2667 3596 2853 3604
rect 3107 3596 3733 3604
rect 4227 3596 4853 3604
rect 1107 3576 1293 3584
rect 1527 3576 1593 3584
rect 1676 3576 1713 3584
rect -24 3556 53 3564
rect 527 3556 733 3564
rect 787 3556 873 3564
rect 1027 3556 1133 3564
rect 1147 3556 1193 3564
rect 1367 3556 1473 3564
rect 1676 3564 1684 3576
rect 2127 3576 2313 3584
rect 2427 3576 2693 3584
rect 2887 3576 3053 3584
rect 3187 3576 3272 3584
rect 3307 3576 3513 3584
rect 3736 3584 3744 3593
rect 3736 3576 3873 3584
rect 4927 3576 5213 3584
rect 5547 3576 5573 3584
rect 1487 3556 1684 3564
rect 1827 3556 1873 3564
rect 2216 3556 2333 3564
rect 2216 3547 2224 3556
rect 2347 3556 2612 3564
rect 2647 3556 2713 3564
rect 2867 3556 3553 3564
rect 5707 3556 5733 3564
rect 147 3536 233 3544
rect 927 3536 953 3544
rect 1167 3544 1180 3547
rect 1167 3533 1184 3544
rect -24 3516 33 3524
rect 607 3516 653 3524
rect 707 3516 793 3524
rect 216 3485 224 3513
rect 987 3520 1104 3524
rect 987 3516 1107 3520
rect 836 3487 844 3512
rect 873 3504 887 3513
rect 1093 3506 1107 3516
rect 873 3500 924 3504
rect 876 3496 924 3500
rect 127 3476 213 3484
rect 267 3476 293 3484
rect 447 3476 493 3484
rect 687 3476 813 3484
rect 836 3476 853 3487
rect 840 3473 853 3476
rect 916 3484 924 3496
rect 916 3476 1033 3484
rect 1176 3485 1184 3533
rect 1216 3536 1273 3544
rect 1216 3485 1224 3536
rect 2207 3536 2224 3547
rect 2207 3533 2220 3536
rect 1267 3516 1293 3524
rect 1606 3513 1607 3520
rect 1416 3487 1424 3513
rect 1456 3485 1464 3513
rect 1593 3504 1607 3513
rect 1496 3500 1607 3504
rect 1493 3496 1603 3500
rect 1493 3487 1507 3496
rect 1616 3484 1624 3513
rect 1653 3504 1667 3513
rect 1653 3500 1704 3504
rect 1656 3496 1704 3500
rect 1596 3480 1624 3484
rect 1593 3476 1624 3480
rect 1696 3484 1704 3496
rect 1776 3486 1784 3533
rect 2073 3524 2087 3533
rect 2073 3520 2253 3524
rect 2076 3516 2253 3520
rect 2267 3516 2393 3524
rect 1793 3504 1807 3513
rect 1793 3500 1884 3504
rect 1796 3496 1884 3500
rect 1696 3476 1733 3484
rect 1593 3467 1607 3476
rect 1876 3484 1884 3496
rect 1956 3487 1964 3513
rect 1993 3504 2007 3513
rect 1976 3500 2007 3504
rect 1976 3496 2004 3500
rect 1876 3476 1932 3484
rect 307 3456 353 3464
rect 627 3456 893 3464
rect 907 3456 1113 3464
rect 1976 3464 1984 3496
rect 2007 3476 2093 3484
rect 2236 3480 2273 3484
rect 2233 3476 2273 3480
rect 2233 3467 2247 3476
rect 2407 3476 2453 3484
rect 2516 3486 2524 3533
rect 2627 3536 2704 3544
rect 2560 3524 2573 3527
rect 2556 3513 2573 3524
rect 2556 3486 2564 3513
rect 2673 3504 2687 3513
rect 2656 3500 2687 3504
rect 2656 3496 2684 3500
rect 2656 3484 2664 3496
rect 2696 3487 2704 3536
rect 2747 3536 2813 3544
rect 2927 3536 2973 3544
rect 2987 3536 3093 3544
rect 3967 3536 4033 3544
rect 4467 3536 4693 3544
rect 4707 3536 4793 3544
rect 4956 3536 5133 3544
rect 2796 3504 2804 3514
rect 2996 3516 3033 3524
rect 2796 3496 2884 3504
rect 2647 3476 2664 3484
rect 2687 3476 2704 3487
rect 2687 3473 2700 3476
rect 2747 3476 2833 3484
rect 2876 3484 2884 3496
rect 2936 3487 2944 3513
rect 2876 3476 2893 3484
rect 1976 3456 2053 3464
rect 2996 3464 3004 3516
rect 3160 3524 3173 3527
rect 3156 3513 3173 3524
rect 3227 3516 3273 3524
rect 3156 3486 3164 3513
rect 3316 3484 3324 3513
rect 3436 3504 3444 3514
rect 3607 3517 3693 3525
rect 3716 3516 3813 3524
rect 3436 3500 3464 3504
rect 3436 3496 3467 3500
rect 3453 3487 3467 3496
rect 3316 3476 3353 3484
rect 3536 3485 3544 3513
rect 3716 3504 3724 3516
rect 3936 3516 4073 3524
rect 3627 3496 3724 3504
rect 3696 3476 3833 3484
rect 2967 3456 3004 3464
rect 3696 3464 3704 3476
rect 3936 3486 3944 3516
rect 4116 3484 4124 3514
rect 4347 3516 4373 3524
rect 4447 3517 4513 3525
rect 4567 3516 4592 3524
rect 4627 3517 4653 3525
rect 4833 3504 4847 3513
rect 4833 3500 4933 3504
rect 4836 3496 4933 3500
rect 4056 3476 4124 3484
rect 4356 3480 4393 3484
rect 4353 3476 4393 3480
rect 4056 3467 4064 3476
rect 3607 3456 3704 3464
rect 3747 3456 3973 3464
rect 4047 3456 4064 3467
rect 4353 3467 4367 3476
rect 4407 3476 4524 3484
rect 4047 3453 4060 3456
rect 4516 3464 4524 3476
rect 4547 3476 4613 3484
rect 4727 3476 4773 3484
rect 4516 3456 4553 3464
rect 4716 3464 4724 3472
rect 4647 3456 4724 3464
rect 67 3436 133 3444
rect 607 3436 673 3444
rect 807 3436 853 3444
rect 1187 3436 1333 3444
rect 1627 3436 1873 3444
rect 1947 3436 2133 3444
rect 2227 3436 2373 3444
rect 2707 3436 2753 3444
rect 3307 3436 3453 3444
rect 4836 3444 4844 3496
rect 4956 3484 4964 3536
rect 5087 3516 5153 3524
rect 5307 3516 5353 3524
rect 5456 3516 5553 3524
rect 5067 3496 5124 3504
rect 5116 3486 5124 3496
rect 4867 3476 4964 3484
rect 5433 3484 5447 3493
rect 5387 3480 5447 3484
rect 5387 3476 5444 3480
rect 5087 3456 5333 3464
rect 5456 3464 5464 3516
rect 5667 3516 5713 3524
rect 5616 3467 5624 3513
rect 5427 3456 5464 3464
rect 5687 3456 5713 3464
rect 4687 3436 4844 3444
rect 796 3424 804 3433
rect 587 3416 804 3424
rect 887 3416 953 3424
rect 1287 3416 1393 3424
rect 1687 3416 1892 3424
rect 1927 3416 2113 3424
rect 2327 3416 2633 3424
rect 2787 3416 2953 3424
rect 3707 3416 3853 3424
rect 3896 3420 4473 3424
rect 3893 3416 4473 3420
rect 3893 3407 3907 3416
rect 5407 3416 5453 3424
rect 5467 3416 5633 3424
rect 487 3396 553 3404
rect 747 3396 773 3404
rect 1367 3396 1684 3404
rect 467 3376 693 3384
rect 1047 3376 1072 3384
rect 1107 3376 1253 3384
rect 1336 3376 1493 3384
rect 1336 3367 1344 3376
rect 1676 3384 1684 3396
rect 1716 3396 1793 3404
rect 1716 3384 1724 3396
rect 2147 3396 2193 3404
rect 2247 3396 2673 3404
rect 3027 3396 3073 3404
rect 3227 3396 3273 3404
rect 3467 3396 3613 3404
rect 3687 3396 3753 3404
rect 4067 3396 4453 3404
rect 4647 3396 4813 3404
rect 4967 3396 5693 3404
rect 1676 3376 1724 3384
rect 1747 3376 1833 3384
rect 2067 3376 2113 3384
rect 2267 3376 2453 3384
rect 2627 3376 2733 3384
rect 2907 3376 2933 3384
rect 2996 3376 3193 3384
rect 47 3356 373 3364
rect 547 3356 833 3364
rect 847 3356 993 3364
rect 1007 3356 1333 3364
rect 1547 3356 1573 3364
rect 1727 3356 1813 3364
rect 1907 3356 2033 3364
rect 2267 3356 2333 3364
rect 2767 3356 2873 3364
rect 2996 3364 3004 3376
rect 3507 3376 3793 3384
rect 3807 3376 3833 3384
rect 3887 3376 4033 3384
rect 4167 3376 4213 3384
rect 4527 3376 4604 3384
rect 2887 3356 3004 3364
rect 3267 3356 3373 3364
rect 3887 3356 3993 3364
rect 4596 3364 4604 3376
rect 4667 3376 4773 3384
rect 4987 3376 5073 3384
rect 4596 3356 4753 3364
rect 4767 3356 4933 3364
rect 4947 3356 5373 3364
rect 107 3336 253 3344
rect 407 3336 513 3344
rect 567 3336 653 3344
rect 747 3336 964 3344
rect 47 3316 73 3324
rect 956 3324 964 3336
rect 987 3336 1133 3344
rect 1387 3336 1553 3344
rect 1767 3336 1793 3344
rect 1907 3336 1933 3344
rect 2067 3336 2353 3344
rect 2467 3336 2693 3344
rect 2867 3336 3353 3344
rect 3567 3336 3713 3344
rect 4107 3336 4233 3344
rect 5007 3336 5233 3344
rect 956 3316 1207 3324
rect 1193 3309 1207 3316
rect 1307 3316 1353 3324
rect 247 3297 333 3305
rect 356 3296 413 3304
rect 356 3284 364 3296
rect 467 3296 524 3304
rect 316 3276 364 3284
rect 516 3284 524 3296
rect 547 3304 560 3307
rect 547 3293 564 3304
rect 587 3296 653 3304
rect 887 3298 933 3306
rect 1047 3304 1060 3307
rect 1047 3293 1064 3304
rect 1087 3296 1124 3304
rect 516 3280 543 3284
rect 516 3276 547 3280
rect 316 3266 324 3276
rect 533 3267 547 3276
rect 27 3256 173 3264
rect 546 3260 547 3267
rect 556 3266 564 3293
rect 607 3256 713 3264
rect 727 3256 773 3264
rect 796 3264 804 3293
rect 1056 3267 1064 3293
rect 796 3256 813 3264
rect 1116 3247 1124 3296
rect 1156 3296 1193 3304
rect 1156 3267 1164 3296
rect 1216 3267 1224 3313
rect 1487 3316 1733 3324
rect 1867 3316 1953 3324
rect 2047 3316 2304 3324
rect 1560 3304 1573 3307
rect 1556 3293 1573 3304
rect 1647 3296 1683 3304
rect 1287 3276 1413 3284
rect 1267 3256 1313 3264
rect 1556 3266 1564 3293
rect 1675 3267 1683 3296
rect 1807 3296 1833 3304
rect 1907 3296 1924 3304
rect 1707 3256 1733 3264
rect 1916 3264 1924 3296
rect 1947 3296 1984 3304
rect 1976 3284 1984 3296
rect 1976 3280 2004 3284
rect 1976 3276 2007 3280
rect 1993 3267 2007 3276
rect 1916 3256 1953 3264
rect 967 3236 1013 3244
rect 1547 3236 1613 3244
rect 1996 3244 2004 3253
rect 1807 3236 2004 3244
rect 287 3216 313 3224
rect 487 3216 653 3224
rect 707 3216 1293 3224
rect 727 3196 973 3204
rect 1367 3196 1433 3204
rect 1707 3196 1953 3204
rect 2016 3204 2024 3295
rect 2176 3296 2212 3304
rect 2076 3267 2084 3293
rect 2176 3284 2184 3296
rect 2156 3276 2184 3284
rect 2156 3267 2164 3276
rect 2067 3256 2084 3267
rect 2067 3253 2080 3256
rect 2147 3256 2164 3267
rect 2236 3264 2244 3293
rect 2296 3267 2304 3316
rect 2727 3316 2933 3324
rect 2447 3296 2544 3304
rect 2536 3284 2544 3296
rect 2567 3296 2733 3304
rect 2336 3280 2544 3284
rect 2333 3276 2544 3280
rect 2333 3267 2347 3276
rect 2536 3267 2544 3276
rect 2596 3267 2604 3296
rect 2827 3296 2844 3304
rect 2176 3260 2244 3264
rect 2173 3256 2244 3260
rect 2147 3253 2160 3256
rect 2173 3247 2187 3256
rect 2387 3256 2473 3264
rect 2647 3256 2673 3264
rect 2476 3244 2484 3253
rect 2836 3247 2844 3296
rect 2856 3267 2864 3316
rect 3487 3316 3653 3324
rect 3987 3324 4000 3327
rect 3987 3313 4004 3324
rect 4027 3316 4053 3324
rect 4747 3316 4793 3324
rect 5547 3316 5613 3324
rect 2987 3296 3113 3304
rect 3327 3296 3444 3304
rect 2896 3267 2904 3293
rect 3273 3284 3287 3293
rect 3273 3280 3304 3284
rect 3276 3276 3307 3280
rect 3293 3267 3307 3276
rect 3436 3266 3444 3296
rect 3687 3297 3732 3305
rect 3867 3297 3933 3305
rect 3996 3304 4004 3313
rect 3996 3296 4053 3304
rect 3516 3267 3524 3293
rect 3633 3284 3647 3293
rect 3556 3280 3647 3284
rect 3556 3276 3644 3280
rect 3556 3267 3564 3276
rect 3547 3256 3564 3267
rect 3547 3253 3560 3256
rect 3587 3255 3653 3263
rect 3756 3264 3764 3293
rect 3836 3284 3844 3294
rect 4176 3296 4213 3304
rect 4176 3284 4184 3296
rect 4307 3296 4373 3304
rect 4627 3297 4693 3305
rect 4767 3304 4780 3307
rect 4767 3293 4784 3304
rect 4836 3296 4893 3304
rect 3836 3276 4184 3284
rect 4396 3280 4573 3284
rect 4393 3276 4573 3280
rect 3756 3256 3893 3264
rect 4076 3266 4084 3276
rect 4393 3267 4407 3276
rect 4776 3284 4784 3293
rect 4816 3284 4824 3294
rect 4776 3276 4824 3284
rect 4836 3267 4844 3296
rect 5167 3296 5233 3304
rect 5247 3296 5333 3304
rect 5507 3296 5693 3304
rect 4956 3267 4964 3293
rect 4267 3256 4353 3264
rect 5367 3256 5393 3264
rect 2476 3236 2573 3244
rect 2587 3236 2713 3244
rect 2836 3246 2860 3247
rect 2836 3236 2853 3246
rect 2840 3233 2853 3236
rect 2967 3236 3453 3244
rect 3627 3236 3673 3244
rect 3687 3236 3813 3244
rect 4627 3236 4913 3244
rect 5487 3236 5593 3244
rect 2147 3216 2213 3224
rect 2287 3216 2413 3224
rect 3167 3216 3393 3224
rect 3527 3216 3593 3224
rect 3907 3216 4153 3224
rect 4247 3216 4953 3224
rect 2016 3196 2084 3204
rect 527 3176 873 3184
rect 1007 3176 1453 3184
rect 1667 3176 1833 3184
rect 2007 3176 2053 3184
rect 2076 3184 2084 3196
rect 2167 3196 2253 3204
rect 2587 3196 2793 3204
rect 2947 3196 3133 3204
rect 3467 3196 3853 3204
rect 4027 3196 4113 3204
rect 4227 3196 5193 3204
rect 5347 3196 5533 3204
rect 2076 3176 2253 3184
rect 3267 3176 3433 3184
rect 3447 3176 3873 3184
rect 3927 3176 4293 3184
rect 4507 3180 5084 3184
rect 4507 3176 5087 3180
rect 247 3156 273 3164
rect 287 3156 2092 3164
rect 2127 3156 2273 3164
rect 2407 3156 2913 3164
rect 3067 3156 3353 3164
rect 3367 3156 3473 3164
rect 3487 3156 3533 3164
rect 3916 3164 3924 3173
rect 3647 3156 3924 3164
rect 5073 3167 5087 3176
rect 5287 3176 5313 3184
rect 307 3136 613 3144
rect 667 3136 733 3144
rect 1027 3136 1793 3144
rect 2276 3144 2284 3153
rect 1847 3136 2164 3144
rect 2276 3136 2633 3144
rect 387 3116 713 3124
rect 987 3116 1693 3124
rect 1907 3116 2004 3124
rect 27 3096 293 3104
rect 427 3096 433 3104
rect 447 3096 673 3104
rect 747 3096 1373 3104
rect 1996 3104 2004 3116
rect 2027 3116 2073 3124
rect 2156 3124 2164 3136
rect 2647 3136 2753 3144
rect 2867 3136 4993 3144
rect 5007 3136 5273 3144
rect 5287 3136 5433 3144
rect 2156 3116 2573 3124
rect 2627 3116 2833 3124
rect 3127 3116 4213 3124
rect 4307 3116 4593 3124
rect 4807 3116 4933 3124
rect 1996 3096 2593 3104
rect 2727 3096 2873 3104
rect 3147 3096 3293 3104
rect 3827 3096 4193 3104
rect 4547 3096 4673 3104
rect 467 3076 593 3084
rect 1227 3076 1253 3084
rect 1987 3076 2173 3084
rect 2187 3076 2313 3084
rect 3367 3076 3553 3084
rect 3567 3076 3693 3084
rect 3927 3076 4233 3084
rect 4487 3076 4973 3084
rect 5127 3076 5493 3084
rect 147 3056 373 3064
rect 447 3056 533 3064
rect 647 3056 713 3064
rect 756 3056 993 3064
rect -24 3036 13 3044
rect 87 3036 113 3044
rect 756 3044 764 3056
rect 1287 3056 1373 3064
rect 1387 3056 1473 3064
rect 1496 3056 1953 3064
rect 607 3036 764 3044
rect 1496 3044 1504 3056
rect 2007 3056 2052 3064
rect 2087 3056 2624 3064
rect 1307 3036 1504 3044
rect 2616 3044 2624 3056
rect 3687 3056 3804 3064
rect 2616 3036 2893 3044
rect 2987 3036 3173 3044
rect 3796 3044 3804 3056
rect 3907 3056 4293 3064
rect 5527 3056 5553 3064
rect 3796 3036 4033 3044
rect 3936 3027 3944 3036
rect 4407 3036 4633 3044
rect 187 3016 233 3024
rect 387 3016 473 3024
rect 527 3016 564 3024
rect -24 2996 13 3004
rect 76 2967 84 2994
rect 420 3004 433 3007
rect 416 2993 433 3004
rect 156 2967 164 2993
rect 67 2956 84 2967
rect 67 2953 80 2956
rect 416 2964 424 2993
rect 407 2956 424 2964
rect 467 2954 533 2962
rect 556 2947 564 3016
rect 887 3016 953 3024
rect 1267 3016 1413 3024
rect 2147 3016 2184 3024
rect 687 2997 733 3005
rect 827 2997 873 3005
rect 576 2967 584 2993
rect 636 2984 644 2994
rect 776 2984 784 2994
rect 1173 3004 1187 3013
rect 1173 3000 1313 3004
rect 1176 2996 1313 3000
rect 1327 2996 1393 3004
rect 636 2980 704 2984
rect 636 2976 707 2980
rect 776 2976 844 2984
rect 693 2967 707 2976
rect 747 2956 793 2964
rect 836 2964 844 2976
rect 836 2956 893 2964
rect 1013 2964 1027 2973
rect 947 2960 1027 2964
rect 947 2956 1024 2960
rect 1187 2954 1353 2962
rect 1376 2947 1384 2996
rect 1447 2996 1653 3004
rect 1836 3000 1893 3004
rect 1833 2996 1893 3000
rect 1833 2986 1847 2996
rect 2046 2994 2047 3008
rect 1427 2956 1853 2964
rect 1867 2956 1893 2964
rect 1956 2964 1964 2993
rect 2036 2984 2044 2994
rect 2067 2996 2153 3004
rect 2036 2976 2104 2984
rect 2096 2964 2104 2976
rect 1956 2956 2024 2964
rect 2096 2956 2133 2964
rect 47 2936 133 2944
rect 627 2936 713 2944
rect 887 2936 913 2944
rect 1647 2936 1913 2944
rect 2016 2944 2024 2956
rect 2176 2947 2184 3016
rect 2387 3016 2473 3024
rect 3927 3016 3944 3027
rect 3927 3013 3940 3016
rect 4987 3016 5093 3024
rect 5200 3024 5213 3027
rect 5196 3013 5213 3024
rect 5547 3016 5673 3024
rect 2687 2996 2784 3004
rect 2216 2967 2224 2993
rect 2436 2964 2444 2994
rect 2367 2956 2444 2964
rect 2567 2956 2713 2964
rect 2776 2964 2784 2996
rect 2807 2996 2833 3004
rect 2847 2996 2873 3004
rect 2927 2996 3053 3004
rect 3127 2997 3233 3005
rect 3056 2984 3064 2994
rect 3056 2976 3124 2984
rect 2776 2956 2853 2964
rect 2907 2956 2952 2964
rect 2987 2955 3033 2963
rect 3116 2964 3124 2976
rect 3116 2956 3144 2964
rect 2016 2936 2073 2944
rect 2167 2936 2184 2947
rect 2167 2933 2180 2936
rect 2247 2936 2293 2944
rect 3136 2944 3144 2956
rect 3307 2955 3353 2963
rect 3376 2964 3384 3013
rect 3447 2996 3493 3004
rect 3727 2997 3753 3005
rect 3827 2996 3944 3004
rect 3716 2984 3724 2994
rect 3696 2976 3724 2984
rect 3696 2966 3704 2976
rect 3936 2966 3944 2996
rect 4196 2996 4293 3004
rect 3376 2956 3453 2964
rect 3507 2954 3533 2962
rect 3787 2955 3873 2963
rect 4196 2965 4204 2996
rect 4316 2996 4393 3004
rect 4316 2966 4324 2996
rect 4447 2996 4533 3004
rect 4576 2947 4584 2994
rect 4607 2956 4633 2964
rect 4647 2956 4673 2964
rect 4847 2956 4873 2964
rect 4887 2956 5033 2964
rect 5047 2956 5093 2964
rect 3136 2936 3173 2944
rect 3567 2936 3593 2944
rect 4267 2936 4413 2944
rect 267 2916 492 2924
rect 616 2924 624 2933
rect 527 2916 624 2924
rect 1567 2916 1613 2924
rect 1627 2916 1993 2924
rect 2107 2916 2633 2924
rect 2867 2916 3093 2924
rect 3427 2916 4133 2924
rect 4387 2916 4473 2924
rect 4727 2916 5113 2924
rect 5127 2916 5153 2924
rect 5196 2924 5204 3013
rect 5216 2996 5313 3004
rect 5216 2966 5224 2996
rect 5467 2996 5804 3004
rect 5247 2936 5413 2944
rect 5196 2916 5272 2924
rect 5307 2916 5513 2924
rect 207 2896 433 2904
rect 547 2896 853 2904
rect 907 2896 1053 2904
rect 1556 2904 1564 2913
rect 1407 2896 1564 2904
rect 2327 2896 2593 2904
rect 4587 2896 4773 2904
rect 4787 2896 4913 2904
rect 4927 2896 5333 2904
rect 427 2876 693 2884
rect 1227 2876 1773 2884
rect 1827 2876 1973 2884
rect 3127 2876 3333 2884
rect 4087 2876 4113 2884
rect 4127 2876 4553 2884
rect 5227 2876 5313 2884
rect 447 2856 653 2864
rect 1447 2856 1713 2864
rect 1807 2856 1873 2864
rect 2187 2856 2353 2864
rect 2847 2856 2913 2864
rect 3087 2856 3493 2864
rect 4147 2856 5233 2864
rect 1087 2836 1173 2844
rect 1467 2836 1633 2844
rect 1927 2836 2113 2844
rect 2607 2836 2753 2844
rect 3107 2836 3453 2844
rect 5127 2836 5273 2844
rect 5367 2836 5533 2844
rect 107 2816 173 2824
rect 227 2816 273 2824
rect 867 2816 1033 2824
rect 1047 2816 1233 2824
rect 1727 2816 1873 2824
rect 2147 2816 2313 2824
rect 2687 2816 2773 2824
rect 3787 2816 3933 2824
rect 3947 2816 4033 2824
rect 4127 2816 4193 2824
rect 4367 2816 4693 2824
rect 5387 2816 5513 2824
rect 47 2796 73 2804
rect 247 2796 313 2804
rect 327 2796 353 2804
rect 1387 2796 1424 2804
rect 140 2784 153 2787
rect 116 2747 124 2775
rect 136 2773 153 2784
rect 336 2776 473 2784
rect 136 2747 144 2773
rect 47 2736 92 2744
rect 196 2744 204 2773
rect 336 2747 344 2776
rect 496 2776 593 2784
rect 496 2764 504 2776
rect 456 2756 504 2764
rect 196 2736 213 2744
rect 136 2724 144 2733
rect 267 2736 333 2744
rect 456 2746 464 2756
rect 636 2747 644 2775
rect 707 2776 733 2784
rect 776 2744 784 2775
rect 927 2777 953 2785
rect 976 2776 993 2784
rect 976 2764 984 2776
rect 1116 2776 1253 2784
rect 1033 2764 1047 2773
rect 896 2760 984 2764
rect 893 2756 984 2760
rect 1016 2760 1047 2764
rect 1016 2756 1044 2760
rect 893 2747 907 2756
rect 667 2736 872 2744
rect 1016 2746 1024 2756
rect 1096 2747 1104 2774
rect 1087 2736 1104 2747
rect 1087 2733 1100 2736
rect 1116 2727 1124 2776
rect 1276 2776 1353 2784
rect 1276 2764 1284 2776
rect 1256 2760 1284 2764
rect 1253 2756 1284 2760
rect 1253 2747 1267 2756
rect 1416 2747 1424 2796
rect 1467 2796 1493 2804
rect 1667 2796 1693 2804
rect 1907 2796 1933 2804
rect 1947 2796 2113 2804
rect 2127 2796 2593 2804
rect 2767 2796 2964 2804
rect 1527 2776 1593 2784
rect 1696 2776 1773 2784
rect 1696 2747 1704 2776
rect 1547 2736 1573 2744
rect 1587 2736 1633 2744
rect 1796 2744 1804 2793
rect 1827 2776 1904 2784
rect 1796 2736 1833 2744
rect 1896 2746 1904 2776
rect 2047 2776 2224 2784
rect 2216 2764 2224 2776
rect 2307 2777 2433 2785
rect 2527 2776 2593 2784
rect 2216 2756 2244 2764
rect 1947 2736 1973 2744
rect 2147 2736 2193 2744
rect 2236 2746 2244 2756
rect 2256 2744 2264 2774
rect 2747 2776 2933 2784
rect 2256 2736 2393 2744
rect 2447 2736 2613 2744
rect 2676 2744 2684 2773
rect 2696 2764 2704 2774
rect 2956 2784 2964 2796
rect 4167 2804 4180 2807
rect 4167 2794 4184 2804
rect 4160 2793 4184 2794
rect 4967 2796 5073 2804
rect 5176 2796 5253 2804
rect 2956 2776 2993 2784
rect 3007 2776 3053 2784
rect 3667 2778 3713 2786
rect 4056 2776 4153 2784
rect 2696 2756 3033 2764
rect 3773 2764 3787 2773
rect 3756 2760 3787 2764
rect 3756 2756 3784 2760
rect 2676 2736 2753 2744
rect 2887 2735 2933 2743
rect 3067 2736 3093 2744
rect 3367 2736 3453 2744
rect 3467 2736 3553 2744
rect 3756 2744 3764 2756
rect 3707 2736 3764 2744
rect 3816 2744 3824 2774
rect 3787 2736 3824 2744
rect 4056 2744 4064 2776
rect 4176 2746 4184 2793
rect 4287 2777 4333 2785
rect 4567 2776 4613 2784
rect 3967 2736 4064 2744
rect 4347 2736 4533 2744
rect 4656 2744 4664 2774
rect 4767 2776 4833 2784
rect 4927 2776 4973 2784
rect 5176 2747 5184 2796
rect 5607 2796 5644 2804
rect 5260 2784 5273 2787
rect 5256 2773 5273 2784
rect 5447 2777 5573 2785
rect 5256 2747 5264 2773
rect 4587 2736 4664 2744
rect 4827 2736 5033 2744
rect 5107 2736 5133 2744
rect 5316 2744 5324 2773
rect 5636 2747 5644 2796
rect 5667 2776 5733 2784
rect 5316 2736 5493 2744
rect 5687 2736 5804 2744
rect 136 2716 373 2724
rect 627 2716 984 2724
rect 976 2707 984 2716
rect 1107 2716 1124 2727
rect 1107 2713 1120 2716
rect 2027 2716 2073 2724
rect 2087 2716 2273 2724
rect 2627 2716 2653 2724
rect 3047 2716 3133 2724
rect 3867 2716 4033 2724
rect 4047 2716 4213 2724
rect 4227 2716 4793 2724
rect 4807 2716 5053 2724
rect 5067 2716 5333 2724
rect 5347 2716 5433 2724
rect 427 2696 493 2704
rect 647 2696 793 2704
rect 987 2696 1113 2704
rect 1427 2696 1673 2704
rect 2667 2696 2813 2704
rect 2827 2696 3213 2704
rect 3227 2696 3253 2704
rect 3767 2696 3993 2704
rect 4627 2696 4713 2704
rect 4787 2696 4853 2704
rect 5007 2696 5152 2704
rect 5187 2696 5373 2704
rect 5627 2696 5673 2704
rect 1287 2676 1933 2684
rect 4896 2676 4953 2684
rect 987 2656 1053 2664
rect 1067 2656 1453 2664
rect 2547 2656 2913 2664
rect 4507 2656 4673 2664
rect 4896 2664 4904 2676
rect 4767 2656 4904 2664
rect 5047 2656 5193 2664
rect 27 2636 933 2644
rect 1127 2636 1213 2644
rect 1267 2636 1373 2644
rect 1507 2636 1713 2644
rect 1727 2636 2553 2644
rect 4027 2636 4313 2644
rect 4927 2636 5533 2644
rect 207 2616 553 2624
rect 967 2616 1073 2624
rect 1087 2616 1593 2624
rect 1807 2616 2153 2624
rect 2327 2616 2453 2624
rect 2467 2616 2653 2624
rect 1147 2596 1253 2604
rect 1347 2596 1493 2604
rect 2147 2596 2713 2604
rect 5436 2596 5593 2604
rect 767 2576 973 2584
rect 1187 2576 3233 2584
rect 3627 2576 4273 2584
rect 4287 2576 4433 2584
rect 4447 2576 4473 2584
rect 5436 2584 5444 2596
rect 4587 2576 5444 2584
rect 47 2556 173 2564
rect 1007 2556 1113 2564
rect 1227 2556 2533 2564
rect 4427 2556 4553 2564
rect 5416 2560 5493 2564
rect 5413 2556 5493 2560
rect 5413 2547 5427 2556
rect 1587 2536 1693 2544
rect 1847 2536 1913 2544
rect 4087 2536 4113 2544
rect 5127 2536 5253 2544
rect 287 2516 413 2524
rect 667 2516 753 2524
rect 767 2516 893 2524
rect 1147 2516 1193 2524
rect 1307 2516 1453 2524
rect 1567 2516 1813 2524
rect 2207 2516 2293 2524
rect 2307 2516 2513 2524
rect 3407 2516 3533 2524
rect 4007 2516 4173 2524
rect 4307 2516 4373 2524
rect 4447 2516 4693 2524
rect 4707 2516 5164 2524
rect 5156 2507 5164 2516
rect 5447 2516 5553 2524
rect 5567 2516 5693 2524
rect 927 2496 1113 2504
rect 1487 2496 1613 2504
rect 1887 2496 1993 2504
rect 2007 2496 2273 2504
rect 2287 2496 2473 2504
rect 2487 2496 2673 2504
rect 3136 2496 3313 2504
rect 80 2484 93 2487
rect 76 2473 93 2484
rect 147 2476 193 2484
rect 387 2476 433 2484
rect 76 2447 84 2473
rect 296 2447 304 2473
rect 316 2464 324 2474
rect 627 2476 793 2484
rect 807 2476 893 2484
rect 1160 2484 1173 2487
rect 1156 2473 1173 2484
rect 1227 2476 1284 2484
rect 316 2456 344 2464
rect 67 2436 84 2447
rect 67 2433 80 2436
rect 127 2436 213 2444
rect 336 2444 344 2456
rect 1156 2447 1164 2473
rect 336 2436 364 2444
rect 356 2427 364 2436
rect 647 2434 693 2442
rect 707 2436 773 2444
rect 927 2435 1053 2443
rect 1276 2446 1284 2476
rect 1427 2477 1553 2485
rect 1356 2447 1364 2474
rect 1687 2476 1713 2484
rect 1940 2484 1953 2487
rect 1787 2476 1844 2484
rect 1836 2447 1844 2476
rect 1936 2473 1953 2484
rect 2016 2476 2053 2484
rect 1247 2436 1273 2444
rect 1347 2436 1364 2447
rect 1347 2433 1360 2436
rect 1547 2435 1633 2443
rect 1647 2436 1692 2444
rect 1727 2435 1753 2443
rect 1936 2445 1944 2473
rect 2016 2464 2024 2476
rect 2167 2477 2232 2485
rect 2267 2477 2333 2485
rect 2347 2476 2433 2484
rect 2456 2476 2573 2484
rect 2456 2464 2464 2476
rect 2767 2476 2793 2484
rect 2916 2476 2993 2484
rect 1987 2456 2024 2464
rect 2416 2456 2464 2464
rect 2087 2436 2233 2444
rect 2416 2446 2424 2456
rect 2916 2447 2924 2476
rect 3136 2487 3144 2496
rect 3387 2504 3400 2507
rect 3387 2493 3404 2504
rect 4067 2496 4133 2504
rect 4347 2496 4444 2504
rect 5156 2496 5173 2507
rect 3107 2476 3132 2484
rect 3167 2477 3193 2485
rect 3216 2476 3293 2484
rect 3036 2447 3044 2473
rect 2247 2436 2353 2444
rect 2367 2436 2413 2444
rect 2527 2436 2813 2444
rect 3216 2446 3224 2476
rect 3356 2444 3364 2473
rect 3396 2464 3404 2493
rect 3627 2477 3653 2485
rect 3727 2477 3753 2485
rect 3947 2476 3973 2484
rect 4047 2476 4224 2484
rect 3396 2456 3424 2464
rect 3416 2446 3424 2456
rect 3267 2436 3364 2444
rect 3847 2436 3913 2444
rect 4216 2445 4224 2476
rect 4247 2476 4364 2484
rect 4356 2445 4364 2476
rect 4436 2447 4444 2496
rect 5160 2493 5173 2496
rect 5187 2500 5404 2504
rect 5187 2496 5407 2500
rect 4767 2477 4813 2485
rect 4516 2464 4524 2474
rect 4947 2476 4973 2484
rect 5247 2477 5273 2485
rect 5393 2487 5407 2496
rect 5433 2464 5447 2473
rect 4516 2456 4704 2464
rect 3987 2434 4013 2442
rect 4107 2434 4133 2442
rect 4696 2444 4704 2456
rect 5356 2460 5447 2464
rect 5456 2476 5513 2484
rect 5356 2456 5444 2460
rect 4696 2436 4733 2444
rect 5356 2446 5364 2456
rect 5456 2447 5464 2476
rect 5607 2476 5713 2484
rect 5727 2476 5753 2484
rect 4947 2435 5053 2443
rect 5447 2436 5464 2447
rect 5447 2433 5460 2436
rect 356 2416 373 2427
rect 360 2413 373 2416
rect 416 2416 553 2424
rect 416 2404 424 2416
rect 887 2416 953 2424
rect 1827 2416 1893 2424
rect 2567 2416 2753 2424
rect 2987 2416 3133 2424
rect 4887 2416 4993 2424
rect 5427 2416 5573 2424
rect 87 2396 424 2404
rect 987 2396 1033 2404
rect 1207 2396 1653 2404
rect 1667 2396 1793 2404
rect 1847 2396 1873 2404
rect 1887 2396 2033 2404
rect 2556 2404 2564 2413
rect 2427 2396 2564 2404
rect 3207 2396 3473 2404
rect 3767 2396 4053 2404
rect 4407 2396 4573 2404
rect 4827 2396 5093 2404
rect 627 2376 733 2384
rect 847 2376 953 2384
rect 1427 2376 1453 2384
rect 2827 2376 3073 2384
rect 3167 2376 3333 2384
rect 47 2356 113 2364
rect 227 2356 413 2364
rect 527 2356 1004 2364
rect 996 2347 1004 2356
rect 1347 2356 1393 2364
rect 2027 2356 2173 2364
rect 2567 2356 2633 2364
rect 1007 2336 1153 2344
rect 1707 2336 1813 2344
rect 2007 2336 2093 2344
rect 2347 2336 2513 2344
rect 2727 2336 2873 2344
rect 3267 2336 3333 2344
rect 4187 2336 4273 2344
rect 5287 2336 5473 2344
rect 267 2316 484 2324
rect 147 2296 293 2304
rect 476 2304 484 2316
rect 527 2316 593 2324
rect 687 2316 973 2324
rect 1027 2316 1313 2324
rect 1367 2316 1573 2324
rect 1807 2316 2133 2324
rect 3356 2316 3773 2324
rect 476 2296 693 2304
rect 867 2296 933 2304
rect 1267 2296 1333 2304
rect 1687 2296 1713 2304
rect 1896 2296 2233 2304
rect 447 2276 733 2284
rect 967 2276 1013 2284
rect 1896 2284 1904 2296
rect 2247 2296 2373 2304
rect 2467 2296 2573 2304
rect 2787 2296 2853 2304
rect 3356 2304 3364 2316
rect 5007 2316 5113 2324
rect 5547 2316 5673 2324
rect 3287 2296 3364 2304
rect 5047 2296 5233 2304
rect 5527 2296 5573 2304
rect 1607 2276 1904 2284
rect 2267 2284 2280 2287
rect 2267 2273 2284 2284
rect 2927 2276 2953 2284
rect 4027 2276 4233 2284
rect 4247 2276 4273 2284
rect 4667 2276 4893 2284
rect 4907 2276 5073 2284
rect 107 2256 173 2264
rect 115 2227 123 2256
rect 227 2256 284 2264
rect 276 2227 284 2256
rect 356 2227 364 2255
rect 427 2256 473 2264
rect 787 2258 913 2266
rect 1167 2257 1293 2265
rect 1427 2257 1553 2265
rect 1687 2264 1700 2267
rect 1687 2253 1704 2264
rect 1727 2256 1773 2264
rect 676 2227 684 2253
rect 1696 2227 1704 2253
rect 47 2216 73 2224
rect 147 2216 193 2224
rect 376 2216 493 2224
rect 376 2204 384 2216
rect 507 2216 593 2224
rect 787 2216 833 2224
rect 927 2216 973 2224
rect 1107 2216 1253 2224
rect 1327 2216 1344 2224
rect 347 2196 384 2204
rect 467 2196 753 2204
rect 1336 2204 1344 2216
rect 1467 2215 1573 2223
rect 1916 2224 1924 2254
rect 2007 2256 2053 2264
rect 2167 2256 2213 2264
rect 2093 2244 2107 2253
rect 2093 2240 2124 2244
rect 2096 2236 2127 2240
rect 2113 2227 2127 2236
rect 1747 2216 1924 2224
rect 1947 2216 2033 2224
rect 2276 2226 2284 2273
rect 2440 2264 2453 2267
rect 2436 2253 2453 2264
rect 2476 2256 2553 2264
rect 2436 2224 2444 2253
rect 2476 2244 2484 2256
rect 2596 2256 2613 2264
rect 2456 2240 2484 2244
rect 2407 2216 2444 2224
rect 2453 2236 2484 2240
rect 2496 2236 2573 2244
rect 2453 2227 2467 2236
rect 2496 2226 2504 2236
rect 2596 2227 2604 2256
rect 2816 2227 2824 2254
rect 2887 2256 3273 2264
rect 3413 2264 3427 2273
rect 3387 2260 3427 2264
rect 3387 2256 3424 2260
rect 3336 2244 3344 2254
rect 3447 2256 3513 2264
rect 3887 2257 3933 2265
rect 3336 2236 3464 2244
rect 2707 2215 2753 2223
rect 2816 2216 2832 2227
rect 2820 2213 2832 2216
rect 2867 2216 3073 2224
rect 3407 2215 3433 2223
rect 3456 2224 3464 2236
rect 3456 2216 3493 2224
rect 3576 2224 3584 2254
rect 4307 2256 4353 2264
rect 4376 2256 4453 2264
rect 4376 2244 4384 2256
rect 4336 2240 4384 2244
rect 4333 2236 4384 2240
rect 4616 2244 4624 2255
rect 4847 2256 4953 2264
rect 5167 2257 5193 2265
rect 5487 2257 5533 2265
rect 5620 2264 5633 2267
rect 4616 2236 4673 2244
rect 4333 2227 4347 2236
rect 5316 2244 5324 2254
rect 5616 2253 5633 2264
rect 5316 2240 5444 2244
rect 5316 2236 5447 2240
rect 5433 2227 5447 2236
rect 5616 2227 5624 2253
rect 3547 2216 3584 2224
rect 3676 2216 3753 2224
rect 1336 2196 1413 2204
rect 1427 2196 1493 2204
rect 2547 2196 2573 2204
rect 2807 2196 2893 2204
rect 3676 2204 3684 2216
rect 3567 2196 3684 2204
rect 3867 2216 3993 2224
rect 4387 2216 4433 2224
rect 4507 2216 4573 2224
rect 4707 2215 4733 2223
rect 4787 2216 4833 2224
rect 4847 2215 4873 2223
rect 5107 2216 5153 2224
rect 3753 2204 3767 2212
rect 5656 2207 5664 2273
rect 5696 2227 5704 2273
rect 3753 2196 4053 2204
rect 4987 2196 5033 2204
rect 5656 2196 5673 2207
rect 5660 2193 5673 2196
rect 727 2176 933 2184
rect 1027 2176 1393 2184
rect 1627 2176 1773 2184
rect 1787 2176 2133 2184
rect 3467 2176 3693 2184
rect 3947 2176 4113 2184
rect 4447 2176 4533 2184
rect 5287 2176 5553 2184
rect 567 2156 873 2164
rect 987 2156 1453 2164
rect 2227 2156 3353 2164
rect 4287 2156 4373 2164
rect 787 2136 1153 2144
rect 1827 2136 1953 2144
rect 2007 2136 2173 2144
rect 2667 2136 3033 2144
rect 3047 2136 3344 2144
rect 3336 2124 3344 2136
rect 5067 2136 5133 2144
rect 5147 2136 5453 2144
rect 3336 2116 3433 2124
rect 4307 2116 4673 2124
rect 4687 2116 4813 2124
rect 4827 2116 5373 2124
rect 5447 2116 5653 2124
rect 1887 2096 2073 2104
rect 3967 2096 4093 2104
rect 5227 2096 5313 2104
rect 267 2076 353 2084
rect 2687 2076 2833 2084
rect 2847 2076 3233 2084
rect 3247 2076 3793 2084
rect 207 2056 453 2064
rect 547 2056 1013 2064
rect 1347 2056 1673 2064
rect 3167 2056 3553 2064
rect 4047 2060 4544 2064
rect 4047 2056 4547 2060
rect 4533 2047 4547 2056
rect 5307 2056 5433 2064
rect 87 2036 113 2044
rect 1007 2036 1133 2044
rect 1307 2036 1773 2044
rect 1867 2036 2013 2044
rect 3667 2036 3993 2044
rect 4667 2036 5013 2044
rect 47 2016 233 2024
rect 527 2016 793 2024
rect 807 2016 2484 2024
rect 2476 2007 2484 2016
rect 2887 2016 3073 2024
rect 3547 2016 3573 2024
rect 4287 2016 4313 2024
rect 4627 2016 4933 2024
rect 5367 2016 5413 2024
rect 27 1996 373 2004
rect 1727 1996 1913 2004
rect 2487 1996 2593 2004
rect 2867 1996 3193 2004
rect 3207 1996 3393 2004
rect 3847 1996 3953 2004
rect 4867 1996 5293 2004
rect 5607 1996 5733 2004
rect 1507 1976 2113 1984
rect 2387 1976 2413 1984
rect 2556 1976 2793 1984
rect -24 1956 13 1964
rect 127 1956 193 1964
rect 327 1957 393 1965
rect 407 1957 433 1965
rect 500 1964 513 1967
rect 496 1953 513 1964
rect 627 1957 653 1965
rect 256 1925 264 1953
rect 496 1926 504 1953
rect 47 1916 93 1924
rect 407 1896 433 1904
rect 556 1904 564 1954
rect 887 1956 913 1964
rect 1167 1957 1233 1965
rect 836 1927 844 1953
rect 827 1916 844 1927
rect 827 1913 840 1916
rect 956 1924 964 1954
rect 1527 1956 1693 1964
rect 2040 1964 2053 1967
rect 1847 1956 1884 1964
rect 1353 1944 1367 1953
rect 1353 1940 1384 1944
rect 1356 1936 1384 1940
rect 867 1916 964 1924
rect 1087 1916 1133 1924
rect 1267 1916 1353 1924
rect 1376 1924 1384 1936
rect 1876 1927 1884 1956
rect 2036 1953 2053 1964
rect 2107 1956 2153 1964
rect 2556 1967 2564 1976
rect 2907 1984 2920 1987
rect 2907 1973 2924 1984
rect 3507 1976 3633 1984
rect 3647 1976 3793 1984
rect 4187 1976 4213 1984
rect 4227 1976 4313 1984
rect 4487 1976 4653 1984
rect 5027 1976 5193 1984
rect 5207 1976 5273 1984
rect 5407 1984 5420 1987
rect 5407 1973 5424 1984
rect 2367 1956 2453 1964
rect 2467 1956 2513 1964
rect 2607 1956 2633 1964
rect 2820 1964 2833 1967
rect 1376 1916 1473 1924
rect 1807 1914 1833 1922
rect 447 1896 564 1904
rect 627 1896 773 1904
rect 1167 1896 1233 1904
rect 2036 1904 2044 1953
rect 2256 1927 2264 1953
rect 2316 1927 2324 1953
rect 2247 1916 2264 1927
rect 2247 1913 2260 1916
rect 2367 1916 2393 1924
rect 2556 1924 2564 1953
rect 2447 1916 2564 1924
rect 2696 1924 2704 1953
rect 2667 1916 2704 1924
rect 2756 1907 2764 1954
rect 2816 1953 2833 1964
rect 2816 1926 2824 1953
rect 2876 1927 2884 1953
rect 2916 1927 2924 1973
rect 3207 1956 3233 1964
rect 3287 1956 3313 1964
rect 3687 1956 3724 1964
rect 2916 1916 2933 1927
rect 2920 1913 2933 1916
rect 3655 1925 3663 1953
rect 3716 1926 3724 1956
rect 3787 1957 3893 1965
rect 4056 1956 4133 1964
rect 3207 1914 3233 1922
rect 3727 1916 3813 1924
rect 4056 1926 4064 1956
rect 4647 1964 4660 1967
rect 4647 1953 4664 1964
rect 4687 1956 4713 1964
rect 4960 1964 4973 1967
rect 4656 1926 4664 1953
rect 3967 1916 4013 1924
rect 4727 1915 4753 1923
rect 4776 1924 4784 1954
rect 4956 1953 4973 1964
rect 5387 1964 5400 1967
rect 5387 1953 5404 1964
rect 4956 1926 4964 1953
rect 5313 1944 5327 1953
rect 5313 1940 5344 1944
rect 5316 1936 5347 1940
rect 5333 1927 5347 1936
rect 4776 1916 4804 1924
rect 4796 1907 4804 1916
rect 5147 1915 5173 1923
rect 5396 1926 5404 1953
rect 5416 1944 5424 1973
rect 5416 1936 5444 1944
rect 1907 1896 2044 1904
rect 2827 1896 2853 1904
rect 2967 1896 3013 1904
rect 4796 1896 4813 1907
rect 4800 1893 4813 1896
rect 4953 1904 4967 1912
rect 5436 1907 5444 1936
rect 5456 1927 5464 1954
rect 5456 1916 5473 1927
rect 5460 1913 5473 1916
rect 5547 1915 5613 1923
rect 5627 1916 5753 1924
rect 4953 1896 5033 1904
rect 5227 1896 5264 1904
rect 107 1876 173 1884
rect 687 1876 773 1884
rect 1847 1876 1933 1884
rect 2787 1876 2873 1884
rect 3807 1876 4053 1884
rect 4427 1876 4453 1884
rect 4796 1876 4853 1884
rect 667 1856 973 1864
rect 1227 1856 1293 1864
rect 1776 1856 1924 1864
rect 1776 1847 1784 1856
rect 1627 1836 1773 1844
rect 1916 1844 1924 1856
rect 1956 1856 2253 1864
rect 1956 1844 1964 1856
rect 2447 1856 2933 1864
rect 3247 1856 3993 1864
rect 4796 1864 4804 1876
rect 5256 1884 5264 1896
rect 5427 1896 5444 1907
rect 5427 1893 5440 1896
rect 5256 1876 5373 1884
rect 4427 1856 4804 1864
rect 5047 1856 5433 1864
rect 1916 1836 1964 1844
rect 2927 1836 3013 1844
rect 3727 1836 3773 1844
rect 5087 1836 5193 1844
rect 387 1816 413 1824
rect 767 1816 913 1824
rect 1367 1816 1413 1824
rect 1427 1816 1553 1824
rect 1567 1816 1633 1824
rect 1767 1816 1913 1824
rect 2047 1816 2844 1824
rect 2187 1796 2233 1804
rect 2836 1804 2844 1816
rect 2867 1816 3313 1824
rect 3327 1816 4173 1824
rect 4187 1816 4333 1824
rect 2836 1796 4493 1804
rect 4927 1796 5173 1804
rect 927 1776 1192 1784
rect 1227 1776 1313 1784
rect 1447 1776 1713 1784
rect 1867 1776 2013 1784
rect 2507 1776 2532 1784
rect 2567 1776 2793 1784
rect 2947 1776 3013 1784
rect 3107 1776 3713 1784
rect 4547 1776 4653 1784
rect 747 1756 813 1764
rect 827 1756 1013 1764
rect 1607 1756 1753 1764
rect 1967 1756 2113 1764
rect 2207 1756 2453 1764
rect 2467 1756 2853 1764
rect 3187 1756 3313 1764
rect 4507 1756 4773 1764
rect 4787 1756 4963 1764
rect 47 1737 113 1745
rect 467 1737 493 1745
rect 593 1744 607 1753
rect 567 1740 607 1744
rect 567 1736 604 1740
rect 647 1737 693 1745
rect 807 1736 993 1744
rect 1096 1736 1153 1744
rect 236 1704 244 1733
rect 927 1720 1064 1724
rect 927 1716 1067 1720
rect 1053 1707 1067 1716
rect 1096 1707 1104 1736
rect 1247 1737 1273 1745
rect 1876 1736 2053 1744
rect 1876 1707 1884 1736
rect 2080 1744 2093 1747
rect 2076 1733 2093 1744
rect 2216 1736 2373 1744
rect 167 1696 244 1704
rect 347 1696 633 1704
rect 727 1695 773 1703
rect 1187 1696 1233 1704
rect 1307 1696 1733 1704
rect 1807 1696 1833 1704
rect 2076 1704 2084 1733
rect 2216 1707 2224 1736
rect 2507 1736 2564 1744
rect 2556 1707 2564 1736
rect 2807 1736 2844 1744
rect 2593 1724 2607 1733
rect 2836 1724 2844 1736
rect 2987 1737 3073 1745
rect 3096 1736 3153 1744
rect 3096 1724 3104 1736
rect 3347 1737 3393 1745
rect 3407 1736 3493 1744
rect 3547 1738 3573 1746
rect 3747 1737 3793 1745
rect 3936 1736 3993 1744
rect 2593 1720 2624 1724
rect 2596 1716 2624 1720
rect 2836 1716 3004 1724
rect 2616 1707 2624 1716
rect 1987 1696 2084 1704
rect 2127 1696 2153 1704
rect 2427 1696 2513 1704
rect 2616 1696 2633 1707
rect 2620 1693 2633 1696
rect 2996 1706 3004 1716
rect 3036 1716 3104 1724
rect 3036 1706 3044 1716
rect 3936 1707 3944 1736
rect 4047 1737 4113 1745
rect 4187 1736 4393 1744
rect 4596 1736 4633 1744
rect 4596 1707 4604 1736
rect 4687 1737 4713 1745
rect 4727 1736 4853 1744
rect 4896 1707 4904 1734
rect 4955 1707 4963 1756
rect 5027 1756 5147 1764
rect 5133 1748 5147 1756
rect 5367 1756 5404 1764
rect 4976 1707 4984 1735
rect 5067 1737 5093 1745
rect 5147 1736 5224 1744
rect 3627 1695 3713 1703
rect 4036 1696 4153 1704
rect 4036 1687 4044 1696
rect 4227 1695 4313 1703
rect 4667 1696 4753 1704
rect 4767 1696 4813 1704
rect 4896 1696 4913 1707
rect 4900 1693 4913 1696
rect 5127 1696 5173 1704
rect 5216 1704 5224 1736
rect 5267 1736 5324 1744
rect 5316 1707 5324 1736
rect 5396 1707 5404 1756
rect 5427 1744 5440 1747
rect 5427 1733 5444 1744
rect 5216 1696 5273 1704
rect 5436 1706 5444 1733
rect 5476 1707 5484 1813
rect 5527 1776 5653 1784
rect 5627 1737 5673 1745
rect 5516 1707 5524 1733
rect 1127 1676 2813 1684
rect 2827 1676 2873 1684
rect 3187 1676 3333 1684
rect 4027 1676 4044 1687
rect 4027 1673 4040 1676
rect 5207 1676 5233 1684
rect 5507 1676 5553 1684
rect 227 1656 273 1664
rect 287 1656 393 1664
rect 407 1656 813 1664
rect 1027 1656 1333 1664
rect 1467 1656 2213 1664
rect 2907 1656 3073 1664
rect 3087 1656 3133 1664
rect 3227 1656 3304 1664
rect 587 1636 633 1644
rect 1016 1644 1024 1653
rect 647 1636 1024 1644
rect 1367 1636 1733 1644
rect 1747 1636 2693 1644
rect 2707 1636 2993 1644
rect 3296 1644 3304 1656
rect 3547 1656 3673 1664
rect 4127 1656 4273 1664
rect 4447 1656 4513 1664
rect 5067 1656 5373 1664
rect 5427 1656 5473 1664
rect 3296 1636 3333 1644
rect 3527 1636 3873 1644
rect 4027 1636 4053 1644
rect 4627 1636 4733 1644
rect 4887 1636 4973 1644
rect 1507 1616 1593 1624
rect 1667 1616 1853 1624
rect 1867 1616 1933 1624
rect 2167 1616 2653 1624
rect 2667 1616 2893 1624
rect 2947 1616 3273 1624
rect 5307 1616 5513 1624
rect 1387 1596 1433 1604
rect 1527 1596 1973 1604
rect 3647 1596 3733 1604
rect 3747 1596 3893 1604
rect 5027 1596 5533 1604
rect 2287 1576 2393 1584
rect 2407 1576 3333 1584
rect 1347 1556 1513 1564
rect 1967 1556 2033 1564
rect 2047 1556 2153 1564
rect 2267 1556 2353 1564
rect 4347 1556 4933 1564
rect 5067 1556 5273 1564
rect 727 1536 1093 1544
rect 1187 1536 1273 1544
rect 1327 1536 2413 1544
rect 2467 1536 2513 1544
rect 2627 1536 2973 1544
rect 3847 1536 3913 1544
rect 4927 1536 5113 1544
rect 5487 1536 5513 1544
rect 5527 1536 5713 1544
rect 827 1516 853 1524
rect 967 1516 1113 1524
rect 1827 1516 2013 1524
rect 2167 1516 2293 1524
rect 3167 1516 3313 1524
rect 3327 1516 3553 1524
rect 4107 1516 4253 1524
rect 467 1496 1273 1504
rect 2127 1496 2233 1504
rect 2387 1496 2613 1504
rect 2807 1496 3433 1504
rect 3727 1496 4073 1504
rect 4467 1496 5013 1504
rect 5287 1496 5313 1504
rect 5447 1496 5673 1504
rect 827 1476 973 1484
rect 1567 1476 1613 1484
rect 2007 1476 2293 1484
rect 2727 1476 2833 1484
rect 1307 1456 1413 1464
rect 2196 1456 2273 1464
rect 167 1436 313 1444
rect 700 1444 713 1447
rect 587 1436 604 1444
rect 596 1407 604 1436
rect 696 1433 713 1444
rect 796 1436 933 1444
rect 487 1396 513 1404
rect 527 1396 553 1404
rect 696 1406 704 1433
rect 796 1406 804 1436
rect 1196 1436 1273 1444
rect 1196 1406 1204 1436
rect 1587 1436 1673 1444
rect 2140 1444 2152 1447
rect 1676 1407 1684 1434
rect 1676 1396 1693 1407
rect 1680 1393 1693 1396
rect 2076 1404 2084 1434
rect 2136 1433 2152 1444
rect 2196 1444 2204 1456
rect 2487 1456 2533 1464
rect 2887 1456 3133 1464
rect 3147 1456 3193 1464
rect 3793 1456 4153 1464
rect 2360 1444 2373 1447
rect 2187 1436 2204 1444
rect 2356 1433 2373 1444
rect 2733 1444 2747 1453
rect 3793 1448 3807 1456
rect 4727 1456 4784 1464
rect 2716 1440 2747 1444
rect 2716 1436 2744 1440
rect 2756 1436 2793 1444
rect 2136 1406 2144 1433
rect 2356 1406 2364 1433
rect 2496 1407 2504 1433
rect 2716 1424 2724 1436
rect 2756 1424 2764 1436
rect 2916 1436 3033 1444
rect 2696 1416 2724 1424
rect 2736 1416 2764 1424
rect 1987 1396 2084 1404
rect 2696 1406 2704 1416
rect 2736 1406 2744 1416
rect 2607 1395 2653 1403
rect 2916 1404 2924 1436
rect 3287 1436 3333 1444
rect 3387 1436 3413 1444
rect 3467 1436 3593 1444
rect 3747 1437 3793 1445
rect 4400 1444 4413 1447
rect 2867 1396 2924 1404
rect 3487 1396 3533 1404
rect 3636 1404 3644 1433
rect 3676 1407 3684 1433
rect 3627 1396 3644 1404
rect 3667 1396 3684 1407
rect 3667 1393 3680 1396
rect 3856 1404 3864 1434
rect 4216 1407 4224 1434
rect 4396 1433 4413 1444
rect 4496 1436 4553 1444
rect 4396 1407 4404 1433
rect 4496 1424 4504 1436
rect 4667 1436 4693 1444
rect 4733 1424 4747 1433
rect 4436 1416 4504 1424
rect 4696 1420 4747 1424
rect 4696 1416 4744 1420
rect 3747 1396 3864 1404
rect 3987 1396 4053 1404
rect 4216 1396 4233 1407
rect 4220 1393 4233 1396
rect 4436 1405 4444 1416
rect 4487 1396 4513 1404
rect 4696 1404 4704 1416
rect 4647 1396 4704 1404
rect 4776 1404 4784 1456
rect 5567 1456 5653 1464
rect 5136 1436 5213 1444
rect 5136 1406 5144 1436
rect 5236 1436 5333 1444
rect 5236 1406 5244 1436
rect 5607 1437 5713 1445
rect 4727 1396 4784 1404
rect 4947 1395 4973 1403
rect 5416 1404 5424 1433
rect 5367 1396 5453 1404
rect 5627 1395 5693 1403
rect 347 1376 413 1384
rect 1507 1376 1713 1384
rect 1727 1376 1953 1384
rect 3347 1376 3433 1384
rect 3447 1376 3573 1384
rect 3587 1376 3693 1384
rect 4347 1376 4373 1384
rect 4547 1376 4613 1384
rect 2707 1356 2893 1364
rect 4067 1356 4653 1364
rect 5207 1356 5393 1364
rect 627 1336 753 1344
rect 767 1336 884 1344
rect 67 1316 113 1324
rect 876 1324 884 1336
rect 2067 1336 2273 1344
rect 2387 1336 2533 1344
rect 2827 1336 2873 1344
rect 2887 1336 3373 1344
rect 3707 1336 3733 1344
rect 4047 1336 4253 1344
rect 876 1316 1213 1324
rect 2507 1316 2553 1324
rect 3947 1316 5093 1324
rect 5307 1316 5433 1324
rect 867 1296 1433 1304
rect 1567 1296 2173 1304
rect 2307 1296 2353 1304
rect 2376 1296 2813 1304
rect 107 1276 193 1284
rect 607 1276 833 1284
rect 847 1276 933 1284
rect 1007 1276 1073 1284
rect 1247 1276 1373 1284
rect 1587 1276 1853 1284
rect 1867 1276 2033 1284
rect 2376 1284 2384 1296
rect 4527 1296 4573 1304
rect 5527 1296 5593 1304
rect 2227 1276 2384 1284
rect 3647 1276 3693 1284
rect 3707 1276 3793 1284
rect 3867 1276 4093 1284
rect 4107 1276 4193 1284
rect 4667 1276 4713 1284
rect 136 1260 444 1264
rect 133 1256 444 1260
rect 133 1247 147 1256
rect 436 1247 444 1256
rect 1607 1256 1893 1264
rect 2487 1256 2513 1264
rect 2647 1256 2864 1264
rect 447 1236 513 1244
rect 587 1236 633 1244
rect 727 1236 753 1244
rect 767 1236 893 1244
rect 1007 1236 1153 1244
rect 1167 1236 1253 1244
rect 1327 1236 1353 1244
rect 1407 1236 1453 1244
rect 1727 1236 2053 1244
rect 2856 1244 2864 1256
rect 4887 1256 4973 1264
rect 5027 1256 5073 1264
rect 5087 1256 5113 1264
rect 5187 1256 5293 1264
rect 2856 1236 2933 1244
rect 3007 1236 3173 1244
rect 4387 1236 4673 1244
rect 5227 1236 5273 1244
rect 227 1217 653 1225
rect 776 1216 833 1224
rect 56 1187 64 1214
rect 47 1176 64 1187
rect 47 1173 60 1176
rect 776 1186 784 1216
rect 1420 1224 1433 1227
rect 1307 1216 1384 1224
rect 1376 1187 1384 1216
rect 1416 1213 1433 1224
rect 1487 1216 1533 1224
rect 1556 1216 1593 1224
rect 1416 1187 1424 1213
rect 1556 1204 1564 1216
rect 1516 1196 1564 1204
rect 1616 1196 1713 1204
rect 227 1176 253 1184
rect 547 1176 633 1184
rect 647 1175 713 1183
rect 827 1175 853 1183
rect 927 1176 993 1184
rect 1127 1176 1173 1184
rect 1227 1176 1273 1184
rect 1516 1186 1524 1196
rect 1616 1186 1624 1196
rect 1796 1184 1804 1214
rect 1867 1216 1924 1224
rect 1916 1187 1924 1216
rect 1987 1216 2033 1224
rect 2367 1217 2433 1225
rect 2527 1217 2613 1225
rect 2076 1187 2084 1214
rect 2747 1216 2793 1224
rect 3387 1216 3533 1224
rect 1796 1176 1873 1184
rect 1967 1176 2013 1184
rect 2076 1176 2093 1187
rect 2080 1173 2093 1176
rect 2147 1176 2193 1184
rect 2207 1176 2533 1184
rect 2656 1184 2664 1213
rect 2656 1176 2673 1184
rect 447 1156 573 1164
rect 587 1156 813 1164
rect 1467 1156 1553 1164
rect 2127 1156 2313 1164
rect 2696 1164 2704 1214
rect 2836 1187 2844 1214
rect 3747 1217 3853 1225
rect 4027 1216 4093 1224
rect 4207 1216 4333 1224
rect 2836 1176 2853 1187
rect 2840 1173 2853 1176
rect 3107 1176 3133 1184
rect 3207 1176 3273 1184
rect 3287 1175 3393 1183
rect 3407 1175 3433 1183
rect 3807 1176 4073 1184
rect 4196 1184 4204 1215
rect 4527 1224 4540 1227
rect 4527 1213 4544 1224
rect 4787 1216 4833 1224
rect 4853 1224 4867 1233
rect 4853 1220 4904 1224
rect 4856 1216 4904 1220
rect 4396 1187 4404 1213
rect 4167 1176 4204 1184
rect 4227 1176 4353 1184
rect 4536 1186 4544 1213
rect 4896 1187 4904 1216
rect 5067 1224 5080 1227
rect 5067 1213 5084 1224
rect 5076 1187 5084 1213
rect 5207 1217 5253 1225
rect 5527 1216 5593 1224
rect 5093 1204 5107 1213
rect 5093 1200 5453 1204
rect 5096 1196 5453 1200
rect 4787 1175 4813 1183
rect 5007 1176 5073 1184
rect 2587 1156 2704 1164
rect 2827 1156 2993 1164
rect 3007 1156 3153 1164
rect 3667 1156 3693 1164
rect 4736 1156 4953 1164
rect 4736 1147 4744 1156
rect 4967 1156 5173 1164
rect 5267 1156 5433 1164
rect 687 1136 793 1144
rect 927 1136 973 1144
rect 1487 1136 1533 1144
rect 1587 1136 1673 1144
rect 1927 1136 2073 1144
rect 2627 1136 2693 1144
rect 4127 1136 4633 1144
rect 4647 1136 4733 1144
rect 4867 1136 4913 1144
rect 4987 1136 5133 1144
rect 5287 1136 5333 1144
rect 1887 1116 2633 1124
rect 3147 1116 3833 1124
rect 5207 1116 5393 1124
rect 347 1096 1033 1104
rect 1987 1096 2153 1104
rect 2247 1096 2624 1104
rect 87 1076 153 1084
rect 167 1076 193 1084
rect 2147 1076 2233 1084
rect 2247 1076 2413 1084
rect 2616 1084 2624 1096
rect 2687 1096 2913 1104
rect 3156 1096 3233 1104
rect 3156 1084 3164 1096
rect 3367 1096 3713 1104
rect 3987 1096 4613 1104
rect 4667 1096 5153 1104
rect 2616 1076 3164 1084
rect 5307 1076 5613 1084
rect 2607 1056 3193 1064
rect 4627 1056 4913 1064
rect 4927 1056 5273 1064
rect 787 1036 1073 1044
rect 2287 1036 3413 1044
rect 3567 1036 4273 1044
rect 4607 1036 4733 1044
rect 2327 1016 2813 1024
rect 4907 1016 5113 1024
rect 887 996 1553 1004
rect 3187 996 3453 1004
rect 3767 996 3913 1004
rect 4047 996 4093 1004
rect 5467 996 5733 1004
rect 1507 976 1613 984
rect 1667 976 1913 984
rect 2367 976 2392 984
rect 2427 976 2673 984
rect 2967 976 3553 984
rect 4487 976 4513 984
rect 4527 976 4653 984
rect 5287 980 5664 984
rect 5287 976 5667 980
rect 5653 967 5667 976
rect 347 956 584 964
rect 107 936 273 944
rect 576 944 584 956
rect 627 956 693 964
rect 1027 956 1393 964
rect 1487 956 2053 964
rect 2067 956 2333 964
rect 2347 956 2713 964
rect 2727 956 2833 964
rect 3407 956 3473 964
rect 3496 956 3533 964
rect 576 936 784 944
rect 227 916 304 924
rect 47 876 73 884
rect 296 884 304 916
rect 447 916 473 924
rect 547 917 653 925
rect 373 904 387 913
rect 776 907 784 936
rect 1056 936 1133 944
rect 827 916 864 924
rect 640 904 653 907
rect 356 900 387 904
rect 356 896 384 900
rect 296 876 313 884
rect 356 867 364 896
rect 636 893 653 904
rect 856 904 864 916
rect 947 917 973 925
rect 1056 904 1064 936
rect 1727 936 1753 944
rect 1807 936 1833 944
rect 1927 936 1953 944
rect 2987 936 3193 944
rect 3287 936 3364 944
rect 856 896 964 904
rect 387 875 513 883
rect 636 884 644 893
rect 956 886 964 896
rect 1016 896 1064 904
rect 536 880 644 884
rect 533 876 644 880
rect 533 867 547 876
rect 1016 884 1024 896
rect 1076 887 1084 914
rect 1307 916 1333 924
rect 1387 916 1413 924
rect 1007 876 1024 884
rect 1067 876 1084 887
rect 1496 886 1504 933
rect 1067 873 1080 876
rect 1267 875 1293 883
rect 1367 880 1404 884
rect 1367 876 1407 880
rect 1393 867 1407 876
rect 167 856 193 864
rect 727 856 893 864
rect 1516 864 1524 914
rect 1736 887 1744 913
rect 1856 887 1864 914
rect 2507 916 2532 924
rect 2567 924 2580 927
rect 2567 913 2584 924
rect 2687 916 2733 924
rect 2947 916 2984 924
rect 1936 887 1944 913
rect 2313 904 2327 913
rect 2313 900 2484 904
rect 2316 896 2484 900
rect 1847 876 1864 887
rect 1847 873 1860 876
rect 2047 875 2073 883
rect 2367 875 2453 883
rect 2476 884 2484 896
rect 2576 887 2584 913
rect 2896 887 2904 913
rect 2476 876 2553 884
rect 2576 876 2593 887
rect 2580 873 2593 876
rect 2887 876 2904 887
rect 2976 884 2984 916
rect 3047 917 3073 925
rect 3313 904 3327 913
rect 3236 900 3327 904
rect 3233 896 3324 900
rect 3233 887 3247 896
rect 2976 876 3093 884
rect 2887 873 2900 876
rect 3356 886 3364 936
rect 3496 944 3504 956
rect 3587 956 3673 964
rect 3907 956 4053 964
rect 4327 956 4453 964
rect 4567 956 4613 964
rect 3387 936 3504 944
rect 4027 936 4213 944
rect 5027 936 5053 944
rect 5067 936 5253 944
rect 5427 936 5533 944
rect 3467 916 3524 924
rect 3516 904 3524 916
rect 3547 917 3573 925
rect 3920 924 3933 927
rect 3516 896 3664 904
rect 3656 886 3664 896
rect 3467 876 3653 884
rect 3676 884 3684 913
rect 3796 887 3804 914
rect 3916 913 3933 924
rect 3987 924 4000 927
rect 3987 913 4004 924
rect 3676 876 3773 884
rect 3796 876 3813 887
rect 3800 873 3813 876
rect 3916 886 3924 913
rect 3996 886 4004 913
rect 4456 887 4464 914
rect 4567 916 4584 924
rect 4516 887 4524 913
rect 4576 887 4584 916
rect 4627 924 4640 927
rect 4627 913 4644 924
rect 4807 917 4833 925
rect 5167 917 5193 925
rect 5327 917 5373 925
rect 5387 916 5444 924
rect 4636 904 4644 913
rect 4636 896 4744 904
rect 4227 876 4433 884
rect 4456 876 4473 887
rect 4460 873 4473 876
rect 4627 876 4693 884
rect 4736 884 4744 896
rect 5436 887 5444 916
rect 5467 924 5480 927
rect 5467 913 5484 924
rect 5567 917 5593 925
rect 4736 876 4813 884
rect 5207 876 5273 884
rect 1487 856 1524 864
rect 1787 856 1953 864
rect 3167 856 3293 864
rect 3407 856 3433 864
rect 3653 864 3667 872
rect 5476 886 5484 913
rect 5656 904 5664 914
rect 5656 900 5684 904
rect 5656 896 5687 900
rect 5673 887 5687 896
rect 3653 856 3973 864
rect 4187 856 4233 864
rect 4507 856 4553 864
rect 4947 856 4973 864
rect 5027 856 5053 864
rect 5067 856 5093 864
rect 5116 856 5253 864
rect 567 836 893 844
rect 956 836 1344 844
rect 47 816 113 824
rect 327 816 413 824
rect 956 824 964 836
rect 867 816 964 824
rect 1336 824 1344 836
rect 1467 836 1553 844
rect 1727 836 2004 844
rect 1336 816 1473 824
rect 1687 816 1713 824
rect 1996 824 2004 836
rect 2087 836 2293 844
rect 2507 836 2593 844
rect 3107 836 3253 844
rect 4207 836 4333 844
rect 4347 836 4413 844
rect 4427 836 4573 844
rect 5116 844 5124 856
rect 5307 856 5393 864
rect 4827 836 5124 844
rect 5356 836 5713 844
rect 1996 816 2053 824
rect 2107 816 2133 824
rect 2387 816 2673 824
rect 2747 816 3033 824
rect 5356 824 5364 836
rect 5267 816 5364 824
rect 5387 816 5533 824
rect 287 796 373 804
rect 487 796 593 804
rect 1307 796 1953 804
rect 2487 796 2573 804
rect 2867 796 2993 804
rect 3207 796 3653 804
rect 3667 796 3813 804
rect 3827 796 4473 804
rect 4487 796 4533 804
rect 5067 796 5133 804
rect 907 776 1193 784
rect 1607 776 1633 784
rect 1827 784 1840 787
rect 1827 773 1844 784
rect 1907 776 1933 784
rect 2067 776 2273 784
rect 2567 776 2693 784
rect 3307 776 3473 784
rect 3847 776 3873 784
rect 4587 776 4633 784
rect 127 756 513 764
rect 527 756 573 764
rect 627 756 673 764
rect 1067 756 1093 764
rect 1836 764 1844 773
rect 1836 756 2204 764
rect 2196 747 2204 756
rect 2347 756 2633 764
rect 2767 756 2813 764
rect 2827 756 3073 764
rect 3647 756 3733 764
rect 3747 756 3773 764
rect 3787 756 3813 764
rect 3827 756 4133 764
rect 4147 756 4393 764
rect 4407 756 4553 764
rect 4567 756 5353 764
rect 247 736 293 744
rect 487 736 533 744
rect 1127 736 1204 744
rect 1196 724 1204 736
rect 1267 736 1413 744
rect 1427 736 1573 744
rect 1587 736 1813 744
rect 2207 736 2513 744
rect 2527 736 2873 744
rect 4067 736 4093 744
rect 4207 736 4333 744
rect 4467 736 4513 744
rect 4667 736 5073 744
rect 667 716 1164 724
rect 1196 716 1293 724
rect 236 684 244 694
rect 327 696 353 704
rect 407 696 424 704
rect 67 676 244 684
rect 416 667 424 696
rect 1156 684 1164 716
rect 1967 716 2253 724
rect 1187 697 1213 705
rect 1367 696 1413 704
rect 1607 704 1620 707
rect 1607 693 1624 704
rect 2373 704 2387 713
rect 2576 716 2733 724
rect 2373 700 2413 704
rect 2376 696 2413 700
rect 2576 704 2584 716
rect 2467 696 2624 704
rect 1156 676 1204 684
rect 1436 680 1573 684
rect 116 656 173 664
rect 116 627 124 656
rect 267 655 313 663
rect 467 656 493 664
rect 547 656 713 664
rect 867 656 933 664
rect 1067 655 1113 663
rect 1196 664 1204 676
rect 1433 676 1573 680
rect 1433 667 1447 676
rect 1196 656 1273 664
rect 1327 655 1353 663
rect 1616 666 1624 693
rect 1807 656 1873 664
rect 1976 664 1984 694
rect 2616 667 2624 696
rect 2807 698 2833 706
rect 2916 704 2924 733
rect 2947 716 2973 724
rect 3107 716 3293 724
rect 3727 716 3953 724
rect 4016 716 4593 724
rect 2916 696 2944 704
rect 1927 656 1984 664
rect 2067 655 2093 663
rect 2267 656 2493 664
rect 2507 656 2533 664
rect 2767 656 2813 664
rect 2936 666 2944 696
rect 3076 696 3193 704
rect 3076 684 3084 696
rect 3547 697 3573 705
rect 3056 676 3084 684
rect 3056 666 3064 676
rect 3436 667 3444 693
rect 3656 684 3664 713
rect 3796 696 3833 704
rect 3636 680 3664 684
rect 3633 676 3664 680
rect 3633 667 3647 676
rect 3676 667 3684 695
rect 3796 684 3804 696
rect 3887 696 3933 704
rect 3756 680 3804 684
rect 3753 676 3804 680
rect 3753 667 3767 676
rect 3096 656 3173 664
rect 3096 647 3104 656
rect 3227 655 3353 663
rect 3827 656 3853 664
rect 4016 666 4024 716
rect 4607 716 4693 724
rect 4707 716 5173 724
rect 5227 716 5313 724
rect 4047 696 4093 704
rect 4116 696 4213 704
rect 4116 684 4124 696
rect 4327 697 4373 705
rect 4396 696 4513 704
rect 4076 680 4124 684
rect 4073 676 4124 680
rect 4073 667 4087 676
rect 4396 666 4404 696
rect 5347 704 5360 707
rect 5347 693 5364 704
rect 4576 667 4584 693
rect 5056 667 5064 693
rect 5096 667 5104 693
rect 5216 684 5224 693
rect 5196 680 5224 684
rect 5193 676 5224 680
rect 5193 667 5207 676
rect 5356 667 5364 693
rect 4807 656 5013 664
rect 5447 655 5573 663
rect 2367 636 2433 644
rect 2987 636 3033 644
rect 3087 636 3104 647
rect 3087 633 3100 636
rect 3216 644 3224 652
rect 3127 636 3224 644
rect 3427 636 3473 644
rect 3487 636 3593 644
rect 4107 636 4192 644
rect 4227 636 4313 644
rect 5087 636 5133 644
rect 5667 636 5693 644
rect 547 616 773 624
rect 787 616 873 624
rect 1007 616 1093 624
rect 1227 616 1393 624
rect 1687 616 1713 624
rect 1727 616 1833 624
rect 1847 616 2153 624
rect 2167 616 2253 624
rect 2267 616 2973 624
rect 1396 604 1404 613
rect 3116 624 3124 633
rect 2987 616 3124 624
rect 3447 616 4073 624
rect 4167 616 4473 624
rect 1396 596 2333 604
rect 2356 596 2513 604
rect 1767 576 2193 584
rect 2356 584 2364 596
rect 2787 596 2893 604
rect 3667 596 3753 604
rect 3847 596 3893 604
rect 4207 596 4353 604
rect 5187 596 5273 604
rect 2207 576 2364 584
rect 2567 576 3464 584
rect 827 556 993 564
rect 1927 556 2393 564
rect 2527 556 3413 564
rect 3456 564 3464 576
rect 3916 576 4173 584
rect 3456 556 3513 564
rect 3916 564 3924 576
rect 4687 576 4893 584
rect 5067 576 5433 584
rect 3627 556 3924 564
rect 3947 556 4153 564
rect 4547 556 4593 564
rect 4607 556 4753 564
rect 5407 556 5493 564
rect 1267 536 1753 544
rect 3107 536 3253 544
rect 3267 536 3293 544
rect 3416 544 3424 553
rect 3416 536 3693 544
rect 5127 536 5193 544
rect 1587 516 2373 524
rect 2667 516 4153 524
rect 4247 516 4293 524
rect 4347 516 4633 524
rect 207 496 293 504
rect 1127 496 1233 504
rect 1247 496 1473 504
rect 1487 496 1553 504
rect 1747 496 1853 504
rect 5027 496 5153 504
rect 5327 496 5393 504
rect 1693 484 1707 493
rect 1607 476 3233 484
rect 3307 476 3953 484
rect 3967 476 3993 484
rect 4207 476 4253 484
rect 87 456 413 464
rect 1827 456 1913 464
rect 2027 456 2253 464
rect 2387 456 2733 464
rect 3207 456 3833 464
rect 4627 456 4653 464
rect 4667 456 4793 464
rect 1647 436 1733 444
rect 1807 436 1953 444
rect 1967 436 1993 444
rect 2007 436 2553 444
rect 2927 436 3053 444
rect 3707 436 3853 444
rect 3867 436 4033 444
rect 4267 436 4393 444
rect 4467 436 4533 444
rect 5087 436 5273 444
rect 5287 436 5673 444
rect 327 416 693 424
rect 707 416 813 424
rect 827 416 1093 424
rect 1107 416 1133 424
rect 1207 416 1353 424
rect 2247 416 2333 424
rect 4187 416 4673 424
rect 127 404 140 407
rect 127 393 144 404
rect 267 396 444 404
rect 136 366 144 393
rect 436 366 444 396
rect 467 397 493 405
rect 727 397 753 405
rect 947 396 1053 404
rect 1387 396 1433 404
rect 1767 404 1780 407
rect 1767 393 1784 404
rect 107 356 133 364
rect 507 356 553 364
rect 576 364 584 393
rect 1456 376 1573 384
rect 576 356 633 364
rect 647 355 853 363
rect 1007 356 1313 364
rect 1456 365 1464 376
rect 1776 366 1784 393
rect 1367 356 1413 364
rect 1527 355 1733 363
rect 1836 364 1844 394
rect 1927 396 2053 404
rect 2147 397 2173 405
rect 1836 356 1933 364
rect 2096 364 2104 393
rect 2196 366 2204 413
rect 2216 384 2224 394
rect 2587 396 2633 404
rect 2216 376 2393 384
rect 2533 384 2547 393
rect 2787 397 2813 405
rect 2993 384 3007 393
rect 2456 376 2784 384
rect 2993 380 3064 384
rect 2996 376 3064 380
rect 2456 366 2464 376
rect 1987 356 2104 364
rect 2607 356 2753 364
rect 2776 364 2784 376
rect 2776 356 2833 364
rect 2987 354 3033 362
rect 407 336 873 344
rect 887 336 1873 344
rect 2707 336 2733 344
rect 3056 344 3064 376
rect 3196 364 3204 394
rect 3387 396 3453 404
rect 3527 397 3653 405
rect 3576 367 3584 397
rect 3807 397 3833 405
rect 4067 396 4093 404
rect 4107 396 4133 404
rect 3716 367 3724 393
rect 4196 367 4204 393
rect 4236 367 4244 393
rect 3127 356 3204 364
rect 3347 355 3373 363
rect 3867 355 3913 363
rect 4027 356 4073 364
rect 4296 366 4304 416
rect 4327 396 4453 404
rect 4476 396 4493 404
rect 4476 367 4484 396
rect 4520 404 4533 407
rect 4467 356 4484 367
rect 4516 393 4533 404
rect 4587 396 4684 404
rect 4516 366 4524 393
rect 4676 384 4684 396
rect 4707 396 4753 404
rect 4887 396 4913 404
rect 4927 396 4953 404
rect 5067 396 5113 404
rect 5187 396 5213 404
rect 5347 397 5373 405
rect 5507 397 5553 405
rect 5013 384 5027 393
rect 4676 376 4784 384
rect 5013 380 5104 384
rect 5016 376 5104 380
rect 4467 353 4480 356
rect 4776 365 4784 376
rect 5096 366 5104 376
rect 4787 356 4853 364
rect 5467 356 5533 364
rect 3056 336 3164 344
rect 3156 327 3164 336
rect 3507 336 3613 344
rect 4107 336 4253 344
rect 5127 336 5233 344
rect 5247 336 5393 344
rect 1087 316 1253 324
rect 1347 316 1413 324
rect 1827 316 1853 324
rect 2407 316 2773 324
rect 3167 316 3473 324
rect 3607 316 3673 324
rect 4247 316 4293 324
rect 4467 316 4633 324
rect 4647 316 4693 324
rect 5396 324 5404 333
rect 5396 316 5673 324
rect 727 296 1033 304
rect 2027 296 2133 304
rect 2616 296 2953 304
rect 2387 276 2453 284
rect 2616 284 2624 296
rect 3007 296 3493 304
rect 3547 296 3833 304
rect 2467 276 2624 284
rect 2647 276 2713 284
rect 2727 276 2933 284
rect 3047 276 3073 284
rect 3307 276 3433 284
rect 4167 276 4993 284
rect 5107 276 5633 284
rect 2247 256 2433 264
rect 3067 256 3253 264
rect 3487 256 3573 264
rect 3727 256 3753 264
rect 4227 256 4353 264
rect 4687 256 4873 264
rect 5387 256 5453 264
rect 1087 236 1593 244
rect 2236 244 2244 253
rect 1987 236 2244 244
rect 2707 236 2753 244
rect 2767 236 3393 244
rect 3967 236 3993 244
rect 367 216 433 224
rect 1747 216 1993 224
rect 2867 216 2993 224
rect 3287 216 3453 224
rect 3607 216 4753 224
rect 4807 216 4993 224
rect 5016 216 5113 224
rect 967 196 1233 204
rect 1247 196 1453 204
rect 1836 196 1873 204
rect 47 177 93 185
rect 107 176 133 184
rect 407 176 484 184
rect 476 164 484 176
rect 507 176 553 184
rect 636 164 644 174
rect 727 176 853 184
rect 876 176 913 184
rect 876 164 884 176
rect 1007 176 1033 184
rect 1327 177 1353 185
rect 1507 176 1553 184
rect 1576 176 1673 184
rect 1576 164 1584 176
rect 476 160 544 164
rect 576 160 884 164
rect 476 156 547 160
rect 533 147 547 156
rect 87 135 193 143
rect 267 136 353 144
rect 467 135 493 143
rect 573 156 884 160
rect 1536 156 1584 164
rect 573 147 587 156
rect 727 135 753 143
rect 867 136 992 144
rect 1027 136 1053 144
rect 1536 146 1544 156
rect 1836 147 1844 196
rect 2273 196 2553 204
rect 2273 188 2287 196
rect 3127 196 3173 204
rect 5016 204 5024 216
rect 5167 216 5404 224
rect 2207 176 2273 184
rect 2356 176 2373 184
rect 1936 164 1944 174
rect 1936 156 1964 164
rect 1207 135 1493 143
rect 1667 136 1793 144
rect 1887 135 1913 143
rect 1956 144 1964 156
rect 2356 147 2364 176
rect 2667 176 2773 184
rect 2787 176 2813 184
rect 3013 164 3027 173
rect 3236 164 3244 193
rect 2447 156 2724 164
rect 1956 136 1992 144
rect 2027 135 2133 143
rect 2467 136 2493 144
rect 2647 135 2693 143
rect 2716 144 2724 156
rect 2936 160 3027 164
rect 2936 156 3024 160
rect 3216 156 3244 164
rect 3347 176 3444 184
rect 3293 164 3307 173
rect 3293 160 3344 164
rect 3296 156 3347 160
rect 2936 146 2944 156
rect 3216 146 3224 156
rect 3333 147 3347 156
rect 2716 136 2873 144
rect 3436 146 3444 176
rect 3476 146 3484 193
rect 3547 176 3773 184
rect 3536 147 3544 174
rect 3873 184 3887 193
rect 4996 196 5024 204
rect 5396 204 5404 216
rect 5447 216 5513 224
rect 5396 196 5533 204
rect 3847 180 3887 184
rect 3847 176 3884 180
rect 3907 177 3953 185
rect 3976 176 3993 184
rect 3976 164 3984 176
rect 4227 176 4413 184
rect 4427 176 4513 184
rect 4687 177 4733 185
rect 4947 177 4973 185
rect 4996 164 5004 196
rect 5087 176 5133 184
rect 5156 176 5193 184
rect 3856 160 3984 164
rect 4816 160 5004 164
rect 3527 136 3544 147
rect 3853 156 3984 160
rect 4813 156 5004 160
rect 3853 147 3867 156
rect 4813 147 4827 156
rect 3527 133 3540 136
rect 3727 135 3753 143
rect 3987 136 4433 144
rect 4447 135 4473 143
rect 4547 136 4593 144
rect 4667 136 4773 144
rect 4907 136 4933 144
rect 327 116 693 124
rect 707 116 813 124
rect 827 116 1133 124
rect 1387 116 1433 124
rect 1587 116 1693 124
rect 2696 124 2704 132
rect 2696 116 2833 124
rect 3473 124 3487 132
rect 3327 116 3487 124
rect 3756 124 3764 132
rect 3756 116 4033 124
rect 4936 124 4944 133
rect 5007 136 5053 144
rect 5156 146 5164 176
rect 5267 176 5333 184
rect 5347 178 5393 186
rect 5436 147 5444 196
rect 5487 136 5513 144
rect 4936 116 5333 124
rect 5507 116 5553 124
rect 1367 96 1553 104
rect 1607 96 1653 104
rect 1967 96 2293 104
rect 2307 96 2413 104
rect 2507 96 2593 104
rect 3407 96 3453 104
rect 3507 96 3593 104
rect 4967 96 5113 104
rect 5307 96 5393 104
rect 5447 96 5593 104
rect 207 76 413 84
rect 1107 76 1233 84
rect 2007 76 2073 84
rect 2756 76 3153 84
rect 2756 64 2764 76
rect 3907 76 4093 84
rect 2407 56 2764 64
rect 3287 56 3653 64
rect 5087 56 5233 64
rect 5247 56 5373 64
rect 2887 36 3053 44
rect 2367 16 2393 24
rect 2507 16 2553 24
use NOR2X1  _723_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726536993
transform 1 0 3870 0 1 790
box -12 -8 92 272
use INVX2  _724_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726533902
transform 1 0 3750 0 -1 790
box -12 -8 72 272
use NOR2X1  _725_
timestamp 1726536993
transform -1 0 3090 0 -1 790
box -12 -8 92 272
use OAI21X1  _726_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726538409
transform 1 0 4390 0 1 790
box -12 -8 112 272
use INVX2  _727_
timestamp 1726533902
transform -1 0 2830 0 -1 790
box -12 -8 72 272
use NOR2X1  _728_
timestamp 1726536993
transform 1 0 2790 0 -1 1310
box -12 -8 92 272
use AOI22X1  _729_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726480912
transform 1 0 3470 0 -1 1830
box -14 -8 132 272
use OAI21X1  _730_
timestamp 1726538409
transform 1 0 3990 0 1 790
box -12 -8 112 272
use INVX1  _731_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726531033
transform 1 0 4530 0 1 790
box -12 -8 72 272
use INVX1  _732_
timestamp 1726531033
transform 1 0 5530 0 1 270
box -12 -8 72 272
use NAND2X1  _733_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726535706
transform 1 0 5350 0 -1 790
box -12 -8 92 272
use OAI21X1  _734_
timestamp 1726538409
transform 1 0 5350 0 1 790
box -12 -8 112 272
use AOI22X1  _735_
timestamp 1726480912
transform 1 0 2910 0 -1 1310
box -14 -8 132 272
use OAI21X1  _736_
timestamp 1726538409
transform -1 0 4350 0 1 790
box -12 -8 112 272
use INVX1  _737_
timestamp 1726531033
transform 1 0 3170 0 1 270
box -12 -8 72 272
use NAND2X1  _738_
timestamp 1726535706
transform 1 0 3850 0 -1 790
box -12 -8 92 272
use OAI21X1  _739_
timestamp 1726538409
transform -1 0 4570 0 -1 790
box -12 -8 112 272
use AOI22X1  _740_
timestamp 1726480912
transform 1 0 2610 0 -1 790
box -14 -8 132 272
use OAI21X1  _741_
timestamp 1726538409
transform -1 0 4430 0 -1 790
box -12 -8 112 272
use NOR2X1  _742_
timestamp 1726536993
transform -1 0 3310 0 1 790
box -12 -8 92 272
use OAI21X1  _743_
timestamp 1726538409
transform 1 0 3730 0 1 790
box -12 -8 112 272
use AOI22X1  _744_
timestamp 1726480912
transform 1 0 2230 0 1 790
box -14 -8 132 272
use OAI21X1  _745_
timestamp 1726538409
transform 1 0 3350 0 1 790
box -12 -8 112 272
use INVX2  _746_
timestamp 1726533902
transform -1 0 3570 0 1 2870
box -12 -8 72 272
use NAND2X1  _747_
timestamp 1726535706
transform -1 0 3150 0 -1 2870
box -12 -8 92 272
use OAI21X1  _748_
timestamp 1726538409
transform -1 0 3470 0 1 2870
box -12 -8 112 272
use INVX1  _749_
timestamp 1726531033
transform 1 0 3710 0 1 4430
box -12 -8 72 272
use NAND2X1  _750_
timestamp 1726535706
transform -1 0 3250 0 -1 3910
box -12 -8 92 272
use OAI21X1  _751_
timestamp 1726538409
transform -1 0 3390 0 -1 3910
box -12 -8 112 272
use INVX2  _752_
timestamp 1726533902
transform 1 0 2810 0 -1 4430
box -12 -8 72 272
use NAND2X1  _753_
timestamp 1726535706
transform -1 0 3230 0 1 3910
box -12 -8 92 272
use OAI21X1  _754_
timestamp 1726538409
transform -1 0 3490 0 1 3910
box -12 -8 112 272
use INVX2  _755_
timestamp 1726533902
transform 1 0 3810 0 1 4430
box -12 -8 72 272
use NAND2X1  _756_
timestamp 1726535706
transform -1 0 3350 0 1 3910
box -12 -8 92 272
use OAI21X1  _757_
timestamp 1726538409
transform 1 0 3530 0 1 3910
box -12 -8 112 272
use NAND2X1  _758_
timestamp 1726535706
transform 1 0 2870 0 1 2870
box -12 -8 92 272
use OAI21X1  _759_
timestamp 1726538409
transform -1 0 3090 0 1 2870
box -12 -8 112 272
use NAND2X1  _760_
timestamp 1726535706
transform 1 0 2610 0 1 3390
box -12 -8 92 272
use OAI21X1  _761_
timestamp 1726538409
transform -1 0 2890 0 -1 3910
box -12 -8 112 272
use NAND2X1  _762_
timestamp 1726535706
transform 1 0 3510 0 1 3390
box -12 -8 92 272
use OAI21X1  _763_
timestamp 1726538409
transform -1 0 3730 0 1 3390
box -12 -8 112 272
use NAND2X1  _764_
timestamp 1726535706
transform 1 0 3290 0 -1 3390
box -12 -8 92 272
use OAI21X1  _765_
timestamp 1726538409
transform -1 0 3510 0 -1 3390
box -12 -8 112 272
use INVX1  _766_
timestamp 1726531033
transform -1 0 2930 0 1 1830
box -12 -8 72 272
use NAND2X1  _767_
timestamp 1726535706
transform 1 0 2730 0 -1 1830
box -12 -8 92 272
use OAI21X1  _768_
timestamp 1726538409
transform -1 0 2830 0 1 1830
box -12 -8 112 272
use INVX1  _769_
timestamp 1726531033
transform 1 0 510 0 -1 1310
box -12 -8 72 272
use NAND2X1  _770_
timestamp 1726535706
transform 1 0 770 0 -1 790
box -12 -8 92 272
use OAI21X1  _771_
timestamp 1726538409
transform 1 0 610 0 -1 1310
box -12 -8 112 272
use INVX1  _772_
timestamp 1726531033
transform -1 0 110 0 1 270
box -12 -8 72 272
use NAND2X1  _773_
timestamp 1726535706
transform 1 0 530 0 1 270
box -12 -8 92 272
use OAI21X1  _774_
timestamp 1726538409
transform 1 0 390 0 1 270
box -12 -8 112 272
use INVX1  _775_
timestamp 1726531033
transform -1 0 110 0 -1 270
box -12 -8 72 272
use NAND2X1  _776_
timestamp 1726535706
transform 1 0 530 0 -1 270
box -12 -8 92 272
use OAI21X1  _777_
timestamp 1726538409
transform 1 0 390 0 -1 270
box -12 -8 112 272
use INVX1  _778_
timestamp 1726531033
transform 1 0 1270 0 1 2350
box -12 -8 72 272
use NAND2X1  _779_
timestamp 1726535706
transform -1 0 1510 0 1 1830
box -12 -8 92 272
use OAI21X1  _780_
timestamp 1726538409
transform 1 0 1290 0 -1 2350
box -12 -8 112 272
use INVX1  _781_
timestamp 1726531033
transform -1 0 2930 0 -1 2350
box -12 -8 72 272
use NAND2X1  _782_
timestamp 1726535706
transform -1 0 2690 0 1 1830
box -12 -8 92 272
use OAI21X1  _783_
timestamp 1726538409
transform -1 0 2830 0 -1 2350
box -12 -8 112 272
use INVX1  _784_
timestamp 1726531033
transform 1 0 1630 0 -1 1830
box -12 -8 72 272
use NAND2X1  _785_
timestamp 1726535706
transform 1 0 1870 0 -1 790
box -12 -8 92 272
use OAI21X1  _786_
timestamp 1726538409
transform -1 0 1970 0 -1 1830
box -12 -8 112 272
use INVX1  _787_
timestamp 1726531033
transform -1 0 710 0 1 1310
box -12 -8 72 272
use NAND2X1  _788_
timestamp 1726535706
transform 1 0 890 0 -1 790
box -12 -8 92 272
use OAI21X1  _789_
timestamp 1726538409
transform 1 0 750 0 1 1310
box -12 -8 112 272
use INVX1  _790_
timestamp 1726531033
transform -1 0 4030 0 -1 2350
box -12 -8 72 272
use NAND2X1  _791_
timestamp 1726535706
transform -1 0 3950 0 -1 1830
box -12 -8 92 272
use OAI21X1  _792_
timestamp 1726538409
transform 1 0 3830 0 -1 2350
box -12 -8 112 272
use INVX1  _793_
timestamp 1726531033
transform 1 0 5590 0 -1 1310
box -12 -8 72 272
use NAND2X1  _794_
timestamp 1726535706
transform -1 0 4750 0 -1 1310
box -12 -8 92 272
use OAI21X1  _795_
timestamp 1726538409
transform -1 0 5310 0 -1 1310
box -12 -8 112 272
use INVX1  _796_
timestamp 1726531033
transform -1 0 4910 0 -1 2350
box -12 -8 72 272
use NAND2X1  _797_
timestamp 1726535706
transform -1 0 4750 0 1 1310
box -12 -8 92 272
use OAI21X1  _798_
timestamp 1726538409
transform -1 0 4810 0 -1 2350
box -12 -8 112 272
use INVX1  _799_
timestamp 1726531033
transform -1 0 4190 0 -1 1830
box -12 -8 72 272
use NAND2X1  _800_
timestamp 1726535706
transform -1 0 4130 0 -1 1310
box -12 -8 92 272
use OAI21X1  _801_
timestamp 1726538409
transform 1 0 3990 0 -1 1830
box -12 -8 112 272
use INVX1  _802_
timestamp 1726531033
transform -1 0 4930 0 -1 790
box -12 -8 72 272
use NAND2X1  _803_
timestamp 1726535706
transform 1 0 3990 0 1 270
box -12 -8 92 272
use OAI21X1  _804_
timestamp 1726538409
transform -1 0 4710 0 -1 790
box -12 -8 112 272
use INVX1  _805_
timestamp 1726531033
transform 1 0 4410 0 -1 270
box -12 -8 72 272
use NAND2X1  _806_
timestamp 1726535706
transform -1 0 3870 0 -1 270
box -12 -8 92 272
use OAI21X1  _807_
timestamp 1726538409
transform -1 0 4010 0 -1 270
box -12 -8 112 272
use INVX1  _808_
timestamp 1726531033
transform -1 0 2850 0 1 270
box -12 -8 72 272
use NAND2X1  _809_
timestamp 1726535706
transform -1 0 2110 0 1 270
box -12 -8 92 272
use OAI21X1  _810_
timestamp 1726538409
transform -1 0 2250 0 1 270
box -12 -8 112 272
use INVX1  _811_
timestamp 1726531033
transform 1 0 2270 0 -1 270
box -12 -8 72 272
use NAND2X1  _812_
timestamp 1726535706
transform -1 0 1850 0 -1 270
box -12 -8 92 272
use OAI21X1  _813_
timestamp 1726538409
transform -1 0 1990 0 -1 270
box -12 -8 112 272
use INVX1  _814_
timestamp 1726531033
transform 1 0 2590 0 -1 2870
box -12 -8 72 272
use NAND3X1  _815_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726536591
transform 1 0 1970 0 -1 2870
box -12 -8 112 272
use OAI21X1  _816_
timestamp 1726538409
transform -1 0 2310 0 -1 2870
box -12 -8 112 272
use INVX8  _817_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726534447
transform 1 0 3210 0 1 1830
box -12 -8 133 272
use NAND2X1  _818_
timestamp 1726535706
transform -1 0 1290 0 -1 2870
box -12 -8 92 272
use NAND2X1  _819_
timestamp 1726535706
transform 1 0 1490 0 -1 2870
box -12 -8 92 272
use XNOR2X1  _820_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726561449
transform -1 0 1110 0 1 2350
box -12 -8 152 272
use NAND2X1  _821_
timestamp 1726535706
transform 1 0 530 0 -1 1830
box -12 -8 92 272
use OAI21X1  _822_
timestamp 1726538409
transform -1 0 750 0 -1 1830
box -12 -8 112 272
use NOR2X1  _823_
timestamp 1726536993
transform -1 0 930 0 1 2350
box -12 -8 92 272
use NAND2X1  _824_
timestamp 1726535706
transform -1 0 1270 0 1 2870
box -12 -8 92 272
use NAND2X1  _825_
timestamp 1726535706
transform 1 0 1170 0 -1 3390
box -12 -8 92 272
use NOR2X1  _826_
timestamp 1726536993
transform 1 0 1090 0 -1 2870
box -12 -8 92 272
use AOI22X1  _827_
timestamp 1726480912
transform 1 0 1330 0 -1 2870
box -14 -8 132 272
use OAI21X1  _828_
timestamp 1726538409
transform 1 0 950 0 -1 2870
box -12 -8 112 272
use INVX1  _829_
timestamp 1726531033
transform 1 0 850 0 -1 2870
box -12 -8 72 272
use AND2X2  _830_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726549440
transform -1 0 1670 0 1 2870
box -12 -8 112 273
use AND2X2  _831_
timestamp 1726549440
transform 1 0 1310 0 1 2870
box -12 -8 112 273
use NAND2X1  _832_
timestamp 1726535706
transform -1 0 1530 0 1 2870
box -12 -8 92 272
use INVX1  _833_
timestamp 1726531033
transform 1 0 1870 0 -1 2870
box -12 -8 72 272
use INVX1  _834_
timestamp 1726531033
transform -1 0 3490 0 -1 4950
box -12 -8 72 272
use NAND2X1  _835_
timestamp 1726535706
transform -1 0 1690 0 -1 2870
box -12 -8 92 272
use OAI21X1  _836_
timestamp 1726538409
transform -1 0 1830 0 -1 2870
box -12 -8 112 272
use NAND3X1  _837_
timestamp 1726536591
transform -1 0 810 0 -1 2870
box -12 -8 112 272
use NAND3X1  _838_
timestamp 1726536591
transform -1 0 810 0 1 2350
box -12 -8 112 272
use INVX1  _839_
timestamp 1726531033
transform -1 0 630 0 -1 2350
box -12 -8 72 272
use AOI21X1  _840_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726549551
transform -1 0 670 0 1 2350
box -12 -8 112 272
use OAI21X1  _841_
timestamp 1726538409
transform -1 0 530 0 -1 2350
box -12 -8 112 272
use INVX1  _842_
timestamp 1726531033
transform 1 0 230 0 -1 790
box -12 -8 72 272
use NAND2X1  _843_
timestamp 1726535706
transform 1 0 390 0 -1 1310
box -12 -8 92 272
use AND2X2  _844_
timestamp 1726549440
transform -1 0 390 0 1 1310
box -12 -8 112 273
use INVX1  _845_
timestamp 1726531033
transform 1 0 50 0 -1 1310
box -12 -8 72 272
use NAND2X1  _846_
timestamp 1726535706
transform 1 0 1970 0 1 3390
box -12 -8 92 272
use AOI21X1  _847_
timestamp 1726549551
transform -1 0 670 0 -1 2870
box -12 -8 112 272
use NAND2X1  _848_
timestamp 1726535706
transform -1 0 1370 0 -1 3390
box -12 -8 92 272
use NAND2X1  _849_
timestamp 1726535706
transform -1 0 750 0 1 4430
box -12 -8 92 272
use NOR2X1  _850_
timestamp 1726536993
transform -1 0 750 0 -1 3390
box -12 -8 92 272
use AOI22X1  _851_
timestamp 1726480912
transform -1 0 1250 0 1 3390
box -14 -8 132 272
use OAI21X1  _852_
timestamp 1726538409
transform -1 0 630 0 -1 3390
box -12 -8 112 272
use INVX1  _853_
timestamp 1726531033
transform -1 0 850 0 -1 3390
box -12 -8 72 272
use AND2X2  _854_
timestamp 1726549440
transform 1 0 1290 0 1 3390
box -12 -8 112 273
use NAND2X1  _855_
timestamp 1726535706
transform 1 0 1430 0 1 3390
box -12 -8 92 272
use INVX1  _856_
timestamp 1726531033
transform 1 0 890 0 1 3390
box -12 -8 72 272
use NAND3X1  _857_
timestamp 1726536591
transform -1 0 850 0 1 3390
box -12 -8 112 272
use NAND3X1  _858_
timestamp 1726536591
transform -1 0 570 0 1 2870
box -12 -8 112 272
use OAI21X1  _859_
timestamp 1726538409
transform -1 0 850 0 1 2870
box -12 -8 112 272
use AOI21X1  _860_
timestamp 1726549551
transform -1 0 710 0 1 3390
box -12 -8 112 272
use INVX2  _861_
timestamp 1726533902
transform -1 0 1850 0 -1 3910
box -12 -8 72 272
use OAI21X1  _862_
timestamp 1726538409
transform -1 0 1790 0 1 3390
box -12 -8 112 272
use INVX2  _863_
timestamp 1726533902
transform -1 0 2630 0 -1 4430
box -12 -8 72 272
use INVX1  _864_
timestamp 1726531033
transform 1 0 970 0 -1 4430
box -12 -8 72 272
use OAI21X1  _865_
timestamp 1726538409
transform -1 0 1930 0 1 3390
box -12 -8 112 272
use AOI21X1  _866_
timestamp 1726549551
transform -1 0 1650 0 1 3390
box -12 -8 112 272
use OAI21X1  _867_
timestamp 1726538409
transform 1 0 610 0 1 2870
box -12 -8 112 272
use NAND3X1  _868_
timestamp 1726536591
transform -1 0 290 0 1 2870
box -12 -8 112 272
use INVX1  _869_
timestamp 1726531033
transform -1 0 210 0 -1 3390
box -12 -8 72 272
use NAND3X1  _870_
timestamp 1726536591
transform -1 0 430 0 1 2870
box -12 -8 112 272
use OAI21X1  _871_
timestamp 1726538409
transform -1 0 530 0 -1 2870
box -12 -8 112 272
use NAND3X1  _872_
timestamp 1726536591
transform -1 0 390 0 -1 2870
box -12 -8 112 272
use AOI21X1  _873_
timestamp 1726549551
transform 1 0 290 0 -1 2350
box -12 -8 112 272
use NAND3X1  _874_
timestamp 1726536591
transform -1 0 250 0 -1 2350
box -12 -8 112 272
use NAND2X1  _875_
timestamp 1726535706
transform -1 0 130 0 1 1830
box -12 -8 92 272
use OAI22X1  _876_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726541006
transform 1 0 170 0 1 1830
box -12 -8 132 272
use INVX1  _877_
timestamp 1726531033
transform -1 0 1010 0 -1 2350
box -12 -8 72 272
use INVX1  _878_
timestamp 1726531033
transform -1 0 110 0 -1 2350
box -12 -8 72 272
use AOI21X1  _879_
timestamp 1726549551
transform -1 0 490 0 -1 3390
box -12 -8 112 272
use OAI21X1  _880_
timestamp 1726538409
transform -1 0 350 0 -1 3390
box -12 -8 112 272
use OAI21X1  _881_
timestamp 1726538409
transform 1 0 990 0 1 3390
box -12 -8 112 272
use AND2X2  _882_
timestamp 1726549440
transform 1 0 950 0 1 4950
box -12 -8 112 273
use NAND2X1  _883_
timestamp 1726535706
transform -1 0 1250 0 1 3910
box -12 -8 92 272
use AOI22X1  _884_
timestamp 1726480912
transform 1 0 790 0 1 4430
box -14 -8 132 272
use INVX1  _885_
timestamp 1726531033
transform -1 0 110 0 1 4430
box -12 -8 72 272
use NAND2X1  _886_
timestamp 1726535706
transform 1 0 1070 0 -1 4430
box -12 -8 92 272
use INVX1  _887_
timestamp 1726531033
transform -1 0 110 0 -1 4430
box -12 -8 72 272
use NAND3X1  _888_
timestamp 1726536591
transform 1 0 470 0 1 3910
box -12 -8 112 272
use NAND2X1  _889_
timestamp 1726535706
transform 1 0 470 0 -1 5470
box -12 -8 92 272
use NOR2X1  _890_
timestamp 1726536993
transform 1 0 310 0 1 4430
box -12 -8 92 272
use OAI21X1  _891_
timestamp 1726538409
transform 1 0 290 0 -1 4430
box -12 -8 112 272
use AOI21X1  _892_
timestamp 1726549551
transform -1 0 530 0 -1 3910
box -12 -8 112 272
use AOI21X1  _893_
timestamp 1726549551
transform -1 0 570 0 1 3390
box -12 -8 112 272
use NAND3X1  _894_
timestamp 1726536591
transform -1 0 430 0 1 3910
box -12 -8 112 272
use OAI21X1  _895_
timestamp 1726538409
transform -1 0 250 0 -1 4430
box -12 -8 112 272
use AOI21X1  _896_
timestamp 1726549551
transform 1 0 190 0 1 3910
box -12 -8 112 272
use NAND2X1  _897_
timestamp 1726535706
transform -1 0 2430 0 1 3390
box -12 -8 92 272
use INVX1  _898_
timestamp 1726531033
transform 1 0 2110 0 -1 2870
box -12 -8 72 272
use INVX2  _899_
timestamp 1726533902
transform -1 0 3490 0 -1 3910
box -12 -8 72 272
use NAND2X1  _900_
timestamp 1726535706
transform -1 0 2310 0 1 3390
box -12 -8 92 272
use OAI21X1  _901_
timestamp 1726538409
transform -1 0 2230 0 -1 3390
box -12 -8 112 272
use OAI21X1  _902_
timestamp 1726538409
transform 1 0 2090 0 1 3390
box -12 -8 112 272
use OAI21X1  _903_
timestamp 1726538409
transform -1 0 390 0 -1 3910
box -12 -8 112 272
use NAND3X1  _904_
timestamp 1726536591
transform -1 0 150 0 1 3910
box -12 -8 112 272
use NAND3X1  _905_
timestamp 1726536591
transform 1 0 570 0 -1 3910
box -12 -8 112 272
use INVX1  _906_
timestamp 1726531033
transform -1 0 110 0 -1 3910
box -12 -8 72 272
use NAND3X1  _907_
timestamp 1726536591
transform 1 0 190 0 1 3390
box -12 -8 112 272
use NAND3X1  _908_
timestamp 1726536591
transform 1 0 330 0 1 3390
box -12 -8 112 272
use INVX1  _909_
timestamp 1726531033
transform -1 0 250 0 -1 2870
box -12 -8 72 272
use AOI21X1  _910_
timestamp 1726549551
transform -1 0 150 0 -1 2870
box -12 -8 112 272
use AOI21X1  _911_
timestamp 1726549551
transform -1 0 150 0 1 3390
box -12 -8 112 272
use INVX1  _912_
timestamp 1726531033
transform -1 0 110 0 -1 3390
box -12 -8 72 272
use OAI21X1  _913_
timestamp 1726538409
transform -1 0 150 0 1 2870
box -12 -8 112 272
use AOI21X1  _914_
timestamp 1726549551
transform 1 0 190 0 1 2350
box -12 -8 112 272
use NAND3X1  _915_
timestamp 1726536591
transform -1 0 150 0 1 2350
box -12 -8 112 272
use NAND2X1  _916_
timestamp 1726535706
transform 1 0 830 0 -1 2350
box -12 -8 92 272
use OAI22X1  _917_
timestamp 1726541006
transform -1 0 790 0 -1 2350
box -12 -8 132 272
use AND2X2  _918_
timestamp 1726549440
transform -1 0 1990 0 -1 3910
box -12 -8 112 273
use NAND2X1  _919_
timestamp 1726535706
transform -1 0 1350 0 -1 3910
box -12 -8 92 272
use INVX1  _920_
timestamp 1726531033
transform 1 0 1290 0 1 3910
box -12 -8 72 272
use AOI21X1  _921_
timestamp 1726549551
transform 1 0 150 0 -1 3910
box -12 -8 112 272
use NAND2X1  _922_
timestamp 1726535706
transform 1 0 2670 0 -1 3910
box -12 -8 92 272
use AND2X2  _923_
timestamp 1726549440
transform 1 0 2030 0 -1 3910
box -12 -8 112 273
use OAI21X1  _924_
timestamp 1726538409
transform 1 0 2170 0 -1 3910
box -12 -8 112 272
use INVX2  _925_
timestamp 1726533902
transform 1 0 3890 0 1 3910
box -12 -8 72 272
use OAI21X1  _926_
timestamp 1726538409
transform -1 0 2430 0 1 3910
box -12 -8 112 272
use NAND3X1  _927_
timestamp 1726536591
transform -1 0 2290 0 1 3910
box -12 -8 112 272
use INVX1  _928_
timestamp 1726531033
transform 1 0 2570 0 -1 3910
box -12 -8 72 272
use NAND2X1  _929_
timestamp 1726535706
transform -1 0 2390 0 -1 3910
box -12 -8 92 272
use OAI21X1  _930_
timestamp 1726538409
transform -1 0 2570 0 1 3390
box -12 -8 112 272
use NAND3X1  _931_
timestamp 1726536591
transform -1 0 2530 0 -1 3910
box -12 -8 112 272
use NAND2X1  _932_
timestamp 1726535706
transform 1 0 850 0 -1 4430
box -12 -8 92 272
use OAI22X1  _933_
timestamp 1726541006
transform -1 0 270 0 1 4430
box -12 -8 132 272
use INVX1  _934_
timestamp 1726531033
transform -1 0 390 0 1 4950
box -12 -8 72 272
use NAND2X1  _935_
timestamp 1726535706
transform 1 0 1030 0 -1 4950
box -12 -8 92 272
use NAND3X1  _936_
timestamp 1726536591
transform -1 0 690 0 -1 5470
box -12 -8 112 272
use NAND2X1  _937_
timestamp 1726535706
transform 1 0 730 0 -1 5470
box -12 -8 92 272
use NAND3X1  _938_
timestamp 1726536591
transform -1 0 430 0 -1 5470
box -12 -8 112 272
use NAND3X1  _939_
timestamp 1726536591
transform 1 0 190 0 -1 5470
box -12 -8 112 272
use INVX1  _940_
timestamp 1726531033
transform 1 0 710 0 1 4950
box -12 -8 72 272
use AND2X2  _941_
timestamp 1726549440
transform 1 0 1110 0 -1 5470
box -12 -8 112 273
use NAND2X1  _942_
timestamp 1726535706
transform 1 0 1090 0 1 4950
box -12 -8 92 272
use OAI21X1  _943_
timestamp 1726538409
transform -1 0 990 0 -1 4950
box -12 -8 112 272
use NAND3X1  _944_
timestamp 1726536591
transform -1 0 670 0 1 4950
box -12 -8 112 272
use NAND3X1  _945_
timestamp 1726536591
transform -1 0 430 0 -1 4950
box -12 -8 112 272
use AOI21X1  _946_
timestamp 1726549551
transform -1 0 530 0 1 4950
box -12 -8 112 272
use AOI21X1  _947_
timestamp 1726549551
transform -1 0 150 0 -1 5470
box -12 -8 112 272
use OAI21X1  _948_
timestamp 1726538409
transform -1 0 150 0 1 4950
box -12 -8 112 272
use NAND3X1  _949_
timestamp 1726536591
transform -1 0 150 0 -1 4950
box -12 -8 112 272
use AND2X2  _950_
timestamp 1726549440
transform -1 0 810 0 -1 4430
box -12 -8 112 273
use NAND3X1  _951_
timestamp 1726536591
transform -1 0 570 0 -1 4950
box -12 -8 112 272
use OAI21X1  _952_
timestamp 1726538409
transform 1 0 190 0 1 4950
box -12 -8 112 272
use NAND3X1  _953_
timestamp 1726536591
transform 1 0 430 0 -1 4430
box -12 -8 112 272
use NAND3X1  _954_
timestamp 1726536591
transform 1 0 610 0 1 3910
box -12 -8 112 272
use OAI21X1  _955_
timestamp 1726538409
transform 1 0 710 0 -1 3910
box -12 -8 112 272
use AOI21X1  _956_
timestamp 1726549551
transform 1 0 570 0 -1 4430
box -12 -8 112 272
use AOI21X1  _957_
timestamp 1726549551
transform 1 0 190 0 -1 4950
box -12 -8 112 272
use OAI21X1  _958_
timestamp 1726538409
transform 1 0 890 0 1 3910
box -12 -8 112 272
use NAND3X1  _959_
timestamp 1726536591
transform -1 0 1130 0 1 3910
box -12 -8 112 272
use NAND3X1  _960_
timestamp 1726536591
transform 1 0 850 0 -1 3910
box -12 -8 112 272
use OAI21X1  _961_
timestamp 1726538409
transform -1 0 850 0 1 3910
box -12 -8 112 272
use NAND3X1  _962_
timestamp 1726536591
transform -1 0 1230 0 -1 3910
box -12 -8 112 272
use NAND2X1  _963_
timestamp 1726535706
transform 1 0 1050 0 -1 3390
box -12 -8 92 272
use NAND2X1  _964_
timestamp 1726535706
transform -1 0 970 0 1 2870
box -12 -8 92 272
use XNOR2X1  _965_
timestamp 1726561449
transform 1 0 1010 0 1 2870
box -12 -8 152 272
use NAND2X1  _966_
timestamp 1726535706
transform 1 0 3310 0 1 2350
box -12 -8 92 272
use OAI21X1  _967_
timestamp 1726538409
transform -1 0 3270 0 1 2350
box -12 -8 112 272
use INVX1  _968_
timestamp 1726531033
transform 1 0 1810 0 -1 2350
box -12 -8 72 272
use AOI22X1  _969_
timestamp 1726480912
transform -1 0 1010 0 -1 3390
box -14 -8 132 272
use AOI21X1  _970_
timestamp 1726549551
transform 1 0 990 0 -1 3910
box -12 -8 112 272
use OAI21X1  _971_
timestamp 1726538409
transform 1 0 1390 0 -1 3910
box -12 -8 112 272
use NAND2X1  _972_
timestamp 1726535706
transform -1 0 2030 0 -1 4430
box -12 -8 92 272
use OAI21X1  _973_
timestamp 1726538409
transform -1 0 2150 0 1 3910
box -12 -8 112 272
use INVX1  _974_
timestamp 1726531033
transform -1 0 1250 0 -1 4430
box -12 -8 72 272
use INVX1  _975_
timestamp 1726531033
transform 1 0 430 0 1 4430
box -12 -8 72 272
use AOI21X1  _976_
timestamp 1726549551
transform 1 0 530 0 1 4430
box -12 -8 112 272
use NAND2X1  _977_
timestamp 1726535706
transform 1 0 2750 0 1 3910
box -12 -8 92 272
use AND2X2  _978_
timestamp 1726549440
transform -1 0 2970 0 1 3910
box -12 -8 112 273
use OAI21X1  _979_
timestamp 1726538409
transform -1 0 2710 0 1 3910
box -12 -8 112 272
use AND2X2  _980_
timestamp 1726549440
transform 1 0 1810 0 -1 4430
box -12 -8 112 273
use OAI21X1  _981_
timestamp 1726538409
transform 1 0 2430 0 -1 4430
box -12 -8 112 272
use NAND3X1  _982_
timestamp 1726536591
transform -1 0 2570 0 1 3910
box -12 -8 112 272
use INVX1  _983_
timestamp 1726531033
transform -1 0 2270 0 -1 4430
box -12 -8 72 272
use NAND2X1  _984_
timestamp 1726535706
transform 1 0 2310 0 -1 4430
box -12 -8 92 272
use OAI21X1  _985_
timestamp 1726538409
transform -1 0 2170 0 -1 4430
box -12 -8 112 272
use NAND3X1  _986_
timestamp 1726536591
transform 1 0 2150 0 1 4430
box -12 -8 112 272
use NAND2X1  _987_
timestamp 1726535706
transform -1 0 1970 0 1 4430
box -12 -8 92 272
use NOR2X1  _988_
timestamp 1726536993
transform 1 0 850 0 -1 5470
box -12 -8 92 272
use AOI21X1  _989_
timestamp 1726549551
transform 1 0 810 0 1 4950
box -12 -8 112 272
use NAND2X1  _990_
timestamp 1726535706
transform 1 0 2210 0 -1 5470
box -12 -8 92 272
use NAND2X1  _991_
timestamp 1726535706
transform -1 0 2550 0 1 4950
box -12 -8 92 272
use NAND3X1  _992_
timestamp 1726536591
transform -1 0 2430 0 1 4950
box -12 -8 112 272
use NAND2X1  _993_
timestamp 1726535706
transform 1 0 2730 0 1 4950
box -12 -8 92 272
use NAND3X1  _994_
timestamp 1726536591
transform -1 0 2690 0 1 4950
box -12 -8 112 272
use NAND3X1  _995_
timestamp 1726536591
transform -1 0 2150 0 1 4950
box -12 -8 112 272
use INVX1  _996_
timestamp 1726531033
transform -1 0 2170 0 -1 5470
box -12 -8 72 272
use AND2X2  _997_
timestamp 1726549440
transform -1 0 2550 0 -1 5470
box -12 -8 112 273
use NAND2X1  _998_
timestamp 1726535706
transform 1 0 1830 0 -1 5470
box -12 -8 92 272
use OAI21X1  _999_
timestamp 1726538409
transform -1 0 2450 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1000_
timestamp 1726536591
transform -1 0 1790 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1001_
timestamp 1726536591
transform -1 0 1730 0 1 4950
box -12 -8 112 272
use AOI22X1  _1002_
timestamp 1726480912
transform -1 0 1370 0 -1 5470
box -14 -8 132 272
use OAI21X1  _1003_
timestamp 1726538409
transform 1 0 1210 0 1 4950
box -12 -8 112 272
use AOI22X1  _1004_
timestamp 1726480912
transform 1 0 1530 0 -1 5470
box -14 -8 132 272
use AOI21X1  _1005_
timestamp 1726549551
transform -1 0 2290 0 1 4950
box -12 -8 112 272
use OAI21X1  _1006_
timestamp 1726538409
transform -1 0 1450 0 1 4950
box -12 -8 112 272
use NAND3X1  _1007_
timestamp 1726536591
transform -1 0 1510 0 -1 4950
box -12 -8 112 272
use AND2X2  _1008_
timestamp 1726549440
transform -1 0 2110 0 1 4430
box -12 -8 112 273
use NAND3X1  _1009_
timestamp 1726536591
transform 1 0 1770 0 1 4950
box -12 -8 112 272
use OAI21X1  _1010_
timestamp 1726538409
transform -1 0 1590 0 1 4950
box -12 -8 112 272
use NAND3X1  _1011_
timestamp 1726536591
transform -1 0 1790 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1012_
timestamp 1726536591
transform -1 0 1170 0 1 4430
box -12 -8 112 272
use AOI21X1  _1013_
timestamp 1726549551
transform 1 0 610 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1014_
timestamp 1726538409
transform -1 0 850 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1015_
timestamp 1726549551
transform -1 0 1930 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1016_
timestamp 1726549551
transform 1 0 1550 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1017_
timestamp 1726538409
transform -1 0 1590 0 1 4430
box -12 -8 112 272
use NAND3X1  _1018_
timestamp 1726536591
transform -1 0 1390 0 -1 4430
box -12 -8 112 272
use NAND3X1  _1019_
timestamp 1726536591
transform 1 0 1210 0 1 4430
box -12 -8 112 272
use OAI21X1  _1020_
timestamp 1726538409
transform -1 0 1730 0 1 4430
box -12 -8 112 272
use NAND3X1  _1021_
timestamp 1726536591
transform -1 0 1730 0 1 3910
box -12 -8 112 272
use NAND2X1  _1022_
timestamp 1726535706
transform 1 0 1670 0 -1 3910
box -12 -8 92 272
use XNOR2X1  _1023_
timestamp 1726561449
transform -1 0 1550 0 -1 3390
box -12 -8 152 272
use NOR2X1  _1024_
timestamp 1726536993
transform -1 0 1950 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1025_
timestamp 1726536591
transform -1 0 1630 0 -1 3910
box -12 -8 112 272
use INVX1  _1026_
timestamp 1726531033
transform 1 0 1530 0 1 3910
box -12 -8 72 272
use AOI21X1  _1027_
timestamp 1726549551
transform 1 0 1390 0 1 3910
box -12 -8 112 272
use AOI21X1  _1028_
timestamp 1726549551
transform 1 0 1910 0 1 3910
box -12 -8 112 272
use AOI21X1  _1029_
timestamp 1726549551
transform 1 0 1430 0 -1 4430
box -12 -8 112 272
use OAI21X1  _1030_
timestamp 1726538409
transform -1 0 1870 0 1 3910
box -12 -8 112 272
use NAND3X1  _1031_
timestamp 1726536591
transform 1 0 1730 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1032_
timestamp 1726535706
transform -1 0 1970 0 1 2870
box -12 -8 92 272
use OAI22X1  _1033_
timestamp 1726541006
transform 1 0 1850 0 1 2350
box -12 -8 132 272
use OAI21X1  _1034_
timestamp 1726538409
transform 1 0 1590 0 -1 3390
box -12 -8 112 272
use INVX1  _1035_
timestamp 1726531033
transform 1 0 1570 0 -1 4430
box -12 -8 72 272
use AOI21X1  _1036_
timestamp 1726549551
transform 1 0 1670 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1037_
timestamp 1726535706
transform -1 0 2370 0 1 4430
box -12 -8 92 272
use INVX1  _1038_
timestamp 1726531033
transform 1 0 3110 0 1 4430
box -12 -8 72 272
use INVX1  _1039_
timestamp 1726531033
transform 1 0 2110 0 -1 4950
box -12 -8 72 272
use AOI21X1  _1040_
timestamp 1726549551
transform 1 0 2210 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1041_
timestamp 1726535706
transform -1 0 3130 0 -1 4430
box -12 -8 92 272
use AND2X2  _1042_
timestamp 1726549440
transform 1 0 3570 0 -1 4430
box -12 -8 112 273
use OAI21X1  _1043_
timestamp 1726538409
transform 1 0 3310 0 -1 4430
box -12 -8 112 272
use AND2X2  _1044_
timestamp 1726549440
transform 1 0 2910 0 -1 4430
box -12 -8 112 273
use OAI21X1  _1045_
timestamp 1726538409
transform -1 0 3110 0 1 3910
box -12 -8 112 272
use NAND3X1  _1046_
timestamp 1726536591
transform -1 0 3270 0 -1 4430
box -12 -8 112 272
use INVX1  _1047_
timestamp 1726531033
transform 1 0 3350 0 1 4430
box -12 -8 72 272
use NAND2X1  _1048_
timestamp 1726535706
transform 1 0 3450 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1049_
timestamp 1726535706
transform 1 0 3670 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1050_
timestamp 1726538409
transform 1 0 3530 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1051_
timestamp 1726536591
transform -1 0 3550 0 1 4430
box -12 -8 112 272
use NAND2X1  _1052_
timestamp 1726535706
transform -1 0 3270 0 -1 4950
box -12 -8 92 272
use AOI22X1  _1053_
timestamp 1726480912
transform 1 0 1950 0 -1 5470
box -14 -8 132 272
use NAND2X1  _1054_
timestamp 1726535706
transform -1 0 4030 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1055_
timestamp 1726535706
transform -1 0 4070 0 1 4950
box -12 -8 92 272
use NOR2X1  _1056_
timestamp 1726536993
transform 1 0 4110 0 1 4950
box -12 -8 92 272
use AOI22X1  _1057_
timestamp 1726480912
transform -1 0 3950 0 1 4950
box -14 -8 132 272
use OAI21X1  _1058_
timestamp 1726538409
transform -1 0 4170 0 -1 5470
box -12 -8 112 272
use INVX1  _1059_
timestamp 1726531033
transform 1 0 4590 0 -1 5470
box -12 -8 72 272
use AND2X2  _1060_
timestamp 1726549440
transform -1 0 3790 0 1 4950
box -12 -8 112 273
use NAND2X1  _1061_
timestamp 1726535706
transform -1 0 4310 0 1 4950
box -12 -8 92 272
use INVX1  _1062_
timestamp 1726531033
transform 1 0 4490 0 -1 5470
box -12 -8 72 272
use NAND3X1  _1063_
timestamp 1726536591
transform -1 0 4450 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1064_
timestamp 1726536591
transform 1 0 3390 0 -1 5470
box -12 -8 112 272
use AOI22X1  _1065_
timestamp 1726480912
transform 1 0 2730 0 -1 5470
box -14 -8 132 272
use OAI21X1  _1066_
timestamp 1726538409
transform 1 0 2590 0 -1 5470
box -12 -8 112 272
use AOI21X1  _1067_
timestamp 1726549551
transform -1 0 4310 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1068_
timestamp 1726538409
transform 1 0 3670 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1069_
timestamp 1726538409
transform 1 0 3530 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1070_
timestamp 1726549551
transform 1 0 3810 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1071_
timestamp 1726538409
transform -1 0 3770 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1072_
timestamp 1726536591
transform -1 0 3510 0 1 4950
box -12 -8 112 272
use AND2X2  _1073_
timestamp 1726549440
transform -1 0 3150 0 -1 4950
box -12 -8 112 273
use NAND3X1  _1074_
timestamp 1726536591
transform -1 0 3350 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1075_
timestamp 1726538409
transform -1 0 3910 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1076_
timestamp 1726536591
transform -1 0 3230 0 1 4950
box -12 -8 112 272
use NAND3X1  _1077_
timestamp 1726536591
transform 1 0 2850 0 1 4950
box -12 -8 112 272
use AOI21X1  _1078_
timestamp 1726549551
transform 1 0 1910 0 1 4950
box -12 -8 112 272
use OAI21X1  _1079_
timestamp 1726538409
transform 1 0 1970 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1080_
timestamp 1726549551
transform -1 0 3090 0 1 4950
box -12 -8 112 272
use AOI21X1  _1081_
timestamp 1726549551
transform -1 0 3370 0 1 4950
box -12 -8 112 272
use OAI21X1  _1082_
timestamp 1726538409
transform 1 0 2630 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1083_
timestamp 1726549551
transform -1 0 2930 0 1 4430
box -12 -8 112 272
use NAND3X1  _1084_
timestamp 1726536591
transform -1 0 2870 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1085_
timestamp 1726538409
transform -1 0 2590 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1086_
timestamp 1726549551
transform 1 0 2690 0 1 4430
box -12 -8 112 272
use OAI21X1  _1087_
timestamp 1726538409
transform -1 0 2770 0 -1 4430
box -12 -8 112 272
use AOI21X1  _1088_
timestamp 1726549551
transform 1 0 1270 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1089_
timestamp 1726538409
transform 1 0 1350 0 1 4430
box -12 -8 112 272
use NAND3X1  _1090_
timestamp 1726536591
transform -1 0 2650 0 1 4430
box -12 -8 112 272
use NAND3X1  _1091_
timestamp 1726536591
transform 1 0 2970 0 1 4430
box -12 -8 112 272
use NAND3X1  _1092_
timestamp 1726536591
transform 1 0 2410 0 1 4430
box -12 -8 112 272
use NAND2X1  _1093_
timestamp 1726535706
transform 1 0 2530 0 -1 3390
box -12 -8 92 272
use XOR2X1  _1094_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726561008
transform 1 0 1710 0 1 2870
box -12 -8 152 272
use NAND2X1  _1095_
timestamp 1726535706
transform -1 0 890 0 1 1830
box -12 -8 92 272
use OAI21X1  _1096_
timestamp 1726538409
transform -1 0 1030 0 1 1830
box -12 -8 112 272
use NAND2X1  _1097_
timestamp 1726535706
transform 1 0 4530 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1098_
timestamp 1726535706
transform -1 0 2350 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1099_
timestamp 1726535706
transform -1 0 2730 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1100_
timestamp 1726538409
transform 1 0 2770 0 -1 3390
box -12 -8 112 272
use AOI21X1  _1101_
timestamp 1726549551
transform 1 0 2910 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1102_
timestamp 1726538409
transform 1 0 3210 0 1 4430
box -12 -8 112 272
use NAND2X1  _1103_
timestamp 1726535706
transform 1 0 3590 0 1 4430
box -12 -8 92 272
use INVX1  _1104_
timestamp 1726531033
transform 1 0 5670 0 1 4950
box -12 -8 72 272
use INVX1  _1105_
timestamp 1726531033
transform 1 0 3010 0 -1 5470
box -12 -8 72 272
use AOI21X1  _1106_
timestamp 1726549551
transform 1 0 3110 0 -1 5470
box -12 -8 112 272
use INVX2  _1107_
timestamp 1726533902
transform 1 0 3790 0 1 3910
box -12 -8 72 272
use NOR2X1  _1108_
timestamp 1726536993
transform 1 0 3670 0 1 3910
box -12 -8 92 272
use AND2X2  _1109_
timestamp 1726549440
transform 1 0 3870 0 -1 4430
box -12 -8 112 273
use AOI22X1  _1110_
timestamp 1726480912
transform 1 0 3710 0 -1 4430
box -14 -8 132 272
use AOI21X1  _1111_
timestamp 1726549551
transform 1 0 4010 0 -1 4430
box -12 -8 112 272
use XNOR2X1  _1112_
timestamp 1726561449
transform 1 0 4150 0 1 4430
box -12 -8 152 272
use AOI21X1  _1113_
timestamp 1726549551
transform 1 0 4690 0 -1 5470
box -12 -8 112 272
use NAND2X1  _1114_
timestamp 1726535706
transform -1 0 4030 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1115_
timestamp 1726535706
transform -1 0 3990 0 1 4430
box -12 -8 92 272
use NAND2X1  _1116_
timestamp 1726535706
transform -1 0 4110 0 1 4430
box -12 -8 92 272
use OAI21X1  _1117_
timestamp 1726538409
transform 1 0 4070 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1118_
timestamp 1726538409
transform 1 0 4210 0 -1 4950
box -12 -8 112 272
use NOR2X1  _1119_
timestamp 1726536993
transform -1 0 4830 0 1 4950
box -12 -8 92 272
use OAI21X1  _1120_
timestamp 1726538409
transform -1 0 4450 0 1 4950
box -12 -8 112 272
use XOR2X1  _1121_
timestamp 1726561008
transform -1 0 4490 0 -1 4950
box -12 -8 152 272
use NOR2X1  _1122_
timestamp 1726536993
transform 1 0 4490 0 1 4950
box -12 -8 92 272
use OAI21X1  _1123_
timestamp 1726538409
transform 1 0 4950 0 -1 4950
box -12 -8 112 272
use XOR2X1  _1124_
timestamp 1726561008
transform 1 0 4470 0 1 4430
box -12 -8 152 272
use OAI21X1  _1125_
timestamp 1726538409
transform -1 0 4710 0 1 4950
box -12 -8 112 272
use NAND2X1  _1126_
timestamp 1726535706
transform 1 0 4870 0 1 4950
box -12 -8 92 272
use NAND3X1  _1127_
timestamp 1726536591
transform 1 0 4990 0 1 4950
box -12 -8 112 272
use NAND3X1  _1128_
timestamp 1726536591
transform 1 0 5130 0 1 4950
box -12 -8 112 272
use AOI21X1  _1129_
timestamp 1726549551
transform 1 0 3530 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1130_
timestamp 1726538409
transform 1 0 3550 0 1 4950
box -12 -8 112 272
use AOI21X1  _1131_
timestamp 1726549551
transform 1 0 4970 0 -1 5470
box -12 -8 112 272
use NAND2X1  _1132_
timestamp 1726535706
transform 1 0 5110 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1133_
timestamp 1726538409
transform 1 0 4830 0 -1 5470
box -12 -8 112 272
use AOI21X1  _1134_
timestamp 1726549551
transform 1 0 5230 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1135_
timestamp 1726538409
transform -1 0 5470 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1136_
timestamp 1726536591
transform 1 0 5530 0 1 4950
box -12 -8 112 272
use NAND3X1  _1137_
timestamp 1726536591
transform 1 0 5230 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1138_
timestamp 1726538409
transform 1 0 5510 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1139_
timestamp 1726536591
transform 1 0 5550 0 1 4430
box -12 -8 112 272
use NAND3X1  _1140_
timestamp 1726536591
transform 1 0 5410 0 1 4430
box -12 -8 112 272
use INVX1  _1141_
timestamp 1726531033
transform -1 0 5370 0 1 4430
box -12 -8 72 272
use AOI21X1  _1142_
timestamp 1726549551
transform -1 0 5610 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1143_
timestamp 1726549551
transform -1 0 5370 0 1 4950
box -12 -8 112 272
use OAI21X1  _1144_
timestamp 1726538409
transform -1 0 5470 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1145_
timestamp 1726535706
transform 1 0 5310 0 -1 3390
box -12 -8 92 272
use XOR2X1  _1146_
timestamp 1726561008
transform 1 0 5010 0 -1 3390
box -12 -8 152 272
use OAI21X1  _1147_
timestamp 1726538409
transform 1 0 4650 0 -1 2870
box -12 -8 112 272
use INVX1  _1148_
timestamp 1726531033
transform -1 0 5630 0 -1 3390
box -12 -8 72 272
use AOI21X1  _1149_
timestamp 1726549551
transform 1 0 5430 0 -1 3390
box -12 -8 112 272
use AOI22X1  _1150_
timestamp 1726480912
transform 1 0 4150 0 -1 4430
box -14 -8 132 272
use INVX1  _1151_
timestamp 1726531033
transform -1 0 4890 0 -1 4430
box -12 -8 72 272
use OAI21X1  _1152_
timestamp 1726538409
transform 1 0 4670 0 -1 4950
box -12 -8 112 272
use NOR2X1  _1153_
timestamp 1726536993
transform -1 0 4250 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1154_
timestamp 1726535706
transform 1 0 3910 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1155_
timestamp 1726535706
transform 1 0 4370 0 1 3390
box -12 -8 92 272
use OR2X2  _1156_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726542447
transform 1 0 4290 0 -1 3910
box -12 -8 112 272
use OAI21X1  _1157_
timestamp 1726538409
transform 1 0 4030 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1158_
timestamp 1726536591
transform 1 0 4430 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1159_
timestamp 1726535706
transform 1 0 4110 0 1 3910
box -12 -8 92 272
use NAND2X1  _1160_
timestamp 1726535706
transform -1 0 4070 0 1 3910
box -12 -8 92 272
use OAI21X1  _1161_
timestamp 1726538409
transform -1 0 4470 0 1 3910
box -12 -8 112 272
use OAI21X1  _1162_
timestamp 1726538409
transform 1 0 4230 0 1 3910
box -12 -8 112 272
use NAND2X1  _1163_
timestamp 1726535706
transform -1 0 4510 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1164_
timestamp 1726538409
transform 1 0 4330 0 1 4430
box -12 -8 112 272
use NOR2X1  _1165_
timestamp 1726536993
transform -1 0 4390 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1166_
timestamp 1726536591
transform 1 0 4550 0 -1 4430
box -12 -8 112 272
use NAND3X1  _1167_
timestamp 1726536591
transform 1 0 4650 0 1 4430
box -12 -8 112 272
use AOI21X1  _1168_
timestamp 1726549551
transform -1 0 4910 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1169_
timestamp 1726549551
transform 1 0 4690 0 -1 4430
box -12 -8 112 272
use INVX1  _1170_
timestamp 1726531033
transform 1 0 5210 0 1 4430
box -12 -8 72 272
use OAI21X1  _1171_
timestamp 1726538409
transform 1 0 5070 0 1 4430
box -12 -8 112 272
use NAND3X1  _1172_
timestamp 1726536591
transform 1 0 5070 0 -1 4430
box -12 -8 112 272
use NAND3X1  _1173_
timestamp 1726536591
transform 1 0 4790 0 1 4430
box -12 -8 112 272
use OAI21X1  _1174_
timestamp 1726538409
transform -1 0 5030 0 1 4430
box -12 -8 112 272
use NAND3X1  _1175_
timestamp 1726536591
transform 1 0 4930 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1176_
timestamp 1726535706
transform -1 0 5410 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1177_
timestamp 1726536591
transform 1 0 5450 0 -1 4430
box -12 -8 112 272
use AOI21X1  _1178_
timestamp 1726549551
transform 1 0 5090 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1179_
timestamp 1726538409
transform 1 0 5650 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1180_
timestamp 1726536591
transform 1 0 5590 0 -1 4430
box -12 -8 112 272
use AND2X2  _1181_
timestamp 1726549440
transform 1 0 5570 0 -1 3910
box -12 -8 112 273
use XOR2X1  _1182_
timestamp 1726561008
transform -1 0 5670 0 1 2870
box -12 -8 152 272
use NAND2X1  _1183_
timestamp 1726535706
transform 1 0 5410 0 1 4950
box -12 -8 92 272
use OAI21X1  _1184_
timestamp 1726538409
transform -1 0 5630 0 1 1830
box -12 -8 112 272
use INVX1  _1185_
timestamp 1726531033
transform -1 0 5010 0 1 2350
box -12 -8 72 272
use NAND2X1  _1186_
timestamp 1726535706
transform 1 0 5330 0 -1 3910
box -12 -8 92 272
use NOR2X1  _1187_
timestamp 1726536993
transform 1 0 5190 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1188_
timestamp 1726535706
transform -1 0 5370 0 1 3910
box -12 -8 92 272
use NAND2X1  _1189_
timestamp 1726535706
transform -1 0 5250 0 1 3910
box -12 -8 92 272
use INVX1  _1190_
timestamp 1726531033
transform 1 0 5330 0 1 3390
box -12 -8 72 272
use AOI21X1  _1191_
timestamp 1726549551
transform 1 0 5270 0 1 2870
box -12 -8 112 272
use NAND2X1  _1192_
timestamp 1726535706
transform 1 0 5210 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1193_
timestamp 1726538409
transform 1 0 4510 0 1 3910
box -12 -8 112 272
use INVX1  _1194_
timestamp 1726531033
transform -1 0 4630 0 -1 3910
box -12 -8 72 272
use OR2X2  _1195_
timestamp 1726542447
transform 1 0 4530 0 -1 4950
box -12 -8 112 272
use NOR2X1  _1196_
timestamp 1726536993
transform 1 0 3790 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1197_
timestamp 1726538409
transform 1 0 4490 0 1 3390
box -12 -8 112 272
use NAND2X1  _1198_
timestamp 1726535706
transform -1 0 4090 0 1 3390
box -12 -8 92 272
use OAI21X1  _1199_
timestamp 1726538409
transform -1 0 4730 0 1 3390
box -12 -8 112 272
use XOR2X1  _1200_
timestamp 1726561008
transform 1 0 4930 0 1 3390
box -12 -8 152 272
use AOI21X1  _1201_
timestamp 1726549551
transform 1 0 4650 0 1 3910
box -12 -8 112 272
use NAND3X1  _1202_
timestamp 1726536591
transform 1 0 4790 0 1 3910
box -12 -8 112 272
use INVX1  _1203_
timestamp 1726531033
transform -1 0 4870 0 -1 3910
box -12 -8 72 272
use OAI21X1  _1204_
timestamp 1726538409
transform -1 0 4770 0 -1 3910
box -12 -8 112 272
use INVX1  _1205_
timestamp 1726531033
transform 1 0 4930 0 1 3910
box -12 -8 72 272
use NAND3X1  _1206_
timestamp 1726536591
transform 1 0 5030 0 1 3910
box -12 -8 112 272
use AND2X2  _1207_
timestamp 1726549440
transform 1 0 5050 0 -1 3910
box -12 -8 112 273
use NAND2X1  _1208_
timestamp 1726535706
transform 1 0 5210 0 1 3390
box -12 -8 92 272
use OR2X2  _1209_
timestamp 1726542447
transform -1 0 5290 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1210_
timestamp 1726535706
transform -1 0 4870 0 1 2870
box -12 -8 92 272
use NAND2X1  _1211_
timestamp 1726535706
transform -1 0 4990 0 1 2870
box -12 -8 92 272
use AND2X2  _1212_
timestamp 1726549440
transform -1 0 2490 0 -1 3390
box -12 -8 112 273
use NAND3X1  _1213_
timestamp 1726536591
transform 1 0 1990 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1214_
timestamp 1726536591
transform 1 0 5610 0 1 3390
box -12 -8 112 272
use AOI21X1  _1215_
timestamp 1726549551
transform 1 0 2910 0 -1 3390
box -12 -8 112 272
use INVX1  _1216_
timestamp 1726531033
transform 1 0 5030 0 1 2870
box -12 -8 72 272
use OAI21X1  _1217_
timestamp 1726538409
transform -1 0 5230 0 1 2870
box -12 -8 112 272
use NAND3X1  _1218_
timestamp 1726536591
transform 1 0 5050 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1219_
timestamp 1726538409
transform 1 0 5050 0 1 2350
box -12 -8 112 272
use NAND2X1  _1220_
timestamp 1726535706
transform 1 0 5550 0 1 2350
box -12 -8 92 272
use AOI21X1  _1221_
timestamp 1726549551
transform -1 0 5010 0 -1 3910
box -12 -8 112 272
use INVX1  _1222_
timestamp 1726531033
transform 1 0 5110 0 1 3390
box -12 -8 72 272
use OAI22X1  _1223_
timestamp 1726541006
transform 1 0 4770 0 1 3390
box -12 -8 132 272
use OAI21X1  _1224_
timestamp 1726538409
transform 1 0 4050 0 -1 3390
box -12 -8 112 272
use NOR2X1  _1225_
timestamp 1726536993
transform 1 0 3790 0 -1 3390
box -12 -8 92 272
use INVX1  _1226_
timestamp 1726531033
transform -1 0 3750 0 -1 3390
box -12 -8 72 272
use OR2X2  _1227_
timestamp 1726542447
transform 1 0 3750 0 1 2870
box -12 -8 112 272
use AND2X2  _1228_
timestamp 1726549440
transform 1 0 4190 0 -1 3390
box -12 -8 112 273
use XNOR2X1  _1229_
timestamp 1726561449
transform 1 0 4450 0 -1 3390
box -12 -8 152 272
use XOR2X1  _1230_
timestamp 1726561008
transform 1 0 5430 0 1 3390
box -12 -8 152 272
use INVX1  _1231_
timestamp 1726531033
transform 1 0 5470 0 -1 2870
box -12 -8 72 272
use NAND3X1  _1232_
timestamp 1726536591
transform 1 0 5190 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1233_
timestamp 1726538409
transform -1 0 4890 0 -1 2870
box -12 -8 112 272
use NAND2X1  _1234_
timestamp 1726535706
transform -1 0 5010 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1235_
timestamp 1726536591
transform 1 0 5330 0 -1 2870
box -12 -8 112 272
use NAND2X1  _1236_
timestamp 1726535706
transform -1 0 5510 0 1 2350
box -12 -8 92 272
use INVX1  _1237_
timestamp 1726531033
transform 1 0 3910 0 1 2350
box -12 -8 72 272
use NOR2X1  _1238_
timestamp 1726536993
transform 1 0 4890 0 -1 3390
box -12 -8 92 272
use AOI21X1  _1239_
timestamp 1726549551
transform -1 0 4850 0 -1 3390
box -12 -8 112 272
use NOR2X1  _1240_
timestamp 1726536993
transform -1 0 4710 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1241_
timestamp 1726536591
transform -1 0 4750 0 1 2870
box -12 -8 112 272
use OAI21X1  _1242_
timestamp 1726538409
transform -1 0 4610 0 1 2870
box -12 -8 112 272
use NAND2X1  _1243_
timestamp 1726535706
transform -1 0 4410 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1244_
timestamp 1726538409
transform 1 0 3550 0 -1 3390
box -12 -8 112 272
use OR2X2  _1245_
timestamp 1726542447
transform 1 0 3910 0 -1 3390
box -12 -8 112 272
use INVX1  _1246_
timestamp 1726531033
transform -1 0 3950 0 1 2870
box -12 -8 72 272
use OAI21X1  _1247_
timestamp 1726538409
transform -1 0 3710 0 1 2870
box -12 -8 112 272
use AND2X2  _1248_
timestamp 1726549440
transform -1 0 3770 0 -1 2870
box -12 -8 112 273
use NOR2X1  _1249_
timestamp 1726536993
transform 1 0 4030 0 -1 2870
box -12 -8 92 272
use INVX1  _1250_
timestamp 1726531033
transform -1 0 4330 0 1 2870
box -12 -8 72 272
use OAI21X1  _1251_
timestamp 1726538409
transform 1 0 4370 0 1 2870
box -12 -8 112 272
use AOI21X1  _1252_
timestamp 1726549551
transform -1 0 4230 0 1 2870
box -12 -8 112 272
use INVX1  _1253_
timestamp 1726531033
transform 1 0 3930 0 -1 2870
box -12 -8 72 272
use OAI21X1  _1254_
timestamp 1726538409
transform 1 0 4150 0 -1 2870
box -12 -8 112 272
use OAI22X1  _1255_
timestamp 1726541006
transform 1 0 4010 0 1 2350
box -12 -8 132 272
use INVX1  _1256_
timestamp 1726531033
transform 1 0 4630 0 1 790
box -12 -8 72 272
use AOI21X1  _1257_
timestamp 1726549551
transform -1 0 4090 0 1 2870
box -12 -8 112 272
use AND2X2  _1258_
timestamp 1726549440
transform 1 0 4170 0 1 2350
box -12 -8 112 273
use AOI22X1  _1259_
timestamp 1726480912
transform -1 0 4430 0 1 2350
box -14 -8 132 272
use NOR2X1  _1260_
timestamp 1726536993
transform -1 0 2450 0 1 1830
box -12 -8 92 272
use INVX1  _1261_
timestamp 1726531033
transform 1 0 2390 0 -1 1830
box -12 -8 72 272
use NAND2X1  _1262_
timestamp 1726535706
transform -1 0 2570 0 1 1830
box -12 -8 92 272
use NAND2X1  _1263_
timestamp 1726535706
transform -1 0 2570 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1264_
timestamp 1726535706
transform -1 0 3190 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1265_
timestamp 1726538409
transform 1 0 2970 0 -1 1830
box -12 -8 112 272
use INVX1  _1266_
timestamp 1726531033
transform 1 0 550 0 1 1310
box -12 -8 72 272
use NOR2X1  _1267_
timestamp 1726536993
transform 1 0 890 0 -1 1310
box -12 -8 92 272
use NOR2X1  _1268_
timestamp 1726536993
transform 1 0 430 0 1 1310
box -12 -8 92 272
use NOR2X1  _1269_
timestamp 1726536993
transform -1 0 1210 0 1 1310
box -12 -8 92 272
use NAND2X1  _1270_
timestamp 1726535706
transform -1 0 1470 0 1 1310
box -12 -8 92 272
use OAI21X1  _1271_
timestamp 1726538409
transform 1 0 1250 0 1 1310
box -12 -8 112 272
use NAND2X1  _1272_
timestamp 1726535706
transform 1 0 1370 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1273_
timestamp 1726535706
transform 1 0 1870 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1274_
timestamp 1726538409
transform -1 0 1590 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1275_
timestamp 1726538409
transform 1 0 750 0 -1 1310
box -12 -8 112 272
use XOR2X1  _1276_
timestamp 1726561008
transform -1 0 190 0 -1 790
box -12 -8 152 272
use XNOR2X1  _1277_
timestamp 1726561449
transform -1 0 730 0 -1 790
box -12 -8 152 272
use NAND2X1  _1278_
timestamp 1726535706
transform 1 0 1390 0 -1 790
box -12 -8 92 272
use OAI21X1  _1279_
timestamp 1726538409
transform 1 0 1250 0 -1 790
box -12 -8 112 272
use NOR2X1  _1280_
timestamp 1726536993
transform -1 0 410 0 -1 790
box -12 -8 92 272
use AOI21X1  _1281_
timestamp 1726549551
transform -1 0 550 0 -1 790
box -12 -8 112 272
use NOR2X1  _1282_
timestamp 1726536993
transform -1 0 130 0 1 790
box -12 -8 92 272
use NOR2X1  _1283_
timestamp 1726536993
transform -1 0 250 0 1 790
box -12 -8 92 272
use NOR2X1  _1284_
timestamp 1726536993
transform -1 0 370 0 1 790
box -12 -8 92 272
use XOR2X1  _1285_
timestamp 1726561008
transform 1 0 650 0 1 790
box -12 -8 152 272
use NAND2X1  _1286_
timestamp 1726535706
transform 1 0 1330 0 1 790
box -12 -8 92 272
use OAI21X1  _1287_
timestamp 1726538409
transform 1 0 950 0 1 790
box -12 -8 112 272
use NAND2X1  _1288_
timestamp 1726535706
transform -1 0 3550 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1289_
timestamp 1726535706
transform -1 0 1510 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1290_
timestamp 1726535706
transform -1 0 1230 0 1 2350
box -12 -8 92 272
use AND2X2  _1291_
timestamp 1726549440
transform 1 0 1610 0 1 2350
box -12 -8 112 273
use INVX1  _1292_
timestamp 1726531033
transform 1 0 1750 0 1 2350
box -12 -8 72 272
use INVX1  _1293_
timestamp 1726531033
transform 1 0 410 0 1 790
box -12 -8 72 272
use OAI21X1  _1294_
timestamp 1726538409
transform 1 0 510 0 1 790
box -12 -8 112 272
use INVX1  _1295_
timestamp 1726531033
transform 1 0 1910 0 -1 2350
box -12 -8 72 272
use NAND2X1  _1296_
timestamp 1726535706
transform -1 0 2090 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1297_
timestamp 1726535706
transform 1 0 1690 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1298_
timestamp 1726535706
transform 1 0 2130 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1299_
timestamp 1726538409
transform 1 0 3330 0 -1 2350
box -12 -8 112 272
use NAND2X1  _1300_
timestamp 1726535706
transform 1 0 2610 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1301_
timestamp 1726538409
transform 1 0 1550 0 -1 2350
box -12 -8 112 272
use OR2X2  _1302_
timestamp 1726542447
transform -1 0 3010 0 1 2350
box -12 -8 112 272
use NAND2X1  _1303_
timestamp 1726535706
transform 1 0 3050 0 1 2350
box -12 -8 92 272
use AND2X2  _1304_
timestamp 1726549440
transform -1 0 2870 0 1 2350
box -12 -8 112 273
use NOR2X1  _1305_
timestamp 1726536993
transform -1 0 2430 0 -1 2350
box -12 -8 92 272
use INVX1  _1306_
timestamp 1726531033
transform 1 0 2250 0 -1 2350
box -12 -8 72 272
use INVX1  _1307_
timestamp 1726531033
transform 1 0 2550 0 1 2350
box -12 -8 72 272
use OAI21X1  _1308_
timestamp 1726538409
transform 1 0 2410 0 1 2350
box -12 -8 112 272
use OAI21X1  _1309_
timestamp 1726538409
transform 1 0 2470 0 -1 2350
box -12 -8 112 272
use NAND2X1  _1310_
timestamp 1726535706
transform -1 0 2010 0 1 1310
box -12 -8 92 272
use OAI21X1  _1311_
timestamp 1726538409
transform -1 0 2370 0 1 2350
box -12 -8 112 272
use XOR2X1  _1312_
timestamp 1726561008
transform 1 0 1550 0 1 1830
box -12 -8 152 272
use NOR2X1  _1313_
timestamp 1726536993
transform 1 0 2270 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1314_
timestamp 1726535706
transform 1 0 2250 0 1 1830
box -12 -8 92 272
use NAND2X1  _1315_
timestamp 1726535706
transform 1 0 2150 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1316_
timestamp 1726538409
transform -1 0 2150 0 1 1310
box -12 -8 112 272
use OAI21X1  _1317_
timestamp 1726538409
transform 1 0 2010 0 -1 1830
box -12 -8 112 272
use NOR2X1  _1318_
timestamp 1726536993
transform 1 0 1150 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1319_
timestamp 1726535706
transform -1 0 1110 0 -1 1830
box -12 -8 92 272
use INVX1  _1320_
timestamp 1726531033
transform 1 0 1070 0 1 1830
box -12 -8 72 272
use NOR2X1  _1321_
timestamp 1726536993
transform 1 0 1270 0 -1 1830
box -12 -8 92 272
use XNOR2X1  _1322_
timestamp 1726561449
transform -1 0 1890 0 1 1310
box -12 -8 152 272
use NAND2X1  _1323_
timestamp 1726535706
transform 1 0 2110 0 1 790
box -12 -8 92 272
use OAI21X1  _1324_
timestamp 1726538409
transform -1 0 1830 0 1 790
box -12 -8 112 272
use NAND2X1  _1325_
timestamp 1726535706
transform 1 0 4410 0 1 1310
box -12 -8 92 272
use OAI21X1  _1326_
timestamp 1726538409
transform 1 0 2130 0 1 2350
box -12 -8 112 272
use NAND2X1  _1327_
timestamp 1726535706
transform -1 0 1390 0 1 1830
box -12 -8 92 272
use OAI21X1  _1328_
timestamp 1726538409
transform -1 0 1270 0 1 1830
box -12 -8 112 272
use AND2X2  _1329_
timestamp 1726549440
transform 1 0 1730 0 -1 1830
box -12 -8 112 273
use AOI21X1  _1330_
timestamp 1726549551
transform -1 0 1830 0 1 1830
box -12 -8 112 272
use NOR2X1  _1331_
timestamp 1726536993
transform -1 0 2090 0 1 2350
box -12 -8 92 272
use NAND3X1  _1332_
timestamp 1726536591
transform -1 0 1970 0 1 1830
box -12 -8 112 272
use NAND2X1  _1333_
timestamp 1726535706
transform 1 0 2010 0 1 1830
box -12 -8 92 272
use OR2X2  _1334_
timestamp 1726542447
transform 1 0 4430 0 -1 2350
box -12 -8 112 272
use NAND2X1  _1335_
timestamp 1726535706
transform -1 0 4390 0 -1 2350
box -12 -8 92 272
use AND2X2  _1336_
timestamp 1726549440
transform 1 0 4570 0 -1 2350
box -12 -8 112 273
use NOR2X1  _1337_
timestamp 1726536993
transform -1 0 4550 0 -1 1830
box -12 -8 92 272
use INVX1  _1338_
timestamp 1726531033
transform -1 0 4790 0 -1 1830
box -12 -8 72 272
use INVX1  _1339_
timestamp 1726531033
transform 1 0 4650 0 1 1830
box -12 -8 72 272
use OAI21X1  _1340_
timestamp 1726538409
transform -1 0 4690 0 -1 1830
box -12 -8 112 272
use OAI21X1  _1341_
timestamp 1726538409
transform -1 0 4630 0 1 1310
box -12 -8 112 272
use OAI21X1  _1342_
timestamp 1726538409
transform 1 0 4750 0 1 1830
box -12 -8 112 272
use NOR2X1  _1343_
timestamp 1726536993
transform 1 0 5530 0 1 3910
box -12 -8 92 272
use NAND2X1  _1344_
timestamp 1726535706
transform -1 0 5490 0 1 1310
box -12 -8 92 272
use INVX1  _1345_
timestamp 1726531033
transform -1 0 5370 0 1 1310
box -12 -8 72 272
use NOR2X1  _1346_
timestamp 1726536993
transform 1 0 5190 0 1 1310
box -12 -8 92 272
use INVX1  _1347_
timestamp 1726531033
transform -1 0 5150 0 1 1310
box -12 -8 72 272
use XOR2X1  _1348_
timestamp 1726561008
transform 1 0 4790 0 1 1310
box -12 -8 152 272
use NAND2X1  _1349_
timestamp 1726535706
transform -1 0 5310 0 1 790
box -12 -8 92 272
use OAI21X1  _1350_
timestamp 1726538409
transform 1 0 5090 0 1 790
box -12 -8 112 272
use NAND2X1  _1351_
timestamp 1726535706
transform 1 0 4750 0 -1 790
box -12 -8 92 272
use NOR2X1  _1352_
timestamp 1726536993
transform -1 0 4910 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1353_
timestamp 1726538409
transform 1 0 5390 0 1 1830
box -12 -8 112 272
use AOI21X1  _1354_
timestamp 1726549551
transform 1 0 4950 0 -1 1830
box -12 -8 112 272
use NOR2X1  _1355_
timestamp 1726536993
transform 1 0 5070 0 -1 2350
box -12 -8 92 272
use NOR2X1  _1356_
timestamp 1726536993
transform 1 0 4950 0 -1 2350
box -12 -8 92 272
use NOR2X1  _1357_
timestamp 1726536993
transform 1 0 5190 0 -1 2350
box -12 -8 92 272
use INVX1  _1358_
timestamp 1726531033
transform 1 0 5350 0 -1 1830
box -12 -8 72 272
use AND2X2  _1359_
timestamp 1726549440
transform 1 0 5070 0 -1 1310
box -12 -8 112 273
use OAI21X1  _1360_
timestamp 1726538409
transform -1 0 5030 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1361_
timestamp 1726538409
transform -1 0 4890 0 -1 1310
box -12 -8 112 272
use NOR2X1  _1362_
timestamp 1726536993
transform 1 0 5090 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1363_
timestamp 1726536993
transform -1 0 4970 0 1 1830
box -12 -8 92 272
use NOR2X1  _1364_
timestamp 1726536993
transform 1 0 5310 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1365_
timestamp 1726535706
transform 1 0 5650 0 -1 2350
box -12 -8 92 272
use INVX1  _1366_
timestamp 1726531033
transform -1 0 5490 0 -1 2350
box -12 -8 72 272
use NOR2X1  _1367_
timestamp 1726536993
transform -1 0 5230 0 1 1830
box -12 -8 92 272
use XOR2X1  _1368_
timestamp 1726561008
transform -1 0 4610 0 1 1830
box -12 -8 152 272
use NAND2X1  _1369_
timestamp 1726535706
transform -1 0 3690 0 1 1830
box -12 -8 92 272
use OAI21X1  _1370_
timestamp 1726538409
transform -1 0 4070 0 1 1830
box -12 -8 112 272
use NAND2X1  _1371_
timestamp 1726535706
transform -1 0 5610 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1372_
timestamp 1726549551
transform 1 0 5010 0 1 1830
box -12 -8 112 272
use NAND2X1  _1373_
timestamp 1726535706
transform 1 0 5270 0 1 1830
box -12 -8 92 272
use OAI21X1  _1374_
timestamp 1726538409
transform -1 0 5310 0 -1 1830
box -12 -8 112 272
use NAND2X1  _1375_
timestamp 1726535706
transform -1 0 4190 0 1 270
box -12 -8 92 272
use NOR2X1  _1376_
timestamp 1726536993
transform -1 0 4310 0 1 270
box -12 -8 92 272
use INVX1  _1377_
timestamp 1726531033
transform 1 0 4850 0 1 270
box -12 -8 72 272
use AND2X2  _1378_
timestamp 1726549440
transform 1 0 4950 0 1 270
box -12 -8 112 273
use NOR2X1  _1379_
timestamp 1726536993
transform 1 0 5630 0 1 270
box -12 -8 92 272
use INVX1  _1380_
timestamp 1726531033
transform -1 0 5250 0 1 270
box -12 -8 72 272
use INVX1  _1381_
timestamp 1726531033
transform 1 0 5090 0 1 270
box -12 -8 72 272
use OAI21X1  _1382_
timestamp 1726538409
transform 1 0 5210 0 -1 790
box -12 -8 112 272
use OAI21X1  _1383_
timestamp 1726538409
transform -1 0 5630 0 1 1310
box -12 -8 112 272
use OAI21X1  _1384_
timestamp 1726538409
transform -1 0 5190 0 -1 270
box -12 -8 112 272
use NOR2X1  _1385_
timestamp 1726536993
transform 1 0 4510 0 -1 270
box -12 -8 92 272
use NOR2X1  _1386_
timestamp 1726536993
transform 1 0 4470 0 1 270
box -12 -8 92 272
use NOR2X1  _1387_
timestamp 1726536993
transform 1 0 4590 0 1 270
box -12 -8 92 272
use INVX1  _1388_
timestamp 1726531033
transform 1 0 4870 0 -1 270
box -12 -8 72 272
use OR2X2  _1389_
timestamp 1726542447
transform 1 0 5230 0 -1 270
box -12 -8 112 272
use AOI21X1  _1390_
timestamp 1726549551
transform 1 0 5370 0 -1 270
box -12 -8 112 272
use AOI22X1  _1391_
timestamp 1726480912
transform 1 0 5510 0 -1 270
box -14 -8 132 272
use AOI21X1  _1392_
timestamp 1726549551
transform -1 0 4810 0 1 270
box -12 -8 112 272
use INVX1  _1393_
timestamp 1726531033
transform -1 0 4690 0 -1 270
box -12 -8 72 272
use NOR2X1  _1394_
timestamp 1726536993
transform 1 0 4970 0 -1 270
box -12 -8 92 272
use AOI21X1  _1395_
timestamp 1726549551
transform -1 0 4830 0 -1 270
box -12 -8 112 272
use INVX1  _1396_
timestamp 1726531033
transform -1 0 2770 0 -1 270
box -12 -8 72 272
use NOR2X1  _1397_
timestamp 1726536993
transform 1 0 2890 0 1 270
box -12 -8 92 272
use OAI21X1  _1398_
timestamp 1726538409
transform 1 0 2810 0 -1 270
box -12 -8 112 272
use OAI22X1  _1399_
timestamp 1726541006
transform -1 0 3130 0 1 270
box -12 -8 132 272
use NAND2X1  _1400_
timestamp 1726535706
transform -1 0 2950 0 1 790
box -12 -8 92 272
use NAND3X1  _1401_
timestamp 1726536591
transform 1 0 2530 0 1 270
box -12 -8 112 272
use OAI21X1  _1402_
timestamp 1726538409
transform -1 0 2670 0 -1 270
box -12 -8 112 272
use NAND2X1  _1403_
timestamp 1726535706
transform 1 0 2670 0 1 270
box -12 -8 92 272
use OAI21X1  _1404_
timestamp 1726538409
transform 1 0 2870 0 -1 790
box -12 -8 112 272
use INVX1  _1405_
timestamp 1726531033
transform 1 0 2370 0 -1 270
box -12 -8 72 272
use NAND3X1  _1406_
timestamp 1726536591
transform 1 0 3610 0 -1 790
box -12 -8 112 272
use NAND2X1  _1407_
timestamp 1726535706
transform -1 0 3710 0 1 270
box -12 -8 92 272
use OAI21X1  _1408_
timestamp 1726538409
transform 1 0 3490 0 1 270
box -12 -8 112 272
use INVX1  _1409_
timestamp 1726531033
transform -1 0 2530 0 -1 270
box -12 -8 72 272
use NAND2X1  _1410_
timestamp 1726535706
transform -1 0 3370 0 -1 270
box -12 -8 92 272
use OAI21X1  _1411_
timestamp 1726538409
transform -1 0 3510 0 -1 270
box -12 -8 112 272
use INVX1  _1412_
timestamp 1726531033
transform -1 0 3450 0 1 270
box -12 -8 72 272
use NAND2X1  _1413_
timestamp 1726535706
transform 1 0 1910 0 1 270
box -12 -8 92 272
use OAI21X1  _1414_
timestamp 1726538409
transform 1 0 1770 0 1 270
box -12 -8 112 272
use INVX1  _1415_
timestamp 1726531033
transform -1 0 3250 0 -1 270
box -12 -8 72 272
use NAND2X1  _1416_
timestamp 1726535706
transform 1 0 1650 0 -1 270
box -12 -8 92 272
use OAI21X1  _1417_
timestamp 1726538409
transform -1 0 1610 0 -1 270
box -12 -8 112 272
use NOR2X1  _1418_
timestamp 1726536993
transform 1 0 4130 0 1 790
box -12 -8 92 272
use NOR2X1  _1419_
timestamp 1726536993
transform -1 0 3630 0 1 1310
box -12 -8 92 272
use AOI21X1  _1420_
timestamp 1726549551
transform 1 0 3410 0 1 1310
box -12 -8 112 272
use NOR2X1  _1421_
timestamp 1726536993
transform -1 0 4390 0 -1 1310
box -12 -8 92 272
use AOI21X1  _1422_
timestamp 1726549551
transform 1 0 4170 0 -1 1310
box -12 -8 112 272
use NOR2X1  _1423_
timestamp 1726536993
transform 1 0 4050 0 1 1310
box -12 -8 92 272
use AOI21X1  _1424_
timestamp 1726549551
transform 1 0 3670 0 1 1310
box -12 -8 112 272
use NOR2X1  _1425_
timestamp 1726536993
transform 1 0 3690 0 -1 1310
box -12 -8 92 272
use AOI21X1  _1426_
timestamp 1726549551
transform 1 0 3310 0 -1 1310
box -12 -8 112 272
use INVX1  _1427_
timestamp 1726531033
transform -1 0 2570 0 -1 790
box -12 -8 72 272
use OAI21X1  _1428_
timestamp 1726538409
transform -1 0 2090 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1429_
timestamp 1726538409
transform -1 0 2230 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1430_
timestamp 1726538409
transform -1 0 2750 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1431_
timestamp 1726538409
transform 1 0 2510 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1432_
timestamp 1726538409
transform -1 0 2470 0 -1 790
box -12 -8 112 272
use OAI21X1  _1433_
timestamp 1726538409
transform 1 0 2230 0 -1 790
box -12 -8 112 272
use OAI21X1  _1434_
timestamp 1726538409
transform 1 0 1450 0 1 790
box -12 -8 112 272
use OAI21X1  _1435_
timestamp 1726538409
transform -1 0 1690 0 1 790
box -12 -8 112 272
use NOR2X1  _1436_
timestamp 1726536993
transform -1 0 2750 0 1 1310
box -12 -8 92 272
use AOI21X1  _1437_
timestamp 1726549551
transform 1 0 2790 0 1 1310
box -12 -8 112 272
use NOR2X1  _1438_
timestamp 1726536993
transform -1 0 1470 0 -1 270
box -12 -8 92 272
use AOI21X1  _1439_
timestamp 1726549551
transform -1 0 1490 0 1 270
box -12 -8 112 272
use NOR2X1  _1440_
timestamp 1726536993
transform -1 0 970 0 1 270
box -12 -8 92 272
use AOI21X1  _1441_
timestamp 1726549551
transform -1 0 1110 0 1 270
box -12 -8 112 272
use NOR2X1  _1442_
timestamp 1726536993
transform -1 0 970 0 -1 270
box -12 -8 92 272
use AOI21X1  _1443_
timestamp 1726549551
transform -1 0 1110 0 -1 270
box -12 -8 112 272
use NAND2X1  _1444_
timestamp 1726535706
transform 1 0 2750 0 1 2870
box -12 -8 92 272
use OAI21X1  _1445_
timestamp 1726538409
transform 1 0 2690 0 -1 2870
box -12 -8 112 272
use NAND2X1  _1446_
timestamp 1726535706
transform 1 0 2270 0 1 2870
box -12 -8 92 272
use OAI21X1  _1447_
timestamp 1726538409
transform 1 0 2130 0 1 2870
box -12 -8 112 272
use NAND2X1  _1448_
timestamp 1726535706
transform 1 0 2870 0 1 3390
box -12 -8 92 272
use OAI21X1  _1449_
timestamp 1726538409
transform 1 0 2730 0 1 3390
box -12 -8 112 272
use NAND2X1  _1450_
timestamp 1726535706
transform -1 0 3330 0 1 3390
box -12 -8 92 272
use OAI21X1  _1451_
timestamp 1726538409
transform 1 0 3370 0 1 3390
box -12 -8 112 272
use DFFPOSX1  _1452_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726550864
transform 1 0 3090 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1453_
timestamp 1726550864
transform 1 0 2890 0 -1 3910
box -13 -8 253 272
use DFFPOSX1  _1454_
timestamp 1726550864
transform 1 0 4090 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1455_
timestamp 1726550864
transform 1 0 3730 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1456_
timestamp 1726550864
transform -1 0 3170 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1457_
timestamp 1726550864
transform -1 0 350 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1458_
timestamp 1726550864
transform -1 0 350 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1459_
timestamp 1726550864
transform -1 0 350 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1460_
timestamp 1726550864
transform 1 0 1010 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1461_
timestamp 1726550864
transform -1 0 3170 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1462_
timestamp 1726550864
transform -1 0 1590 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1463_
timestamp 1726550864
transform 1 0 850 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1464_
timestamp 1726550864
transform 1 0 4030 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1465_
timestamp 1726550864
transform 1 0 5310 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1466_
timestamp 1726550864
transform 1 0 4430 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1467_
timestamp 1726550864
transform 1 0 4190 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1468_
timestamp 1726550864
transform -1 0 5170 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1469_
timestamp 1726550864
transform 1 0 4010 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1470_
timestamp 1726550864
transform 1 0 2250 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1471_
timestamp 1726550864
transform 1 0 1990 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1472_
timestamp 1726550864
transform 1 0 2310 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1473_
timestamp 1726550864
transform 1 0 250 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1474_
timestamp 1726550864
transform -1 0 250 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1475_
timestamp 1726550864
transform -1 0 250 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1476_
timestamp 1726550864
transform 1 0 290 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1477_
timestamp 1726550864
transform -1 0 3630 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1478_
timestamp 1726550864
transform 1 0 1330 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1479_
timestamp 1726550864
transform 1 0 530 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1480_
timestamp 1726550864
transform -1 0 4490 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1481_
timestamp 1726550864
transform 1 0 5410 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1482_
timestamp 1726550864
transform 1 0 4670 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1483_
timestamp 1726550864
transform 1 0 5150 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1484_
timestamp 1726550864
transform 1 0 3630 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1485_
timestamp 1726550864
transform 1 0 4190 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1486_
timestamp 1726550864
transform 1 0 3190 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1487_
timestamp 1726550864
transform 1 0 1590 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1488_
timestamp 1726550864
transform 1 0 970 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1489_
timestamp 1726550864
transform 1 0 1050 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1490_
timestamp 1726550864
transform -1 0 3790 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1491_
timestamp 1726550864
transform 1 0 2150 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1492_
timestamp 1726550864
transform 1 0 2230 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1493_
timestamp 1726550864
transform 1 0 1830 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1494_
timestamp 1726550864
transform -1 0 4630 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1495_
timestamp 1726550864
transform -1 0 5670 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1496_
timestamp 1726550864
transform -1 0 4930 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1497_
timestamp 1726550864
transform -1 0 3930 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1498_
timestamp 1726550864
transform -1 0 5690 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1499_
timestamp 1726550864
transform 1 0 5250 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1500_
timestamp 1726550864
transform 1 0 2910 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1501_
timestamp 1726550864
transform 1 0 3090 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1502_
timestamp 1726550864
transform 1 0 3710 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1503_
timestamp 1726550864
transform -1 0 3750 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1504_
timestamp 1726550864
transform -1 0 1730 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1505_
timestamp 1726550864
transform 1 0 1110 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1506_
timestamp 1726550864
transform 1 0 3590 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1507_
timestamp 1726550864
transform 1 0 4130 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1508_
timestamp 1726550864
transform 1 0 3770 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1509_
timestamp 1726550864
transform 1 0 3410 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1510_
timestamp 1726550864
transform -1 0 1710 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1511_
timestamp 1726550864
transform 1 0 2390 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1512_
timestamp 1726550864
transform -1 0 2190 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1513_
timestamp 1726550864
transform -1 0 1710 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1514_
timestamp 1726550864
transform -1 0 3130 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1515_
timestamp 1726550864
transform 1 0 1110 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1516_
timestamp 1726550864
transform -1 0 850 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1517_
timestamp 1726550864
transform -1 0 850 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1518_
timestamp 1726550864
transform 1 0 2790 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1519_
timestamp 1726550864
transform 1 0 2350 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1520_
timestamp 1726550864
transform 1 0 2950 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1521_
timestamp 1726550864
transform -1 0 3250 0 -1 3390
box -13 -8 253 272
use DFFPOSX1  _1522_
timestamp 1726550864
transform 1 0 290 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1523_
timestamp 1726550864
transform 1 0 2590 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1524_
timestamp 1726550864
transform 1 0 2950 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1525_
timestamp 1726550864
transform 1 0 3330 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1526_
timestamp 1726550864
transform 1 0 3450 0 1 790
box -13 -8 253 272
use BUFX2  _1527_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726549730
transform 1 0 5570 0 -1 2870
box -12 -8 92 272
use BUFX2  _1528_
timestamp 1726549730
transform 1 0 5410 0 1 2870
box -12 -8 92 272
use BUFX2  _1529_
timestamp 1726549730
transform 1 0 5450 0 -1 3910
box -12 -8 92 272
use BUFX2  _1530_
timestamp 1726549730
transform 1 0 5650 0 1 3910
box -12 -8 92 272
use BUFX2  _1531_
timestamp 1726549730
transform 1 0 5410 0 1 3910
box -12 -8 92 272
use BUFX2  _1532_
timestamp 1726549730
transform 1 0 4090 0 -1 790
box -12 -8 92 272
use BUFX2  _1533_
timestamp 1726549730
transform 1 0 4290 0 -1 270
box -12 -8 92 272
use BUFX2  _1534_
timestamp 1726549730
transform 1 0 4350 0 1 270
box -12 -8 92 272
use BUFX2  _1535_
timestamp 1726549730
transform 1 0 4210 0 -1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert0
timestamp 1726549730
transform 1 0 1750 0 -1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert1
timestamp 1726549730
transform -1 0 2730 0 1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert2
timestamp 1726549730
transform -1 0 1330 0 -1 1310
box -12 -8 92 272
use BUFX2  BUFX2_insert3
timestamp 1726549730
transform -1 0 3350 0 1 270
box -12 -8 92 272
use BUFX2  BUFX2_insert4
timestamp 1726549730
transform 1 0 3810 0 -1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert5
timestamp 1726549730
transform 1 0 3970 0 -1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert6
timestamp 1726549730
transform -1 0 3290 0 -1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert15
timestamp 1726549730
transform -1 0 1490 0 -1 5470
box -12 -8 92 272
use BUFX2  BUFX2_insert16
timestamp 1726549730
transform 1 0 1770 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert17
timestamp 1726549730
transform -1 0 1030 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert18
timestamp 1726549730
transform -1 0 2970 0 -1 5470
box -12 -8 92 272
use BUFX2  BUFX2_insert19
timestamp 1726549730
transform 1 0 4970 0 1 1310
box -12 -8 92 272
use BUFX2  BUFX2_insert20
timestamp 1726549730
transform -1 0 2590 0 1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert21
timestamp 1726549730
transform 1 0 2850 0 -1 1830
box -12 -8 92 272
use BUFX2  BUFX2_insert22
timestamp 1726549730
transform 1 0 4970 0 1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert23
timestamp 1726549730
transform -1 0 4190 0 1 1830
box -12 -8 92 272
use BUFX2  BUFX2_insert24
timestamp 1726549730
transform -1 0 2210 0 1 1830
box -12 -8 92 272
use BUFX2  BUFX2_insert25
timestamp 1726549730
transform -1 0 2470 0 1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert26
timestamp 1726549730
transform -1 0 2090 0 1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert27
timestamp 1726549730
transform 1 0 830 0 1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert28
timestamp 1726549730
transform 1 0 2630 0 1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert29
timestamp 1726549730
transform 1 0 2610 0 -1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert30
timestamp 1726549730
transform 1 0 1150 0 -1 4950
box -12 -8 92 272
use BUFX2  BUFX2_insert31
timestamp 1726549730
transform -1 0 2410 0 -1 5470
box -12 -8 92 272
use BUFX2  BUFX2_insert32
timestamp 1726549730
transform 1 0 3310 0 -1 4950
box -12 -8 92 272
use BUFX2  BUFX2_insert33
timestamp 1726549730
transform -1 0 1070 0 -1 5470
box -12 -8 92 272
use CLKBUF1  CLKBUF1_insert7 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726549955
transform 1 0 3810 0 -1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert8
timestamp 1726549955
transform 1 0 3070 0 -1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert9
timestamp 1726549955
transform 1 0 3170 0 1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert10
timestamp 1726549955
transform -1 0 3390 0 -1 2870
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert11
timestamp 1726549955
transform 1 0 3370 0 1 1830
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert12
timestamp 1726549955
transform -1 0 1210 0 -1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert13
timestamp 1726549955
transform 1 0 3430 0 -1 2870
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert14
timestamp 1726549955
transform -1 0 990 0 -1 1830
box -12 -8 212 272
use FILL  FILL84150x78150 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1700315010
transform -1 0 5630 0 -1 5470
box -12 -8 32 272
use FILL  FILL84450x150
timestamp 1700315010
transform -1 0 5650 0 -1 270
box -12 -8 32 272
use FILL  FILL84450x19650
timestamp 1700315010
transform 1 0 5630 0 1 1310
box -12 -8 32 272
use FILL  FILL84450x27450
timestamp 1700315010
transform 1 0 5630 0 1 1830
box -12 -8 32 272
use FILL  FILL84450x35250
timestamp 1700315010
transform 1 0 5630 0 1 2350
box -12 -8 32 272
use FILL  FILL84450x46950
timestamp 1700315010
transform -1 0 5650 0 -1 3390
box -12 -8 32 272
use FILL  FILL84450x78150
timestamp 1700315010
transform -1 0 5650 0 -1 5470
box -12 -8 32 272
use FILL  FILL84750x150
timestamp 1700315010
transform -1 0 5670 0 -1 270
box -12 -8 32 272
use FILL  FILL84750x15750
timestamp 1700315010
transform -1 0 5670 0 -1 1310
box -12 -8 32 272
use FILL  FILL84750x19650
timestamp 1700315010
transform 1 0 5650 0 1 1310
box -12 -8 32 272
use FILL  FILL84750x23550
timestamp 1700315010
transform -1 0 5670 0 -1 1830
box -12 -8 32 272
use FILL  FILL84750x27450
timestamp 1700315010
transform 1 0 5650 0 1 1830
box -12 -8 32 272
use FILL  FILL84750x35250
timestamp 1700315010
transform 1 0 5650 0 1 2350
box -12 -8 32 272
use FILL  FILL84750x39150
timestamp 1700315010
transform -1 0 5670 0 -1 2870
box -12 -8 32 272
use FILL  FILL84750x46950
timestamp 1700315010
transform -1 0 5670 0 -1 3390
box -12 -8 32 272
use FILL  FILL84750x66450
timestamp 1700315010
transform 1 0 5650 0 1 4430
box -12 -8 32 272
use FILL  FILL84750x78150
timestamp 1700315010
transform -1 0 5670 0 -1 5470
box -12 -8 32 272
use FILL  FILL85050x150
timestamp 1700315010
transform -1 0 5690 0 -1 270
box -12 -8 32 272
use FILL  FILL85050x7950
timestamp 1700315010
transform -1 0 5690 0 -1 790
box -12 -8 32 272
use FILL  FILL85050x15750
timestamp 1700315010
transform -1 0 5690 0 -1 1310
box -12 -8 32 272
use FILL  FILL85050x19650
timestamp 1700315010
transform 1 0 5670 0 1 1310
box -12 -8 32 272
use FILL  FILL85050x23550
timestamp 1700315010
transform -1 0 5690 0 -1 1830
box -12 -8 32 272
use FILL  FILL85050x27450
timestamp 1700315010
transform 1 0 5670 0 1 1830
box -12 -8 32 272
use FILL  FILL85050x35250
timestamp 1700315010
transform 1 0 5670 0 1 2350
box -12 -8 32 272
use FILL  FILL85050x39150
timestamp 1700315010
transform -1 0 5690 0 -1 2870
box -12 -8 32 272
use FILL  FILL85050x43050
timestamp 1700315010
transform 1 0 5670 0 1 2870
box -12 -8 32 272
use FILL  FILL85050x46950
timestamp 1700315010
transform -1 0 5690 0 -1 3390
box -12 -8 32 272
use FILL  FILL85050x54750
timestamp 1700315010
transform -1 0 5690 0 -1 3910
box -12 -8 32 272
use FILL  FILL85050x66450
timestamp 1700315010
transform 1 0 5670 0 1 4430
box -12 -8 32 272
use FILL  FILL85050x78150
timestamp 1700315010
transform -1 0 5690 0 -1 5470
box -12 -8 32 272
use FILL  FILL85350x150
timestamp 1700315010
transform -1 0 5710 0 -1 270
box -12 -8 32 272
use FILL  FILL85350x7950
timestamp 1700315010
transform -1 0 5710 0 -1 790
box -12 -8 32 272
use FILL  FILL85350x11850
timestamp 1700315010
transform 1 0 5690 0 1 790
box -12 -8 32 272
use FILL  FILL85350x15750
timestamp 1700315010
transform -1 0 5710 0 -1 1310
box -12 -8 32 272
use FILL  FILL85350x19650
timestamp 1700315010
transform 1 0 5690 0 1 1310
box -12 -8 32 272
use FILL  FILL85350x23550
timestamp 1700315010
transform -1 0 5710 0 -1 1830
box -12 -8 32 272
use FILL  FILL85350x27450
timestamp 1700315010
transform 1 0 5690 0 1 1830
box -12 -8 32 272
use FILL  FILL85350x35250
timestamp 1700315010
transform 1 0 5690 0 1 2350
box -12 -8 32 272
use FILL  FILL85350x39150
timestamp 1700315010
transform -1 0 5710 0 -1 2870
box -12 -8 32 272
use FILL  FILL85350x43050
timestamp 1700315010
transform 1 0 5690 0 1 2870
box -12 -8 32 272
use FILL  FILL85350x46950
timestamp 1700315010
transform -1 0 5710 0 -1 3390
box -12 -8 32 272
use FILL  FILL85350x54750
timestamp 1700315010
transform -1 0 5710 0 -1 3910
box -12 -8 32 272
use FILL  FILL85350x62550
timestamp 1700315010
transform -1 0 5710 0 -1 4430
box -12 -8 32 272
use FILL  FILL85350x66450
timestamp 1700315010
transform 1 0 5690 0 1 4430
box -12 -8 32 272
use FILL  FILL85350x78150
timestamp 1700315010
transform -1 0 5710 0 -1 5470
box -12 -8 32 272
use FILL  FILL85650x150
timestamp 1700315010
transform -1 0 5730 0 -1 270
box -12 -8 32 272
use FILL  FILL85650x4050
timestamp 1700315010
transform 1 0 5710 0 1 270
box -12 -8 32 272
use FILL  FILL85650x7950
timestamp 1700315010
transform -1 0 5730 0 -1 790
box -12 -8 32 272
use FILL  FILL85650x11850
timestamp 1700315010
transform 1 0 5710 0 1 790
box -12 -8 32 272
use FILL  FILL85650x15750
timestamp 1700315010
transform -1 0 5730 0 -1 1310
box -12 -8 32 272
use FILL  FILL85650x19650
timestamp 1700315010
transform 1 0 5710 0 1 1310
box -12 -8 32 272
use FILL  FILL85650x23550
timestamp 1700315010
transform -1 0 5730 0 -1 1830
box -12 -8 32 272
use FILL  FILL85650x27450
timestamp 1700315010
transform 1 0 5710 0 1 1830
box -12 -8 32 272
use FILL  FILL85650x35250
timestamp 1700315010
transform 1 0 5710 0 1 2350
box -12 -8 32 272
use FILL  FILL85650x39150
timestamp 1700315010
transform -1 0 5730 0 -1 2870
box -12 -8 32 272
use FILL  FILL85650x43050
timestamp 1700315010
transform 1 0 5710 0 1 2870
box -12 -8 32 272
use FILL  FILL85650x46950
timestamp 1700315010
transform -1 0 5730 0 -1 3390
box -12 -8 32 272
use FILL  FILL85650x50850
timestamp 1700315010
transform 1 0 5710 0 1 3390
box -12 -8 32 272
use FILL  FILL85650x54750
timestamp 1700315010
transform -1 0 5730 0 -1 3910
box -12 -8 32 272
use FILL  FILL85650x62550
timestamp 1700315010
transform -1 0 5730 0 -1 4430
box -12 -8 32 272
use FILL  FILL85650x66450
timestamp 1700315010
transform 1 0 5710 0 1 4430
box -12 -8 32 272
use FILL  FILL85650x78150
timestamp 1700315010
transform -1 0 5730 0 -1 5470
box -12 -8 32 272
use FILL  FILL85950x150
timestamp 1700315010
transform -1 0 5750 0 -1 270
box -12 -8 32 272
use FILL  FILL85950x4050
timestamp 1700315010
transform 1 0 5730 0 1 270
box -12 -8 32 272
use FILL  FILL85950x7950
timestamp 1700315010
transform -1 0 5750 0 -1 790
box -12 -8 32 272
use FILL  FILL85950x11850
timestamp 1700315010
transform 1 0 5730 0 1 790
box -12 -8 32 272
use FILL  FILL85950x15750
timestamp 1700315010
transform -1 0 5750 0 -1 1310
box -12 -8 32 272
use FILL  FILL85950x19650
timestamp 1700315010
transform 1 0 5730 0 1 1310
box -12 -8 32 272
use FILL  FILL85950x23550
timestamp 1700315010
transform -1 0 5750 0 -1 1830
box -12 -8 32 272
use FILL  FILL85950x27450
timestamp 1700315010
transform 1 0 5730 0 1 1830
box -12 -8 32 272
use FILL  FILL85950x31350
timestamp 1700315010
transform -1 0 5750 0 -1 2350
box -12 -8 32 272
use FILL  FILL85950x35250
timestamp 1700315010
transform 1 0 5730 0 1 2350
box -12 -8 32 272
use FILL  FILL85950x39150
timestamp 1700315010
transform -1 0 5750 0 -1 2870
box -12 -8 32 272
use FILL  FILL85950x43050
timestamp 1700315010
transform 1 0 5730 0 1 2870
box -12 -8 32 272
use FILL  FILL85950x46950
timestamp 1700315010
transform -1 0 5750 0 -1 3390
box -12 -8 32 272
use FILL  FILL85950x50850
timestamp 1700315010
transform 1 0 5730 0 1 3390
box -12 -8 32 272
use FILL  FILL85950x54750
timestamp 1700315010
transform -1 0 5750 0 -1 3910
box -12 -8 32 272
use FILL  FILL85950x58650
timestamp 1700315010
transform 1 0 5730 0 1 3910
box -12 -8 32 272
use FILL  FILL85950x62550
timestamp 1700315010
transform -1 0 5750 0 -1 4430
box -12 -8 32 272
use FILL  FILL85950x66450
timestamp 1700315010
transform 1 0 5730 0 1 4430
box -12 -8 32 272
use FILL  FILL85950x74250
timestamp 1700315010
transform 1 0 5730 0 1 4950
box -12 -8 32 272
use FILL  FILL85950x78150
timestamp 1700315010
transform -1 0 5750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__723_
timestamp 1700315010
transform 1 0 3830 0 1 790
box -12 -8 32 272
use FILL  FILL_0__724_
timestamp 1700315010
transform 1 0 3710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__725_
timestamp 1700315010
transform -1 0 2990 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__726_
timestamp 1700315010
transform 1 0 4350 0 1 790
box -12 -8 32 272
use FILL  FILL_0__727_
timestamp 1700315010
transform -1 0 2750 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__728_
timestamp 1700315010
transform 1 0 2750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__729_
timestamp 1700315010
transform 1 0 3430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__730_
timestamp 1700315010
transform 1 0 3950 0 1 790
box -12 -8 32 272
use FILL  FILL_0__731_
timestamp 1700315010
transform 1 0 4490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__732_
timestamp 1700315010
transform 1 0 5490 0 1 270
box -12 -8 32 272
use FILL  FILL_0__733_
timestamp 1700315010
transform 1 0 5310 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__734_
timestamp 1700315010
transform 1 0 5310 0 1 790
box -12 -8 32 272
use FILL  FILL_0__735_
timestamp 1700315010
transform 1 0 2870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__736_
timestamp 1700315010
transform -1 0 4230 0 1 790
box -12 -8 32 272
use FILL  FILL_0__737_
timestamp 1700315010
transform 1 0 3130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__738_
timestamp 1700315010
transform 1 0 3810 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__739_
timestamp 1700315010
transform -1 0 4450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__740_
timestamp 1700315010
transform 1 0 2570 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__741_
timestamp 1700315010
transform -1 0 4310 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__742_
timestamp 1700315010
transform -1 0 3210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__743_
timestamp 1700315010
transform 1 0 3690 0 1 790
box -12 -8 32 272
use FILL  FILL_0__744_
timestamp 1700315010
transform 1 0 2190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__745_
timestamp 1700315010
transform 1 0 3310 0 1 790
box -12 -8 32 272
use FILL  FILL_0__746_
timestamp 1700315010
transform -1 0 3490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__747_
timestamp 1700315010
transform -1 0 3050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__748_
timestamp 1700315010
transform -1 0 3350 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__749_
timestamp 1700315010
transform 1 0 3670 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__750_
timestamp 1700315010
transform -1 0 3150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__751_
timestamp 1700315010
transform -1 0 3270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__752_
timestamp 1700315010
transform 1 0 2770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__753_
timestamp 1700315010
transform -1 0 3130 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__754_
timestamp 1700315010
transform -1 0 3370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__755_
timestamp 1700315010
transform 1 0 3770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__756_
timestamp 1700315010
transform -1 0 3250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__757_
timestamp 1700315010
transform 1 0 3490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__758_
timestamp 1700315010
transform 1 0 2830 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__759_
timestamp 1700315010
transform -1 0 2970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__760_
timestamp 1700315010
transform 1 0 2570 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__761_
timestamp 1700315010
transform -1 0 2770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__762_
timestamp 1700315010
transform 1 0 3470 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__763_
timestamp 1700315010
transform -1 0 3610 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__764_
timestamp 1700315010
transform 1 0 3250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__765_
timestamp 1700315010
transform -1 0 3390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__766_
timestamp 1700315010
transform -1 0 2850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__767_
timestamp 1700315010
transform 1 0 2690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__768_
timestamp 1700315010
transform -1 0 2710 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__769_
timestamp 1700315010
transform 1 0 470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__770_
timestamp 1700315010
transform 1 0 730 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__771_
timestamp 1700315010
transform 1 0 570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__772_
timestamp 1700315010
transform -1 0 30 0 1 270
box -12 -8 32 272
use FILL  FILL_0__773_
timestamp 1700315010
transform 1 0 490 0 1 270
box -12 -8 32 272
use FILL  FILL_0__774_
timestamp 1700315010
transform 1 0 350 0 1 270
box -12 -8 32 272
use FILL  FILL_0__775_
timestamp 1700315010
transform -1 0 30 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__776_
timestamp 1700315010
transform 1 0 490 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__777_
timestamp 1700315010
transform 1 0 350 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__778_
timestamp 1700315010
transform 1 0 1230 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__779_
timestamp 1700315010
transform -1 0 1410 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__780_
timestamp 1700315010
transform 1 0 1250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__781_
timestamp 1700315010
transform -1 0 2850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__782_
timestamp 1700315010
transform -1 0 2590 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__783_
timestamp 1700315010
transform -1 0 2710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__784_
timestamp 1700315010
transform 1 0 1590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__785_
timestamp 1700315010
transform 1 0 1830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__786_
timestamp 1700315010
transform -1 0 1850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__787_
timestamp 1700315010
transform -1 0 630 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__788_
timestamp 1700315010
transform 1 0 850 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__789_
timestamp 1700315010
transform 1 0 710 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__790_
timestamp 1700315010
transform -1 0 3950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__791_
timestamp 1700315010
transform -1 0 3850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__792_
timestamp 1700315010
transform 1 0 3790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__793_
timestamp 1700315010
transform 1 0 5550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__794_
timestamp 1700315010
transform -1 0 4650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__795_
timestamp 1700315010
transform -1 0 5190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__796_
timestamp 1700315010
transform -1 0 4830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__797_
timestamp 1700315010
transform -1 0 4650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__798_
timestamp 1700315010
transform -1 0 4690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__799_
timestamp 1700315010
transform -1 0 4110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__800_
timestamp 1700315010
transform -1 0 4030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__801_
timestamp 1700315010
transform 1 0 3950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__802_
timestamp 1700315010
transform -1 0 4850 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__803_
timestamp 1700315010
transform 1 0 3950 0 1 270
box -12 -8 32 272
use FILL  FILL_0__804_
timestamp 1700315010
transform -1 0 4590 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__805_
timestamp 1700315010
transform 1 0 4370 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__806_
timestamp 1700315010
transform -1 0 3770 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__807_
timestamp 1700315010
transform -1 0 3890 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__808_
timestamp 1700315010
transform -1 0 2770 0 1 270
box -12 -8 32 272
use FILL  FILL_0__809_
timestamp 1700315010
transform -1 0 2010 0 1 270
box -12 -8 32 272
use FILL  FILL_0__810_
timestamp 1700315010
transform -1 0 2130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__811_
timestamp 1700315010
transform 1 0 2230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__812_
timestamp 1700315010
transform -1 0 1750 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__813_
timestamp 1700315010
transform -1 0 1870 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__814_
timestamp 1700315010
transform 1 0 2550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__815_
timestamp 1700315010
transform 1 0 1930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__816_
timestamp 1700315010
transform -1 0 2190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__817_
timestamp 1700315010
transform 1 0 3170 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__818_
timestamp 1700315010
transform -1 0 1190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__819_
timestamp 1700315010
transform 1 0 1450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__820_
timestamp 1700315010
transform -1 0 950 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__821_
timestamp 1700315010
transform 1 0 490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__822_
timestamp 1700315010
transform -1 0 630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__823_
timestamp 1700315010
transform -1 0 830 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__824_
timestamp 1700315010
transform -1 0 1170 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__825_
timestamp 1700315010
transform 1 0 1130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__826_
timestamp 1700315010
transform 1 0 1050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__827_
timestamp 1700315010
transform 1 0 1290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__828_
timestamp 1700315010
transform 1 0 910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__829_
timestamp 1700315010
transform 1 0 810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__830_
timestamp 1700315010
transform -1 0 1550 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__831_
timestamp 1700315010
transform 1 0 1270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__832_
timestamp 1700315010
transform -1 0 1430 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__833_
timestamp 1700315010
transform 1 0 1830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__834_
timestamp 1700315010
transform -1 0 3410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__835_
timestamp 1700315010
transform -1 0 1590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__836_
timestamp 1700315010
transform -1 0 1710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__837_
timestamp 1700315010
transform -1 0 690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__838_
timestamp 1700315010
transform -1 0 690 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__839_
timestamp 1700315010
transform -1 0 550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__840_
timestamp 1700315010
transform -1 0 550 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__841_
timestamp 1700315010
transform -1 0 410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__842_
timestamp 1700315010
transform 1 0 190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__843_
timestamp 1700315010
transform 1 0 350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__844_
timestamp 1700315010
transform -1 0 270 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__845_
timestamp 1700315010
transform 1 0 10 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__846_
timestamp 1700315010
transform 1 0 1930 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__847_
timestamp 1700315010
transform -1 0 550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__848_
timestamp 1700315010
transform -1 0 1270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__849_
timestamp 1700315010
transform -1 0 650 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__850_
timestamp 1700315010
transform -1 0 650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__851_
timestamp 1700315010
transform -1 0 1110 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__852_
timestamp 1700315010
transform -1 0 510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__853_
timestamp 1700315010
transform -1 0 770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__854_
timestamp 1700315010
transform 1 0 1250 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__855_
timestamp 1700315010
transform 1 0 1390 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__856_
timestamp 1700315010
transform 1 0 850 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__857_
timestamp 1700315010
transform -1 0 730 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__858_
timestamp 1700315010
transform -1 0 450 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__859_
timestamp 1700315010
transform -1 0 730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__860_
timestamp 1700315010
transform -1 0 590 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__861_
timestamp 1700315010
transform -1 0 1770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__862_
timestamp 1700315010
transform -1 0 1670 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__863_
timestamp 1700315010
transform -1 0 2550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__864_
timestamp 1700315010
transform 1 0 930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__865_
timestamp 1700315010
transform -1 0 1810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__866_
timestamp 1700315010
transform -1 0 1530 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__867_
timestamp 1700315010
transform 1 0 570 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__868_
timestamp 1700315010
transform -1 0 170 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__869_
timestamp 1700315010
transform -1 0 130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__870_
timestamp 1700315010
transform -1 0 310 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__871_
timestamp 1700315010
transform -1 0 410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__872_
timestamp 1700315010
transform -1 0 270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__873_
timestamp 1700315010
transform 1 0 250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__874_
timestamp 1700315010
transform -1 0 130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__875_
timestamp 1700315010
transform -1 0 30 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__876_
timestamp 1700315010
transform 1 0 130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__877_
timestamp 1700315010
transform -1 0 930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__878_
timestamp 1700315010
transform -1 0 30 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__879_
timestamp 1700315010
transform -1 0 370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__880_
timestamp 1700315010
transform -1 0 230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__881_
timestamp 1700315010
transform 1 0 950 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__882_
timestamp 1700315010
transform 1 0 910 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__883_
timestamp 1700315010
transform -1 0 1150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__884_
timestamp 1700315010
transform 1 0 750 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__885_
timestamp 1700315010
transform -1 0 30 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__886_
timestamp 1700315010
transform 1 0 1030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__887_
timestamp 1700315010
transform -1 0 30 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__888_
timestamp 1700315010
transform 1 0 430 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__889_
timestamp 1700315010
transform 1 0 430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__890_
timestamp 1700315010
transform 1 0 270 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__891_
timestamp 1700315010
transform 1 0 250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__892_
timestamp 1700315010
transform -1 0 410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__893_
timestamp 1700315010
transform -1 0 450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__894_
timestamp 1700315010
transform -1 0 310 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__895_
timestamp 1700315010
transform -1 0 130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__896_
timestamp 1700315010
transform 1 0 150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__897_
timestamp 1700315010
transform -1 0 2330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__898_
timestamp 1700315010
transform 1 0 2070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__899_
timestamp 1700315010
transform -1 0 3410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__900_
timestamp 1700315010
transform -1 0 2210 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__901_
timestamp 1700315010
transform -1 0 2110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__902_
timestamp 1700315010
transform 1 0 2050 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__903_
timestamp 1700315010
transform -1 0 270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__904_
timestamp 1700315010
transform -1 0 30 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__905_
timestamp 1700315010
transform 1 0 530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__906_
timestamp 1700315010
transform -1 0 30 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__907_
timestamp 1700315010
transform 1 0 150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__908_
timestamp 1700315010
transform 1 0 290 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__909_
timestamp 1700315010
transform -1 0 170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__910_
timestamp 1700315010
transform -1 0 30 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__911_
timestamp 1700315010
transform -1 0 30 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__912_
timestamp 1700315010
transform -1 0 30 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__913_
timestamp 1700315010
transform -1 0 30 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__914_
timestamp 1700315010
transform 1 0 150 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__915_
timestamp 1700315010
transform -1 0 30 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__916_
timestamp 1700315010
transform 1 0 790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__917_
timestamp 1700315010
transform -1 0 650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__918_
timestamp 1700315010
transform -1 0 1870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__919_
timestamp 1700315010
transform -1 0 1250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__920_
timestamp 1700315010
transform 1 0 1250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__921_
timestamp 1700315010
transform 1 0 110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__922_
timestamp 1700315010
transform 1 0 2630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__923_
timestamp 1700315010
transform 1 0 1990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__924_
timestamp 1700315010
transform 1 0 2130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__925_
timestamp 1700315010
transform 1 0 3850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__926_
timestamp 1700315010
transform -1 0 2310 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__927_
timestamp 1700315010
transform -1 0 2170 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__928_
timestamp 1700315010
transform 1 0 2530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__929_
timestamp 1700315010
transform -1 0 2290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__930_
timestamp 1700315010
transform -1 0 2450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__931_
timestamp 1700315010
transform -1 0 2410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__932_
timestamp 1700315010
transform 1 0 810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__933_
timestamp 1700315010
transform -1 0 130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__934_
timestamp 1700315010
transform -1 0 310 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__935_
timestamp 1700315010
transform 1 0 990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__936_
timestamp 1700315010
transform -1 0 570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__937_
timestamp 1700315010
transform 1 0 690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__938_
timestamp 1700315010
transform -1 0 310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__939_
timestamp 1700315010
transform 1 0 150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__940_
timestamp 1700315010
transform 1 0 670 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__941_
timestamp 1700315010
transform 1 0 1070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__942_
timestamp 1700315010
transform 1 0 1050 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__943_
timestamp 1700315010
transform -1 0 870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__944_
timestamp 1700315010
transform -1 0 550 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__945_
timestamp 1700315010
transform -1 0 310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__946_
timestamp 1700315010
transform -1 0 410 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__947_
timestamp 1700315010
transform -1 0 30 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__948_
timestamp 1700315010
transform -1 0 30 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__949_
timestamp 1700315010
transform -1 0 30 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__950_
timestamp 1700315010
transform -1 0 690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__951_
timestamp 1700315010
transform -1 0 450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__952_
timestamp 1700315010
transform 1 0 150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__953_
timestamp 1700315010
transform 1 0 390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__954_
timestamp 1700315010
transform 1 0 570 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__955_
timestamp 1700315010
transform 1 0 670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__956_
timestamp 1700315010
transform 1 0 530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__957_
timestamp 1700315010
transform 1 0 150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__958_
timestamp 1700315010
transform 1 0 850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__959_
timestamp 1700315010
transform -1 0 1010 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__960_
timestamp 1700315010
transform 1 0 810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__961_
timestamp 1700315010
transform -1 0 730 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__962_
timestamp 1700315010
transform -1 0 1110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__963_
timestamp 1700315010
transform 1 0 1010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__964_
timestamp 1700315010
transform -1 0 870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__965_
timestamp 1700315010
transform 1 0 970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__966_
timestamp 1700315010
transform 1 0 3270 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__967_
timestamp 1700315010
transform -1 0 3150 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__968_
timestamp 1700315010
transform 1 0 1770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__969_
timestamp 1700315010
transform -1 0 870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__970_
timestamp 1700315010
transform 1 0 950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__971_
timestamp 1700315010
transform 1 0 1350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__972_
timestamp 1700315010
transform -1 0 1930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__973_
timestamp 1700315010
transform -1 0 2030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__974_
timestamp 1700315010
transform -1 0 1170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__975_
timestamp 1700315010
transform 1 0 390 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__976_
timestamp 1700315010
transform 1 0 490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__977_
timestamp 1700315010
transform 1 0 2710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__978_
timestamp 1700315010
transform -1 0 2850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__979_
timestamp 1700315010
transform -1 0 2590 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__980_
timestamp 1700315010
transform 1 0 1770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__981_
timestamp 1700315010
transform 1 0 2390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__982_
timestamp 1700315010
transform -1 0 2450 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__983_
timestamp 1700315010
transform -1 0 2190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__984_
timestamp 1700315010
transform 1 0 2270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__985_
timestamp 1700315010
transform -1 0 2050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__986_
timestamp 1700315010
transform 1 0 2110 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__987_
timestamp 1700315010
transform -1 0 1870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__988_
timestamp 1700315010
transform 1 0 810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__989_
timestamp 1700315010
transform 1 0 770 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__990_
timestamp 1700315010
transform 1 0 2170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__991_
timestamp 1700315010
transform -1 0 2450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__992_
timestamp 1700315010
transform -1 0 2310 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__993_
timestamp 1700315010
transform 1 0 2690 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__994_
timestamp 1700315010
transform -1 0 2570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__995_
timestamp 1700315010
transform -1 0 2030 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__996_
timestamp 1700315010
transform -1 0 2090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__997_
timestamp 1700315010
transform -1 0 2430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__998_
timestamp 1700315010
transform 1 0 1790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__999_
timestamp 1700315010
transform -1 0 2330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1000_
timestamp 1700315010
transform -1 0 1670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1001_
timestamp 1700315010
transform -1 0 1610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1002_
timestamp 1700315010
transform -1 0 1230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1003_
timestamp 1700315010
transform 1 0 1170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1004_
timestamp 1700315010
transform 1 0 1490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1005_
timestamp 1700315010
transform -1 0 2170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1006_
timestamp 1700315010
transform -1 0 1330 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1007_
timestamp 1700315010
transform -1 0 1390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1008_
timestamp 1700315010
transform -1 0 1990 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1009_
timestamp 1700315010
transform 1 0 1730 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1010_
timestamp 1700315010
transform -1 0 1470 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1011_
timestamp 1700315010
transform -1 0 1670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1012_
timestamp 1700315010
transform -1 0 1050 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1013_
timestamp 1700315010
transform 1 0 570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1014_
timestamp 1700315010
transform -1 0 730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1015_
timestamp 1700315010
transform -1 0 1810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1016_
timestamp 1700315010
transform 1 0 1510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1017_
timestamp 1700315010
transform -1 0 1470 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1018_
timestamp 1700315010
transform -1 0 1270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1019_
timestamp 1700315010
transform 1 0 1170 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1020_
timestamp 1700315010
transform -1 0 1610 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1021_
timestamp 1700315010
transform -1 0 1610 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1022_
timestamp 1700315010
transform 1 0 1630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1023_
timestamp 1700315010
transform -1 0 1390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1024_
timestamp 1700315010
transform -1 0 1850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1025_
timestamp 1700315010
transform -1 0 1510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1026_
timestamp 1700315010
transform 1 0 1490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1027_
timestamp 1700315010
transform 1 0 1350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1028_
timestamp 1700315010
transform 1 0 1870 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1029_
timestamp 1700315010
transform 1 0 1390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1030_
timestamp 1700315010
transform -1 0 1750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1031_
timestamp 1700315010
transform 1 0 1690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1032_
timestamp 1700315010
transform -1 0 1870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1033_
timestamp 1700315010
transform 1 0 1810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1034_
timestamp 1700315010
transform 1 0 1550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1035_
timestamp 1700315010
transform 1 0 1530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1036_
timestamp 1700315010
transform 1 0 1630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1037_
timestamp 1700315010
transform -1 0 2270 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1038_
timestamp 1700315010
transform 1 0 3070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1039_
timestamp 1700315010
transform 1 0 2070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1040_
timestamp 1700315010
transform 1 0 2170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1041_
timestamp 1700315010
transform -1 0 3030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1042_
timestamp 1700315010
transform 1 0 3530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1043_
timestamp 1700315010
transform 1 0 3270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1044_
timestamp 1700315010
transform 1 0 2870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1045_
timestamp 1700315010
transform -1 0 2990 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1046_
timestamp 1700315010
transform -1 0 3150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1047_
timestamp 1700315010
transform 1 0 3310 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1048_
timestamp 1700315010
transform 1 0 3410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1049_
timestamp 1700315010
transform 1 0 3630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1050_
timestamp 1700315010
transform 1 0 3490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1051_
timestamp 1700315010
transform -1 0 3430 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1052_
timestamp 1700315010
transform -1 0 3170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1053_
timestamp 1700315010
transform 1 0 1910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1054_
timestamp 1700315010
transform -1 0 3930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1055_
timestamp 1700315010
transform -1 0 3970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1056_
timestamp 1700315010
transform 1 0 4070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1057_
timestamp 1700315010
transform -1 0 3810 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1058_
timestamp 1700315010
transform -1 0 4050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1059_
timestamp 1700315010
transform 1 0 4550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1060_
timestamp 1700315010
transform -1 0 3670 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1061_
timestamp 1700315010
transform -1 0 4210 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1062_
timestamp 1700315010
transform 1 0 4450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1063_
timestamp 1700315010
transform -1 0 4330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1064_
timestamp 1700315010
transform 1 0 3350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1065_
timestamp 1700315010
transform 1 0 2690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1066_
timestamp 1700315010
transform 1 0 2550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1067_
timestamp 1700315010
transform -1 0 4190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1068_
timestamp 1700315010
transform 1 0 3630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1069_
timestamp 1700315010
transform 1 0 3490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1070_
timestamp 1700315010
transform 1 0 3770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1071_
timestamp 1700315010
transform -1 0 3650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1072_
timestamp 1700315010
transform -1 0 3390 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1073_
timestamp 1700315010
transform -1 0 3030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1074_
timestamp 1700315010
transform -1 0 3230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1075_
timestamp 1700315010
transform -1 0 3790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1076_
timestamp 1700315010
transform -1 0 3110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1077_
timestamp 1700315010
transform 1 0 2810 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1078_
timestamp 1700315010
transform 1 0 1870 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1079_
timestamp 1700315010
transform 1 0 1930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1080_
timestamp 1700315010
transform -1 0 2970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1081_
timestamp 1700315010
transform -1 0 3250 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1082_
timestamp 1700315010
transform 1 0 2590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1083_
timestamp 1700315010
transform -1 0 2810 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1084_
timestamp 1700315010
transform -1 0 2750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1085_
timestamp 1700315010
transform -1 0 2470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1086_
timestamp 1700315010
transform 1 0 2650 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1087_
timestamp 1700315010
transform -1 0 2650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1088_
timestamp 1700315010
transform 1 0 1230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1089_
timestamp 1700315010
transform 1 0 1310 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1090_
timestamp 1700315010
transform -1 0 2530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1091_
timestamp 1700315010
transform 1 0 2930 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1092_
timestamp 1700315010
transform 1 0 2370 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1093_
timestamp 1700315010
transform 1 0 2490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1094_
timestamp 1700315010
transform 1 0 1670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1095_
timestamp 1700315010
transform -1 0 790 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1096_
timestamp 1700315010
transform -1 0 910 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1097_
timestamp 1700315010
transform 1 0 4490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1098_
timestamp 1700315010
transform -1 0 2250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1099_
timestamp 1700315010
transform -1 0 2630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1100_
timestamp 1700315010
transform 1 0 2730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1101_
timestamp 1700315010
transform 1 0 2870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1102_
timestamp 1700315010
transform 1 0 3170 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1103_
timestamp 1700315010
transform 1 0 3550 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1104_
timestamp 1700315010
transform 1 0 5630 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1105_
timestamp 1700315010
transform 1 0 2970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1106_
timestamp 1700315010
transform 1 0 3070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1107_
timestamp 1700315010
transform 1 0 3750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1108_
timestamp 1700315010
transform 1 0 3630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1109_
timestamp 1700315010
transform 1 0 3830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1110_
timestamp 1700315010
transform 1 0 3670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1111_
timestamp 1700315010
transform 1 0 3970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1112_
timestamp 1700315010
transform 1 0 4110 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1113_
timestamp 1700315010
transform 1 0 4650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1114_
timestamp 1700315010
transform -1 0 3930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1115_
timestamp 1700315010
transform -1 0 3890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1116_
timestamp 1700315010
transform -1 0 4010 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1117_
timestamp 1700315010
transform 1 0 4030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1118_
timestamp 1700315010
transform 1 0 4170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1119_
timestamp 1700315010
transform -1 0 4730 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1120_
timestamp 1700315010
transform -1 0 4330 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1121_
timestamp 1700315010
transform -1 0 4330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1122_
timestamp 1700315010
transform 1 0 4450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1123_
timestamp 1700315010
transform 1 0 4910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1124_
timestamp 1700315010
transform 1 0 4430 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1125_
timestamp 1700315010
transform -1 0 4590 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1126_
timestamp 1700315010
transform 1 0 4830 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1127_
timestamp 1700315010
transform 1 0 4950 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1128_
timestamp 1700315010
transform 1 0 5090 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1129_
timestamp 1700315010
transform 1 0 3490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1130_
timestamp 1700315010
transform 1 0 3510 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1131_
timestamp 1700315010
transform 1 0 4930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1132_
timestamp 1700315010
transform 1 0 5070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1133_
timestamp 1700315010
transform 1 0 4790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1134_
timestamp 1700315010
transform 1 0 5190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1135_
timestamp 1700315010
transform -1 0 5350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1136_
timestamp 1700315010
transform 1 0 5490 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1137_
timestamp 1700315010
transform 1 0 5190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1138_
timestamp 1700315010
transform 1 0 5470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1139_
timestamp 1700315010
transform 1 0 5510 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1140_
timestamp 1700315010
transform 1 0 5370 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1141_
timestamp 1700315010
transform -1 0 5290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1142_
timestamp 1700315010
transform -1 0 5490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1143_
timestamp 1700315010
transform -1 0 5250 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1144_
timestamp 1700315010
transform -1 0 5350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1145_
timestamp 1700315010
transform 1 0 5270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1146_
timestamp 1700315010
transform 1 0 4970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1147_
timestamp 1700315010
transform 1 0 4610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1148_
timestamp 1700315010
transform -1 0 5550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1149_
timestamp 1700315010
transform 1 0 5390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1150_
timestamp 1700315010
transform 1 0 4110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1151_
timestamp 1700315010
transform -1 0 4810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1152_
timestamp 1700315010
transform 1 0 4630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1153_
timestamp 1700315010
transform -1 0 4150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1154_
timestamp 1700315010
transform 1 0 3870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1155_
timestamp 1700315010
transform 1 0 4330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1156_
timestamp 1700315010
transform 1 0 4250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1157_
timestamp 1700315010
transform 1 0 3990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1158_
timestamp 1700315010
transform 1 0 4390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1159_
timestamp 1700315010
transform 1 0 4070 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1160_
timestamp 1700315010
transform -1 0 3970 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1161_
timestamp 1700315010
transform -1 0 4350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1162_
timestamp 1700315010
transform 1 0 4190 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1163_
timestamp 1700315010
transform -1 0 4410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1164_
timestamp 1700315010
transform 1 0 4290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1165_
timestamp 1700315010
transform -1 0 4290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1166_
timestamp 1700315010
transform 1 0 4510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1167_
timestamp 1700315010
transform 1 0 4610 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1168_
timestamp 1700315010
transform -1 0 4790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1169_
timestamp 1700315010
transform 1 0 4650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1170_
timestamp 1700315010
transform 1 0 5170 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1171_
timestamp 1700315010
transform 1 0 5030 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1172_
timestamp 1700315010
transform 1 0 5030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1173_
timestamp 1700315010
transform 1 0 4750 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1174_
timestamp 1700315010
transform -1 0 4910 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1175_
timestamp 1700315010
transform 1 0 4890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1176_
timestamp 1700315010
transform -1 0 5310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1177_
timestamp 1700315010
transform 1 0 5410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1178_
timestamp 1700315010
transform 1 0 5050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1179_
timestamp 1700315010
transform 1 0 5610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1180_
timestamp 1700315010
transform 1 0 5550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1181_
timestamp 1700315010
transform 1 0 5530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1182_
timestamp 1700315010
transform -1 0 5510 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1183_
timestamp 1700315010
transform 1 0 5370 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1184_
timestamp 1700315010
transform -1 0 5510 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1185_
timestamp 1700315010
transform -1 0 4930 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1186_
timestamp 1700315010
transform 1 0 5290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1187_
timestamp 1700315010
transform 1 0 5150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1188_
timestamp 1700315010
transform -1 0 5270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1189_
timestamp 1700315010
transform -1 0 5150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1190_
timestamp 1700315010
transform 1 0 5290 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1191_
timestamp 1700315010
transform 1 0 5230 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1192_
timestamp 1700315010
transform 1 0 5170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1193_
timestamp 1700315010
transform 1 0 4470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1194_
timestamp 1700315010
transform -1 0 4550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1195_
timestamp 1700315010
transform 1 0 4490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1196_
timestamp 1700315010
transform 1 0 3750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1197_
timestamp 1700315010
transform 1 0 4450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1198_
timestamp 1700315010
transform -1 0 3990 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1199_
timestamp 1700315010
transform -1 0 4610 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1200_
timestamp 1700315010
transform 1 0 4890 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1201_
timestamp 1700315010
transform 1 0 4610 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1202_
timestamp 1700315010
transform 1 0 4750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1203_
timestamp 1700315010
transform -1 0 4790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1204_
timestamp 1700315010
transform -1 0 4650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1205_
timestamp 1700315010
transform 1 0 4890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1206_
timestamp 1700315010
transform 1 0 4990 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1207_
timestamp 1700315010
transform 1 0 5010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1208_
timestamp 1700315010
transform 1 0 5170 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1209_
timestamp 1700315010
transform -1 0 5170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1210_
timestamp 1700315010
transform -1 0 4770 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1211_
timestamp 1700315010
transform -1 0 4890 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1212_
timestamp 1700315010
transform -1 0 2370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1213_
timestamp 1700315010
transform 1 0 1950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1214_
timestamp 1700315010
transform 1 0 5570 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1215_
timestamp 1700315010
transform 1 0 2870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1216_
timestamp 1700315010
transform 1 0 4990 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1217_
timestamp 1700315010
transform -1 0 5110 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1218_
timestamp 1700315010
transform 1 0 5010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1219_
timestamp 1700315010
transform 1 0 5010 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1220_
timestamp 1700315010
transform 1 0 5510 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1221_
timestamp 1700315010
transform -1 0 4890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1222_
timestamp 1700315010
transform 1 0 5070 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1223_
timestamp 1700315010
transform 1 0 4730 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1224_
timestamp 1700315010
transform 1 0 4010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1225_
timestamp 1700315010
transform 1 0 3750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1226_
timestamp 1700315010
transform -1 0 3670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1227_
timestamp 1700315010
transform 1 0 3710 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1228_
timestamp 1700315010
transform 1 0 4150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1229_
timestamp 1700315010
transform 1 0 4410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1230_
timestamp 1700315010
transform 1 0 5390 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1231_
timestamp 1700315010
transform 1 0 5430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1232_
timestamp 1700315010
transform 1 0 5150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1233_
timestamp 1700315010
transform -1 0 4770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1234_
timestamp 1700315010
transform -1 0 4910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1235_
timestamp 1700315010
transform 1 0 5290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1236_
timestamp 1700315010
transform -1 0 5410 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1237_
timestamp 1700315010
transform 1 0 3870 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1238_
timestamp 1700315010
transform 1 0 4850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1239_
timestamp 1700315010
transform -1 0 4730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1240_
timestamp 1700315010
transform -1 0 4610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1241_
timestamp 1700315010
transform -1 0 4630 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1242_
timestamp 1700315010
transform -1 0 4490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1243_
timestamp 1700315010
transform -1 0 4310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1244_
timestamp 1700315010
transform 1 0 3510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1245_
timestamp 1700315010
transform 1 0 3870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1246_
timestamp 1700315010
transform -1 0 3870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1247_
timestamp 1700315010
transform -1 0 3590 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1248_
timestamp 1700315010
transform -1 0 3650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1249_
timestamp 1700315010
transform 1 0 3990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1250_
timestamp 1700315010
transform -1 0 4250 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1251_
timestamp 1700315010
transform 1 0 4330 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1252_
timestamp 1700315010
transform -1 0 4110 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1253_
timestamp 1700315010
transform 1 0 3890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1254_
timestamp 1700315010
transform 1 0 4110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1255_
timestamp 1700315010
transform 1 0 3970 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1256_
timestamp 1700315010
transform 1 0 4590 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1257_
timestamp 1700315010
transform -1 0 3970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1258_
timestamp 1700315010
transform 1 0 4130 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1259_
timestamp 1700315010
transform -1 0 4290 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1260_
timestamp 1700315010
transform -1 0 2350 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1261_
timestamp 1700315010
transform 1 0 2350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1262_
timestamp 1700315010
transform -1 0 2470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1263_
timestamp 1700315010
transform -1 0 2470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1264_
timestamp 1700315010
transform -1 0 3090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1265_
timestamp 1700315010
transform 1 0 2930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1266_
timestamp 1700315010
transform 1 0 510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1267_
timestamp 1700315010
transform 1 0 850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1268_
timestamp 1700315010
transform 1 0 390 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1269_
timestamp 1700315010
transform -1 0 1110 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1270_
timestamp 1700315010
transform -1 0 1370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1271_
timestamp 1700315010
transform 1 0 1210 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1272_
timestamp 1700315010
transform 1 0 1330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1273_
timestamp 1700315010
transform 1 0 1830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1274_
timestamp 1700315010
transform -1 0 1470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1275_
timestamp 1700315010
transform 1 0 710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1276_
timestamp 1700315010
transform -1 0 30 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1277_
timestamp 1700315010
transform -1 0 570 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1278_
timestamp 1700315010
transform 1 0 1350 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1279_
timestamp 1700315010
transform 1 0 1210 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1280_
timestamp 1700315010
transform -1 0 310 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1281_
timestamp 1700315010
transform -1 0 430 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1282_
timestamp 1700315010
transform -1 0 30 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1283_
timestamp 1700315010
transform -1 0 150 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1284_
timestamp 1700315010
transform -1 0 270 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1285_
timestamp 1700315010
transform 1 0 610 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1286_
timestamp 1700315010
transform 1 0 1290 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1287_
timestamp 1700315010
transform 1 0 910 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1288_
timestamp 1700315010
transform -1 0 3450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1289_
timestamp 1700315010
transform -1 0 1410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1290_
timestamp 1700315010
transform -1 0 1130 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1291_
timestamp 1700315010
transform 1 0 1570 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1292_
timestamp 1700315010
transform 1 0 1710 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1293_
timestamp 1700315010
transform 1 0 370 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1294_
timestamp 1700315010
transform 1 0 470 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1295_
timestamp 1700315010
transform 1 0 1870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1296_
timestamp 1700315010
transform -1 0 1990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1297_
timestamp 1700315010
transform 1 0 1650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1298_
timestamp 1700315010
transform 1 0 2090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1299_
timestamp 1700315010
transform 1 0 3290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1300_
timestamp 1700315010
transform 1 0 2570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1301_
timestamp 1700315010
transform 1 0 1510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1302_
timestamp 1700315010
transform -1 0 2890 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1303_
timestamp 1700315010
transform 1 0 3010 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1304_
timestamp 1700315010
transform -1 0 2750 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1305_
timestamp 1700315010
transform -1 0 2330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1306_
timestamp 1700315010
transform 1 0 2210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1307_
timestamp 1700315010
transform 1 0 2510 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1308_
timestamp 1700315010
transform 1 0 2370 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1309_
timestamp 1700315010
transform 1 0 2430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1310_
timestamp 1700315010
transform -1 0 1910 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1311_
timestamp 1700315010
transform -1 0 2250 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1312_
timestamp 1700315010
transform 1 0 1510 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1313_
timestamp 1700315010
transform 1 0 2230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1314_
timestamp 1700315010
transform 1 0 2210 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1315_
timestamp 1700315010
transform 1 0 2110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1316_
timestamp 1700315010
transform -1 0 2030 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1317_
timestamp 1700315010
transform 1 0 1970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1318_
timestamp 1700315010
transform 1 0 1110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1319_
timestamp 1700315010
transform -1 0 1010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1320_
timestamp 1700315010
transform 1 0 1030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1321_
timestamp 1700315010
transform 1 0 1230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1322_
timestamp 1700315010
transform -1 0 1730 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1323_
timestamp 1700315010
transform 1 0 2070 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1324_
timestamp 1700315010
transform -1 0 1710 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1325_
timestamp 1700315010
transform 1 0 4370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1326_
timestamp 1700315010
transform 1 0 2090 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1327_
timestamp 1700315010
transform -1 0 1290 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1328_
timestamp 1700315010
transform -1 0 1150 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1329_
timestamp 1700315010
transform 1 0 1690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1330_
timestamp 1700315010
transform -1 0 1710 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1331_
timestamp 1700315010
transform -1 0 1990 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1332_
timestamp 1700315010
transform -1 0 1850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1333_
timestamp 1700315010
transform 1 0 1970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1334_
timestamp 1700315010
transform 1 0 4390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1335_
timestamp 1700315010
transform -1 0 4290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1336_
timestamp 1700315010
transform 1 0 4530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1337_
timestamp 1700315010
transform -1 0 4450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1338_
timestamp 1700315010
transform -1 0 4710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1339_
timestamp 1700315010
transform 1 0 4610 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1340_
timestamp 1700315010
transform -1 0 4570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1341_
timestamp 1700315010
transform -1 0 4510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1342_
timestamp 1700315010
transform 1 0 4710 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1343_
timestamp 1700315010
transform 1 0 5490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1344_
timestamp 1700315010
transform -1 0 5390 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1345_
timestamp 1700315010
transform -1 0 5290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1346_
timestamp 1700315010
transform 1 0 5150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1347_
timestamp 1700315010
transform -1 0 5070 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1348_
timestamp 1700315010
transform 1 0 4750 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1349_
timestamp 1700315010
transform -1 0 5210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1350_
timestamp 1700315010
transform 1 0 5050 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1351_
timestamp 1700315010
transform 1 0 4710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1352_
timestamp 1700315010
transform -1 0 4810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1353_
timestamp 1700315010
transform 1 0 5350 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1354_
timestamp 1700315010
transform 1 0 4910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1355_
timestamp 1700315010
transform 1 0 5030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1356_
timestamp 1700315010
transform 1 0 4910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1357_
timestamp 1700315010
transform 1 0 5150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1358_
timestamp 1700315010
transform 1 0 5310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1359_
timestamp 1700315010
transform 1 0 5030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1360_
timestamp 1700315010
transform -1 0 4910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1361_
timestamp 1700315010
transform -1 0 4770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1362_
timestamp 1700315010
transform 1 0 5050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1363_
timestamp 1700315010
transform -1 0 4870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1364_
timestamp 1700315010
transform 1 0 5270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1365_
timestamp 1700315010
transform 1 0 5610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1366_
timestamp 1700315010
transform -1 0 5410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1367_
timestamp 1700315010
transform -1 0 5130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1368_
timestamp 1700315010
transform -1 0 4450 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1369_
timestamp 1700315010
transform -1 0 3590 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1370_
timestamp 1700315010
transform -1 0 3950 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1371_
timestamp 1700315010
transform -1 0 5510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1372_
timestamp 1700315010
transform 1 0 4970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1373_
timestamp 1700315010
transform 1 0 5230 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1374_
timestamp 1700315010
transform -1 0 5190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1375_
timestamp 1700315010
transform -1 0 4090 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1376_
timestamp 1700315010
transform -1 0 4210 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1377_
timestamp 1700315010
transform 1 0 4810 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1378_
timestamp 1700315010
transform 1 0 4910 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1379_
timestamp 1700315010
transform 1 0 5590 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1380_
timestamp 1700315010
transform -1 0 5170 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1381_
timestamp 1700315010
transform 1 0 5050 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1382_
timestamp 1700315010
transform 1 0 5170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1383_
timestamp 1700315010
transform -1 0 5510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1384_
timestamp 1700315010
transform -1 0 5070 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1385_
timestamp 1700315010
transform 1 0 4470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1386_
timestamp 1700315010
transform 1 0 4430 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1387_
timestamp 1700315010
transform 1 0 4550 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1388_
timestamp 1700315010
transform 1 0 4830 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1389_
timestamp 1700315010
transform 1 0 5190 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1390_
timestamp 1700315010
transform 1 0 5330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1391_
timestamp 1700315010
transform 1 0 5470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1392_
timestamp 1700315010
transform -1 0 4690 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1393_
timestamp 1700315010
transform -1 0 4610 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1394_
timestamp 1700315010
transform 1 0 4930 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1395_
timestamp 1700315010
transform -1 0 4710 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1396_
timestamp 1700315010
transform -1 0 2690 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1397_
timestamp 1700315010
transform 1 0 2850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1398_
timestamp 1700315010
transform 1 0 2770 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1399_
timestamp 1700315010
transform -1 0 2990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1400_
timestamp 1700315010
transform -1 0 2850 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1401_
timestamp 1700315010
transform 1 0 2490 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1402_
timestamp 1700315010
transform -1 0 2550 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1403_
timestamp 1700315010
transform 1 0 2630 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1404_
timestamp 1700315010
transform 1 0 2830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1405_
timestamp 1700315010
transform 1 0 2330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1406_
timestamp 1700315010
transform 1 0 3570 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1407_
timestamp 1700315010
transform -1 0 3610 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1408_
timestamp 1700315010
transform 1 0 3450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1409_
timestamp 1700315010
transform -1 0 2450 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1410_
timestamp 1700315010
transform -1 0 3270 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1411_
timestamp 1700315010
transform -1 0 3390 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1412_
timestamp 1700315010
transform -1 0 3370 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1413_
timestamp 1700315010
transform 1 0 1870 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1414_
timestamp 1700315010
transform 1 0 1730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1415_
timestamp 1700315010
transform -1 0 3170 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1416_
timestamp 1700315010
transform 1 0 1610 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1417_
timestamp 1700315010
transform -1 0 1490 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1418_
timestamp 1700315010
transform 1 0 4090 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1419_
timestamp 1700315010
transform -1 0 3530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1420_
timestamp 1700315010
transform 1 0 3370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1421_
timestamp 1700315010
transform -1 0 4290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1422_
timestamp 1700315010
transform 1 0 4130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1423_
timestamp 1700315010
transform 1 0 4010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1424_
timestamp 1700315010
transform 1 0 3630 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1425_
timestamp 1700315010
transform 1 0 3650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1426_
timestamp 1700315010
transform 1 0 3270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1427_
timestamp 1700315010
transform -1 0 2490 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1428_
timestamp 1700315010
transform -1 0 1970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1429_
timestamp 1700315010
transform -1 0 2110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1430_
timestamp 1700315010
transform -1 0 2630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1431_
timestamp 1700315010
transform 1 0 2470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1432_
timestamp 1700315010
transform -1 0 2350 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1433_
timestamp 1700315010
transform 1 0 2190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1434_
timestamp 1700315010
transform 1 0 1410 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1435_
timestamp 1700315010
transform -1 0 1570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1436_
timestamp 1700315010
transform -1 0 2650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1437_
timestamp 1700315010
transform 1 0 2750 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1438_
timestamp 1700315010
transform -1 0 1370 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1439_
timestamp 1700315010
transform -1 0 1370 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1440_
timestamp 1700315010
transform -1 0 870 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1441_
timestamp 1700315010
transform -1 0 990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1442_
timestamp 1700315010
transform -1 0 870 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1443_
timestamp 1700315010
transform -1 0 990 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1444_
timestamp 1700315010
transform 1 0 2710 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1445_
timestamp 1700315010
transform 1 0 2650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1446_
timestamp 1700315010
transform 1 0 2230 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1447_
timestamp 1700315010
transform 1 0 2090 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1448_
timestamp 1700315010
transform 1 0 2830 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1449_
timestamp 1700315010
transform 1 0 2690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1450_
timestamp 1700315010
transform -1 0 3210 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1451_
timestamp 1700315010
transform 1 0 3330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1527_
timestamp 1700315010
transform 1 0 5530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1528_
timestamp 1700315010
transform 1 0 5370 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1529_
timestamp 1700315010
transform 1 0 5410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1530_
timestamp 1700315010
transform 1 0 5610 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1531_
timestamp 1700315010
transform 1 0 5370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1532_
timestamp 1700315010
transform 1 0 4050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1533_
timestamp 1700315010
transform 1 0 4250 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1534_
timestamp 1700315010
transform 1 0 4310 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1535_
timestamp 1700315010
transform 1 0 4170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1700315010
transform 1 0 1710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1700315010
transform -1 0 2630 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1700315010
transform -1 0 1230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1700315010
transform -1 0 3250 0 1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1700315010
transform 1 0 3770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1700315010
transform 1 0 3930 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1700315010
transform -1 0 3190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert15
timestamp 1700315010
transform -1 0 1390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1700315010
transform 1 0 1730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1700315010
transform -1 0 930 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1700315010
transform -1 0 2870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1700315010
transform 1 0 4930 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1700315010
transform -1 0 2490 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1700315010
transform 1 0 2810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1700315010
transform 1 0 4930 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1700315010
transform -1 0 4090 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1700315010
transform -1 0 2110 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1700315010
transform -1 0 2370 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1700315010
transform -1 0 1990 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1700315010
transform 1 0 790 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1700315010
transform 1 0 2590 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1700315010
transform 1 0 2570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1700315010
transform 1 0 1110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1700315010
transform -1 0 2310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1700315010
transform 1 0 3270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert33
timestamp 1700315010
transform -1 0 950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert7
timestamp 1700315010
transform 1 0 3770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1700315010
transform 1 0 3030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1700315010
transform 1 0 3130 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 3170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1700315010
transform 1 0 3330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert13
timestamp 1700315010
transform 1 0 3390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert14
timestamp 1700315010
transform -1 0 770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__723_
timestamp 1700315010
transform 1 0 3850 0 1 790
box -12 -8 32 272
use FILL  FILL_1__724_
timestamp 1700315010
transform 1 0 3730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__725_
timestamp 1700315010
transform -1 0 3010 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__726_
timestamp 1700315010
transform 1 0 4370 0 1 790
box -12 -8 32 272
use FILL  FILL_1__727_
timestamp 1700315010
transform -1 0 2770 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__728_
timestamp 1700315010
transform 1 0 2770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__729_
timestamp 1700315010
transform 1 0 3450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__730_
timestamp 1700315010
transform 1 0 3970 0 1 790
box -12 -8 32 272
use FILL  FILL_1__731_
timestamp 1700315010
transform 1 0 4510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__732_
timestamp 1700315010
transform 1 0 5510 0 1 270
box -12 -8 32 272
use FILL  FILL_1__733_
timestamp 1700315010
transform 1 0 5330 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__734_
timestamp 1700315010
transform 1 0 5330 0 1 790
box -12 -8 32 272
use FILL  FILL_1__735_
timestamp 1700315010
transform 1 0 2890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__736_
timestamp 1700315010
transform -1 0 4250 0 1 790
box -12 -8 32 272
use FILL  FILL_1__737_
timestamp 1700315010
transform 1 0 3150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__738_
timestamp 1700315010
transform 1 0 3830 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__739_
timestamp 1700315010
transform -1 0 4470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__740_
timestamp 1700315010
transform 1 0 2590 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__741_
timestamp 1700315010
transform -1 0 4330 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__742_
timestamp 1700315010
transform -1 0 3230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__743_
timestamp 1700315010
transform 1 0 3710 0 1 790
box -12 -8 32 272
use FILL  FILL_1__744_
timestamp 1700315010
transform 1 0 2210 0 1 790
box -12 -8 32 272
use FILL  FILL_1__745_
timestamp 1700315010
transform 1 0 3330 0 1 790
box -12 -8 32 272
use FILL  FILL_1__746_
timestamp 1700315010
transform -1 0 3510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__747_
timestamp 1700315010
transform -1 0 3070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__748_
timestamp 1700315010
transform -1 0 3370 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__749_
timestamp 1700315010
transform 1 0 3690 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__750_
timestamp 1700315010
transform -1 0 3170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__751_
timestamp 1700315010
transform -1 0 3290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__752_
timestamp 1700315010
transform 1 0 2790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__753_
timestamp 1700315010
transform -1 0 3150 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__754_
timestamp 1700315010
transform -1 0 3390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__755_
timestamp 1700315010
transform 1 0 3790 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__756_
timestamp 1700315010
transform -1 0 3270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__757_
timestamp 1700315010
transform 1 0 3510 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__758_
timestamp 1700315010
transform 1 0 2850 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__759_
timestamp 1700315010
transform -1 0 2990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__760_
timestamp 1700315010
transform 1 0 2590 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__761_
timestamp 1700315010
transform -1 0 2790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__762_
timestamp 1700315010
transform 1 0 3490 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__763_
timestamp 1700315010
transform -1 0 3630 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__764_
timestamp 1700315010
transform 1 0 3270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__765_
timestamp 1700315010
transform -1 0 3410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__766_
timestamp 1700315010
transform -1 0 2870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__767_
timestamp 1700315010
transform 1 0 2710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__768_
timestamp 1700315010
transform -1 0 2730 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__769_
timestamp 1700315010
transform 1 0 490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__770_
timestamp 1700315010
transform 1 0 750 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__771_
timestamp 1700315010
transform 1 0 590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__772_
timestamp 1700315010
transform -1 0 50 0 1 270
box -12 -8 32 272
use FILL  FILL_1__773_
timestamp 1700315010
transform 1 0 510 0 1 270
box -12 -8 32 272
use FILL  FILL_1__774_
timestamp 1700315010
transform 1 0 370 0 1 270
box -12 -8 32 272
use FILL  FILL_1__775_
timestamp 1700315010
transform -1 0 50 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__776_
timestamp 1700315010
transform 1 0 510 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__777_
timestamp 1700315010
transform 1 0 370 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__778_
timestamp 1700315010
transform 1 0 1250 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__779_
timestamp 1700315010
transform -1 0 1430 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__780_
timestamp 1700315010
transform 1 0 1270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__781_
timestamp 1700315010
transform -1 0 2870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__782_
timestamp 1700315010
transform -1 0 2610 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__783_
timestamp 1700315010
transform -1 0 2730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__784_
timestamp 1700315010
transform 1 0 1610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__785_
timestamp 1700315010
transform 1 0 1850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__786_
timestamp 1700315010
transform -1 0 1870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__787_
timestamp 1700315010
transform -1 0 650 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__788_
timestamp 1700315010
transform 1 0 870 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__789_
timestamp 1700315010
transform 1 0 730 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__790_
timestamp 1700315010
transform -1 0 3970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__791_
timestamp 1700315010
transform -1 0 3870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__792_
timestamp 1700315010
transform 1 0 3810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__793_
timestamp 1700315010
transform 1 0 5570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__794_
timestamp 1700315010
transform -1 0 4670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__795_
timestamp 1700315010
transform -1 0 5210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__796_
timestamp 1700315010
transform -1 0 4850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__797_
timestamp 1700315010
transform -1 0 4670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__798_
timestamp 1700315010
transform -1 0 4710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__799_
timestamp 1700315010
transform -1 0 4130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__800_
timestamp 1700315010
transform -1 0 4050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__801_
timestamp 1700315010
transform 1 0 3970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__802_
timestamp 1700315010
transform -1 0 4870 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__803_
timestamp 1700315010
transform 1 0 3970 0 1 270
box -12 -8 32 272
use FILL  FILL_1__804_
timestamp 1700315010
transform -1 0 4610 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__805_
timestamp 1700315010
transform 1 0 4390 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__806_
timestamp 1700315010
transform -1 0 3790 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__807_
timestamp 1700315010
transform -1 0 3910 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__808_
timestamp 1700315010
transform -1 0 2790 0 1 270
box -12 -8 32 272
use FILL  FILL_1__809_
timestamp 1700315010
transform -1 0 2030 0 1 270
box -12 -8 32 272
use FILL  FILL_1__810_
timestamp 1700315010
transform -1 0 2150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__811_
timestamp 1700315010
transform 1 0 2250 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__812_
timestamp 1700315010
transform -1 0 1770 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__813_
timestamp 1700315010
transform -1 0 1890 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__814_
timestamp 1700315010
transform 1 0 2570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__815_
timestamp 1700315010
transform 1 0 1950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__816_
timestamp 1700315010
transform -1 0 2210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__817_
timestamp 1700315010
transform 1 0 3190 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__818_
timestamp 1700315010
transform -1 0 1210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__819_
timestamp 1700315010
transform 1 0 1470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__820_
timestamp 1700315010
transform -1 0 970 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__821_
timestamp 1700315010
transform 1 0 510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__822_
timestamp 1700315010
transform -1 0 650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__823_
timestamp 1700315010
transform -1 0 850 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__824_
timestamp 1700315010
transform -1 0 1190 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__825_
timestamp 1700315010
transform 1 0 1150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__826_
timestamp 1700315010
transform 1 0 1070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__827_
timestamp 1700315010
transform 1 0 1310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__828_
timestamp 1700315010
transform 1 0 930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__829_
timestamp 1700315010
transform 1 0 830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__830_
timestamp 1700315010
transform -1 0 1570 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__831_
timestamp 1700315010
transform 1 0 1290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__832_
timestamp 1700315010
transform -1 0 1450 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__833_
timestamp 1700315010
transform 1 0 1850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__834_
timestamp 1700315010
transform -1 0 3430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__835_
timestamp 1700315010
transform -1 0 1610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__836_
timestamp 1700315010
transform -1 0 1730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__837_
timestamp 1700315010
transform -1 0 710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__838_
timestamp 1700315010
transform -1 0 710 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__839_
timestamp 1700315010
transform -1 0 570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__840_
timestamp 1700315010
transform -1 0 570 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__841_
timestamp 1700315010
transform -1 0 430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__842_
timestamp 1700315010
transform 1 0 210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__843_
timestamp 1700315010
transform 1 0 370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__844_
timestamp 1700315010
transform -1 0 290 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__845_
timestamp 1700315010
transform 1 0 30 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__846_
timestamp 1700315010
transform 1 0 1950 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__847_
timestamp 1700315010
transform -1 0 570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__848_
timestamp 1700315010
transform -1 0 1290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__849_
timestamp 1700315010
transform -1 0 670 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__850_
timestamp 1700315010
transform -1 0 670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__851_
timestamp 1700315010
transform -1 0 1130 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__852_
timestamp 1700315010
transform -1 0 530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__853_
timestamp 1700315010
transform -1 0 790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__854_
timestamp 1700315010
transform 1 0 1270 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__855_
timestamp 1700315010
transform 1 0 1410 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__856_
timestamp 1700315010
transform 1 0 870 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__857_
timestamp 1700315010
transform -1 0 750 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__858_
timestamp 1700315010
transform -1 0 470 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__859_
timestamp 1700315010
transform -1 0 750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__860_
timestamp 1700315010
transform -1 0 610 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__861_
timestamp 1700315010
transform -1 0 1790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__862_
timestamp 1700315010
transform -1 0 1690 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__863_
timestamp 1700315010
transform -1 0 2570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__864_
timestamp 1700315010
transform 1 0 950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__865_
timestamp 1700315010
transform -1 0 1830 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__866_
timestamp 1700315010
transform -1 0 1550 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__867_
timestamp 1700315010
transform 1 0 590 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__868_
timestamp 1700315010
transform -1 0 190 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__869_
timestamp 1700315010
transform -1 0 150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__870_
timestamp 1700315010
transform -1 0 330 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__871_
timestamp 1700315010
transform -1 0 430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__872_
timestamp 1700315010
transform -1 0 290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__873_
timestamp 1700315010
transform 1 0 270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__874_
timestamp 1700315010
transform -1 0 150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__875_
timestamp 1700315010
transform -1 0 50 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__876_
timestamp 1700315010
transform 1 0 150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__877_
timestamp 1700315010
transform -1 0 950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__878_
timestamp 1700315010
transform -1 0 50 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__879_
timestamp 1700315010
transform -1 0 390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__880_
timestamp 1700315010
transform -1 0 250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__881_
timestamp 1700315010
transform 1 0 970 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__882_
timestamp 1700315010
transform 1 0 930 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__883_
timestamp 1700315010
transform -1 0 1170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__884_
timestamp 1700315010
transform 1 0 770 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__885_
timestamp 1700315010
transform -1 0 50 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__886_
timestamp 1700315010
transform 1 0 1050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__887_
timestamp 1700315010
transform -1 0 50 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__888_
timestamp 1700315010
transform 1 0 450 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__889_
timestamp 1700315010
transform 1 0 450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__890_
timestamp 1700315010
transform 1 0 290 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__891_
timestamp 1700315010
transform 1 0 270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__892_
timestamp 1700315010
transform -1 0 430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__893_
timestamp 1700315010
transform -1 0 470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__894_
timestamp 1700315010
transform -1 0 330 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__895_
timestamp 1700315010
transform -1 0 150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__896_
timestamp 1700315010
transform 1 0 170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__897_
timestamp 1700315010
transform -1 0 2350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__898_
timestamp 1700315010
transform 1 0 2090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__899_
timestamp 1700315010
transform -1 0 3430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__900_
timestamp 1700315010
transform -1 0 2230 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__901_
timestamp 1700315010
transform -1 0 2130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__902_
timestamp 1700315010
transform 1 0 2070 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__903_
timestamp 1700315010
transform -1 0 290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__904_
timestamp 1700315010
transform -1 0 50 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__905_
timestamp 1700315010
transform 1 0 550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__906_
timestamp 1700315010
transform -1 0 50 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__907_
timestamp 1700315010
transform 1 0 170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__908_
timestamp 1700315010
transform 1 0 310 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__909_
timestamp 1700315010
transform -1 0 190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__910_
timestamp 1700315010
transform -1 0 50 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__911_
timestamp 1700315010
transform -1 0 50 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__912_
timestamp 1700315010
transform -1 0 50 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__913_
timestamp 1700315010
transform -1 0 50 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__914_
timestamp 1700315010
transform 1 0 170 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__915_
timestamp 1700315010
transform -1 0 50 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__916_
timestamp 1700315010
transform 1 0 810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__917_
timestamp 1700315010
transform -1 0 670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__918_
timestamp 1700315010
transform -1 0 1890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__919_
timestamp 1700315010
transform -1 0 1270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__920_
timestamp 1700315010
transform 1 0 1270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__921_
timestamp 1700315010
transform 1 0 130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__922_
timestamp 1700315010
transform 1 0 2650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__923_
timestamp 1700315010
transform 1 0 2010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__924_
timestamp 1700315010
transform 1 0 2150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__925_
timestamp 1700315010
transform 1 0 3870 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__926_
timestamp 1700315010
transform -1 0 2330 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__927_
timestamp 1700315010
transform -1 0 2190 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__928_
timestamp 1700315010
transform 1 0 2550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__929_
timestamp 1700315010
transform -1 0 2310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__930_
timestamp 1700315010
transform -1 0 2470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__931_
timestamp 1700315010
transform -1 0 2430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__932_
timestamp 1700315010
transform 1 0 830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__933_
timestamp 1700315010
transform -1 0 150 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__934_
timestamp 1700315010
transform -1 0 330 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__935_
timestamp 1700315010
transform 1 0 1010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__936_
timestamp 1700315010
transform -1 0 590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__937_
timestamp 1700315010
transform 1 0 710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__938_
timestamp 1700315010
transform -1 0 330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__939_
timestamp 1700315010
transform 1 0 170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__940_
timestamp 1700315010
transform 1 0 690 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__941_
timestamp 1700315010
transform 1 0 1090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__942_
timestamp 1700315010
transform 1 0 1070 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__943_
timestamp 1700315010
transform -1 0 890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__944_
timestamp 1700315010
transform -1 0 570 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__945_
timestamp 1700315010
transform -1 0 330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__946_
timestamp 1700315010
transform -1 0 430 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__947_
timestamp 1700315010
transform -1 0 50 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__948_
timestamp 1700315010
transform -1 0 50 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__949_
timestamp 1700315010
transform -1 0 50 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__950_
timestamp 1700315010
transform -1 0 710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__951_
timestamp 1700315010
transform -1 0 470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__952_
timestamp 1700315010
transform 1 0 170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__953_
timestamp 1700315010
transform 1 0 410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__954_
timestamp 1700315010
transform 1 0 590 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__955_
timestamp 1700315010
transform 1 0 690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__956_
timestamp 1700315010
transform 1 0 550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__957_
timestamp 1700315010
transform 1 0 170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__958_
timestamp 1700315010
transform 1 0 870 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__959_
timestamp 1700315010
transform -1 0 1030 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__960_
timestamp 1700315010
transform 1 0 830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__961_
timestamp 1700315010
transform -1 0 750 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__962_
timestamp 1700315010
transform -1 0 1130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__963_
timestamp 1700315010
transform 1 0 1030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__964_
timestamp 1700315010
transform -1 0 890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__965_
timestamp 1700315010
transform 1 0 990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__966_
timestamp 1700315010
transform 1 0 3290 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__967_
timestamp 1700315010
transform -1 0 3170 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__968_
timestamp 1700315010
transform 1 0 1790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__969_
timestamp 1700315010
transform -1 0 890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__970_
timestamp 1700315010
transform 1 0 970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__971_
timestamp 1700315010
transform 1 0 1370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__972_
timestamp 1700315010
transform -1 0 1950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__973_
timestamp 1700315010
transform -1 0 2050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__974_
timestamp 1700315010
transform -1 0 1190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__975_
timestamp 1700315010
transform 1 0 410 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__976_
timestamp 1700315010
transform 1 0 510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__977_
timestamp 1700315010
transform 1 0 2730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__978_
timestamp 1700315010
transform -1 0 2870 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__979_
timestamp 1700315010
transform -1 0 2610 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__980_
timestamp 1700315010
transform 1 0 1790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__981_
timestamp 1700315010
transform 1 0 2410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__982_
timestamp 1700315010
transform -1 0 2470 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__983_
timestamp 1700315010
transform -1 0 2210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__984_
timestamp 1700315010
transform 1 0 2290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__985_
timestamp 1700315010
transform -1 0 2070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__986_
timestamp 1700315010
transform 1 0 2130 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__987_
timestamp 1700315010
transform -1 0 1890 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__988_
timestamp 1700315010
transform 1 0 830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__989_
timestamp 1700315010
transform 1 0 790 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__990_
timestamp 1700315010
transform 1 0 2190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__991_
timestamp 1700315010
transform -1 0 2470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__992_
timestamp 1700315010
transform -1 0 2330 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__993_
timestamp 1700315010
transform 1 0 2710 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__994_
timestamp 1700315010
transform -1 0 2590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__995_
timestamp 1700315010
transform -1 0 2050 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__996_
timestamp 1700315010
transform -1 0 2110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__997_
timestamp 1700315010
transform -1 0 2450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__998_
timestamp 1700315010
transform 1 0 1810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__999_
timestamp 1700315010
transform -1 0 2350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1000_
timestamp 1700315010
transform -1 0 1690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1001_
timestamp 1700315010
transform -1 0 1630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1002_
timestamp 1700315010
transform -1 0 1250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1003_
timestamp 1700315010
transform 1 0 1190 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1004_
timestamp 1700315010
transform 1 0 1510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1005_
timestamp 1700315010
transform -1 0 2190 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1006_
timestamp 1700315010
transform -1 0 1350 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1007_
timestamp 1700315010
transform -1 0 1410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1008_
timestamp 1700315010
transform -1 0 2010 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1009_
timestamp 1700315010
transform 1 0 1750 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1010_
timestamp 1700315010
transform -1 0 1490 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1011_
timestamp 1700315010
transform -1 0 1690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1012_
timestamp 1700315010
transform -1 0 1070 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1013_
timestamp 1700315010
transform 1 0 590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1014_
timestamp 1700315010
transform -1 0 750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1015_
timestamp 1700315010
transform -1 0 1830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1016_
timestamp 1700315010
transform 1 0 1530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1017_
timestamp 1700315010
transform -1 0 1490 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1018_
timestamp 1700315010
transform -1 0 1290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1019_
timestamp 1700315010
transform 1 0 1190 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1020_
timestamp 1700315010
transform -1 0 1630 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1021_
timestamp 1700315010
transform -1 0 1630 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1022_
timestamp 1700315010
transform 1 0 1650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1023_
timestamp 1700315010
transform -1 0 1410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1024_
timestamp 1700315010
transform -1 0 1870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1025_
timestamp 1700315010
transform -1 0 1530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1026_
timestamp 1700315010
transform 1 0 1510 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1027_
timestamp 1700315010
transform 1 0 1370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1028_
timestamp 1700315010
transform 1 0 1890 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1029_
timestamp 1700315010
transform 1 0 1410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1030_
timestamp 1700315010
transform -1 0 1770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1031_
timestamp 1700315010
transform 1 0 1710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1032_
timestamp 1700315010
transform -1 0 1890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1033_
timestamp 1700315010
transform 1 0 1830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1034_
timestamp 1700315010
transform 1 0 1570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1035_
timestamp 1700315010
transform 1 0 1550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1036_
timestamp 1700315010
transform 1 0 1650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1037_
timestamp 1700315010
transform -1 0 2290 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1038_
timestamp 1700315010
transform 1 0 3090 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1039_
timestamp 1700315010
transform 1 0 2090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1040_
timestamp 1700315010
transform 1 0 2190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1041_
timestamp 1700315010
transform -1 0 3050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1042_
timestamp 1700315010
transform 1 0 3550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1043_
timestamp 1700315010
transform 1 0 3290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1044_
timestamp 1700315010
transform 1 0 2890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1045_
timestamp 1700315010
transform -1 0 3010 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1046_
timestamp 1700315010
transform -1 0 3170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1047_
timestamp 1700315010
transform 1 0 3330 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1048_
timestamp 1700315010
transform 1 0 3430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1049_
timestamp 1700315010
transform 1 0 3650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1050_
timestamp 1700315010
transform 1 0 3510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1051_
timestamp 1700315010
transform -1 0 3450 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1052_
timestamp 1700315010
transform -1 0 3190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1053_
timestamp 1700315010
transform 1 0 1930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1054_
timestamp 1700315010
transform -1 0 3950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1055_
timestamp 1700315010
transform -1 0 3990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1056_
timestamp 1700315010
transform 1 0 4090 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1057_
timestamp 1700315010
transform -1 0 3830 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1058_
timestamp 1700315010
transform -1 0 4070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1059_
timestamp 1700315010
transform 1 0 4570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1060_
timestamp 1700315010
transform -1 0 3690 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1061_
timestamp 1700315010
transform -1 0 4230 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1062_
timestamp 1700315010
transform 1 0 4470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1063_
timestamp 1700315010
transform -1 0 4350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1064_
timestamp 1700315010
transform 1 0 3370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1065_
timestamp 1700315010
transform 1 0 2710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1066_
timestamp 1700315010
transform 1 0 2570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1067_
timestamp 1700315010
transform -1 0 4210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1068_
timestamp 1700315010
transform 1 0 3650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1069_
timestamp 1700315010
transform 1 0 3510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1070_
timestamp 1700315010
transform 1 0 3790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1071_
timestamp 1700315010
transform -1 0 3670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1072_
timestamp 1700315010
transform -1 0 3410 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1073_
timestamp 1700315010
transform -1 0 3050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1074_
timestamp 1700315010
transform -1 0 3250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1075_
timestamp 1700315010
transform -1 0 3810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1076_
timestamp 1700315010
transform -1 0 3130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1077_
timestamp 1700315010
transform 1 0 2830 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1078_
timestamp 1700315010
transform 1 0 1890 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1079_
timestamp 1700315010
transform 1 0 1950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1080_
timestamp 1700315010
transform -1 0 2990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1081_
timestamp 1700315010
transform -1 0 3270 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1082_
timestamp 1700315010
transform 1 0 2610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1083_
timestamp 1700315010
transform -1 0 2830 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1084_
timestamp 1700315010
transform -1 0 2770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1085_
timestamp 1700315010
transform -1 0 2490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1086_
timestamp 1700315010
transform 1 0 2670 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1087_
timestamp 1700315010
transform -1 0 2670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1088_
timestamp 1700315010
transform 1 0 1250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1089_
timestamp 1700315010
transform 1 0 1330 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1090_
timestamp 1700315010
transform -1 0 2550 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1091_
timestamp 1700315010
transform 1 0 2950 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1092_
timestamp 1700315010
transform 1 0 2390 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1093_
timestamp 1700315010
transform 1 0 2510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1094_
timestamp 1700315010
transform 1 0 1690 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1095_
timestamp 1700315010
transform -1 0 810 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1096_
timestamp 1700315010
transform -1 0 930 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1097_
timestamp 1700315010
transform 1 0 4510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1098_
timestamp 1700315010
transform -1 0 2270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1099_
timestamp 1700315010
transform -1 0 2650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1100_
timestamp 1700315010
transform 1 0 2750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1101_
timestamp 1700315010
transform 1 0 2890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1102_
timestamp 1700315010
transform 1 0 3190 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1103_
timestamp 1700315010
transform 1 0 3570 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1104_
timestamp 1700315010
transform 1 0 5650 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1105_
timestamp 1700315010
transform 1 0 2990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1106_
timestamp 1700315010
transform 1 0 3090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1107_
timestamp 1700315010
transform 1 0 3770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1108_
timestamp 1700315010
transform 1 0 3650 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1109_
timestamp 1700315010
transform 1 0 3850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1110_
timestamp 1700315010
transform 1 0 3690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1111_
timestamp 1700315010
transform 1 0 3990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1112_
timestamp 1700315010
transform 1 0 4130 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1113_
timestamp 1700315010
transform 1 0 4670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1114_
timestamp 1700315010
transform -1 0 3950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1115_
timestamp 1700315010
transform -1 0 3910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1116_
timestamp 1700315010
transform -1 0 4030 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1117_
timestamp 1700315010
transform 1 0 4050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1118_
timestamp 1700315010
transform 1 0 4190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1119_
timestamp 1700315010
transform -1 0 4750 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1120_
timestamp 1700315010
transform -1 0 4350 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1121_
timestamp 1700315010
transform -1 0 4350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1122_
timestamp 1700315010
transform 1 0 4470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1123_
timestamp 1700315010
transform 1 0 4930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1124_
timestamp 1700315010
transform 1 0 4450 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1125_
timestamp 1700315010
transform -1 0 4610 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1126_
timestamp 1700315010
transform 1 0 4850 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1127_
timestamp 1700315010
transform 1 0 4970 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1128_
timestamp 1700315010
transform 1 0 5110 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1129_
timestamp 1700315010
transform 1 0 3510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1130_
timestamp 1700315010
transform 1 0 3530 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1131_
timestamp 1700315010
transform 1 0 4950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1132_
timestamp 1700315010
transform 1 0 5090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1133_
timestamp 1700315010
transform 1 0 4810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1134_
timestamp 1700315010
transform 1 0 5210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1135_
timestamp 1700315010
transform -1 0 5370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1136_
timestamp 1700315010
transform 1 0 5510 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1137_
timestamp 1700315010
transform 1 0 5210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1138_
timestamp 1700315010
transform 1 0 5490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1139_
timestamp 1700315010
transform 1 0 5530 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1140_
timestamp 1700315010
transform 1 0 5390 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1141_
timestamp 1700315010
transform -1 0 5310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1142_
timestamp 1700315010
transform -1 0 5510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1143_
timestamp 1700315010
transform -1 0 5270 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1144_
timestamp 1700315010
transform -1 0 5370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1145_
timestamp 1700315010
transform 1 0 5290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1146_
timestamp 1700315010
transform 1 0 4990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1147_
timestamp 1700315010
transform 1 0 4630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1148_
timestamp 1700315010
transform -1 0 5570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1149_
timestamp 1700315010
transform 1 0 5410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1150_
timestamp 1700315010
transform 1 0 4130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1151_
timestamp 1700315010
transform -1 0 4830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1152_
timestamp 1700315010
transform 1 0 4650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1153_
timestamp 1700315010
transform -1 0 4170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1154_
timestamp 1700315010
transform 1 0 3890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1155_
timestamp 1700315010
transform 1 0 4350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1156_
timestamp 1700315010
transform 1 0 4270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1157_
timestamp 1700315010
transform 1 0 4010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1158_
timestamp 1700315010
transform 1 0 4410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1159_
timestamp 1700315010
transform 1 0 4090 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1160_
timestamp 1700315010
transform -1 0 3990 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1161_
timestamp 1700315010
transform -1 0 4370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1162_
timestamp 1700315010
transform 1 0 4210 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1163_
timestamp 1700315010
transform -1 0 4430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1164_
timestamp 1700315010
transform 1 0 4310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1165_
timestamp 1700315010
transform -1 0 4310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1166_
timestamp 1700315010
transform 1 0 4530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1167_
timestamp 1700315010
transform 1 0 4630 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1168_
timestamp 1700315010
transform -1 0 4810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1169_
timestamp 1700315010
transform 1 0 4670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1170_
timestamp 1700315010
transform 1 0 5190 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1171_
timestamp 1700315010
transform 1 0 5050 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1172_
timestamp 1700315010
transform 1 0 5050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1173_
timestamp 1700315010
transform 1 0 4770 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1174_
timestamp 1700315010
transform -1 0 4930 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1175_
timestamp 1700315010
transform 1 0 4910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1176_
timestamp 1700315010
transform -1 0 5330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1177_
timestamp 1700315010
transform 1 0 5430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1178_
timestamp 1700315010
transform 1 0 5070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1179_
timestamp 1700315010
transform 1 0 5630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1180_
timestamp 1700315010
transform 1 0 5570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1181_
timestamp 1700315010
transform 1 0 5550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1182_
timestamp 1700315010
transform -1 0 5530 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1183_
timestamp 1700315010
transform 1 0 5390 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1184_
timestamp 1700315010
transform -1 0 5530 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1185_
timestamp 1700315010
transform -1 0 4950 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1186_
timestamp 1700315010
transform 1 0 5310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1187_
timestamp 1700315010
transform 1 0 5170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1188_
timestamp 1700315010
transform -1 0 5290 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1189_
timestamp 1700315010
transform -1 0 5170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1190_
timestamp 1700315010
transform 1 0 5310 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1191_
timestamp 1700315010
transform 1 0 5250 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1192_
timestamp 1700315010
transform 1 0 5190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1193_
timestamp 1700315010
transform 1 0 4490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1194_
timestamp 1700315010
transform -1 0 4570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1195_
timestamp 1700315010
transform 1 0 4510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1196_
timestamp 1700315010
transform 1 0 3770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1197_
timestamp 1700315010
transform 1 0 4470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1198_
timestamp 1700315010
transform -1 0 4010 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1199_
timestamp 1700315010
transform -1 0 4630 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1200_
timestamp 1700315010
transform 1 0 4910 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1201_
timestamp 1700315010
transform 1 0 4630 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1202_
timestamp 1700315010
transform 1 0 4770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1203_
timestamp 1700315010
transform -1 0 4810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1204_
timestamp 1700315010
transform -1 0 4670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1205_
timestamp 1700315010
transform 1 0 4910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1206_
timestamp 1700315010
transform 1 0 5010 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1207_
timestamp 1700315010
transform 1 0 5030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1208_
timestamp 1700315010
transform 1 0 5190 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1209_
timestamp 1700315010
transform -1 0 5190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1210_
timestamp 1700315010
transform -1 0 4790 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1211_
timestamp 1700315010
transform -1 0 4910 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1212_
timestamp 1700315010
transform -1 0 2390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1213_
timestamp 1700315010
transform 1 0 1970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1214_
timestamp 1700315010
transform 1 0 5590 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1215_
timestamp 1700315010
transform 1 0 2890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1216_
timestamp 1700315010
transform 1 0 5010 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1217_
timestamp 1700315010
transform -1 0 5130 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1218_
timestamp 1700315010
transform 1 0 5030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1219_
timestamp 1700315010
transform 1 0 5030 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1220_
timestamp 1700315010
transform 1 0 5530 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1221_
timestamp 1700315010
transform -1 0 4910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1222_
timestamp 1700315010
transform 1 0 5090 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1223_
timestamp 1700315010
transform 1 0 4750 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1224_
timestamp 1700315010
transform 1 0 4030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1225_
timestamp 1700315010
transform 1 0 3770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1226_
timestamp 1700315010
transform -1 0 3690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1227_
timestamp 1700315010
transform 1 0 3730 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1228_
timestamp 1700315010
transform 1 0 4170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1229_
timestamp 1700315010
transform 1 0 4430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1230_
timestamp 1700315010
transform 1 0 5410 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1231_
timestamp 1700315010
transform 1 0 5450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1232_
timestamp 1700315010
transform 1 0 5170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1233_
timestamp 1700315010
transform -1 0 4790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1234_
timestamp 1700315010
transform -1 0 4930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1235_
timestamp 1700315010
transform 1 0 5310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1236_
timestamp 1700315010
transform -1 0 5430 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1237_
timestamp 1700315010
transform 1 0 3890 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1238_
timestamp 1700315010
transform 1 0 4870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1239_
timestamp 1700315010
transform -1 0 4750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1240_
timestamp 1700315010
transform -1 0 4630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1241_
timestamp 1700315010
transform -1 0 4650 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1242_
timestamp 1700315010
transform -1 0 4510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1243_
timestamp 1700315010
transform -1 0 4330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1244_
timestamp 1700315010
transform 1 0 3530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1245_
timestamp 1700315010
transform 1 0 3890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1246_
timestamp 1700315010
transform -1 0 3890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1247_
timestamp 1700315010
transform -1 0 3610 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1248_
timestamp 1700315010
transform -1 0 3670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1249_
timestamp 1700315010
transform 1 0 4010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1250_
timestamp 1700315010
transform -1 0 4270 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1251_
timestamp 1700315010
transform 1 0 4350 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1252_
timestamp 1700315010
transform -1 0 4130 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1253_
timestamp 1700315010
transform 1 0 3910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1254_
timestamp 1700315010
transform 1 0 4130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1255_
timestamp 1700315010
transform 1 0 3990 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1256_
timestamp 1700315010
transform 1 0 4610 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1257_
timestamp 1700315010
transform -1 0 3990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1258_
timestamp 1700315010
transform 1 0 4150 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1259_
timestamp 1700315010
transform -1 0 4310 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1260_
timestamp 1700315010
transform -1 0 2370 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1261_
timestamp 1700315010
transform 1 0 2370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1262_
timestamp 1700315010
transform -1 0 2490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1263_
timestamp 1700315010
transform -1 0 2490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1264_
timestamp 1700315010
transform -1 0 3110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1265_
timestamp 1700315010
transform 1 0 2950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1266_
timestamp 1700315010
transform 1 0 530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1267_
timestamp 1700315010
transform 1 0 870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1268_
timestamp 1700315010
transform 1 0 410 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1269_
timestamp 1700315010
transform -1 0 1130 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1270_
timestamp 1700315010
transform -1 0 1390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1271_
timestamp 1700315010
transform 1 0 1230 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1272_
timestamp 1700315010
transform 1 0 1350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1273_
timestamp 1700315010
transform 1 0 1850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1274_
timestamp 1700315010
transform -1 0 1490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1275_
timestamp 1700315010
transform 1 0 730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1276_
timestamp 1700315010
transform -1 0 50 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1277_
timestamp 1700315010
transform -1 0 590 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1278_
timestamp 1700315010
transform 1 0 1370 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1279_
timestamp 1700315010
transform 1 0 1230 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1280_
timestamp 1700315010
transform -1 0 330 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1281_
timestamp 1700315010
transform -1 0 450 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1282_
timestamp 1700315010
transform -1 0 50 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1283_
timestamp 1700315010
transform -1 0 170 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1284_
timestamp 1700315010
transform -1 0 290 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1285_
timestamp 1700315010
transform 1 0 630 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1286_
timestamp 1700315010
transform 1 0 1310 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1287_
timestamp 1700315010
transform 1 0 930 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1288_
timestamp 1700315010
transform -1 0 3470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1289_
timestamp 1700315010
transform -1 0 1430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1290_
timestamp 1700315010
transform -1 0 1150 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1291_
timestamp 1700315010
transform 1 0 1590 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1292_
timestamp 1700315010
transform 1 0 1730 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1293_
timestamp 1700315010
transform 1 0 390 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1294_
timestamp 1700315010
transform 1 0 490 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1295_
timestamp 1700315010
transform 1 0 1890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1296_
timestamp 1700315010
transform -1 0 2010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1297_
timestamp 1700315010
transform 1 0 1670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1298_
timestamp 1700315010
transform 1 0 2110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1299_
timestamp 1700315010
transform 1 0 3310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1300_
timestamp 1700315010
transform 1 0 2590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1301_
timestamp 1700315010
transform 1 0 1530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1302_
timestamp 1700315010
transform -1 0 2910 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1303_
timestamp 1700315010
transform 1 0 3030 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1304_
timestamp 1700315010
transform -1 0 2770 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1305_
timestamp 1700315010
transform -1 0 2350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1306_
timestamp 1700315010
transform 1 0 2230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1307_
timestamp 1700315010
transform 1 0 2530 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1308_
timestamp 1700315010
transform 1 0 2390 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1309_
timestamp 1700315010
transform 1 0 2450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1310_
timestamp 1700315010
transform -1 0 1930 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1311_
timestamp 1700315010
transform -1 0 2270 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1312_
timestamp 1700315010
transform 1 0 1530 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1313_
timestamp 1700315010
transform 1 0 2250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1314_
timestamp 1700315010
transform 1 0 2230 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1315_
timestamp 1700315010
transform 1 0 2130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1316_
timestamp 1700315010
transform -1 0 2050 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1317_
timestamp 1700315010
transform 1 0 1990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1318_
timestamp 1700315010
transform 1 0 1130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1319_
timestamp 1700315010
transform -1 0 1030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1320_
timestamp 1700315010
transform 1 0 1050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1321_
timestamp 1700315010
transform 1 0 1250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1322_
timestamp 1700315010
transform -1 0 1750 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1323_
timestamp 1700315010
transform 1 0 2090 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1324_
timestamp 1700315010
transform -1 0 1730 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1325_
timestamp 1700315010
transform 1 0 4390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1326_
timestamp 1700315010
transform 1 0 2110 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1327_
timestamp 1700315010
transform -1 0 1310 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1328_
timestamp 1700315010
transform -1 0 1170 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1329_
timestamp 1700315010
transform 1 0 1710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1330_
timestamp 1700315010
transform -1 0 1730 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1331_
timestamp 1700315010
transform -1 0 2010 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1332_
timestamp 1700315010
transform -1 0 1870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1333_
timestamp 1700315010
transform 1 0 1990 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1334_
timestamp 1700315010
transform 1 0 4410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1335_
timestamp 1700315010
transform -1 0 4310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1336_
timestamp 1700315010
transform 1 0 4550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1337_
timestamp 1700315010
transform -1 0 4470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1338_
timestamp 1700315010
transform -1 0 4730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1339_
timestamp 1700315010
transform 1 0 4630 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1340_
timestamp 1700315010
transform -1 0 4590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1341_
timestamp 1700315010
transform -1 0 4530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1342_
timestamp 1700315010
transform 1 0 4730 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1343_
timestamp 1700315010
transform 1 0 5510 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1344_
timestamp 1700315010
transform -1 0 5410 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1345_
timestamp 1700315010
transform -1 0 5310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1346_
timestamp 1700315010
transform 1 0 5170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1347_
timestamp 1700315010
transform -1 0 5090 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1348_
timestamp 1700315010
transform 1 0 4770 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1349_
timestamp 1700315010
transform -1 0 5230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1350_
timestamp 1700315010
transform 1 0 5070 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1351_
timestamp 1700315010
transform 1 0 4730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1352_
timestamp 1700315010
transform -1 0 4830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1353_
timestamp 1700315010
transform 1 0 5370 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1354_
timestamp 1700315010
transform 1 0 4930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1355_
timestamp 1700315010
transform 1 0 5050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1356_
timestamp 1700315010
transform 1 0 4930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1357_
timestamp 1700315010
transform 1 0 5170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1358_
timestamp 1700315010
transform 1 0 5330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1359_
timestamp 1700315010
transform 1 0 5050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1360_
timestamp 1700315010
transform -1 0 4930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1361_
timestamp 1700315010
transform -1 0 4790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1362_
timestamp 1700315010
transform 1 0 5070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1363_
timestamp 1700315010
transform -1 0 4890 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1364_
timestamp 1700315010
transform 1 0 5290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1365_
timestamp 1700315010
transform 1 0 5630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1366_
timestamp 1700315010
transform -1 0 5430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1367_
timestamp 1700315010
transform -1 0 5150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1368_
timestamp 1700315010
transform -1 0 4470 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1369_
timestamp 1700315010
transform -1 0 3610 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1370_
timestamp 1700315010
transform -1 0 3970 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1371_
timestamp 1700315010
transform -1 0 5530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1372_
timestamp 1700315010
transform 1 0 4990 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1373_
timestamp 1700315010
transform 1 0 5250 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1374_
timestamp 1700315010
transform -1 0 5210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1375_
timestamp 1700315010
transform -1 0 4110 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1376_
timestamp 1700315010
transform -1 0 4230 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1377_
timestamp 1700315010
transform 1 0 4830 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1378_
timestamp 1700315010
transform 1 0 4930 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1379_
timestamp 1700315010
transform 1 0 5610 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1380_
timestamp 1700315010
transform -1 0 5190 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1381_
timestamp 1700315010
transform 1 0 5070 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1382_
timestamp 1700315010
transform 1 0 5190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1383_
timestamp 1700315010
transform -1 0 5530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1384_
timestamp 1700315010
transform -1 0 5090 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1385_
timestamp 1700315010
transform 1 0 4490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1386_
timestamp 1700315010
transform 1 0 4450 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1387_
timestamp 1700315010
transform 1 0 4570 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1388_
timestamp 1700315010
transform 1 0 4850 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1389_
timestamp 1700315010
transform 1 0 5210 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1390_
timestamp 1700315010
transform 1 0 5350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1391_
timestamp 1700315010
transform 1 0 5490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1392_
timestamp 1700315010
transform -1 0 4710 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1393_
timestamp 1700315010
transform -1 0 4630 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1394_
timestamp 1700315010
transform 1 0 4950 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1395_
timestamp 1700315010
transform -1 0 4730 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1396_
timestamp 1700315010
transform -1 0 2710 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1397_
timestamp 1700315010
transform 1 0 2870 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1398_
timestamp 1700315010
transform 1 0 2790 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1399_
timestamp 1700315010
transform -1 0 3010 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1400_
timestamp 1700315010
transform -1 0 2870 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1401_
timestamp 1700315010
transform 1 0 2510 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1402_
timestamp 1700315010
transform -1 0 2570 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1403_
timestamp 1700315010
transform 1 0 2650 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1404_
timestamp 1700315010
transform 1 0 2850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1405_
timestamp 1700315010
transform 1 0 2350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1406_
timestamp 1700315010
transform 1 0 3590 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1407_
timestamp 1700315010
transform -1 0 3630 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1408_
timestamp 1700315010
transform 1 0 3470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1409_
timestamp 1700315010
transform -1 0 2470 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1410_
timestamp 1700315010
transform -1 0 3290 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1411_
timestamp 1700315010
transform -1 0 3410 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1412_
timestamp 1700315010
transform -1 0 3390 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1413_
timestamp 1700315010
transform 1 0 1890 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1414_
timestamp 1700315010
transform 1 0 1750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1415_
timestamp 1700315010
transform -1 0 3190 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1416_
timestamp 1700315010
transform 1 0 1630 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1417_
timestamp 1700315010
transform -1 0 1510 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1418_
timestamp 1700315010
transform 1 0 4110 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1419_
timestamp 1700315010
transform -1 0 3550 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1420_
timestamp 1700315010
transform 1 0 3390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1421_
timestamp 1700315010
transform -1 0 4310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1422_
timestamp 1700315010
transform 1 0 4150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1423_
timestamp 1700315010
transform 1 0 4030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1424_
timestamp 1700315010
transform 1 0 3650 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1425_
timestamp 1700315010
transform 1 0 3670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1426_
timestamp 1700315010
transform 1 0 3290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1427_
timestamp 1700315010
transform -1 0 2510 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1428_
timestamp 1700315010
transform -1 0 1990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1429_
timestamp 1700315010
transform -1 0 2130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1430_
timestamp 1700315010
transform -1 0 2650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1431_
timestamp 1700315010
transform 1 0 2490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1432_
timestamp 1700315010
transform -1 0 2370 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1433_
timestamp 1700315010
transform 1 0 2210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1434_
timestamp 1700315010
transform 1 0 1430 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1435_
timestamp 1700315010
transform -1 0 1590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1436_
timestamp 1700315010
transform -1 0 2670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1437_
timestamp 1700315010
transform 1 0 2770 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1438_
timestamp 1700315010
transform -1 0 1390 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1439_
timestamp 1700315010
transform -1 0 1390 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1440_
timestamp 1700315010
transform -1 0 890 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1441_
timestamp 1700315010
transform -1 0 1010 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1442_
timestamp 1700315010
transform -1 0 890 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1443_
timestamp 1700315010
transform -1 0 1010 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1444_
timestamp 1700315010
transform 1 0 2730 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1445_
timestamp 1700315010
transform 1 0 2670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1446_
timestamp 1700315010
transform 1 0 2250 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1447_
timestamp 1700315010
transform 1 0 2110 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1448_
timestamp 1700315010
transform 1 0 2850 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1449_
timestamp 1700315010
transform 1 0 2710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1450_
timestamp 1700315010
transform -1 0 3230 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1451_
timestamp 1700315010
transform 1 0 3350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1527_
timestamp 1700315010
transform 1 0 5550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1528_
timestamp 1700315010
transform 1 0 5390 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1529_
timestamp 1700315010
transform 1 0 5430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1530_
timestamp 1700315010
transform 1 0 5630 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1531_
timestamp 1700315010
transform 1 0 5390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1532_
timestamp 1700315010
transform 1 0 4070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1533_
timestamp 1700315010
transform 1 0 4270 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1534_
timestamp 1700315010
transform 1 0 4330 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1535_
timestamp 1700315010
transform 1 0 4190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1700315010
transform 1 0 1730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1700315010
transform -1 0 2650 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1700315010
transform -1 0 1250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1700315010
transform -1 0 3270 0 1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1700315010
transform 1 0 3790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1700315010
transform 1 0 3950 0 -1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert6
timestamp 1700315010
transform -1 0 3210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert15
timestamp 1700315010
transform -1 0 1410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1700315010
transform 1 0 1750 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1700315010
transform -1 0 950 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1700315010
transform -1 0 2890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1700315010
transform 1 0 4950 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1700315010
transform -1 0 2510 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1700315010
transform 1 0 2830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1700315010
transform 1 0 4950 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1700315010
transform -1 0 4110 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1700315010
transform -1 0 2130 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1700315010
transform -1 0 2390 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1700315010
transform -1 0 2010 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert27
timestamp 1700315010
transform 1 0 810 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1700315010
transform 1 0 2610 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert29
timestamp 1700315010
transform 1 0 2590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1700315010
transform 1 0 1130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert31
timestamp 1700315010
transform -1 0 2330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1700315010
transform 1 0 3290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert33
timestamp 1700315010
transform -1 0 970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert7
timestamp 1700315010
transform 1 0 3790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1700315010
transform 1 0 3050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1700315010
transform 1 0 3150 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 3190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1700315010
transform 1 0 3350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 1010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert13
timestamp 1700315010
transform 1 0 3410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert14
timestamp 1700315010
transform -1 0 790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1450_
timestamp 1700315010
transform -1 0 3250 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert33
timestamp 1700315010
transform -1 0 990 0 -1 5470
box -12 -8 32 272
<< labels >>
flabel metal1 s 5763 2 5823 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 3877 5517 3883 5523 3 FreeSans 16 90 0 0 Cin[5]
port 2 nsew
flabel metal2 s 3417 5517 3423 5523 3 FreeSans 16 90 0 0 Cin[2]
port 5 nsew
flabel metal3 s -24 1956 -16 1964 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal3 s 5796 2736 5804 2744 3 FreeSans 16 0 0 0 Vld
port 9 nsew
flabel metal3 s -24 3556 -16 3564 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s -24 3516 -16 3524 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal3 s -24 3036 -16 3044 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal3 s 5796 4076 5804 4084 3 FreeSans 16 0 0 0 Xout[3]
port 14 nsew
flabel metal3 s 5796 4036 5804 4044 3 FreeSans 16 0 0 0 Xout[2]
port 15 nsew
flabel metal3 s 5796 3776 5804 3784 3 FreeSans 16 0 0 0 Xout[1]
port 16 nsew
flabel metal3 s 5796 2996 5804 3004 3 FreeSans 16 0 0 0 Xout[0]
port 17 nsew
flabel metal2 s 2497 -23 2503 -17 7 FreeSans 16 270 0 0 Yin[1]
port 20 nsew
flabel metal2 s 2397 -23 2403 -17 7 FreeSans 16 270 0 0 Yin[0]
port 21 nsew
flabel metal2 s 4337 -23 4343 -17 7 FreeSans 16 270 0 0 Yout[1]
port 24 nsew
flabel metal2 s 3057 5517 3063 5523 3 FreeSans 16 90 0 0 clk
port 26 nsew
flabel metal2 s 2897 5517 2903 5523 3 FreeSans 16 90 0 0 Cin[0]
port 7 nsew
flabel metal2 s 3217 5517 3223 5523 3 FreeSans 16 90 0 0 Cin[1]
port 6 nsew
flabel metal2 s 4177 5517 4183 5523 3 FreeSans 16 90 0 0 Cin[4]
port 3 nsew
flabel metal2 s 3917 5517 3923 5523 3 FreeSans 16 90 0 0 Cin[3]
port 4 nsew
flabel metal2 s 4257 -23 4263 -17 7 FreeSans 16 270 0 0 Yout[2]
port 23 nsew
flabel metal2 s 4117 -23 4123 -17 7 FreeSans 16 270 0 0 Yout[0]
port 25 nsew
flabel metal2 s 4157 -23 4163 -17 7 FreeSans 16 270 0 0 Yout[3]
port 22 nsew
flabel metal2 s 3297 -23 3303 -17 7 FreeSans 16 270 0 0 Yin[3]
port 18 nsew
flabel metal2 s 3337 -23 3343 -17 7 FreeSans 16 270 0 0 Yin[2]
port 19 nsew
<< properties >>
string FIXED_BBOX -40 -40 5800 5520
<< end >>
