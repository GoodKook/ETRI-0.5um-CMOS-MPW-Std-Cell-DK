magic
tech scmos
magscale 1 2
timestamp 1726828718
<< nwell >>
rect -13 154 313 272
rect 60 150 247 154
rect 160 136 247 150
rect 188 135 222 136
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
rect 90 14 94 54
rect 110 14 114 54
rect 130 14 134 54
rect 150 14 154 54
rect 170 14 174 54
rect 192 14 196 54
rect 202 14 206 54
rect 212 14 216 54
rect 232 14 236 34
rect 276 14 280 34
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
rect 80 166 84 246
rect 90 166 94 246
rect 110 166 114 246
rect 130 174 134 246
rect 150 174 154 246
rect 170 174 174 246
rect 192 150 196 246
rect 202 150 206 246
rect 212 150 216 246
rect 232 206 236 246
rect 276 206 280 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 42 40 54
rect 24 14 26 42
rect 38 14 40 42
rect 44 48 60 54
rect 44 14 46 48
rect 58 14 60 48
rect 64 46 80 54
rect 64 14 66 46
rect 78 14 80 46
rect 84 14 90 54
rect 94 50 110 54
rect 94 18 96 50
rect 108 18 110 50
rect 94 14 110 18
rect 114 52 130 54
rect 114 14 116 52
rect 128 14 130 52
rect 134 40 150 54
rect 134 18 136 40
rect 148 18 150 40
rect 134 14 150 18
rect 154 52 170 54
rect 154 14 156 52
rect 168 14 170 52
rect 174 44 192 54
rect 174 14 177 44
rect 189 14 192 44
rect 196 14 202 54
rect 206 14 212 54
rect 216 34 226 54
rect 216 14 218 34
rect 230 14 232 34
rect 236 14 238 34
rect 274 14 276 34
rect 280 14 282 34
<< pdiffusion >>
rect 18 166 20 246
rect 24 180 26 246
rect 38 180 40 246
rect 24 166 40 180
rect 44 180 46 246
rect 58 180 60 246
rect 44 166 60 180
rect 64 176 66 246
rect 78 176 80 246
rect 64 166 80 176
rect 84 166 90 246
rect 94 166 96 246
rect 108 166 110 246
rect 114 174 116 246
rect 128 174 130 246
rect 134 186 136 246
rect 148 186 150 246
rect 134 174 150 186
rect 154 176 156 246
rect 168 176 170 246
rect 154 174 170 176
rect 174 174 177 246
rect 189 174 192 246
rect 114 166 124 174
rect 180 150 192 174
rect 196 150 202 246
rect 206 150 212 246
rect 216 206 218 246
rect 230 206 232 246
rect 236 206 238 246
rect 274 206 276 246
rect 280 206 282 246
rect 216 150 227 206
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 42
rect 46 14 58 48
rect 66 14 78 46
rect 96 18 108 50
rect 116 14 128 52
rect 136 18 148 40
rect 156 14 168 52
rect 177 14 189 44
rect 218 14 230 34
rect 238 14 250 34
rect 262 14 274 34
rect 282 14 294 34
<< pdcontact >>
rect 6 166 18 246
rect 26 180 38 246
rect 46 180 58 246
rect 66 176 78 246
rect 96 166 108 246
rect 116 174 128 246
rect 136 186 148 246
rect 156 176 168 246
rect 177 174 189 246
rect 218 206 230 246
rect 238 206 250 246
rect 262 206 274 246
rect 282 206 294 246
<< psubstratepcontact >>
rect -6 -6 306 6
<< nsubstratencontact >>
rect -6 254 306 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 90 246 94 250
rect 110 246 114 250
rect 130 246 134 250
rect 150 246 154 250
rect 170 246 174 250
rect 192 246 196 250
rect 202 246 206 250
rect 212 246 216 250
rect 232 246 236 250
rect 276 246 280 250
rect 20 129 24 166
rect 20 54 24 117
rect 40 97 44 166
rect 60 117 64 166
rect 40 54 44 84
rect 60 54 64 105
rect 80 97 84 166
rect 90 162 94 166
rect 110 162 114 166
rect 130 162 134 174
rect 150 170 154 174
rect 170 170 174 174
rect 90 158 114 162
rect 120 158 134 162
rect 138 166 154 170
rect 159 166 174 170
rect 80 54 84 84
rect 96 78 100 158
rect 120 97 124 158
rect 138 154 142 166
rect 132 150 142 154
rect 132 122 137 150
rect 159 142 164 166
rect 158 130 164 142
rect 192 135 196 150
rect 96 62 108 66
rect 120 62 124 84
rect 140 62 144 110
rect 159 62 164 130
rect 179 131 196 135
rect 179 123 184 131
rect 202 123 206 150
rect 204 110 206 123
rect 180 72 184 110
rect 180 68 196 72
rect 90 58 114 62
rect 120 58 134 62
rect 140 58 154 62
rect 159 58 174 62
rect 90 54 94 58
rect 110 54 114 58
rect 130 54 134 58
rect 150 54 154 58
rect 170 54 174 58
rect 192 54 196 68
rect 202 54 206 110
rect 212 78 216 150
rect 232 141 236 206
rect 212 65 214 78
rect 212 54 216 65
rect 235 56 240 129
rect 232 51 240 56
rect 232 34 236 51
rect 276 34 280 206
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
rect 90 10 94 14
rect 110 10 114 14
rect 130 10 134 14
rect 150 10 154 14
rect 170 10 174 14
rect 192 10 196 14
rect 202 10 206 14
rect 212 10 216 14
rect 232 10 236 14
rect 276 10 280 14
<< polycontact >>
rect 20 117 32 129
rect 57 105 69 117
rect 40 84 52 97
rect 76 84 88 97
rect 146 130 158 142
rect 132 110 144 122
rect 116 84 128 97
rect 96 66 108 78
rect 172 110 184 123
rect 192 110 204 123
rect 264 164 276 176
rect 230 129 242 141
rect 214 65 226 78
<< metal1 >>
rect -6 266 306 268
rect -6 252 306 254
rect 26 246 38 252
rect 96 246 108 252
rect 136 246 148 252
rect 218 246 230 252
rect 262 246 274 252
rect 46 172 55 180
rect 66 174 78 176
rect 18 166 55 172
rect 128 176 156 180
rect 128 174 168 176
rect 176 174 177 246
rect 236 206 238 215
rect 176 160 189 174
rect 177 146 189 160
rect 236 156 242 206
rect 282 156 290 206
rect 236 150 255 156
rect 146 142 157 146
rect 183 141 189 146
rect 183 135 230 141
rect 69 110 132 117
rect 144 110 172 118
rect 249 117 255 150
rect 263 148 290 156
rect 263 117 271 148
rect 192 104 203 110
rect 116 103 203 104
rect 24 78 34 103
rect 116 97 217 103
rect 52 84 76 91
rect 88 84 116 91
rect 147 78 198 84
rect 24 72 96 78
rect 108 72 155 78
rect 190 72 214 78
rect 18 48 54 54
rect 177 58 183 72
rect 66 46 77 52
rect 26 8 38 14
rect 96 8 108 18
rect 128 46 156 52
rect 136 8 148 18
rect 176 44 183 58
rect 249 48 255 103
rect 176 14 177 44
rect 240 40 255 48
rect 240 34 246 40
rect 263 34 270 103
rect 218 8 226 14
rect 282 8 294 14
rect -6 6 306 8
rect -6 -8 306 -6
<< m2contact >>
rect 63 160 77 174
rect 143 146 157 160
rect 163 146 177 160
rect 250 163 264 177
rect 23 103 37 117
rect 43 103 57 117
rect 203 110 204 117
rect 204 110 217 117
rect 203 103 217 110
rect 243 103 257 117
rect 263 103 277 117
rect 63 52 77 66
rect 163 58 177 72
<< metal2 >>
rect 77 168 250 174
rect 143 160 157 168
rect 46 117 54 134
rect 26 86 34 103
rect 67 66 73 160
rect 167 72 175 146
rect 266 117 274 134
rect 206 86 214 103
rect 246 86 254 103
<< m1p >>
rect -6 252 306 268
rect -6 -8 306 8
<< m2p >>
rect 46 119 54 134
rect 266 119 274 134
rect 26 86 34 101
rect 206 86 214 101
rect 246 86 254 101
<< labels >>
rlabel metal1 -6 252 306 268 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -6 -8 306 8 0 gnd
port 7 nsew ground bidirectional abutment
rlabel metal2 30 90 30 90 3 A
port 1 n signal input
rlabel metal2 50 131 50 131 1 C
port 3 n signal input
rlabel metal2 250 88 250 88 7 YS
port 4 n signal output
rlabel metal2 210 89 210 89 3 B
port 2 n signal input
rlabel metal2 270 127 270 127 5 YC
port 5 n signal output
<< properties >>
string FIXED_BBOX 0 0 300 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
