/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module cpu(
    inout vdd,
    inout gnd,
    output [15:0] AB,
    input [7:0] DI,
    output [7:0] DO,
    input IRQ,
    input NMI,
    input RDY,
    output WE,
    input clk,
    input reset
);

wire C ;
wire D ;
wire I ;
wire N ;
wire V ;
wire Z ;
wire _1677_ ;
wire _1257_ ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _1295_ ;
wire _703_ ;
wire _1389_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _1198_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _929_ ;
wire _509_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire _16_ ;
wire _1195_ ;
wire _54_ ;
wire _603_ ;
wire _1289_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _1098_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _926_ ;
wire _506_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire IRQ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _1727_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1__bF$buf10 ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire WE ;
wire _1383_ ;
wire _294_ ;
wire _13_ ;
wire _1439_ ;
wire _1019_ ;
wire php ;
wire _1192_ ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _1095_ ;
wire _7_ ;
wire RDY ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire adc_sbc ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _1724_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _10_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _1283_ ;
wire _194_ ;
wire _1339_ ;
wire _1092_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire write_back ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _1721_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _902__bF$buf0 ;
wire _902__bF$buf1 ;
wire _902__bF$buf2 ;
wire _902__bF$buf3 ;
wire _1718_ ;
wire _629_ ;
wire _209_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _1374_ ;
wire _285_ ;
wire _1_ ;
wire index_y ;
wire _1183_ ;
wire _1659_ ;
wire _1239_ ;
wire _42_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire clc ;
wire cld ;
wire cli ;
wire clk ;
wire clv ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _1715_ ;
wire _626_ ;
wire _206_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1371_ ;
wire _282_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _1319__bF$buf0 ;
wire _1319__bF$buf1 ;
wire _1319__bF$buf2 ;
wire _1319__bF$buf3 ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _1083_ ;
wire _1559_ ;
wire _1139_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _1027__bF$buf0 ;
wire _1027__bF$buf1 ;
wire _1027__bF$buf2 ;
wire _1027__bF$buf3 ;
wire _1027__bF$buf4 ;
wire _1712_ ;
wire _623_ ;
wire _203_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _1709_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire HC ;
wire _33_ ;
wire _1459_ ;
wire _1039_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire [7:0] ADD ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _1706_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _1609_ ;
wire _1362_ ;
wire RDY_bF$buf0 ;
wire RDY_bF$buf1 ;
wire RDY_bF$buf2 ;
wire RDY_bF$buf3 ;
wire RDY_bF$buf4 ;
wire RDY_bF$buf5 ;
wire RDY_bF$buf6 ;
wire RDY_bF$buf7 ;
wire RDY_bF$buf8 ;
wire RDY_bF$buf9 ;
wire _693_ ;
wire _273_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _1456_ ;
wire _1036_ ;
wire res ;
wire _787_ ;
wire _367_ ;
wire rotate ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire [3:0] alu_op ;
wire _1359_ ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire [1:0] dst_reg ;
wire \u_ALU8.BI7  ;
wire _805_ ;
wire [7:0] DIHOLD ;
wire _65_ ;
wire _1703_ ;
wire _614_ ;
wire _903__bF$buf0 ;
wire _903__bF$buf1 ;
wire _903__bF$buf2 ;
wire _903__bF$buf3 ;
wire [5:0] _1512_ ;
wire _843_ ;
wire _423_ ;
wire [15:0] _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _1738_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _24_ ;
wire _1679_ ;
wire _1259_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _1700_ ;
wire _611_ ;
wire _1714__bF$buf0 ;
wire _1714__bF$buf1 ;
wire _1714__bF$buf2 ;
wire _1714__bF$buf3 ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire \u_ALU8.BCD  ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _21_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire [7:0] \AXYS[1]  ;
wire _1579_ ;
wire _1159_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _928_ ;
wire _508_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _1729_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _1194_ ;
wire _53_ ;
wire _1479_ ;
wire _1059_ ;
wire store ;
wire _602_ ;
wire _1288_ ;
wire _199_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire IRHOLD_valid ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _1726_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _12_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _1285_ ;
wire _196_ ;
wire _1094_ ;
wire _1379_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire _1188_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _1723_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _1__bF$buf0 ;
wire _1__bF$buf1 ;
wire _1__bF$buf2 ;
wire _1__bF$buf3 ;
wire _1__bF$buf4 ;
wire _1__bF$buf5 ;
wire _1__bF$buf6 ;
wire _1__bF$buf7 ;
wire _1__bF$buf8 ;
wire _1__bF$buf9 ;
wire _919_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire backwards ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _44_ ;
wire _1699_ ;
wire _1279_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1720_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire [15:0] PC ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _1717_ ;
wire _628_ ;
wire _208_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _1373_ ;
wire _284_ ;
wire _0_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire adj_bcd ;
wire _41_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire _913_ ;
wire [7:0] \AXYS[3]  ;
wire _1599_ ;
wire _1179_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire compare ;
wire _816_ ;
wire _76_ ;
wire _1714_ ;
wire _625_ ;
wire _205_ ;
wire load_only ;
wire clk_bF$buf10 ;
wire shift ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1370_ ;
wire _281_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire [1:0] src_reg ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _1329_ ;
wire _1082_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire _35_ ;
wire _1149__bF$buf0 ;
wire _1149__bF$buf1 ;
wire _1149__bF$buf2 ;
wire _1149__bF$buf3 ;
wire _1149__bF$buf4 ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _1711_ ;
wire _622_ ;
wire _202_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _1708_ ;
wire _619_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _1593_ ;
wire _1173_ ;
wire _1649_ ;
wire _1229_ ;
wire _32_ ;
wire _1458_ ;
wire _1038_ ;
wire [2:0] cond_code ;
wire _789_ ;
wire _369_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _904_ ;
wire _713_ ;
wire _1399_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _1705_ ;
wire _616_ ;
wire [5:0] state ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire bit_ins ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire [7:0] DI ;
wire [7:0] DO ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _1493_ ;
wire _1073_ ;
wire _1549_ ;
wire _1129_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _1702_ ;
wire _613_ ;
wire _1299_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire [15:0] AB ;
wire [7:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _1737_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _1393_ ;
wire _23_ ;
wire _1449_ ;
wire _1029_ ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire _886__bF$buf0 ;
wire _886__bF$buf1 ;
wire _886__bF$buf2 ;
wire _886__bF$buf3 ;
wire _886__bF$buf4 ;
wire _886__bF$buf5 ;
wire _886__bF$buf6 ;
wire _704_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _1199_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire NMI ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _20_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _1293_ ;
wire _1349_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire plp ;
wire _1196_ ;
wire _55_ ;
wire _604_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _1099_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _1728_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire _295_ ;
wire _14_ ;
wire _1193_ ;
wire _1669_ ;
wire _1249_ ;
wire _52_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _1096_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _1725_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _11_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _1093_ ;
wire [7:0] \AXYS[0]  ;
wire _1569_ ;
wire _1149_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _1722_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _1719_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _1528_ ;
wire _1108_ ;
wire shift_right ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _914__bF$buf0 ;
wire _914__bF$buf1 ;
wire _914__bF$buf2 ;
wire _914__bF$buf3 ;
wire _914__bF$buf4 ;
wire _43_ ;
wire _1469_ ;
wire _1049_ ;
wire [7:0] DIMUX ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _1150__bF$buf0 ;
wire _1150__bF$buf1 ;
wire _1150__bF$buf2 ;
wire _1150__bF$buf3 ;
wire _1150__bF$buf4 ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire [3:0] op ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _1716_ ;
wire _627_ ;
wire _207_ ;
wire _720__bF$buf0 ;
wire _720__bF$buf1 ;
wire _720__bF$buf2 ;
wire _720__bF$buf3 ;
wire _380_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _1619_ ;
wire _1372_ ;
wire _283_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire sec ;
wire sed ;
wire sei ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire [7:0] IRHOLD ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire alu_shift_right ;
wire _1084_ ;
wire _1369_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _1713_ ;
wire _624_ ;
wire _204_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _1519_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire _34_ ;
wire _1689_ ;
wire _1269_ ;
wire NMI_1 ;
wire _812_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _1710_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire adc_bcd ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _1707_ ;
wire _618_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _931__bF$buf0 ;
wire _931__bF$buf1 ;
wire _931__bF$buf2 ;
wire _931__bF$buf3 ;
wire _931__bF$buf4 ;
wire _903_ ;
wire [7:0] \AXYS[2]  ;
wire _1589_ ;
wire _1169_ ;
wire _712_ ;
wire [7:0] ABH ;
wire [7:0] ABL ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire NMI_edge ;
wire _806_ ;
wire _66_ ;
wire _1704_ ;
wire _615_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire [7:0] _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire load_reg ;
wire _709_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire CI ;
wire CO ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _1739_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire inc ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _1701_ ;
wire _612_ ;
wire _1298_ ;
wire reset ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _22_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert83 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319_),
    .Y(_1319__bF$buf0)
);

BUFX2 BUFX2_insert82 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319_),
    .Y(_1319__bF$buf1)
);

BUFX2 BUFX2_insert81 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319_),
    .Y(_1319__bF$buf2)
);

BUFX2 BUFX2_insert80 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319_),
    .Y(_1319__bF$buf3)
);

BUFX2 BUFX2_insert79 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903_),
    .Y(_903__bF$buf0)
);

BUFX2 BUFX2_insert78 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903_),
    .Y(_903__bF$buf1)
);

BUFX2 BUFX2_insert77 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903_),
    .Y(_903__bF$buf2)
);

BUFX2 BUFX2_insert76 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903_),
    .Y(_903__bF$buf3)
);

BUFX2 BUFX2_insert75 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149_),
    .Y(_1149__bF$buf0)
);

BUFX2 BUFX2_insert74 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149_),
    .Y(_1149__bF$buf1)
);

BUFX2 BUFX2_insert73 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149_),
    .Y(_1149__bF$buf2)
);

BUFX2 BUFX2_insert72 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149_),
    .Y(_1149__bF$buf3)
);

BUFX2 BUFX2_insert71 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149_),
    .Y(_1149__bF$buf4)
);

BUFX2 BUFX2_insert70 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .Y(_886__bF$buf0)
);

BUFX2 BUFX2_insert69 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .Y(_886__bF$buf1)
);

BUFX2 BUFX2_insert68 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .Y(_886__bF$buf2)
);

BUFX2 BUFX2_insert67 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .Y(_886__bF$buf3)
);

BUFX2 BUFX2_insert66 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .Y(_886__bF$buf4)
);

BUFX2 BUFX2_insert65 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .Y(_886__bF$buf5)
);

BUFX2 BUFX2_insert64 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886_),
    .Y(_886__bF$buf6)
);

BUFX2 BUFX2_insert63 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714_),
    .Y(_1714__bF$buf0)
);

BUFX2 BUFX2_insert62 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714_),
    .Y(_1714__bF$buf1)
);

BUFX2 BUFX2_insert61 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714_),
    .Y(_1714__bF$buf2)
);

BUFX2 BUFX2_insert60 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714_),
    .Y(_1714__bF$buf3)
);

BUFX2 BUFX2_insert59 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150_),
    .Y(_1150__bF$buf0)
);

BUFX2 BUFX2_insert58 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150_),
    .Y(_1150__bF$buf1)
);

BUFX2 BUFX2_insert57 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150_),
    .Y(_1150__bF$buf2)
);

BUFX2 BUFX2_insert56 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150_),
    .Y(_1150__bF$buf3)
);

BUFX2 BUFX2_insert55 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150_),
    .Y(_1150__bF$buf4)
);

BUFX2 BUFX2_insert54 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931_),
    .Y(_931__bF$buf0)
);

BUFX2 BUFX2_insert53 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931_),
    .Y(_931__bF$buf1)
);

BUFX2 BUFX2_insert52 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931_),
    .Y(_931__bF$buf2)
);

BUFX2 BUFX2_insert51 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931_),
    .Y(_931__bF$buf3)
);

BUFX2 BUFX2_insert50 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931_),
    .Y(_931__bF$buf4)
);

BUFX2 BUFX2_insert49 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027_),
    .Y(_1027__bF$buf0)
);

BUFX2 BUFX2_insert48 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027_),
    .Y(_1027__bF$buf1)
);

BUFX2 BUFX2_insert47 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027_),
    .Y(_1027__bF$buf2)
);

BUFX2 BUFX2_insert46 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027_),
    .Y(_1027__bF$buf3)
);

BUFX2 BUFX2_insert45 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027_),
    .Y(_1027__bF$buf4)
);

BUFX2 BUFX2_insert44 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902_),
    .Y(_902__bF$buf0)
);

BUFX2 BUFX2_insert43 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902_),
    .Y(_902__bF$buf1)
);

BUFX2 BUFX2_insert42 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902_),
    .Y(_902__bF$buf2)
);

BUFX2 BUFX2_insert41 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902_),
    .Y(_902__bF$buf3)
);

BUFX2 BUFX2_insert40 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .Y(_720__bF$buf0)
);

BUFX2 BUFX2_insert39 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .Y(_720__bF$buf1)
);

BUFX2 BUFX2_insert38 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .Y(_720__bF$buf2)
);

BUFX2 BUFX2_insert37 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .Y(_720__bF$buf3)
);

CLKBUF1 CLKBUF1_insert36 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert35 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert34 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert33 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert32 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert31 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert30 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert29 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert28 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert27 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert26 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf10)
);

BUFX2 BUFX2_insert25 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914_),
    .Y(_914__bF$buf0)
);

BUFX2 BUFX2_insert24 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914_),
    .Y(_914__bF$buf1)
);

BUFX2 BUFX2_insert23 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914_),
    .Y(_914__bF$buf2)
);

BUFX2 BUFX2_insert22 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914_),
    .Y(_914__bF$buf3)
);

BUFX2 BUFX2_insert21 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914_),
    .Y(_914__bF$buf4)
);

BUFX2 BUFX2_insert20 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf4)
);

BUFX2 BUFX2_insert15 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf5)
);

BUFX2 BUFX2_insert14 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf6)
);

BUFX2 BUFX2_insert13 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf7)
);

BUFX2 BUFX2_insert12 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf8)
);

BUFX2 BUFX2_insert11 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf9)
);

BUFX2 BUFX2_insert10 (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1_),
    .Y(_1__bF$buf10)
);

BUFX2 BUFX2_insert9 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf0)
);

BUFX2 BUFX2_insert8 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf3)
);

BUFX2 BUFX2_insert5 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf4)
);

BUFX2 BUFX2_insert4 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf5)
);

BUFX2 BUFX2_insert3 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf6)
);

BUFX2 BUFX2_insert2 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf7)
);

BUFX2 BUFX2_insert1 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf8)
);

BUFX2 BUFX2_insert0 (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY),
    .Y(RDY_bF$buf9)
);

INVX1 _1744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIHOLD[0]),
    .Y(_878_)
);

NAND2X1 _1745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DI[0]),
    .B(RDY_bF$buf9),
    .Y(_879_)
);

OAI21X1 _1746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_878_),
    .C(_879_),
    .Y(DIMUX[0])
);

INVX1 _1747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIHOLD[1]),
    .Y(_880_)
);

NAND2X1 _1748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf7),
    .B(DI[1]),
    .Y(_881_)
);

OAI21X1 _1749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf6),
    .B(_880_),
    .C(_881_),
    .Y(DIMUX[1])
);

INVX1 _1750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIHOLD[2]),
    .Y(_882_)
);

NAND2X1 _1751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf5),
    .B(DI[2]),
    .Y(_883_)
);

OAI21X1 _1752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_882_),
    .C(_883_),
    .Y(DIMUX[2])
);

INVX1 _1753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIHOLD[3]),
    .Y(_884_)
);

NAND2X1 _1754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf3),
    .B(DI[3]),
    .Y(_885_)
);

OAI21X1 _1755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_884_),
    .C(_885_),
    .Y(DIMUX[3])
);

INVX8 _1756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf1),
    .Y(_886_)
);

OR2X2 _1757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf0),
    .B(DIHOLD[4]),
    .Y(_887_)
);

OAI21X1 _1758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf6),
    .B(DI[4]),
    .C(_887_),
    .Y(_888_)
);

INVX1 _1759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_888_),
    .Y(DIMUX[4])
);

INVX1 _1760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIHOLD[5]),
    .Y(_889_)
);

NAND2X1 _1761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf9),
    .B(DI[5]),
    .Y(_890_)
);

OAI21X1 _1762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_889_),
    .C(_890_),
    .Y(DIMUX[5])
);

INVX1 _1763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIHOLD[6]),
    .Y(_891_)
);

NAND2X1 _1764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf7),
    .B(DI[6]),
    .Y(_892_)
);

OAI21X1 _1765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf6),
    .B(_891_),
    .C(_892_),
    .Y(DIMUX[6])
);

MUX2X1 _1766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DI[7]),
    .B(DIHOLD[7]),
    .S(RDY_bF$buf5),
    .Y(_893_)
);

INVX1 _1767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .Y(DIMUX[7])
);

INVX1 _1768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(C),
    .Y(_894_)
);

INVX1 _1769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shift),
    .Y(_895_)
);

INVX1 _1770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[2]),
    .Y(_896_)
);

INVX1 _1771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[3]),
    .Y(_897_)
);

NAND2X1 _1772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_896_),
    .B(_897_),
    .Y(_898_)
);

NAND2X1 _1773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[1]),
    .B(state[0]),
    .Y(_899_)
);

NOR2X1 _1774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_899_),
    .B(_898_),
    .Y(_900_)
);

INVX2 _1775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[4]),
    .Y(_901_)
);

NAND2X1 _1776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .B(_901_),
    .Y(_902_)
);

INVX4 _1777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf3),
    .Y(_903_)
);

NAND2X1 _1778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[2]),
    .B(_897_),
    .Y(_904_)
);

INVX1 _1779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[1]),
    .Y(_905_)
);

INVX1 _1780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[0]),
    .Y(_906_)
);

NAND2X1 _1781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_905_),
    .B(_906_),
    .Y(_907_)
);

NOR2X1 _1782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_904_),
    .B(_907_),
    .Y(_908_)
);

OAI21X1 _1783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_900_),
    .B(_908_),
    .C(_903__bF$buf3),
    .Y(_909_)
);

AND2X2 _1784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[2]),
    .B(state[3]),
    .Y(_910_)
);

NOR2X1 _1785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[1]),
    .B(_906_),
    .Y(_911_)
);

NAND2X1 _1786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_910_),
    .B(_911_),
    .Y(_912_)
);

INVX2 _1787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .Y(_913_)
);

NAND2X1 _1788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_913_),
    .B(_901_),
    .Y(_914_)
);

OAI21X1 _1789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_912_),
    .B(_914__bF$buf4),
    .C(_909_),
    .Y(_915_)
);

NOR2X1 _1790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf3),
    .B(_912_),
    .Y(_916_)
);

INVX1 _1791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_916_),
    .Y(_917_)
);

NOR2X1 _1792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(load_only),
    .B(_917_),
    .Y(_918_)
);

AOI22X1 _1793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(rotate),
    .B(_915_),
    .C(_918_),
    .D(_895_),
    .Y(_919_)
);

INVX1 _1794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(rotate),
    .Y(_920_)
);

INVX1 _1795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(compare),
    .Y(_921_)
);

NAND2X1 _1796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(inc),
    .B(_895_),
    .Y(_922_)
);

OAI22X1 _1797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_909_),
    .B(_922_),
    .C(_921_),
    .D(_917_),
    .Y(_923_)
);

NAND2X1 _1798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[1]),
    .B(_906_),
    .Y(_924_)
);

NOR3X1 _1799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_904_),
    .B(_914__bF$buf2),
    .C(_924_),
    .Y(_925_)
);

NOR2X1 _1800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[3]),
    .B(_896_),
    .Y(_926_)
);

NOR2X1 _1801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[1]),
    .B(state[0]),
    .Y(_927_)
);

NAND2X1 _1802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_927_),
    .B(_926_),
    .Y(_928_)
);

NOR2X1 _1803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .B(state[4]),
    .Y(_929_)
);

NAND2X1 _1804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_900_),
    .Y(_930_)
);

NAND2X1 _1805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[4]),
    .B(_913_),
    .Y(_931_)
);

OAI21X1 _1806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_928_),
    .B(_931__bF$buf4),
    .C(_930_),
    .Y(_932_)
);

OAI21X1 _1807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_925_),
    .B(_932_),
    .C(CO),
    .Y(_933_)
);

NAND2X1 _1808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[3]),
    .B(_896_),
    .Y(_934_)
);

NOR2X1 _1809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_924_),
    .B(_934_),
    .Y(_935_)
);

NAND2X1 _1810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf2),
    .B(_935_),
    .Y(_936_)
);

AND2X2 _1811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[1]),
    .B(state[0]),
    .Y(_937_)
);

NAND2X1 _1812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_937_),
    .B(_910_),
    .Y(_938_)
);

INVX1 _1813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_938_),
    .Y(_939_)
);

NAND2X1 _1814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_939_),
    .Y(_940_)
);

NOR2X1 _1815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_924_),
    .B(_898_),
    .Y(_941_)
);

INVX2 _1816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_941_),
    .Y(_942_)
);

NOR2X1 _1817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf3),
    .B(_942_),
    .Y(_943_)
);

INVX1 _1818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_943_),
    .Y(_944_)
);

NAND3X1 _1819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_940_),
    .B(_936_),
    .C(_944_),
    .Y(_945_)
);

NAND2X1 _1820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_926_),
    .B(_911_),
    .Y(_946_)
);

NOR2X1 _1821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf2),
    .B(_946_),
    .Y(_947_)
);

NOR2X1 _1822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[0]),
    .B(_905_),
    .Y(_948_)
);

NAND2X1 _1823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_910_),
    .B(_948_),
    .Y(_949_)
);

NOR2X1 _1824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf2),
    .B(_949_),
    .Y(_950_)
);

NOR2X1 _1825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_950_),
    .B(_947_),
    .Y(_951_)
);

NOR2X1 _1826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_904_),
    .B(_924_),
    .Y(_952_)
);

NAND2X1 _1827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf1),
    .B(_952_),
    .Y(_953_)
);

NAND3X1 _1828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[2]),
    .B(_897_),
    .C(_937_),
    .Y(_954_)
);

INVX1 _1829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_954_),
    .Y(_955_)
);

NAND2X1 _1830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf0),
    .B(_955_),
    .Y(_956_)
);

NOR2X1 _1831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[2]),
    .B(_897_),
    .Y(_957_)
);

NAND2X1 _1832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_937_),
    .B(_957_),
    .Y(_958_)
);

OAI21X1 _1833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf1),
    .B(_958_),
    .C(_956_),
    .Y(_959_)
);

INVX1 _1834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_959_),
    .Y(_960_)
);

NAND3X1 _1835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_953_),
    .B(_951_),
    .C(_960_),
    .Y(_961_)
);

NOR2X1 _1836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_961_),
    .B(_945_),
    .Y(_962_)
);

NAND2X1 _1837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_933_),
    .B(_962_),
    .Y(_963_)
);

AOI21X1 _1838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_920_),
    .B(_923_),
    .C(_963_),
    .Y(_964_)
);

OAI21X1 _1839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_894_),
    .B(_919_),
    .C(_964_),
    .Y(CI)
);

INVX1 _1840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[0]),
    .Y(_965_)
);

INVX2 _1841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[0]),
    .Y(_966_)
);

NOR2X1 _1842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf1),
    .B(_946_),
    .Y(_967_)
);

INVX2 _1843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_967_),
    .Y(_968_)
);

INVX4 _1844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf1),
    .Y(_969_)
);

NAND2X1 _1845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[2]),
    .B(state[3]),
    .Y(_970_)
);

NOR2X1 _1846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_970_),
    .B(_924_),
    .Y(_971_)
);

NAND2X1 _1847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_971_),
    .Y(_972_)
);

NOR2X1 _1848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[2]),
    .B(state[3]),
    .Y(_973_)
);

NAND2X1 _1849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_973_),
    .B(_911_),
    .Y(_974_)
);

OAI21X1 _1850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf0),
    .B(_974_),
    .C(_972_),
    .Y(_975_)
);

NAND2X1 _1851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[0]),
    .B(_905_),
    .Y(_976_)
);

NOR2X1 _1852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_904_),
    .B(_976_),
    .Y(_977_)
);

NAND2X1 _1853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf3),
    .B(_977_),
    .Y(_978_)
);

OAI21X1 _1854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf0),
    .B(_974_),
    .C(_978_),
    .Y(_979_)
);

NOR2X1 _1855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_975_),
    .B(_979_),
    .Y(_980_)
);

INVX1 _1856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_900_),
    .Y(_981_)
);

NOR2X1 _1857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf3),
    .B(_981_),
    .Y(_982_)
);

NOR2X1 _1858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_967_),
    .B(_982_),
    .Y(_983_)
);

NAND2X1 _1859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_911_),
    .B(_957_),
    .Y(_984_)
);

OAI21X1 _1860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf4),
    .B(_984_),
    .C(_983_),
    .Y(_985_)
);

INVX1 _1861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_985_),
    .Y(_986_)
);

NAND2X1 _1862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_913_),
    .B(_935_),
    .Y(_987_)
);

NOR2X1 _1863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf2),
    .B(_928_),
    .Y(_988_)
);

NAND2X1 _1864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_927_),
    .B(_910_),
    .Y(_989_)
);

NOR2X1 _1865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf0),
    .B(_989_),
    .Y(_990_)
);

NOR2X1 _1866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_990_),
    .B(_988_),
    .Y(_991_)
);

INVX1 _1867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_989_),
    .Y(_992_)
);

NOR2X1 _1868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_934_),
    .B(_907_),
    .Y(_993_)
);

OAI21X1 _1869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_993_),
    .B(_992_),
    .C(_929_),
    .Y(_994_)
);

NAND3X1 _1870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_987_),
    .B(_994_),
    .C(_991_),
    .Y(_995_)
);

NAND2X1 _1871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_952_),
    .Y(_996_)
);

OAI21X1 _1872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_935_),
    .B(_941_),
    .C(_903__bF$buf2),
    .Y(_997_)
);

INVX1 _1873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_940_),
    .Y(_998_)
);

OAI21X1 _1874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf4),
    .B(_958_),
    .C(_960_),
    .Y(_999_)
);

OR2X2 _1875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_999_),
    .B(_998_),
    .Y(_1000_)
);

INVX1 _1876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1000_),
    .Y(_1001_)
);

NAND3X1 _1877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_996_),
    .B(_997_),
    .C(_1001_),
    .Y(_1002_)
);

NOR2X1 _1878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_995_),
    .B(_1002_),
    .Y(_1003_)
);

NAND3X1 _1879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_980_),
    .B(_986_),
    .C(_1003_),
    .Y(_1004_)
);

OAI22X1 _1880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_965_),
    .B(_968_),
    .C(_966_),
    .D(_1004_),
    .Y(BI[0])
);

INVX1 _1881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[1]),
    .Y(_1005_)
);

INVX2 _1882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[1]),
    .Y(_1006_)
);

OAI22X1 _1883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1005_),
    .B(_968_),
    .C(_1006_),
    .D(_1004_),
    .Y(BI[1])
);

INVX2 _1884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[2]),
    .Y(_1007_)
);

INVX1 _1885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[2]),
    .Y(_1008_)
);

OAI22X1 _1886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1007_),
    .B(_968_),
    .C(_1008_),
    .D(_1004_),
    .Y(BI[2])
);

INVX2 _1887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[3]),
    .Y(_1009_)
);

INVX2 _1888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[3]),
    .Y(_1010_)
);

OAI22X1 _1889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1009_),
    .B(_968_),
    .C(_1010_),
    .D(_1004_),
    .Y(BI[3])
);

INVX1 _1890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[4]),
    .Y(_1011_)
);

OAI22X1 _1891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1011_),
    .B(_968_),
    .C(_888_),
    .D(_1004_),
    .Y(BI[4])
);

INVX2 _1892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[5]),
    .Y(_1012_)
);

INVX2 _1893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[5]),
    .Y(_1013_)
);

OAI22X1 _1894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1012_),
    .B(_968_),
    .C(_1013_),
    .D(_1004_),
    .Y(BI[5])
);

INVX2 _1895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[6]),
    .Y(_1014_)
);

INVX2 _1896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[6]),
    .Y(_1015_)
);

OAI22X1 _1897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1014_),
    .B(_968_),
    .C(_1015_),
    .D(_1004_),
    .Y(BI[6])
);

INVX2 _1898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[7]),
    .Y(_1016_)
);

OAI22X1 _1899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1016_),
    .B(_968_),
    .C(_893_),
    .D(_1004_),
    .Y(BI[7])
);

INVX1 _1900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(src_reg[1]),
    .Y(_1017_)
);

NAND2X1 _1901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_935_),
    .Y(_1018_)
);

OAI21X1 _1902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf1),
    .B(_969_),
    .C(_992_),
    .Y(_1019_)
);

NOR2X1 _1903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf3),
    .B(_938_),
    .Y(_1020_)
);

NOR2X1 _1904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf3),
    .B(_958_),
    .Y(_1021_)
);

NOR2X1 _1905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1020_),
    .B(_1021_),
    .Y(_1022_)
);

NAND3X1 _1906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1018_),
    .B(_1019_),
    .C(_1022_),
    .Y(_1023_)
);

NAND2X1 _1907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_993_),
    .Y(_1024_)
);

NAND3X1 _1908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_997_),
    .B(_1024_),
    .C(_951_),
    .Y(_1025_)
);

NOR2X1 _1909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1023_),
    .B(_1025_),
    .Y(_1026_)
);

NAND3X1 _1910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_927_),
    .B(_910_),
    .C(_929_),
    .Y(_1027_)
);

NAND2X1 _1911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_900_),
    .Y(_1028_)
);

OAI21X1 _1912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf2),
    .B(_949_),
    .C(_1028_),
    .Y(_1029_)
);

NOR2X1 _1913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_913_),
    .B(_901_),
    .Y(_1030_)
);

NOR2X1 _1914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_898_),
    .B(_907_),
    .Y(_1031_)
);

NAND2X1 _1915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1030_),
    .B(_1031_),
    .Y(_1032_)
);

OAI21X1 _1916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf1),
    .B(_942_),
    .C(_1032_),
    .Y(_1033_)
);

NOR2X1 _1917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1029_),
    .B(_1033_),
    .Y(_1034_)
);

AND2X2 _1918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1034_),
    .B(_1027__bF$buf4),
    .Y(_1035_)
);

NAND2X1 _1919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1035_),
    .B(_1026_),
    .Y(_1036_)
);

INVX1 _1920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf3),
    .Y(_1037_)
);

INVX1 _1921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1034_),
    .Y(_1038_)
);

AOI21X1 _1922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(dst_reg[1]),
    .B(_1037_),
    .C(_1038_),
    .Y(_1039_)
);

OAI21X1 _1923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1017_),
    .B(_1036_),
    .C(_1039_),
    .Y(_1040_)
);

OAI21X1 _1924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1029_),
    .B(_1033_),
    .C(index_y),
    .Y(_1041_)
);

INVX1 _1925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(dst_reg[0]),
    .Y(_1042_)
);

NOR2X1 _1926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1042_),
    .B(_1027__bF$buf2),
    .Y(_1043_)
);

NOR3X1 _1927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1043_),
    .B(_1023_),
    .C(_1025_),
    .Y(_1044_)
);

AND2X2 _1928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1044_),
    .B(_1041_),
    .Y(_1045_)
);

NAND3X1 _1929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(src_reg[0]),
    .B(_1035_),
    .C(_1026_),
    .Y(_1046_)
);

AOI21X1 _1930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1045_),
    .B(_1046_),
    .C(_1040_),
    .Y(_1047_)
);

NAND3X1 _1931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(src_reg[1]),
    .B(_1035_),
    .C(_1026_),
    .Y(_1048_)
);

AOI22X1 _1932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1048_),
    .B(_1039_),
    .C(_1045_),
    .D(_1046_),
    .Y(_1049_)
);

AOI22X1 _1933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[3] [0]),
    .B(_1049_),
    .C(_1047_),
    .D(\AXYS[1] [0]),
    .Y(_1050_)
);

AND2X2 _1934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1048_),
    .B(_1039_),
    .Y(_1051_)
);

NAND3X1 _1935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1041_),
    .B(_1044_),
    .C(_1036_),
    .Y(_1052_)
);

OAI21X1 _1936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(src_reg[0]),
    .B(_1036_),
    .C(_1052_),
    .Y(_1053_)
);

NAND3X1 _1937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [0]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1054_)
);

INVX1 _1938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(src_reg[0]),
    .Y(_1055_)
);

NAND3X1 _1939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1055_),
    .B(_1035_),
    .C(_1026_),
    .Y(_1056_)
);

AOI22X1 _1940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1048_),
    .B(_1039_),
    .C(_1052_),
    .D(_1056_),
    .Y(_1057_)
);

NAND2X1 _1941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [0]),
    .B(_1057_),
    .Y(_1058_)
);

NAND3X1 _1942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1054_),
    .B(_1058_),
    .C(_1050_),
    .Y(_1059_)
);

INVX1 _1943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1059_),
    .Y(_1060_)
);

AOI21X1 _1944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_941_),
    .C(_988_),
    .Y(_1061_)
);

INVX1 _1945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1061_),
    .Y(_1062_)
);

NOR2X1 _1946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf1),
    .B(_974_),
    .Y(_1063_)
);

NOR2X1 _1947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_990_),
    .B(_1063_),
    .Y(_1064_)
);

NAND2X1 _1948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1064_),
    .B(_951_),
    .Y(_1065_)
);

NOR2X1 _1949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1062_),
    .B(_1065_),
    .Y(_1066_)
);

OAI21X1 _1950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf0),
    .B(_969_),
    .C(_935_),
    .Y(_1067_)
);

INVX1 _1951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1067_),
    .Y(_1068_)
);

INVX2 _1952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_993_),
    .Y(_1069_)
);

OAI21X1 _1953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf0),
    .B(_1069_),
    .C(_1032_),
    .Y(_1070_)
);

NOR2X1 _1954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1068_),
    .B(_1070_),
    .Y(_1071_)
);

NOR2X1 _1955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1029_),
    .B(_918_),
    .Y(_1072_)
);

NAND3X1 _1956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1071_),
    .B(_1072_),
    .C(_1066_),
    .Y(_1073_)
);

INVX2 _1957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1073_),
    .Y(_1074_)
);

NAND2X1 _1958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_948_),
    .B(_957_),
    .Y(_1075_)
);

OAI21X1 _1959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf4),
    .B(_1075_),
    .C(_953_),
    .Y(_1076_)
);

INVX1 _1960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1076_),
    .Y(_1077_)
);

NOR2X1 _1961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_899_),
    .B(_934_),
    .Y(_1078_)
);

NAND2X1 _1962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_1078_),
    .Y(_1079_)
);

OAI21X1 _1963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf3),
    .B(_984_),
    .C(_1079_),
    .Y(_1080_)
);

NOR2X1 _1964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1080_),
    .B(_959_),
    .Y(_1081_)
);

NAND3X1 _1965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_940_),
    .B(_1077_),
    .C(_1081_),
    .Y(_1082_)
);

NAND2X1 _1966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[0]),
    .B(_925_),
    .Y(_1083_)
);

OAI21X1 _1967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_966_),
    .B(_983_),
    .C(_1083_),
    .Y(_1084_)
);

AOI21X1 _1968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(ADD[0]),
    .C(_1084_),
    .Y(_1085_)
);

OAI21X1 _1969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1060_),
    .C(_1085_),
    .Y(AI[0])
);

NAND2X1 _1970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[1] [1]),
    .B(_1047_),
    .Y(_1086_)
);

AOI22X1 _1971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .B(\AXYS[3] [1]),
    .C(\AXYS[2] [1]),
    .D(_1057_),
    .Y(_1087_)
);

NAND3X1 _1972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [1]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1088_)
);

NAND3X1 _1973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1088_),
    .B(_1086_),
    .C(_1087_),
    .Y(_1089_)
);

INVX1 _1974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1089_),
    .Y(_1090_)
);

INVX1 _1975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[1]),
    .Y(_1091_)
);

NAND2X1 _1976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_952_),
    .Y(_1092_)
);

NOR2X1 _1977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1091_),
    .B(_1092_),
    .Y(_1093_)
);

INVX1 _1978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1093_),
    .Y(_1094_)
);

OAI21X1 _1979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1006_),
    .B(_983_),
    .C(_1094_),
    .Y(_1095_)
);

AOI21X1 _1980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(ADD[1]),
    .C(_1095_),
    .Y(_1096_)
);

OAI21X1 _1981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1090_),
    .C(_1096_),
    .Y(AI[1])
);

NAND2X1 _1982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[1] [2]),
    .B(_1047_),
    .Y(_1097_)
);

AOI22X1 _1983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .B(\AXYS[3] [2]),
    .C(\AXYS[2] [2]),
    .D(_1057_),
    .Y(_1098_)
);

NAND3X1 _1984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [2]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1099_)
);

NAND3X1 _1985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1099_),
    .B(_1097_),
    .C(_1098_),
    .Y(_1100_)
);

INVX1 _1986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1100_),
    .Y(_1101_)
);

INVX1 _1987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[2]),
    .Y(_1102_)
);

OAI22X1 _1988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1102_),
    .B(_1092_),
    .C(_1008_),
    .D(_983_),
    .Y(_1103_)
);

AOI21X1 _1989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(ADD[2]),
    .C(_1103_),
    .Y(_1104_)
);

OAI21X1 _1990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1101_),
    .C(_1104_),
    .Y(AI[2])
);

NAND2X1 _1991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[1] [3]),
    .B(_1047_),
    .Y(_1105_)
);

AOI22X1 _1992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .B(\AXYS[3] [3]),
    .C(\AXYS[2] [3]),
    .D(_1057_),
    .Y(_1106_)
);

NAND3X1 _1993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [3]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1107_)
);

NAND3X1 _1994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1107_),
    .B(_1105_),
    .C(_1106_),
    .Y(_1108_)
);

INVX1 _1995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1108_),
    .Y(_1109_)
);

NAND2X1 _1996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[3]),
    .B(_925_),
    .Y(_1110_)
);

OAI21X1 _1997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1010_),
    .B(_983_),
    .C(_1110_),
    .Y(_1111_)
);

AOI21X1 _1998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(ADD[3]),
    .C(_1111_),
    .Y(_1112_)
);

OAI21X1 _1999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1109_),
    .C(_1112_),
    .Y(AI[3])
);

NAND2X1 _2000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[1] [4]),
    .B(_1047_),
    .Y(_1113_)
);

AOI22X1 _2001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .B(\AXYS[3] [4]),
    .C(\AXYS[2] [4]),
    .D(_1057_),
    .Y(_1114_)
);

NAND3X1 _2002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [4]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1115_)
);

NAND3X1 _2003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1115_),
    .B(_1113_),
    .C(_1114_),
    .Y(_1116_)
);

INVX1 _2004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1116_),
    .Y(_1117_)
);

NAND2X1 _2005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[4]),
    .B(_925_),
    .Y(_1118_)
);

OAI21X1 _2006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_888_),
    .B(_983_),
    .C(_1118_),
    .Y(_1119_)
);

AOI21X1 _2007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(ADD[4]),
    .C(_1119_),
    .Y(_1120_)
);

OAI21X1 _2008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1117_),
    .C(_1120_),
    .Y(AI[4])
);

NAND2X1 _2009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[1] [5]),
    .B(_1047_),
    .Y(_1121_)
);

AOI22X1 _2010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .B(\AXYS[3] [5]),
    .C(\AXYS[2] [5]),
    .D(_1057_),
    .Y(_1122_)
);

NAND3X1 _2011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [5]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1123_)
);

NAND3X1 _2012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1123_),
    .B(_1121_),
    .C(_1122_),
    .Y(_1124_)
);

INVX1 _2013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1124_),
    .Y(_1125_)
);

NAND2X1 _2014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[5]),
    .B(_925_),
    .Y(_1126_)
);

OAI21X1 _2015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1013_),
    .B(_983_),
    .C(_1126_),
    .Y(_1127_)
);

AOI21X1 _2016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(ADD[5]),
    .C(_1127_),
    .Y(_1128_)
);

OAI21X1 _2017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1125_),
    .C(_1128_),
    .Y(AI[5])
);

NAND2X1 _2018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[1] [6]),
    .B(_1047_),
    .Y(_1129_)
);

AOI22X1 _2019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .B(\AXYS[3] [6]),
    .C(\AXYS[2] [6]),
    .D(_1057_),
    .Y(_1130_)
);

NAND3X1 _2020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [6]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1131_)
);

NAND3X1 _2021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1131_),
    .B(_1129_),
    .C(_1130_),
    .Y(_1132_)
);

INVX1 _2022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1132_),
    .Y(_1133_)
);

INVX1 _2023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[6]),
    .Y(_1134_)
);

NOR2X1 _2024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1134_),
    .B(_1092_),
    .Y(_1135_)
);

INVX1 _2025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1135_),
    .Y(_1136_)
);

OAI21X1 _2026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1015_),
    .B(_983_),
    .C(_1136_),
    .Y(_1137_)
);

AOI21X1 _2027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(ADD[6]),
    .C(_1137_),
    .Y(_1138_)
);

OAI21X1 _2028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1133_),
    .C(_1138_),
    .Y(AI[6])
);

NAND2X1 _2029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[1] [7]),
    .B(_1047_),
    .Y(_1139_)
);

AOI22X1 _2030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .B(\AXYS[3] [7]),
    .C(\AXYS[2] [7]),
    .D(_1057_),
    .Y(_1140_)
);

NAND3X1 _2031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [7]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1141_)
);

NAND3X1 _2032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1141_),
    .B(_1139_),
    .C(_1140_),
    .Y(_1142_)
);

INVX1 _2033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1142_),
    .Y(_1143_)
);

INVX1 _2034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[7]),
    .Y(_1144_)
);

NOR2X1 _2035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1144_),
    .B(_1092_),
    .Y(_1145_)
);

INVX1 _2036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1145_),
    .Y(_1146_)
);

OAI21X1 _2037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .B(_983_),
    .C(_1146_),
    .Y(_1147_)
);

AOI21X1 _2038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1082_),
    .B(AN),
    .C(_1147_),
    .Y(_1148_)
);

OAI21X1 _2039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1074_),
    .B(_1143_),
    .C(_1148_),
    .Y(AI[7])
);

NAND2X1 _2040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_1037_),
    .Y(_1149_)
);

INVX8 _2041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf4),
    .Y(_1150_)
);

INVX1 _2042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD[1]),
    .Y(_1151_)
);

INVX1 _2043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRQ),
    .Y(_1152_)
);

INVX1 _2044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(NMI_edge),
    .Y(_1153_)
);

OAI21X1 _2045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(I),
    .B(_1152_),
    .C(_1153_),
    .Y(_1154_)
);

AOI21X1 _2046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(_1151_),
    .C(_1154_),
    .Y(_1155_)
);

OAI21X1 _2047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(DIMUX[1]),
    .C(_1155_),
    .Y(_1156_)
);

INVX1 _2048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD[0]),
    .Y(_1157_)
);

AOI21X1 _2049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1157_),
    .B(IRHOLD_valid),
    .C(_1154_),
    .Y(_1158_)
);

OAI21X1 _2050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(DIMUX[0]),
    .C(_1158_),
    .Y(_1159_)
);

NAND2X1 _2051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1156_),
    .B(_1159_),
    .Y(_1160_)
);

INVX1 _2052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1160_),
    .Y(_1161_)
);

INVX1 _2053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD[3]),
    .Y(_1162_)
);

AOI21X1 _2054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(_1162_),
    .C(_1154_),
    .Y(_1163_)
);

OAI21X1 _2055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(DIMUX[3]),
    .C(_1163_),
    .Y(_1164_)
);

INVX1 _2056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(I),
    .Y(_1165_)
);

NAND2X1 _2057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1152_),
    .B(_1153_),
    .Y(_1166_)
);

OAI21X1 _2058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1165_),
    .B(NMI_edge),
    .C(_1166_),
    .Y(_1167_)
);

INVX2 _2059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .Y(_1168_)
);

INVX1 _2060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD[2]),
    .Y(_1169_)
);

NAND2X1 _2061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1168_),
    .B(DIMUX[2]),
    .Y(_1170_)
);

OAI21X1 _2062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1168_),
    .B(_1169_),
    .C(_1170_),
    .Y(_1171_)
);

NAND2X1 _2063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1167_),
    .B(_1171_),
    .Y(_1172_)
);

NAND2X1 _2064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1164_),
    .B(_1172_),
    .Y(_1173_)
);

INVX1 _2065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1173_),
    .Y(_1174_)
);

NAND2X1 _2066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1161_),
    .B(_1174_),
    .Y(_1175_)
);

NAND2X1 _2067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(IRHOLD[4]),
    .Y(_1176_)
);

OAI21X1 _2068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(_888_),
    .C(_1176_),
    .Y(_1177_)
);

NAND2X1 _2069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1167_),
    .B(_1177_),
    .Y(_1178_)
);

INVX2 _2070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1178_),
    .Y(_1179_)
);

OAI21X1 _2071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1168_),
    .B(IRHOLD[5]),
    .C(_1167_),
    .Y(_1180_)
);

AOI21X1 _2072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1168_),
    .B(_1013_),
    .C(_1180_),
    .Y(_1181_)
);

NOR2X1 _2073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_1179_),
    .Y(_1182_)
);

NAND2X1 _2074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(IRHOLD[7]),
    .Y(_1183_)
);

OAI21X1 _2075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(IRHOLD_valid),
    .B(_893_),
    .C(_1183_),
    .Y(_1184_)
);

NAND2X1 _2076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1167_),
    .B(_1184_),
    .Y(_1185_)
);

MUX2X1 _2077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[6]),
    .B(IRHOLD[6]),
    .S(_1168_),
    .Y(_1186_)
);

NOR2X1 _2078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1154_),
    .B(_1186_),
    .Y(_1187_)
);

NAND2X1 _2079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .B(_1187_),
    .Y(_1188_)
);

INVX1 _2080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1188_),
    .Y(_1189_)
);

NAND2X1 _2081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1189_),
    .B(_1182_),
    .Y(_1190_)
);

NOR2X1 _2082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1175_),
    .B(_1190_),
    .Y(_1191_)
);

AOI22X1 _2083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf5),
    .B(_947_),
    .C(_1191_),
    .D(_1150__bF$buf4),
    .Y(_1192_)
);

NOR2X1 _2084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf2),
    .B(_928_),
    .Y(_1193_)
);

OAI21X1 _2085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(store),
    .C(_1193_),
    .Y(_1194_)
);

NAND2X1 _2086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf3),
    .B(_1194_),
    .Y(_1195_)
);

NOR2X1 _2087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf1),
    .B(_946_),
    .Y(_1196_)
);

OAI21X1 _2088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_1196_),
    .C(_1195_),
    .Y(_1197_)
);

NAND2X1 _2089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1197_),
    .B(_1192_),
    .Y(_1198_)
);

NOR2X1 _2090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_974_),
    .Y(_1199_)
);

INVX1 _2091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1199_),
    .Y(_1200_)
);

NOR2X1 _2092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf0),
    .B(_938_),
    .Y(_1201_)
);

NAND2X1 _2093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_908_),
    .Y(_1202_)
);

OAI21X1 _2094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf2),
    .B(_974_),
    .C(_1202_),
    .Y(_1203_)
);

NOR2X1 _2095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1201_),
    .B(_1203_),
    .Y(_1204_)
);

OAI21X1 _2096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_913_),
    .B(_1200_),
    .C(_1204_),
    .Y(_1205_)
);

INVX1 _2097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1205_),
    .Y(_1206_)
);

INVX1 _2098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(write_back),
    .Y(_1207_)
);

NAND2X1 _2099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf1),
    .B(_1207_),
    .Y(_1208_)
);

NOR2X1 _2100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1208_),
    .B(_1206_),
    .Y(_1209_)
);

INVX1 _2101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1209_),
    .Y(_1210_)
);

OAI21X1 _2102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1168_),
    .B(IRHOLD[3]),
    .C(_1167_),
    .Y(_1211_)
);

AOI21X1 _2103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1168_),
    .B(_1010_),
    .C(_1211_),
    .Y(_1212_)
);

NAND2X1 _2104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1172_),
    .B(_1212_),
    .Y(_1213_)
);

INVX1 _2105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1159_),
    .Y(_1214_)
);

NAND2X1 _2106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1156_),
    .B(_1214_),
    .Y(_1215_)
);

NAND2X1 _2107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1159_),
    .B(_1164_),
    .Y(_1216_)
);

INVX2 _2108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .Y(_1217_)
);

NAND2X1 _2109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1172_),
    .B(_1217_),
    .Y(_1218_)
);

OAI22X1 _2110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1216_),
    .B(_1218_),
    .C(_1213_),
    .D(_1215_),
    .Y(_1219_)
);

NAND3X1 _2111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf3),
    .B(_1178_),
    .C(_1219_),
    .Y(_1220_)
);

NOR2X1 _2112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_970_),
    .B(_976_),
    .Y(_1221_)
);

NAND2X1 _2113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_1221_),
    .Y(_1222_)
);

OAI21X1 _2114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf3),
    .B(_912_),
    .C(_1222_),
    .Y(_1223_)
);

INVX1 _2115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1196_),
    .Y(_1224_)
);

INVX1 _2116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_974_),
    .Y(_1225_)
);

NAND2X1 _2117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_1225_),
    .Y(_1226_)
);

NAND2X1 _2118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf3),
    .B(_971_),
    .Y(_1227_)
);

NAND3X1 _2119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1227_),
    .B(_1224_),
    .C(_1226_),
    .Y(_1228_)
);

NOR2X1 _2120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1223_),
    .B(_1228_),
    .Y(_1229_)
);

INVX1 _2121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1229_),
    .Y(_1230_)
);

NOR2X1 _2122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf4),
    .B(_1205_),
    .Y(_1231_)
);

NAND2X1 _2123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf3),
    .B(_916_),
    .Y(_1232_)
);

NOR2X1 _2124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf2),
    .B(_989_),
    .Y(_1233_)
);

INVX1 _2125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1233_),
    .Y(_1234_)
);

NOR2X1 _2126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf1),
    .B(_912_),
    .Y(_1235_)
);

NAND2X1 _2127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf2),
    .B(_1235_),
    .Y(_1236_)
);

OAI21X1 _2128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf1),
    .B(_1234_),
    .C(_1236_),
    .Y(_1237_)
);

NAND2X1 _2129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf0),
    .B(_990_),
    .Y(_1238_)
);

OAI21X1 _2130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf9),
    .B(_1222_),
    .C(_1238_),
    .Y(_1239_)
);

NOR2X1 _2131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1239_),
    .B(_1237_),
    .Y(_1240_)
);

OR2X2 _2132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(store),
    .Y(_1241_)
);

NOR2X1 _2133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(write_back),
    .B(_1241_),
    .Y(_1242_)
);

NOR2X1 _2134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf0),
    .B(_930_),
    .Y(_1243_)
);

NOR2X1 _2135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf6),
    .B(_1241_),
    .Y(_1244_)
);

AOI22X1 _2136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1193_),
    .B(_1244_),
    .C(_1243_),
    .D(_1242_),
    .Y(_1245_)
);

NAND3X1 _2137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1232_),
    .B(_1245_),
    .C(_1240_),
    .Y(_1246_)
);

AOI21X1 _2138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1231_),
    .B(_1230_),
    .C(_1246_),
    .Y(_1247_)
);

NAND3X1 _2139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1220_),
    .B(_1247_),
    .C(_1210_),
    .Y(_1248_)
);

OR2X2 _2140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1198_),
    .B(_1248_),
    .Y(_1249_)
);

INVX1 _2141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1249_),
    .Y(_1250_)
);

NOR2X1 _2142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1160_),
    .B(_1213_),
    .Y(_1251_)
);

NAND3X1 _2143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1182_),
    .B(_1185_),
    .C(_1251_),
    .Y(_1252_)
);

INVX1 _2144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1252_),
    .Y(_1253_)
);

AOI22X1 _2145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf5),
    .B(_1063_),
    .C(_1253_),
    .D(_1150__bF$buf2),
    .Y(_1254_)
);

NOR2X1 _2146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1178_),
    .B(_1175_),
    .Y(_1255_)
);

AOI22X1 _2147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf4),
    .B(_967_),
    .C(_1255_),
    .D(_1150__bF$buf1),
    .Y(_1256_)
);

NOR2X1 _2148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf0),
    .B(_1069_),
    .Y(_1257_)
);

OAI21X1 _2149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf3),
    .B(_984_),
    .C(_886__bF$buf3),
    .Y(_1258_)
);

OAI21X1 _2150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf2),
    .B(_1257_),
    .C(_1258_),
    .Y(_1259_)
);

NOR2X1 _2151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf0),
    .B(_1069_),
    .Y(_1260_)
);

OAI21X1 _2152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf4),
    .B(_984_),
    .C(_886__bF$buf1),
    .Y(_1261_)
);

OAI21X1 _2153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf0),
    .B(_1260_),
    .C(_1261_),
    .Y(_1262_)
);

NOR2X1 _2154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf1),
    .B(_1069_),
    .Y(_1263_)
);

OAI21X1 _2155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf0),
    .B(_984_),
    .C(_886__bF$buf6),
    .Y(_1264_)
);

OAI21X1 _2156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf5),
    .B(_1263_),
    .C(_1264_),
    .Y(_1265_)
);

NAND3X1 _2157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1262_),
    .B(_1265_),
    .C(_1259_),
    .Y(_1266_)
);

NAND2X1 _2158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1030_),
    .B(_1225_),
    .Y(_1267_)
);

INVX1 _2159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1032_),
    .Y(_1268_)
);

NAND2X1 _2160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_1268_),
    .Y(_1269_)
);

OAI21X1 _2161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf7),
    .B(_1267_),
    .C(_1269_),
    .Y(_1270_)
);

OAI21X1 _2162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf3),
    .B(_974_),
    .C(_886__bF$buf4),
    .Y(_1271_)
);

INVX2 _2163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1031_),
    .Y(_1272_)
);

OAI21X1 _2164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf2),
    .B(_1272_),
    .C(RDY_bF$buf6),
    .Y(_1273_)
);

AOI21X1 _2165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1271_),
    .B(_1273_),
    .C(_1270_),
    .Y(_1274_)
);

NOR2X1 _2166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf4),
    .B(_974_),
    .Y(_1275_)
);

OAI21X1 _2167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf3),
    .B(_1272_),
    .C(RDY_bF$buf5),
    .Y(_1276_)
);

OAI21X1 _2168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_1275_),
    .C(_1276_),
    .Y(_1277_)
);

NAND2X1 _2169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1277_),
    .B(_1274_),
    .Y(_1278_)
);

NOR2X1 _2170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1266_),
    .B(_1278_),
    .Y(_1279_)
);

NAND3X1 _2171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1256_),
    .B(_1279_),
    .C(_1254_),
    .Y(_1280_)
);

OAI21X1 _2172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1207_),
    .B(_1206_),
    .C(RDY_bF$buf3),
    .Y(_1281_)
);

OAI21X1 _2173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_982_),
    .C(_1281_),
    .Y(_1282_)
);

NOR2X1 _2174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1172_),
    .B(_1212_),
    .Y(_1283_)
);

NOR2X1 _2175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf3),
    .B(_1179_),
    .Y(_1284_)
);

AOI22X1 _2176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf3),
    .B(_1201_),
    .C(_1284_),
    .D(_1283_),
    .Y(_1285_)
);

OAI21X1 _2177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf2),
    .B(_949_),
    .C(RDY_bF$buf1),
    .Y(_1286_)
);

OAI21X1 _2178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf0),
    .B(_998_),
    .C(_1286_),
    .Y(_1287_)
);

NAND2X1 _2179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1287_),
    .B(_1285_),
    .Y(_1288_)
);

MUX2X1 _2180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_956_),
    .B(_953_),
    .S(_886__bF$buf2),
    .Y(_1289_)
);

NAND2X1 _2181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_969_),
    .B(_952_),
    .Y(_1290_)
);

NOR2X1 _2182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf1),
    .B(_954_),
    .Y(_1291_)
);

NAND2X1 _2183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf1),
    .B(_1291_),
    .Y(_1292_)
);

OAI21X1 _2184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf0),
    .B(_1290_),
    .C(_1292_),
    .Y(_1293_)
);

NOR2X1 _2185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1289_),
    .B(_1293_),
    .Y(_1294_)
);

NAND2X1 _2186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(backwards),
    .Y(_1295_)
);

OR2X2 _2187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(backwards),
    .Y(_1296_)
);

NAND2X1 _2188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1295_),
    .B(_1296_),
    .Y(_1297_)
);

OAI21X1 _2189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1297_),
    .B(_1092_),
    .C(RDY_bF$buf9),
    .Y(_1298_)
);

NOR2X1 _2190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf1),
    .B(_954_),
    .Y(_1299_)
);

OAI21X1 _2191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_1299_),
    .C(_1298_),
    .Y(_1300_)
);

NAND2X1 _2192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1300_),
    .B(_1294_),
    .Y(_1301_)
);

NOR2X1 _2193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1301_),
    .B(_1288_),
    .Y(_1302_)
);

NAND2X1 _2194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_941_),
    .Y(_1303_)
);

INVX1 _2195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1303_),
    .Y(_1304_)
);

OAI21X1 _2196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf0),
    .B(_981_),
    .C(_886__bF$buf6),
    .Y(_1305_)
);

OAI21X1 _2197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf5),
    .B(_1304_),
    .C(_1305_),
    .Y(_1306_)
);

OAI21X1 _2198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf0),
    .B(_949_),
    .C(RDY_bF$buf7),
    .Y(_1307_)
);

OAI21X1 _2199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf6),
    .B(_1020_),
    .C(_1307_),
    .Y(_1308_)
);

INVX1 _2200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1028_),
    .Y(_1309_)
);

OAI21X1 _2201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf4),
    .B(_942_),
    .C(RDY_bF$buf5),
    .Y(_1310_)
);

OAI21X1 _2202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_1309_),
    .C(_1310_),
    .Y(_1311_)
);

NAND3X1 _2203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1308_),
    .B(_1306_),
    .C(_1311_),
    .Y(_1312_)
);

OAI21X1 _2204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf4),
    .B(_1075_),
    .C(RDY_bF$buf3),
    .Y(_1313_)
);

OAI21X1 _2205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_1021_),
    .C(_1313_),
    .Y(_1314_)
);

OAI21X1 _2206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf2),
    .B(_1075_),
    .C(RDY_bF$buf1),
    .Y(_1315_)
);

OAI21X1 _2207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf1),
    .B(_958_),
    .C(_886__bF$buf4),
    .Y(_1316_)
);

AND2X2 _2208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1315_),
    .B(_1316_),
    .Y(_1317_)
);

INVX1 _2209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1317_),
    .Y(_1318_)
);

INVX4 _2210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1018_),
    .Y(_1319_)
);

OAI21X1 _2211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf3),
    .B(_958_),
    .C(_886__bF$buf3),
    .Y(_1320_)
);

OAI21X1 _2212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf2),
    .B(_1319__bF$buf3),
    .C(_1320_),
    .Y(_1321_)
);

NAND3X1 _2213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1314_),
    .B(_1321_),
    .C(_1318_),
    .Y(_1322_)
);

NOR2X1 _2214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1312_),
    .B(_1322_),
    .Y(_1323_)
);

NAND3X1 _2215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1323_),
    .B(_1282_),
    .C(_1302_),
    .Y(_1324_)
);

NOR2X1 _2216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1280_),
    .B(_1324_),
    .Y(_1325_)
);

NAND2X1 _2217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1325_),
    .B(_1250_),
    .Y(_1512_[0])
);

NOR2X1 _2218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1213_),
    .B(_1215_),
    .Y(_1326_)
);

AND2X2 _2219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1171_),
    .B(_1167_),
    .Y(_1327_)
);

NAND2X1 _2220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1212_),
    .B(_1327_),
    .Y(_1328_)
);

INVX1 _2221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1328_),
    .Y(_1329_)
);

NOR2X1 _2222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf2),
    .B(_1178_),
    .Y(_1330_)
);

OAI21X1 _2223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1329_),
    .B(_1326_),
    .C(_1330_),
    .Y(_1331_)
);

NOR2X1 _2224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1173_),
    .B(_1215_),
    .Y(_1332_)
);

AOI22X1 _2225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf1),
    .B(_943_),
    .C(_1332_),
    .D(_1330_),
    .Y(_1333_)
);

NOR2X1 _2226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf3),
    .B(_1075_),
    .Y(_1334_)
);

OAI21X1 _2227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf2),
    .B(_984_),
    .C(RDY_bF$buf0),
    .Y(_1335_)
);

OAI21X1 _2228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf9),
    .B(_1334_),
    .C(_1335_),
    .Y(_1336_)
);

NAND2X1 _2229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf2),
    .B(_941_),
    .Y(_1337_)
);

NAND2X1 _2230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_1063_),
    .Y(_1338_)
);

OAI21X1 _2231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf7),
    .B(_1337_),
    .C(_1338_),
    .Y(_1339_)
);

AOI21X1 _2232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf0),
    .B(_1304_),
    .C(_1339_),
    .Y(_1340_)
);

AND2X2 _2233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1340_),
    .B(_1336_),
    .Y(_1341_)
);

NAND3X1 _2234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1331_),
    .B(_1333_),
    .C(_1341_),
    .Y(_1342_)
);

INVX1 _2235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1342_),
    .Y(_1343_)
);

NAND2X1 _2236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_1078_),
    .Y(_1344_)
);

OAI21X1 _2237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf2),
    .B(_984_),
    .C(_1344_),
    .Y(_1345_)
);

NAND3X1 _2238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1229_),
    .B(_1345_),
    .C(_1231_),
    .Y(_1346_)
);

OR2X2 _2239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1290_),
    .B(RDY_bF$buf6),
    .Y(_1347_)
);

INVX1 _2240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .Y(_1348_)
);

NAND2X1 _2241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1178_),
    .B(_1348_),
    .Y(_1349_)
);

NOR2X1 _2242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1188_),
    .B(_1349_),
    .Y(_1350_)
);

NOR2X1 _2243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1160_),
    .B(_1328_),
    .Y(_1351_)
);

NAND3X1 _2244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf0),
    .B(_1351_),
    .C(_1350_),
    .Y(_1352_)
);

NAND3X1 _2245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1347_),
    .B(_1352_),
    .C(_1346_),
    .Y(_1353_)
);

INVX1 _2246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1353_),
    .Y(_1354_)
);

NAND2X1 _2247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1178_),
    .B(_1181_),
    .Y(_1355_)
);

NOR2X1 _2248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1217_),
    .B(_1355_),
    .Y(_1356_)
);

NAND2X1 _2249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1356_),
    .B(_1251_),
    .Y(_1357_)
);

OAI22X1 _2250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf5),
    .B(_972_),
    .C(_1149__bF$buf1),
    .D(_1357_),
    .Y(_1358_)
);

NAND2X1 _2251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_982_),
    .Y(_1359_)
);

NOR2X1 _2252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[4]),
    .B(_949_),
    .Y(_1360_)
);

NAND2X1 _2253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf6),
    .B(_1360_),
    .Y(_1361_)
);

NAND2X1 _2254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1284_),
    .B(_1332_),
    .Y(_1362_)
);

NAND3X1 _2255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1359_),
    .B(_1361_),
    .C(_1362_),
    .Y(_1363_)
);

NOR2X1 _2256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1363_),
    .B(_1358_),
    .Y(_1364_)
);

NOR2X1 _2257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1160_),
    .B(_1173_),
    .Y(_1365_)
);

OAI21X1 _2258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1154_),
    .B(_1186_),
    .C(_1185_),
    .Y(_1366_)
);

NOR2X1 _2259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1366_),
    .B(_1355_),
    .Y(_1367_)
);

NAND3X1 _2260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf4),
    .B(_1365_),
    .C(_1367_),
    .Y(_1368_)
);

OAI21X1 _2261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf3),
    .B(_1018_),
    .C(_1368_),
    .Y(_1369_)
);

NOR2X1 _2262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1188_),
    .B(_1355_),
    .Y(_1370_)
);

NAND3X1 _2263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf3),
    .B(_1365_),
    .C(_1370_),
    .Y(_1371_)
);

OAI21X1 _2264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_936_),
    .C(_1371_),
    .Y(_1372_)
);

INVX1 _2265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(cond_code[0]),
    .Y(_1373_)
);

INVX1 _2266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(V),
    .Y(_1374_)
);

NAND2X1 _2267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(cond_code[2]),
    .B(Z),
    .Y(_1375_)
);

OAI21X1 _2268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(cond_code[2]),
    .B(_1374_),
    .C(_1375_),
    .Y(_1376_)
);

INVX1 _2269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(N),
    .Y(_1377_)
);

NAND2X1 _2270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(C),
    .B(cond_code[2]),
    .Y(_1378_)
);

OAI21X1 _2271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(cond_code[2]),
    .B(_1377_),
    .C(_1378_),
    .Y(_1379_)
);

MUX2X1 _2272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1376_),
    .B(_1379_),
    .S(cond_code[1]),
    .Y(_1380_)
);

OR2X2 _2273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1380_),
    .B(_1373_),
    .Y(_1381_)
);

NAND2X1 _2274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1373_),
    .B(_1380_),
    .Y(_1382_)
);

NAND2X1 _2275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1382_),
    .B(_1381_),
    .Y(_1383_)
);

NOR2X1 _2276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf5),
    .B(_968_),
    .Y(_1384_)
);

NOR2X1 _2277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf4),
    .B(_978_),
    .Y(_1385_)
);

INVX1 _2278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1385_),
    .Y(_1386_)
);

OAI21X1 _2279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf1),
    .B(_953_),
    .C(_1386_),
    .Y(_1387_)
);

AOI21X1 _2280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1383_),
    .B(_1384_),
    .C(_1387_),
    .Y(_1388_)
);

OAI21X1 _2281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf0),
    .B(_1092_),
    .C(_1388_),
    .Y(_1389_)
);

NOR3X1 _2282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1369_),
    .B(_1372_),
    .C(_1389_),
    .Y(_1390_)
);

NAND3X1 _2283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1364_),
    .B(_1390_),
    .C(_1354_),
    .Y(_1391_)
);

NOR2X1 _2284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1324_),
    .B(_1391_),
    .Y(_1392_)
);

NAND2X1 _2285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1343_),
    .B(_1392_),
    .Y(_1512_[1])
);

OAI21X1 _2286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1184_),
    .B(_1177_),
    .C(_1167_),
    .Y(_1393_)
);

INVX1 _2287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1393_),
    .Y(_1394_)
);

NOR2X1 _2288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1156_),
    .B(_1214_),
    .Y(_1395_)
);

INVX1 _2289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1395_),
    .Y(_1396_)
);

NOR2X1 _2290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1213_),
    .B(_1396_),
    .Y(_1397_)
);

AOI21X1 _2291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1394_),
    .B(_1251_),
    .C(_1397_),
    .Y(_1398_)
);

OAI21X1 _2292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1213_),
    .B(_1215_),
    .C(_1328_),
    .Y(_1399_)
);

MUX2X1 _2293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1219_),
    .B(_1399_),
    .S(_1178_),
    .Y(_1400_)
);

NAND2X1 _2294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1400_),
    .B(_1398_),
    .Y(_1401_)
);

NOR2X1 _2295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .B(_1179_),
    .Y(_1402_)
);

OAI21X1 _2296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1367_),
    .B(_1402_),
    .C(_1351_),
    .Y(_1403_)
);

INVX1 _2297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1156_),
    .Y(_1404_)
);

NOR2X1 _2298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1159_),
    .B(_1404_),
    .Y(_1405_)
);

NOR2X1 _2299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1179_),
    .B(_1328_),
    .Y(_1406_)
);

OAI21X1 _2300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1405_),
    .B(_1395_),
    .C(_1406_),
    .Y(_1407_)
);

AND2X2 _2301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1403_),
    .B(_1407_),
    .Y(_1408_)
);

INVX1 _2302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1351_),
    .Y(_1409_)
);

OAI21X1 _2303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1190_),
    .B(_1409_),
    .C(_1252_),
    .Y(_1410_)
);

NAND2X1 _2304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1370_),
    .B(_1351_),
    .Y(_1411_)
);

INVX2 _2305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1187_),
    .Y(_1412_)
);

OAI21X1 _2306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_1412_),
    .C(_1393_),
    .Y(_1413_)
);

OAI21X1 _2307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1175_),
    .B(_1413_),
    .C(_1411_),
    .Y(_1414_)
);

NOR2X1 _2308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1414_),
    .B(_1410_),
    .Y(_1415_)
);

NAND2X1 _2309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1365_),
    .B(_1350_),
    .Y(_1416_)
);

OAI21X1 _2310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1172_),
    .B(_1212_),
    .C(_1150__bF$buf2),
    .Y(_1417_)
);

NOR2X1 _2311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1417_),
    .B(_1332_),
    .Y(_1418_)
);

AND2X2 _2312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1416_),
    .B(_1418_),
    .Y(_1419_)
);

AOI21X1 _2313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1251_),
    .B(_1356_),
    .C(_1255_),
    .Y(_1420_)
);

AND2X2 _2314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1419_),
    .B(_1420_),
    .Y(_1421_)
);

NAND3X1 _2315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1408_),
    .B(_1415_),
    .C(_1421_),
    .Y(_1422_)
);

AND2X2 _2316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1231_),
    .B(_1229_),
    .Y(_1423_)
);

NOR2X1 _2317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .B(_954_),
    .Y(_1424_)
);

NOR2X1 _2318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1424_),
    .B(_916_),
    .Y(_1425_)
);

OAI21X1 _2319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_908_),
    .B(_1031_),
    .C(_903__bF$buf1),
    .Y(_1426_)
);

NOR2X1 _2320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_976_),
    .B(_934_),
    .Y(_1427_)
);

OAI21X1 _2321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_941_),
    .B(_1427_),
    .C(_903__bF$buf0),
    .Y(_1428_)
);

NAND3X1 _2322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1426_),
    .B(_1428_),
    .C(_1425_),
    .Y(_1429_)
);

INVX1 _2323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1384_),
    .Y(_1430_)
);

NOR2X1 _2324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1383_),
    .B(_1430_),
    .Y(_1431_)
);

NAND2X1 _2325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1297_),
    .B(_925_),
    .Y(_1432_)
);

NAND2X1 _2326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf3),
    .B(_990_),
    .Y(_1433_)
);

OAI21X1 _2327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf2),
    .B(_1079_),
    .C(_1433_),
    .Y(_1434_)
);

OAI21X1 _2328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf0),
    .B(_958_),
    .C(RDY_bF$buf9),
    .Y(_1435_)
);

OAI21X1 _2329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_1233_),
    .C(_1435_),
    .Y(_1436_)
);

OAI21X1 _2330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf7),
    .B(_1027__bF$buf1),
    .C(_1436_),
    .Y(_1437_)
);

NOR2X1 _2331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1434_),
    .B(_1437_),
    .Y(_1438_)
);

OAI21X1 _2332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf1),
    .B(_1432_),
    .C(_1438_),
    .Y(_1439_)
);

OR2X2 _2333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1431_),
    .B(_1439_),
    .Y(_1440_)
);

AOI21X1 _2334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1423_),
    .B(_1429_),
    .C(_1440_),
    .Y(_1441_)
);

OAI21X1 _2335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1401_),
    .B(_1422_),
    .C(_1441_),
    .Y(_1442_)
);

INVX1 _2336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1442_),
    .Y(_1443_)
);

INVX1 _2337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_988_),
    .Y(_1444_)
);

OAI22X1 _2338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf6),
    .B(_1444_),
    .C(_1149__bF$buf0),
    .D(_1398_),
    .Y(_1445_)
);

OAI21X1 _2339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(write_back),
    .B(_1241_),
    .C(_1243_),
    .Y(_1446_)
);

OAI21X1 _2340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf1),
    .B(_928_),
    .C(_886__bF$buf0),
    .Y(_1447_)
);

OAI21X1 _2341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf6),
    .B(_1309_),
    .C(_1447_),
    .Y(_1448_)
);

OR2X2 _2342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1202_),
    .B(RDY_bF$buf5),
    .Y(_1449_)
);

NAND3X1 _2343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1448_),
    .B(_1449_),
    .C(_1446_),
    .Y(_1450_)
);

NOR2X1 _2344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1450_),
    .B(_1445_),
    .Y(_1451_)
);

OR2X2 _2345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1358_),
    .B(_1363_),
    .Y(_1452_)
);

NOR2X1 _2346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1389_),
    .B(_1452_),
    .Y(_1453_)
);

NAND2X1 _2347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1354_),
    .B(_1453_),
    .Y(_1454_)
);

NAND3X1 _2348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1308_),
    .B(_1256_),
    .C(_1302_),
    .Y(_1455_)
);

NOR3X1 _2349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1455_),
    .B(_1249_),
    .C(_1454_),
    .Y(_1456_)
);

NAND3X1 _2350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1451_),
    .B(_1443_),
    .C(_1456_),
    .Y(_1512_[2])
);

INVX1 _2351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1401_),
    .Y(_1457_)
);

OR2X2 _2352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1410_),
    .B(_1414_),
    .Y(_1458_)
);

NAND2X1 _2353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1420_),
    .B(_1419_),
    .Y(_1459_)
);

NOR2X1 _2354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1459_),
    .B(_1458_),
    .Y(_1460_)
);

NAND3X1 _2355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1457_),
    .B(_1408_),
    .C(_1460_),
    .Y(_1461_)
);

NAND3X1 _2356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1441_),
    .B(_1451_),
    .C(_1461_),
    .Y(_1462_)
);

AOI22X1 _2357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf5),
    .B(_1268_),
    .C(_1283_),
    .D(_1330_),
    .Y(_1463_)
);

NOR2X1 _2358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf0),
    .B(_1272_),
    .Y(_1464_)
);

MUX2X1 _2359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1464_),
    .B(_998_),
    .S(_886__bF$buf4),
    .Y(_1465_)
);

AND2X2 _2360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1463_),
    .B(_1465_),
    .Y(_1466_)
);

NAND2X1 _2361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf3),
    .B(_1031_),
    .Y(_1467_)
);

NAND2X1 _2362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_1020_),
    .Y(_1468_)
);

OAI21X1 _2363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf3),
    .B(_1467_),
    .C(_1468_),
    .Y(_1469_)
);

NAND2X1 _2364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_1031_),
    .Y(_1470_)
);

NOR2X1 _2365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_1470_),
    .Y(_1471_)
);

NOR2X1 _2366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1471_),
    .B(_1469_),
    .Y(_1472_)
);

NAND2X1 _2367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1472_),
    .B(_1466_),
    .Y(_1473_)
);

NOR2X1 _2368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1473_),
    .B(_1342_),
    .Y(_1474_)
);

NAND2X1 _2369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf3),
    .B(_1260_),
    .Y(_1475_)
);

NAND3X1 _2370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf1),
    .B(_1370_),
    .C(_1351_),
    .Y(_1476_)
);

OAI21X1 _2371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf3),
    .B(_954_),
    .C(RDY_bF$buf1),
    .Y(_1477_)
);

OAI21X1 _2372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf0),
    .B(_1257_),
    .C(_1477_),
    .Y(_1478_)
);

NAND3X1 _2373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1475_),
    .B(_1478_),
    .C(_1476_),
    .Y(_1479_)
);

INVX1 _2374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1479_),
    .Y(_1480_)
);

OR2X2 _2375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1408_),
    .B(_1149__bF$buf4),
    .Y(_1481_)
);

NAND3X1 _2376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1474_),
    .B(_1480_),
    .C(_1481_),
    .Y(_1482_)
);

NOR2X1 _2377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1391_),
    .B(_1482_),
    .Y(_1483_)
);

NAND3X1 _2378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1325_),
    .B(_1250_),
    .C(_1483_),
    .Y(_1484_)
);

INVX1 _2379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1248_),
    .Y(_1485_)
);

NOR2X1 _2380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1479_),
    .B(_1452_),
    .Y(_1486_)
);

NOR2X1 _2381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1369_),
    .B(_1372_),
    .Y(_1487_)
);

INVX1 _2382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1266_),
    .Y(_1488_)
);

NAND3X1 _2383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1308_),
    .B(_1336_),
    .C(_1488_),
    .Y(_1489_)
);

NOR3X1 _2384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1288_),
    .B(_1322_),
    .C(_1489_),
    .Y(_1490_)
);

AND2X2 _2385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1490_),
    .B(_1487_),
    .Y(_1491_)
);

NAND3X1 _2386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1485_),
    .B(_1486_),
    .C(_1491_),
    .Y(_1492_)
);

NOR2X1 _2387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1492_),
    .B(_1442_),
    .Y(_1493_)
);

OAI21X1 _2388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1462_),
    .B(_1484_),
    .C(_1493_),
    .Y(_1512_[3])
);

NAND3X1 _2389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1475_),
    .B(_1476_),
    .C(_1333_),
    .Y(_1494_)
);

NOR2X1 _2390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1494_),
    .B(_1353_),
    .Y(_1495_)
);

NOR2X1 _2391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1239_),
    .B(_1434_),
    .Y(_1496_)
);

INVX1 _2392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1293_),
    .Y(_1497_)
);

AND2X2 _2393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1311_),
    .B(_1321_),
    .Y(_1498_)
);

NAND3X1 _2394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1197_),
    .B(_1497_),
    .C(_1498_),
    .Y(_1499_)
);

NAND3X1 _2395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1262_),
    .B(_1308_),
    .C(_1274_),
    .Y(_1500_)
);

NOR2X1 _2396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1499_),
    .B(_1500_),
    .Y(_1501_)
);

NAND3X1 _2397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1448_),
    .B(_1496_),
    .C(_1501_),
    .Y(_1502_)
);

NOR2X1 _2398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1369_),
    .B(_1502_),
    .Y(_1503_)
);

INVX1 _2399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1466_),
    .Y(_1504_)
);

NOR2X1 _2400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1358_),
    .B(_1504_),
    .Y(_1505_)
);

NAND3X1 _2401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1495_),
    .B(_1505_),
    .C(_1503_),
    .Y(_1512_[4])
);

INVX1 _2402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1192_),
    .Y(_1506_)
);

NOR2X1 _2403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1372_),
    .B(_1506_),
    .Y(_1507_)
);

INVX1 _2404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1478_),
    .Y(_1508_)
);

NOR2X1 _2405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1469_),
    .B(_1508_),
    .Y(_1509_)
);

AND2X2 _2406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1509_),
    .B(_1436_),
    .Y(_1510_)
);

AND2X2 _2407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1510_),
    .B(_1463_),
    .Y(_1511_)
);

AND2X2 _2408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1511_),
    .B(_1285_),
    .Y(_117_)
);

AND2X2 _2409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_117_),
    .B(_1254_),
    .Y(_118_)
);

NOR2X1 _2410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1237_),
    .B(_1339_),
    .Y(_119_)
);

NOR2X1 _2411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1289_),
    .B(_1270_),
    .Y(_120_)
);

NAND2X1 _2412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_119_),
    .B(_120_),
    .Y(_121_)
);

OAI21X1 _2413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf9),
    .B(_1227_),
    .C(_1359_),
    .Y(_122_)
);

NOR2X1 _2414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_122_),
    .B(_1387_),
    .Y(_123_)
);

NAND3X1 _2415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1259_),
    .B(_1318_),
    .C(_123_),
    .Y(_124_)
);

NOR2X1 _2416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_121_),
    .B(_124_),
    .Y(_125_)
);

NAND2X1 _2417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1282_),
    .B(_125_),
    .Y(_126_)
);

NOR2X1 _2418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1445_),
    .B(_126_),
    .Y(_127_)
);

NAND3X1 _2419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1507_),
    .B(_127_),
    .C(_118_),
    .Y(_1512_[5])
);

INVX1 _2420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(op[0]),
    .Y(_128_)
);

INVX2 _2421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_915_),
    .Y(_129_)
);

INVX1 _2422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1275_),
    .Y(_130_)
);

NAND3X1 _2423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf0),
    .B(_130_),
    .C(_129_),
    .Y(_131_)
);

OAI21X1 _2424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_129_),
    .C(_131_),
    .Y(alu_op[0])
);

INVX1 _2425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(op[1]),
    .Y(_132_)
);

OAI21X1 _2426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_132_),
    .B(_129_),
    .C(_131_),
    .Y(alu_op[1])
);

INVX1 _2427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1337_),
    .Y(_133_)
);

NOR2X1 _2428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_133_),
    .B(_1263_),
    .Y(_134_)
);

INVX1 _2429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_134_),
    .Y(_135_)
);

INVX2 _2430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1080_),
    .Y(_136_)
);

OAI21X1 _2431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .B(_1075_),
    .C(_136_),
    .Y(_137_)
);

NOR2X1 _2432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_135_),
    .B(_137_),
    .Y(_138_)
);

AOI22X1 _2433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(backwards),
    .B(_925_),
    .C(_915_),
    .D(op[2]),
    .Y(_139_)
);

NAND2X1 _2434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_139_),
    .B(_138_),
    .Y(alu_op[2])
);

INVX1 _2435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(op[3]),
    .Y(_140_)
);

NOR2X1 _2436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_140_),
    .B(_129_),
    .Y(alu_op[3])
);

OAI21X1 _2437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf4),
    .B(_946_),
    .C(_1204_),
    .Y(_141_)
);

OAI21X1 _2438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1199_),
    .B(_141_),
    .C(store),
    .Y(_142_)
);

NAND3X1 _2439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1227_),
    .B(_142_),
    .C(_138_),
    .Y(_1743_)
);

OAI21X1 _2440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf2),
    .B(_949_),
    .C(_138_),
    .Y(_143_)
);

OAI21X1 _2441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(php),
    .B(_1337_),
    .C(_1227_),
    .Y(_144_)
);

NAND2X1 _2442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[0]),
    .B(_144_),
    .Y(_145_)
);

OAI21X1 _2443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf2),
    .B(_1263_),
    .C(PC[8]),
    .Y(_146_)
);

INVX1 _2444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(php),
    .Y(_147_)
);

NAND2X1 _2445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_935_),
    .Y(_148_)
);

OAI21X1 _2446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_147_),
    .B(_1337_),
    .C(_148_),
    .Y(_149_)
);

AOI22X1 _2447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[0]),
    .B(_1080_),
    .C(_149_),
    .D(C),
    .Y(_150_)
);

NAND3X1 _2448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_145_),
    .B(_146_),
    .C(_150_),
    .Y(_151_)
);

INVX1 _2449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_151_),
    .Y(_152_)
);

OAI21X1 _2450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1060_),
    .C(_152_),
    .Y(_1742_[0])
);

OAI21X1 _2451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf1),
    .B(_1263_),
    .C(PC[9]),
    .Y(_153_)
);

NOR2X1 _2452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_147_),
    .B(_1337_),
    .Y(_154_)
);

OAI21X1 _2453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1334_),
    .B(_154_),
    .C(Z),
    .Y(_155_)
);

AOI22X1 _2454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[1]),
    .B(_1080_),
    .C(_144_),
    .D(ADD[1]),
    .Y(_156_)
);

NAND3X1 _2455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_153_),
    .B(_156_),
    .C(_155_),
    .Y(_157_)
);

INVX1 _2456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_157_),
    .Y(_158_)
);

OAI21X1 _2457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1090_),
    .C(_158_),
    .Y(_1742_[1])
);

NAND2X1 _2458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[2]),
    .B(_144_),
    .Y(_159_)
);

OAI21X1 _2459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf0),
    .B(_1263_),
    .C(PC[10]),
    .Y(_160_)
);

AOI22X1 _2460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[2]),
    .B(_1080_),
    .C(_149_),
    .D(I),
    .Y(_161_)
);

NAND3X1 _2461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_159_),
    .B(_160_),
    .C(_161_),
    .Y(_162_)
);

INVX1 _2462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_162_),
    .Y(_163_)
);

OAI21X1 _2463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1101_),
    .C(_163_),
    .Y(_1742_[2])
);

INVX1 _2464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(D),
    .Y(_164_)
);

INVX1 _2465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_149_),
    .Y(_165_)
);

OAI21X1 _2466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf3),
    .B(_1263_),
    .C(PC[11]),
    .Y(_166_)
);

OAI21X1 _2467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1009_),
    .B(_136_),
    .C(_166_),
    .Y(_167_)
);

AOI21X1 _2468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[3]),
    .B(_144_),
    .C(_167_),
    .Y(_168_)
);

OAI21X1 _2469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_164_),
    .B(_165_),
    .C(_168_),
    .Y(_169_)
);

INVX1 _2470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_169_),
    .Y(_170_)
);

OAI21X1 _2471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1109_),
    .C(_170_),
    .Y(_1742_[3])
);

AOI21X1 _2472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[4]),
    .B(_1080_),
    .C(_154_),
    .Y(_171_)
);

OAI21X1 _2473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .B(_1166_),
    .C(_171_),
    .Y(_172_)
);

INVX1 _2474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[4]),
    .Y(_173_)
);

OAI21X1 _2475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_971_),
    .B(_941_),
    .C(_903__bF$buf2),
    .Y(_174_)
);

OAI21X1 _2476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf2),
    .B(_1263_),
    .C(PC[12]),
    .Y(_175_)
);

OAI21X1 _2477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_173_),
    .B(_174_),
    .C(_175_),
    .Y(_176_)
);

NOR2X1 _2478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_176_),
    .B(_172_),
    .Y(_177_)
);

OAI21X1 _2479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1117_),
    .C(_177_),
    .Y(_1742_[4])
);

OAI21X1 _2480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1012_),
    .B(_136_),
    .C(_165_),
    .Y(_178_)
);

INVX1 _2481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[5]),
    .Y(_179_)
);

OAI21X1 _2482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf1),
    .B(_1263_),
    .C(PC[13]),
    .Y(_180_)
);

OAI21X1 _2483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_179_),
    .B(_174_),
    .C(_180_),
    .Y(_181_)
);

NOR2X1 _2484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_178_),
    .B(_181_),
    .Y(_182_)
);

OAI21X1 _2485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1125_),
    .C(_182_),
    .Y(_1742_[5])
);

OAI21X1 _2486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf0),
    .B(_1263_),
    .C(PC[14]),
    .Y(_183_)
);

OAI21X1 _2487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1014_),
    .B(_136_),
    .C(_183_),
    .Y(_184_)
);

AOI21X1 _2488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[6]),
    .B(_144_),
    .C(_184_),
    .Y(_185_)
);

OAI21X1 _2489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1374_),
    .B(_165_),
    .C(_185_),
    .Y(_186_)
);

INVX1 _2490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_186_),
    .Y(_187_)
);

OAI21X1 _2491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1133_),
    .C(_187_),
    .Y(_1742_[6])
);

OAI21X1 _2492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf3),
    .B(_1263_),
    .C(PC[15]),
    .Y(_188_)
);

OAI21X1 _2493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1016_),
    .B(_136_),
    .C(_188_),
    .Y(_189_)
);

AOI21X1 _2494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .B(_144_),
    .C(_189_),
    .Y(_190_)
);

OAI21X1 _2495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1377_),
    .B(_165_),
    .C(_190_),
    .Y(_191_)
);

INVX1 _2496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_191_),
    .Y(_192_)
);

OAI21X1 _2497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_143_),
    .B(_1143_),
    .C(_192_),
    .Y(_1742_[7])
);

OAI21X1 _2498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf1),
    .B(_946_),
    .C(_1067_),
    .Y(_193_)
);

NOR2X1 _2499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_193_),
    .B(_135_),
    .Y(_194_)
);

INVX2 _2500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_194_),
    .Y(_195_)
);

OAI21X1 _2501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf0),
    .B(_949_),
    .C(_909_),
    .Y(_196_)
);

NAND2X1 _2502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_955_),
    .Y(_197_)
);

NAND3X1 _2503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1202_),
    .B(_197_),
    .C(_1224_),
    .Y(_198_)
);

NOR2X1 _2504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_196_),
    .B(_198_),
    .Y(_199_)
);

INVX2 _2505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_199_),
    .Y(_200_)
);

NOR2X1 _2506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1201_),
    .B(_943_),
    .Y(_201_)
);

NAND2X1 _2507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_201_),
    .B(_194_),
    .Y(_202_)
);

NOR2X1 _2508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_200_),
    .B(_202_),
    .Y(_203_)
);

OAI21X1 _2509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_993_),
    .B(_992_),
    .C(_903__bF$buf1),
    .Y(_204_)
);

NAND3X1 _2510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1077_),
    .B(_204_),
    .C(_1081_),
    .Y(_205_)
);

NOR2X1 _2511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1020_),
    .B(_205_),
    .Y(_206_)
);

NAND3X1 _2512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_940_),
    .B(_1028_),
    .C(_1267_),
    .Y(_207_)
);

NOR2X1 _2513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1464_),
    .B(_207_),
    .Y(_208_)
);

NAND2X1 _2514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_208_),
    .B(_206_),
    .Y(_209_)
);

NAND2X1 _2515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf0),
    .B(_1427_),
    .Y(_210_)
);

INVX1 _2516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1291_),
    .Y(_211_)
);

NAND3X1 _2517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_210_),
    .B(_211_),
    .C(_1226_),
    .Y(_212_)
);

OAI22X1 _2518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf1),
    .B(_974_),
    .C(_931__bF$buf3),
    .D(_984_),
    .Y(_213_)
);

OR2X2 _2519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_932_),
    .B(_213_),
    .Y(_214_)
);

NOR2X1 _2520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_212_),
    .B(_214_),
    .Y(_215_)
);

OAI21X1 _2521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .B(_996_),
    .C(_215_),
    .Y(_216_)
);

NOR2X1 _2522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(_209_),
    .Y(_217_)
);

NAND2X1 _2523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_203_),
    .B(_217_),
    .Y(_218_)
);

NAND2X1 _2524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[0]),
    .B(_209_),
    .Y(_219_)
);

OAI21X1 _2525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_196_),
    .B(_198_),
    .C(ABL[0]),
    .Y(_220_)
);

OAI21X1 _2526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_966_),
    .B(_201_),
    .C(_220_),
    .Y(_221_)
);

AOI21X1 _2527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(ADD[0]),
    .C(_221_),
    .Y(_222_)
);

AND2X2 _2528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_219_),
    .B(_222_),
    .Y(_223_)
);

OAI21X1 _2529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_965_),
    .B(_218_),
    .C(_223_),
    .Y(_224_)
);

AOI21X1 _2530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1059_),
    .B(_195_),
    .C(_224_),
    .Y(_225_)
);

INVX1 _2531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_225_),
    .Y(_1741_[0])
);

OAI21X1 _2532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(_209_),
    .C(ADD[1]),
    .Y(_226_)
);

INVX1 _2533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_201_),
    .Y(_227_)
);

AOI22X1 _2534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[1]),
    .B(_227_),
    .C(_200_),
    .D(ABL[1]),
    .Y(_228_)
);

AND2X2 _2535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_226_),
    .B(_228_),
    .Y(_229_)
);

OAI21X1 _2536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1005_),
    .B(_218_),
    .C(_229_),
    .Y(_230_)
);

AOI21X1 _2537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1089_),
    .B(_195_),
    .C(_230_),
    .Y(_231_)
);

INVX1 _2538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_231_),
    .Y(_1741_[1])
);

OAI21X1 _2539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(_209_),
    .C(ADD[2]),
    .Y(_232_)
);

AOI22X1 _2540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[2]),
    .B(_227_),
    .C(_200_),
    .D(ABL[2]),
    .Y(_233_)
);

AND2X2 _2541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_232_),
    .B(_233_),
    .Y(_234_)
);

OAI21X1 _2542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1007_),
    .B(_218_),
    .C(_234_),
    .Y(_235_)
);

AOI21X1 _2543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1100_),
    .B(_195_),
    .C(_235_),
    .Y(_236_)
);

INVX1 _2544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_236_),
    .Y(_1741_[2])
);

OR2X2 _2545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_209_),
    .B(_216_),
    .Y(_237_)
);

INVX1 _2546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[3]),
    .Y(_238_)
);

OAI22X1 _2547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1010_),
    .B(_201_),
    .C(_238_),
    .D(_199_),
    .Y(_239_)
);

AOI21X1 _2548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_237_),
    .B(ADD[3]),
    .C(_239_),
    .Y(_240_)
);

OAI21X1 _2549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1009_),
    .B(_218_),
    .C(_240_),
    .Y(_241_)
);

AOI21X1 _2550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1108_),
    .B(_195_),
    .C(_241_),
    .Y(_242_)
);

INVX1 _2551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_242_),
    .Y(_1741_[3])
);

NAND2X1 _2552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[4]),
    .B(_209_),
    .Y(_243_)
);

INVX1 _2553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[4]),
    .Y(_244_)
);

OAI22X1 _2554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_888_),
    .B(_201_),
    .C(_244_),
    .D(_199_),
    .Y(_245_)
);

AOI21X1 _2555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(ADD[4]),
    .C(_245_),
    .Y(_246_)
);

AND2X2 _2556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_243_),
    .B(_246_),
    .Y(_247_)
);

OAI21X1 _2557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1011_),
    .B(_218_),
    .C(_247_),
    .Y(_248_)
);

AOI21X1 _2558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1116_),
    .B(_195_),
    .C(_248_),
    .Y(_249_)
);

INVX1 _2559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_249_),
    .Y(_1741_[4])
);

NAND2X1 _2560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[5]),
    .B(_209_),
    .Y(_250_)
);

INVX1 _2561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[5]),
    .Y(_251_)
);

OAI22X1 _2562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1013_),
    .B(_201_),
    .C(_251_),
    .D(_199_),
    .Y(_252_)
);

AOI21X1 _2563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(ADD[5]),
    .C(_252_),
    .Y(_253_)
);

NAND2X1 _2564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_253_),
    .B(_250_),
    .Y(_254_)
);

INVX1 _2565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_254_),
    .Y(_255_)
);

OAI21X1 _2566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1012_),
    .B(_218_),
    .C(_255_),
    .Y(_256_)
);

AOI21X1 _2567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1124_),
    .B(_195_),
    .C(_256_),
    .Y(_257_)
);

INVX1 _2568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_257_),
    .Y(_1741_[5])
);

OAI21X1 _2569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(_209_),
    .C(ADD[6]),
    .Y(_258_)
);

AOI22X1 _2570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[6]),
    .B(_227_),
    .C(_200_),
    .D(ABL[6]),
    .Y(_259_)
);

AND2X2 _2571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_258_),
    .B(_259_),
    .Y(_260_)
);

OAI21X1 _2572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1014_),
    .B(_218_),
    .C(_260_),
    .Y(_261_)
);

AOI21X1 _2573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1132_),
    .B(_195_),
    .C(_261_),
    .Y(_262_)
);

INVX1 _2574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_262_),
    .Y(_1741_[6])
);

OAI21X1 _2575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_216_),
    .B(_209_),
    .C(AN),
    .Y(_263_)
);

AOI22X1 _2576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[7]),
    .B(_227_),
    .C(_200_),
    .D(ABL[7]),
    .Y(_264_)
);

AND2X2 _2577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_263_),
    .B(_264_),
    .Y(_265_)
);

OAI21X1 _2578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1016_),
    .B(_218_),
    .C(_265_),
    .Y(_266_)
);

AOI21X1 _2579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1142_),
    .B(_195_),
    .C(_266_),
    .Y(_267_)
);

INVX1 _2580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_267_),
    .Y(_1741_[7])
);

INVX2 _2581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[8]),
    .Y(_268_)
);

INVX1 _2582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[0]),
    .Y(_269_)
);

INVX2 _2583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_196_),
    .Y(_270_)
);

OAI21X1 _2584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_269_),
    .B(_270_),
    .C(_206_),
    .Y(_271_)
);

INVX2 _2585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_215_),
    .Y(_272_)
);

AOI22X1 _2586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[0]),
    .B(_198_),
    .C(_272_),
    .D(DIMUX[0]),
    .Y(_273_)
);

NAND3X1 _2587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1083_),
    .B(_194_),
    .C(_273_),
    .Y(_274_)
);

NOR2X1 _2588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_274_),
    .Y(_275_)
);

OAI21X1 _2589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_268_),
    .B(_218_),
    .C(_275_),
    .Y(_1741_[8])
);

INVX1 _2590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[9]),
    .Y(_276_)
);

AOI21X1 _2591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_198_),
    .B(ADD[1]),
    .C(_1093_),
    .Y(_277_)
);

OAI21X1 _2592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1091_),
    .B(_270_),
    .C(_277_),
    .Y(_278_)
);

AOI21X1 _2593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_272_),
    .B(DIMUX[1]),
    .C(_278_),
    .Y(_279_)
);

OAI21X1 _2594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_276_),
    .B(_218_),
    .C(_279_),
    .Y(_1741_[9])
);

INVX1 _2595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[10]),
    .Y(_280_)
);

AOI22X1 _2596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[2]),
    .B(_198_),
    .C(_272_),
    .D(DIMUX[2]),
    .Y(_281_)
);

OAI21X1 _2597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_925_),
    .B(_196_),
    .C(ABH[2]),
    .Y(_282_)
);

NAND2X1 _2598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_282_),
    .B(_281_),
    .Y(_283_)
);

INVX1 _2599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_283_),
    .Y(_284_)
);

OAI21X1 _2600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_280_),
    .B(_218_),
    .C(_284_),
    .Y(_1741_[10])
);

INVX2 _2601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[11]),
    .Y(_285_)
);

AOI22X1 _2602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[3]),
    .B(_198_),
    .C(_272_),
    .D(DIMUX[3]),
    .Y(_286_)
);

OAI21X1 _2603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_925_),
    .B(_196_),
    .C(ABH[3]),
    .Y(_287_)
);

NAND2X1 _2604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_287_),
    .B(_286_),
    .Y(_288_)
);

INVX1 _2605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_288_),
    .Y(_289_)
);

OAI21X1 _2606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_285_),
    .B(_218_),
    .C(_289_),
    .Y(_1741_[11])
);

INVX1 _2607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[12]),
    .Y(_290_)
);

INVX1 _2608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[4]),
    .Y(_291_)
);

AOI22X1 _2609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[4]),
    .B(_925_),
    .C(_198_),
    .D(ADD[4]),
    .Y(_292_)
);

OAI21X1 _2610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_291_),
    .B(_270_),
    .C(_292_),
    .Y(_293_)
);

AOI21X1 _2611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_272_),
    .B(DIMUX[4]),
    .C(_293_),
    .Y(_294_)
);

OAI21X1 _2612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_290_),
    .B(_218_),
    .C(_294_),
    .Y(_1741_[12])
);

INVX1 _2613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[13]),
    .Y(_295_)
);

INVX1 _2614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[5]),
    .Y(_296_)
);

AOI22X1 _2615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[5]),
    .B(_925_),
    .C(_198_),
    .D(ADD[5]),
    .Y(_297_)
);

OAI21X1 _2616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_296_),
    .B(_270_),
    .C(_297_),
    .Y(_298_)
);

AOI21X1 _2617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_272_),
    .B(DIMUX[5]),
    .C(_298_),
    .Y(_299_)
);

OAI21X1 _2618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_295_),
    .B(_218_),
    .C(_299_),
    .Y(_1741_[13])
);

INVX1 _2619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[14]),
    .Y(_300_)
);

AOI21X1 _2620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_198_),
    .B(ADD[6]),
    .C(_1135_),
    .Y(_301_)
);

OAI21X1 _2621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1134_),
    .B(_270_),
    .C(_301_),
    .Y(_302_)
);

AOI21X1 _2622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_272_),
    .B(DIMUX[6]),
    .C(_302_),
    .Y(_303_)
);

OAI21X1 _2623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_300_),
    .B(_218_),
    .C(_303_),
    .Y(_1741_[14])
);

INVX1 _2624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[15]),
    .Y(_304_)
);

AOI21X1 _2625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_198_),
    .B(AN),
    .C(_1145_),
    .Y(_305_)
);

OAI21X1 _2626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1144_),
    .B(_270_),
    .C(_305_),
    .Y(_306_)
);

AOI21X1 _2627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_272_),
    .B(DIMUX[7]),
    .C(_306_),
    .Y(_307_)
);

OAI21X1 _2628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_304_),
    .B(_218_),
    .C(_307_),
    .Y(_1741_[15])
);

INVX1 _2629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(adc_sbc),
    .Y(_308_)
);

NOR2X1 _2630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_308_),
    .B(_164_),
    .Y(_0_)
);

INVX1 _2631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(adc_bcd),
    .Y(_309_)
);

NOR2X1 _2632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_309_),
    .B(_917_),
    .Y(\u_ALU8.BCD )
);

INVX1 _2633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shift_right),
    .Y(_310_)
);

NOR2X1 _2634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_310_),
    .B(_129_),
    .Y(alu_shift_right)
);

INVX8 _2635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .Y(_1_)
);

OAI21X1 _2636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf0),
    .B(_942_),
    .C(_1470_),
    .Y(_311_)
);

NOR2X1 _2637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1154_),
    .B(_1027__bF$buf4),
    .Y(_312_)
);

INVX1 _2638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_312_),
    .Y(_313_)
);

OAI21X1 _2639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_913_),
    .B(_901_),
    .C(_1427_),
    .Y(_314_)
);

OAI21X1 _2640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_314_),
    .C(_313_),
    .Y(_315_)
);

NOR2X1 _2641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_311_),
    .B(_315_),
    .Y(_316_)
);

AOI21X1 _2642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_1221_),
    .C(_967_),
    .Y(_317_)
);

NOR2X1 _2643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1424_),
    .B(_1021_),
    .Y(_318_)
);

AND2X2 _2644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_317_),
    .B(_318_),
    .Y(_319_)
);

NAND3X1 _2645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1432_),
    .B(_316_),
    .C(_319_),
    .Y(_320_)
);

OAI22X1 _2646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf3),
    .B(_969_),
    .C(_1221_),
    .D(_1427_),
    .Y(_321_)
);

NAND3X1 _2647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1092_),
    .B(_321_),
    .C(_211_),
    .Y(_322_)
);

NOR2X1 _2648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf3),
    .B(_1167_),
    .Y(_323_)
);

AOI22X1 _2649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[0]),
    .B(_323_),
    .C(_322_),
    .D(ADD[0]),
    .Y(_324_)
);

AOI22X1 _2650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf3),
    .B(_931__bF$buf2),
    .C(_984_),
    .D(_912_),
    .Y(_325_)
);

NOR3X1 _2651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_925_),
    .B(_1291_),
    .C(_325_),
    .Y(_326_)
);

OAI21X1 _2652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf4),
    .B(_954_),
    .C(_1027__bF$buf2),
    .Y(_327_)
);

AOI21X1 _2653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_929_),
    .B(_935_),
    .C(_327_),
    .Y(_328_)
);

OAI21X1 _2654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf1),
    .B(_1154_),
    .C(_197_),
    .Y(_329_)
);

AOI21X1 _2655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_326_),
    .B(_328_),
    .C(_329_),
    .Y(_330_)
);

OAI21X1 _2656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_965_),
    .B(_330_),
    .C(_324_),
    .Y(_331_)
);

NOR2X1 _2657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_320_),
    .B(_331_),
    .Y(_332_)
);

AND2X2 _2658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_331_),
    .B(_320_),
    .Y(_333_)
);

OR2X2 _2659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_333_),
    .B(_886__bF$buf2),
    .Y(_334_)
);

OAI22X1 _2660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_965_),
    .C(_332_),
    .D(_334_),
    .Y(_2_)
);

NAND2X1 _2661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[1]),
    .B(_323_),
    .Y(_335_)
);

OAI21X1 _2662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(res),
    .B(_148_),
    .C(_335_),
    .Y(_336_)
);

AOI21X1 _2663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(ADD[1]),
    .C(_336_),
    .Y(_337_)
);

OAI21X1 _2664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1005_),
    .B(_330_),
    .C(_337_),
    .Y(_338_)
);

NOR2X1 _2665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_338_),
    .B(_333_),
    .Y(_339_)
);

NAND3X1 _2666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_320_),
    .B(_331_),
    .C(_338_),
    .Y(_340_)
);

NAND2X1 _2667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf7),
    .B(_340_),
    .Y(_341_)
);

OAI22X1 _2668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf6),
    .B(_1005_),
    .C(_341_),
    .D(_339_),
    .Y(_3_)
);

INVX1 _2669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_340_),
    .Y(_342_)
);

OAI21X1 _2670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1153_),
    .B(res),
    .C(_1334_),
    .Y(_343_)
);

AOI22X1 _2671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[2]),
    .B(_323_),
    .C(_322_),
    .D(ADD[2]),
    .Y(_344_)
);

NAND2X1 _2672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_343_),
    .B(_344_),
    .Y(_345_)
);

INVX1 _2673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_345_),
    .Y(_346_)
);

OAI21X1 _2674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1007_),
    .B(_330_),
    .C(_346_),
    .Y(_347_)
);

NOR2X1 _2675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_347_),
    .B(_342_),
    .Y(_348_)
);

INVX1 _2676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_347_),
    .Y(_349_)
);

OAI21X1 _2677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_340_),
    .B(_349_),
    .C(RDY_bF$buf5),
    .Y(_350_)
);

OAI22X1 _2678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_1007_),
    .C(_350_),
    .D(_348_),
    .Y(_4_)
);

NOR2X1 _2679_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1291_),
    .B(_325_),
    .Y(_351_)
);

NAND3X1 _2680_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1092_),
    .B(_328_),
    .C(_351_),
    .Y(_352_)
);

INVX2 _2681_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .Y(_353_)
);

AOI21X1 _2682_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_352_),
    .B(_353_),
    .C(_1009_),
    .Y(_354_)
);

INVX1 _2683_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[3]),
    .Y(_355_)
);

AOI21X1 _2684_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[3]),
    .B(_323_),
    .C(_1334_),
    .Y(_356_)
);

OAI21X1 _2685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_355_),
    .B(_326_),
    .C(_356_),
    .Y(_357_)
);

NOR2X1 _2686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_357_),
    .B(_354_),
    .Y(_358_)
);

INVX1 _2687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_358_),
    .Y(_359_)
);

AOI21X1 _2688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_342_),
    .B(_347_),
    .C(_359_),
    .Y(_360_)
);

AOI21X1 _2689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_352_),
    .B(_353_),
    .C(_1007_),
    .Y(_361_)
);

OAI22X1 _2690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_345_),
    .B(_361_),
    .C(_354_),
    .D(_357_),
    .Y(_362_)
);

OAI21X1 _2691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_362_),
    .B(_340_),
    .C(RDY_bF$buf3),
    .Y(_363_)
);

OAI22X1 _2692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_1009_),
    .C(_363_),
    .D(_360_),
    .Y(_5_)
);

NAND3X1 _2693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf0),
    .B(_148_),
    .C(_197_),
    .Y(_364_)
);

NOR2X1 _2694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_364_),
    .B(_322_),
    .Y(_365_)
);

OAI21X1 _2695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .B(_365_),
    .C(PC[2]),
    .Y(_366_)
);

OAI21X1 _2696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .B(_365_),
    .C(PC[3]),
    .Y(_367_)
);

INVX1 _2697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_357_),
    .Y(_368_)
);

AOI22X1 _2698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_367_),
    .B(_368_),
    .C(_346_),
    .D(_366_),
    .Y(_369_)
);

NAND3X1 _2699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_338_),
    .B(_369_),
    .C(_333_),
    .Y(_370_)
);

OAI21X1 _2700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_364_),
    .B(_322_),
    .C(_353_),
    .Y(_371_)
);

AOI21X1 _2701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[4]),
    .B(_323_),
    .C(_1334_),
    .Y(_372_)
);

OAI21X1 _2702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_173_),
    .B(_326_),
    .C(_372_),
    .Y(_373_)
);

AOI21X1 _2703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[4]),
    .B(_371_),
    .C(_373_),
    .Y(_374_)
);

AND2X2 _2704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_370_),
    .B(_374_),
    .Y(_375_)
);

OAI21X1 _2705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_374_),
    .B(_370_),
    .C(RDY_bF$buf1),
    .Y(_376_)
);

OAI22X1 _2706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf0),
    .B(_1011_),
    .C(_376_),
    .D(_375_),
    .Y(_6_)
);

AOI21X1 _2707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_352_),
    .B(_353_),
    .C(_1012_),
    .Y(_377_)
);

INVX2 _2708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_323_),
    .Y(_378_)
);

OAI21X1 _2709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_251_),
    .B(_378_),
    .C(_148_),
    .Y(_379_)
);

INVX1 _2710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_379_),
    .Y(_380_)
);

OAI21X1 _2711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_179_),
    .B(_326_),
    .C(_380_),
    .Y(_381_)
);

NOR2X1 _2712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_377_),
    .B(_381_),
    .Y(_382_)
);

OAI21X1 _2713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_374_),
    .B(_370_),
    .C(_382_),
    .Y(_383_)
);

AOI21X1 _2714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_352_),
    .B(_353_),
    .C(_1011_),
    .Y(_384_)
);

OAI22X1 _2715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_373_),
    .B(_384_),
    .C(_377_),
    .D(_381_),
    .Y(_385_)
);

NOR3X1 _2716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_362_),
    .B(_385_),
    .C(_340_),
    .Y(_386_)
);

INVX1 _2717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_386_),
    .Y(_387_)
);

NAND3X1 _2718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf9),
    .B(_387_),
    .C(_383_),
    .Y(_388_)
);

OAI21X1 _2719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_1012_),
    .C(_388_),
    .Y(_7_)
);

INVX1 _2720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[6]),
    .Y(_389_)
);

OAI21X1 _2721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_389_),
    .B(_378_),
    .C(_148_),
    .Y(_390_)
);

AOI21X1 _2722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(ADD[6]),
    .C(_390_),
    .Y(_391_)
);

OAI21X1 _2723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1014_),
    .B(_330_),
    .C(_391_),
    .Y(_392_)
);

NOR2X1 _2724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_392_),
    .B(_386_),
    .Y(_393_)
);

INVX1 _2725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_392_),
    .Y(_394_)
);

OAI21X1 _2726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_394_),
    .B(_387_),
    .C(RDY_bF$buf7),
    .Y(_395_)
);

OAI22X1 _2727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf6),
    .B(_1014_),
    .C(_393_),
    .D(_395_),
    .Y(_8_)
);

INVX1 _2728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[7]),
    .Y(_396_)
);

OAI21X1 _2729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_396_),
    .B(_378_),
    .C(_148_),
    .Y(_397_)
);

AOI21X1 _2730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(AN),
    .C(_397_),
    .Y(_398_)
);

OAI21X1 _2731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1016_),
    .B(_330_),
    .C(_398_),
    .Y(_399_)
);

AOI21X1 _2732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_386_),
    .B(_392_),
    .C(_399_),
    .Y(_400_)
);

NAND3X1 _2733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_392_),
    .B(_399_),
    .C(_386_),
    .Y(_401_)
);

NAND2X1 _2734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf5),
    .B(_401_),
    .Y(_402_)
);

OAI22X1 _2735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_1016_),
    .C(_400_),
    .D(_402_),
    .Y(_9_)
);

AOI21X1 _2736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_211_),
    .B(_321_),
    .C(_966_),
    .Y(_403_)
);

OAI21X1 _2737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_268_),
    .B(_313_),
    .C(_1083_),
    .Y(_404_)
);

NAND2X1 _2738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[0]),
    .B(_1299_),
    .Y(_405_)
);

NAND2X1 _2739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[0]),
    .B(_323_),
    .Y(_406_)
);

NAND3X1 _2740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .B(_405_),
    .C(_406_),
    .Y(_407_)
);

NOR3X1 _2741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_403_),
    .B(_404_),
    .C(_407_),
    .Y(_408_)
);

OAI21X1 _2742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_268_),
    .B(_352_),
    .C(_408_),
    .Y(_409_)
);

INVX1 _2743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_409_),
    .Y(_410_)
);

AND2X2 _2744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_401_),
    .B(_410_),
    .Y(_411_)
);

OAI21X1 _2745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_410_),
    .B(_401_),
    .C(RDY_bF$buf3),
    .Y(_412_)
);

OAI22X1 _2746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_268_),
    .C(_412_),
    .D(_411_),
    .Y(_10_)
);

OAI21X1 _2747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .B(_365_),
    .C(PC[5]),
    .Y(_413_)
);

AOI21X1 _2748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(ADD[5]),
    .C(_379_),
    .Y(_414_)
);

AOI21X1 _2749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_413_),
    .B(_414_),
    .C(_374_),
    .Y(_415_)
);

NAND3X1 _2750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_392_),
    .B(_399_),
    .C(_415_),
    .Y(_416_)
);

NOR2X1 _2751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_416_),
    .B(_370_),
    .Y(_417_)
);

NOR2X1 _2752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_312_),
    .B(_365_),
    .Y(_418_)
);

INVX1 _2753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_351_),
    .Y(_419_)
);

AOI22X1 _2754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[1]),
    .B(_1299_),
    .C(_323_),
    .D(ABH[1]),
    .Y(_420_)
);

NAND3X1 _2755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .B(_420_),
    .C(_1094_),
    .Y(_421_)
);

AOI21X1 _2756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[1]),
    .B(_419_),
    .C(_421_),
    .Y(_422_)
);

OAI21X1 _2757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_276_),
    .B(_418_),
    .C(_422_),
    .Y(_423_)
);

AOI21X1 _2758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_409_),
    .C(_423_),
    .Y(_424_)
);

NOR2X1 _2759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_404_),
    .B(_407_),
    .Y(_425_)
);

OAI21X1 _2760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_966_),
    .B(_351_),
    .C(_425_),
    .Y(_426_)
);

NOR2X1 _2761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_268_),
    .B(_352_),
    .Y(_427_)
);

OAI21X1 _2762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_426_),
    .B(_427_),
    .C(_423_),
    .Y(_428_)
);

OAI21X1 _2763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_428_),
    .B(_401_),
    .C(RDY_bF$buf1),
    .Y(_429_)
);

OAI22X1 _2764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf0),
    .B(_276_),
    .C(_424_),
    .D(_429_),
    .Y(_11_)
);

NOR2X1 _2765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_428_),
    .B(_401_),
    .Y(_430_)
);

INVX1 _2766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[2]),
    .Y(_431_)
);

OAI21X1 _2767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_431_),
    .B(_197_),
    .C(_148_),
    .Y(_432_)
);

AOI21X1 _2768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[2]),
    .B(_323_),
    .C(_432_),
    .Y(_433_)
);

OAI21X1 _2769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1291_),
    .B(_325_),
    .C(DIMUX[2]),
    .Y(_434_)
);

AOI22X1 _2770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_925_),
    .B(ABH[2]),
    .C(PC[10]),
    .D(_312_),
    .Y(_435_)
);

AND2X2 _2771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_434_),
    .B(_435_),
    .Y(_436_)
);

AND2X2 _2772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_436_),
    .B(_433_),
    .Y(_437_)
);

MUX2X1 _2773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_437_),
    .B(_280_),
    .S(_352_),
    .Y(_438_)
);

NOR2X1 _2774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_438_),
    .B(_430_),
    .Y(_439_)
);

NAND3X1 _2775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_409_),
    .B(_423_),
    .C(_417_),
    .Y(_440_)
);

NAND2X1 _2776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_280_),
    .B(_365_),
    .Y(_441_)
);

NAND2X1 _2777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_433_),
    .B(_436_),
    .Y(_442_)
);

OAI21X1 _2778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_365_),
    .B(_442_),
    .C(_441_),
    .Y(_443_)
);

OAI21X1 _2779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_443_),
    .B(_440_),
    .C(RDY_bF$buf9),
    .Y(_444_)
);

OAI22X1 _2780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_280_),
    .C(_444_),
    .D(_439_),
    .Y(_12_)
);

OAI21X1 _2781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1291_),
    .B(_325_),
    .C(DIMUX[3]),
    .Y(_445_)
);

AOI21X1 _2782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[3]),
    .B(_1299_),
    .C(_1334_),
    .Y(_446_)
);

NAND3X1 _2783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1110_),
    .B(_445_),
    .C(_446_),
    .Y(_447_)
);

INVX1 _2784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[3]),
    .Y(_448_)
);

MUX2X1 _2785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_448_),
    .B(_285_),
    .S(_1154_),
    .Y(_449_)
);

AOI21X1 _2786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1037_),
    .B(_449_),
    .C(_447_),
    .Y(_450_)
);

OAI21X1 _2787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_285_),
    .B(_352_),
    .C(_450_),
    .Y(_451_)
);

AOI21X1 _2788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_430_),
    .B(_438_),
    .C(_451_),
    .Y(_452_)
);

NAND2X1 _2789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[8]),
    .B(_365_),
    .Y(_453_)
);

NAND2X1 _2790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[11]),
    .B(_365_),
    .Y(_454_)
);

AOI22X1 _2791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_408_),
    .B(_453_),
    .C(_450_),
    .D(_454_),
    .Y(_455_)
);

NAND3X1 _2792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_455_),
    .B(_423_),
    .C(_438_),
    .Y(_456_)
);

OAI21X1 _2793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_456_),
    .B(_401_),
    .C(RDY_bF$buf7),
    .Y(_457_)
);

OAI22X1 _2794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf6),
    .B(_285_),
    .C(_457_),
    .D(_452_),
    .Y(_13_)
);

NAND2X1 _2795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[12]),
    .B(_886__bF$buf1),
    .Y(_458_)
);

OAI21X1 _2796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_290_),
    .B(_313_),
    .C(_1118_),
    .Y(_459_)
);

AOI21X1 _2797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[4]),
    .B(_1299_),
    .C(_1334_),
    .Y(_460_)
);

OAI21X1 _2798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_291_),
    .B(_378_),
    .C(_460_),
    .Y(_461_)
);

NOR2X1 _2799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_459_),
    .B(_461_),
    .Y(_462_)
);

OAI21X1 _2800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_888_),
    .B(_351_),
    .C(_462_),
    .Y(_463_)
);

NOR2X1 _2801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_290_),
    .B(_352_),
    .Y(_464_)
);

NOR2X1 _2802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_464_),
    .B(_463_),
    .Y(_465_)
);

NOR3X1 _2803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_456_),
    .B(_416_),
    .C(_370_),
    .Y(_466_)
);

NAND2X1 _2804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_465_),
    .B(_466_),
    .Y(_467_)
);

NOR2X1 _2805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_362_),
    .B(_340_),
    .Y(_468_)
);

NAND2X1 _2806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_392_),
    .B(_399_),
    .Y(_469_)
);

NOR2X1 _2807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_385_),
    .B(_469_),
    .Y(_470_)
);

NAND2X1 _2808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_276_),
    .B(_365_),
    .Y(_471_)
);

OAI21X1 _2809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1291_),
    .B(_325_),
    .C(DIMUX[1]),
    .Y(_472_)
);

INVX1 _2810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[1]),
    .Y(_473_)
);

OAI21X1 _2811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_197_),
    .C(_148_),
    .Y(_474_)
);

AOI21X1 _2812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABH[1]),
    .B(_323_),
    .C(_474_),
    .Y(_475_)
);

AOI21X1 _2813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(PC[9]),
    .B(_312_),
    .C(_1093_),
    .Y(_476_)
);

NAND3X1 _2814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_472_),
    .B(_476_),
    .C(_475_),
    .Y(_477_)
);

OAI21X1 _2815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_365_),
    .B(_477_),
    .C(_471_),
    .Y(_478_)
);

AND2X2 _2816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_445_),
    .B(_1110_),
    .Y(_479_)
);

NAND2X1 _2817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1037_),
    .B(_449_),
    .Y(_480_)
);

NAND3X1 _2818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_446_),
    .B(_480_),
    .C(_479_),
    .Y(_481_)
);

NOR2X1 _2819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_285_),
    .B(_352_),
    .Y(_482_)
);

OAI22X1 _2820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_481_),
    .B(_482_),
    .C(_427_),
    .D(_426_),
    .Y(_483_)
);

NOR3X1 _2821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_478_),
    .B(_443_),
    .C(_483_),
    .Y(_484_)
);

NAND3X1 _2822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_468_),
    .B(_470_),
    .C(_484_),
    .Y(_485_)
);

OAI21X1 _2823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_463_),
    .B(_464_),
    .C(_485_),
    .Y(_486_)
);

AND2X2 _2824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_467_),
    .B(_486_),
    .Y(_487_)
);

OAI21X1 _2825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf0),
    .B(_487_),
    .C(_458_),
    .Y(_14_)
);

INVX1 _2826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_465_),
    .Y(_488_)
);

OAI21X1 _2827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_295_),
    .B(_313_),
    .C(_1126_),
    .Y(_489_)
);

AOI21X1 _2828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[5]),
    .B(_1299_),
    .C(_1334_),
    .Y(_490_)
);

OAI21X1 _2829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_296_),
    .B(_378_),
    .C(_490_),
    .Y(_491_)
);

NOR2X1 _2830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_489_),
    .B(_491_),
    .Y(_492_)
);

OAI21X1 _2831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1013_),
    .B(_351_),
    .C(_492_),
    .Y(_493_)
);

NOR2X1 _2832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_295_),
    .B(_352_),
    .Y(_494_)
);

NOR2X1 _2833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_494_),
    .B(_493_),
    .Y(_495_)
);

AOI21X1 _2834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_466_),
    .B(_488_),
    .C(_495_),
    .Y(_496_)
);

INVX1 _2835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_495_),
    .Y(_497_)
);

NOR3X1 _2836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_465_),
    .B(_497_),
    .C(_485_),
    .Y(_498_)
);

OAI21X1 _2837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_498_),
    .B(_496_),
    .C(RDY_bF$buf5),
    .Y(_499_)
);

OAI21X1 _2838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .B(_295_),
    .C(_499_),
    .Y(_15_)
);

NOR2X1 _2839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_465_),
    .B(_495_),
    .Y(_500_)
);

NOR2X1 _2840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_300_),
    .B(_418_),
    .Y(_501_)
);

NOR2X1 _2841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1334_),
    .B(_1135_),
    .Y(_502_)
);

AOI22X1 _2842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[6]),
    .B(_1299_),
    .C(_323_),
    .D(ABH[6]),
    .Y(_503_)
);

AND2X2 _2843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_502_),
    .B(_503_),
    .Y(_504_)
);

OAI21X1 _2844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1015_),
    .B(_351_),
    .C(_504_),
    .Y(_505_)
);

NOR2X1 _2845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_505_),
    .B(_501_),
    .Y(_506_)
);

NAND3X1 _2846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_500_),
    .B(_506_),
    .C(_466_),
    .Y(_507_)
);

OAI21X1 _2847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_493_),
    .B(_494_),
    .C(_488_),
    .Y(_508_)
);

INVX1 _2848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_506_),
    .Y(_509_)
);

OAI21X1 _2849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_508_),
    .B(_485_),
    .C(_509_),
    .Y(_510_)
);

NAND3X1 _2850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf3),
    .B(_510_),
    .C(_507_),
    .Y(_511_)
);

NAND2X1 _2851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf6),
    .B(_300_),
    .Y(_512_)
);

AND2X2 _2852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_511_),
    .B(_512_),
    .Y(_16_)
);

NOR3X1 _2853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_456_),
    .B(_508_),
    .C(_401_),
    .Y(_513_)
);

NOR2X1 _2854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_304_),
    .B(_418_),
    .Y(_514_)
);

NOR2X1 _2855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1334_),
    .B(_1145_),
    .Y(_515_)
);

AOI22X1 _2856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .B(_1299_),
    .C(_323_),
    .D(ABH[7]),
    .Y(_516_)
);

AND2X2 _2857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_515_),
    .B(_516_),
    .Y(_517_)
);

OAI21X1 _2858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .B(_351_),
    .C(_517_),
    .Y(_518_)
);

NOR2X1 _2859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_518_),
    .B(_514_),
    .Y(_519_)
);

NAND3X1 _2860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_509_),
    .B(_519_),
    .C(_513_),
    .Y(_520_)
);

INVX1 _2861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_519_),
    .Y(_521_)
);

NAND3X1 _2862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_500_),
    .B(_509_),
    .C(_466_),
    .Y(_522_)
);

AOI21X1 _2863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_522_),
    .B(_521_),
    .C(_886__bF$buf5),
    .Y(_523_)
);

AOI22X1 _2864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf4),
    .B(_304_),
    .C(_520_),
    .D(_523_),
    .Y(_17_)
);

INVX1 _2865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(NMI_1),
    .Y(_524_)
);

NAND3X1 _2866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(NMI),
    .B(_524_),
    .C(_1153_),
    .Y(_525_)
);

OAI21X1 _2867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1153_),
    .B(_1021_),
    .C(_525_),
    .Y(_18_)
);

NAND2X1 _2868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf2),
    .B(_1181_),
    .Y(_526_)
);

OAI21X1 _2869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf1),
    .B(_1373_),
    .C(_526_),
    .Y(_19_)
);

NAND2X1 _2870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(cond_code[1]),
    .B(_886__bF$buf3),
    .Y(_527_)
);

OAI21X1 _2871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf2),
    .B(_1412_),
    .C(_527_),
    .Y(_20_)
);

NAND2X1 _2872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(cond_code[2]),
    .B(_886__bF$buf1),
    .Y(_528_)
);

OAI21X1 _2873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf0),
    .B(_1185_),
    .C(_528_),
    .Y(_21_)
);

INVX1 _2874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(plp),
    .Y(_529_)
);

INVX2 _2875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1251_),
    .Y(_530_)
);

NOR2X1 _2876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf3),
    .B(_530_),
    .Y(_531_)
);

NAND2X1 _2877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1367_),
    .B(_531_),
    .Y(_532_)
);

OAI21X1 _2878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_529_),
    .B(_1150__bF$buf0),
    .C(_532_),
    .Y(_22_)
);

INVX1 _2879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_531_),
    .Y(_533_)
);

NOR2X1 _2880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1187_),
    .B(_1181_),
    .Y(_534_)
);

NAND2X1 _2881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1393_),
    .B(_534_),
    .Y(_535_)
);

OAI22X1 _2882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_147_),
    .B(_1150__bF$buf4),
    .C(_535_),
    .D(_533_),
    .Y(_23_)
);

OAI21X1 _2883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf6),
    .B(_1027__bF$buf4),
    .C(clc),
    .Y(_536_)
);

NAND2X1 _2884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1348_),
    .B(_1330_),
    .Y(_537_)
);

OR2X2 _2885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_530_),
    .B(_1366_),
    .Y(_538_)
);

OAI21X1 _2886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_537_),
    .B(_538_),
    .C(_536_),
    .Y(_24_)
);

INVX1 _2887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(sec),
    .Y(_539_)
);

NOR2X1 _2888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf3),
    .B(_526_),
    .Y(_540_)
);

NAND2X1 _2889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1179_),
    .B(_540_),
    .Y(_541_)
);

OAI22X1 _2890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_539_),
    .B(_1150__bF$buf3),
    .C(_541_),
    .D(_538_),
    .Y(_25_)
);

OAI21X1 _2891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf5),
    .B(_1027__bF$buf2),
    .C(cld),
    .Y(_542_)
);

NOR2X1 _2892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .B(_1412_),
    .Y(_543_)
);

NAND2X1 _2893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_1251_),
    .Y(_544_)
);

OAI21X1 _2894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_537_),
    .B(_544_),
    .C(_542_),
    .Y(_26_)
);

INVX1 _2895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(sed),
    .Y(_545_)
);

OAI22X1 _2896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_545_),
    .B(_1150__bF$buf2),
    .C(_541_),
    .D(_544_),
    .Y(_27_)
);

OAI21X1 _2897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf4),
    .B(_1027__bF$buf1),
    .C(cli),
    .Y(_546_)
);

NAND2X1 _2898_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1189_),
    .B(_1251_),
    .Y(_547_)
);

OAI21X1 _2899_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_537_),
    .B(_547_),
    .C(_546_),
    .Y(_28_)
);

INVX1 _2900_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(sei),
    .Y(_548_)
);

OAI22X1 _2901_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_548_),
    .B(_1150__bF$buf1),
    .C(_541_),
    .D(_547_),
    .Y(_29_)
);

OAI21X1 _2902_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf3),
    .B(_1027__bF$buf0),
    .C(clv),
    .Y(_549_)
);

NOR2X1 _2903_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .B(_1187_),
    .Y(_550_)
);

NAND2X1 _2904_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_550_),
    .Y(_551_)
);

NOR2X1 _2905_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1178_),
    .B(_551_),
    .Y(_552_)
);

INVX1 _2906_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_552_),
    .Y(_553_)
);

OAI21X1 _2907_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_553_),
    .B(_533_),
    .C(_549_),
    .Y(_30_)
);

NAND3X1 _2908_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1327_),
    .B(_1178_),
    .C(_1161_),
    .Y(_554_)
);

NAND3X1 _2909_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .B(_1412_),
    .C(_1181_),
    .Y(_555_)
);

NOR2X1 _2910_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_555_),
    .B(_554_),
    .Y(_556_)
);

INVX1 _2911_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_556_),
    .Y(_557_)
);

OAI21X1 _2912_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf2),
    .B(_1027__bF$buf4),
    .C(bit_ins),
    .Y(_558_)
);

OAI21X1 _2913_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf2),
    .B(_557_),
    .C(_558_),
    .Y(_31_)
);

NOR2X1 _2914_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1412_),
    .B(_1348_),
    .Y(_559_)
);

NOR2X1 _2915_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1217_),
    .B(_559_),
    .Y(_560_)
);

AND2X2 _2916_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_560_),
    .B(_1405_),
    .Y(_561_)
);

OAI21X1 _2917_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1217_),
    .B(_1396_),
    .C(_557_),
    .Y(_562_)
);

AOI21X1 _2918_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_561_),
    .C(_562_),
    .Y(_563_)
);

NOR2X1 _2919_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1217_),
    .B(_1396_),
    .Y(_564_)
);

INVX1 _2920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_564_),
    .Y(_565_)
);

NOR2X1 _2921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_556_),
    .B(_561_),
    .Y(_566_)
);

AOI21X1 _2922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_566_),
    .B(_565_),
    .C(_1149__bF$buf1),
    .Y(_567_)
);

AOI22X1 _2923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_1149__bF$buf0),
    .C(_567_),
    .D(_563_),
    .Y(_32_)
);

NAND2X1 _2924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1187_),
    .B(_1348_),
    .Y(_568_)
);

NOR2X1 _2925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1215_),
    .B(_568_),
    .Y(_569_)
);

OAI21X1 _2926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1395_),
    .B(_569_),
    .C(_1185_),
    .Y(_570_)
);

AOI22X1 _2927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_132_),
    .B(_1149__bF$buf4),
    .C(_567_),
    .D(_570_),
    .Y(_33_)
);

INVX1 _2928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(op[2]),
    .Y(_571_)
);

AND2X2 _2929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_1178_),
    .Y(_572_)
);

NAND2X1 _2930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1164_),
    .B(_1178_),
    .Y(_573_)
);

NOR2X1 _2931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1160_),
    .B(_573_),
    .Y(_574_)
);

AOI22X1 _2932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_574_),
    .C(_572_),
    .D(_1351_),
    .Y(_575_)
);

NAND2X1 _2933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1327_),
    .B(_1395_),
    .Y(_576_)
);

OAI21X1 _2934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_576_),
    .C(_1215_),
    .Y(_577_)
);

INVX2 _2935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1397_),
    .Y(_578_)
);

NAND2X1 _2936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_1182_),
    .Y(_579_)
);

OR2X2 _2937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_578_),
    .B(_579_),
    .Y(_580_)
);

NAND2X1 _2938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_550_),
    .B(_1182_),
    .Y(_581_)
);

OAI21X1 _2939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_530_),
    .B(_581_),
    .C(_580_),
    .Y(_582_)
);

AOI21X1 _2940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_577_),
    .C(_582_),
    .Y(_583_)
);

AND2X2 _2941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_583_),
    .B(_575_),
    .Y(_584_)
);

AOI21X1 _2942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1395_),
    .B(_1189_),
    .C(_1149__bF$buf3),
    .Y(_585_)
);

AND2X2 _2943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_566_),
    .B(_585_),
    .Y(_586_)
);

AOI22X1 _2944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_571_),
    .B(_1149__bF$buf2),
    .C(_584_),
    .D(_586_),
    .Y(_34_)
);

INVX1 _2945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_567_),
    .Y(_587_)
);

OAI21X1 _2946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_140_),
    .B(_1150__bF$buf0),
    .C(_587_),
    .Y(_35_)
);

OAI21X1 _2947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1212_),
    .B(_1327_),
    .C(_540_),
    .Y(_588_)
);

OAI22X1 _2948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_920_),
    .B(_1150__bF$buf4),
    .C(_588_),
    .D(_565_),
    .Y(_36_)
);

AOI21X1 _2949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_310_),
    .B(_1149__bF$buf1),
    .C(_585_),
    .Y(_37_)
);

NOR2X1 _2950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1185_),
    .B(_1149__bF$buf0),
    .Y(_589_)
);

AOI22X1 _2951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(compare),
    .B(_1149__bF$buf4),
    .C(_569_),
    .D(_589_),
    .Y(_590_)
);

OAI21X1 _2952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf3),
    .B(_575_),
    .C(_590_),
    .Y(_38_)
);

NAND2X1 _2953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf3),
    .B(_564_),
    .Y(_591_)
);

OAI22X1 _2954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_895_),
    .B(_1150__bF$buf2),
    .C(_1174_),
    .D(_591_),
    .Y(_39_)
);

OAI21X1 _2955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1037_),
    .B(_1263_),
    .C(RDY_bF$buf0),
    .Y(_592_)
);

INVX1 _2956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_592_),
    .Y(_593_)
);

NAND2X1 _2957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(D),
    .B(_1185_),
    .Y(_594_)
);

NAND3X1 _2958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_559_),
    .B(_1405_),
    .C(_593_),
    .Y(_595_)
);

OAI22X1 _2959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_309_),
    .B(_593_),
    .C(_594_),
    .D(_595_),
    .Y(_40_)
);

OAI21X1 _2960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_308_),
    .B(_593_),
    .C(_595_),
    .Y(_41_)
);

INVX1 _2961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_576_),
    .Y(_596_)
);

NAND3X1 _2962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_543_),
    .C(_596_),
    .Y(_597_)
);

AOI22X1 _2963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(inc),
    .B(_1149__bF$buf2),
    .C(_531_),
    .D(_572_),
    .Y(_598_)
);

OAI21X1 _2964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf1),
    .B(_597_),
    .C(_598_),
    .Y(_42_)
);

OAI21X1 _2965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf1),
    .B(_1027__bF$buf3),
    .C(load_only),
    .Y(_599_)
);

OAI21X1 _2966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf0),
    .B(_551_),
    .C(_599_),
    .Y(_43_)
);

NAND2X1 _2967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf1),
    .B(_596_),
    .Y(_600_)
);

OAI22X1 _2968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1207_),
    .B(_1150__bF$buf0),
    .C(_550_),
    .D(_600_),
    .Y(_44_)
);

INVX1 _2969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_589_),
    .Y(_601_)
);

OAI21X1 _2970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_886__bF$buf0),
    .B(_1027__bF$buf2),
    .C(store),
    .Y(_602_)
);

NOR2X1 _2971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1172_),
    .B(_1214_),
    .Y(_603_)
);

OAI21X1 _2972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1405_),
    .B(_603_),
    .C(_534_),
    .Y(_604_)
);

OAI21X1 _2973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_601_),
    .B(_604_),
    .C(_602_),
    .Y(_45_)
);

INVX1 _2974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_550_),
    .Y(_605_)
);

NOR2X1 _2975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1178_),
    .B(_605_),
    .Y(_606_)
);

AOI21X1 _2976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_596_),
    .B(_606_),
    .C(_1326_),
    .Y(_607_)
);

AOI22X1 _2977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(index_y),
    .B(_1149__bF$buf4),
    .C(_1332_),
    .D(_1330_),
    .Y(_608_)
);

OAI21X1 _2978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1149__bF$buf3),
    .B(_607_),
    .C(_608_),
    .Y(_46_)
);

NOR2X1 _2979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_605_),
    .Y(_609_)
);

INVX1 _2980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_609_),
    .Y(_610_)
);

OAI21X1 _2981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1172_),
    .B(_610_),
    .C(_579_),
    .Y(_611_)
);

NAND2X1 _2982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1348_),
    .B(_606_),
    .Y(_612_)
);

NAND2X1 _2983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1217_),
    .B(_1182_),
    .Y(_613_)
);

NOR2X1 _2984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_613_),
    .B(_530_),
    .Y(_614_)
);

INVX1 _2985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_614_),
    .Y(_615_)
);

OAI21X1 _2986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_530_),
    .B(_612_),
    .C(_615_),
    .Y(_616_)
);

AOI21X1 _2987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1161_),
    .B(_611_),
    .C(_616_),
    .Y(_617_)
);

OAI21X1 _2988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_578_),
    .B(_553_),
    .C(_617_),
    .Y(_618_)
);

NAND2X1 _2989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1150__bF$buf4),
    .B(_618_),
    .Y(_619_)
);

OAI21X1 _2990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1055_),
    .B(_1150__bF$buf3),
    .C(_619_),
    .Y(_47_)
);

OAI21X1 _2991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_579_),
    .B(_578_),
    .C(_1150__bF$buf2),
    .Y(_620_)
);

NAND2X1 _2992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1402_),
    .B(_559_),
    .Y(_621_)
);

OAI21X1 _2993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_596_),
    .B(_1397_),
    .C(_609_),
    .Y(_622_)
);

OAI21X1 _2994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1160_),
    .B(_621_),
    .C(_622_),
    .Y(_623_)
);

NOR2X1 _2995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_620_),
    .B(_623_),
    .Y(_624_)
);

AOI22X1 _2996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1017_),
    .B(_1149__bF$buf2),
    .C(_617_),
    .D(_624_),
    .Y(_48_)
);

OAI21X1 _2997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1327_),
    .B(_1178_),
    .C(_1161_),
    .Y(_625_)
);

OAI21X1 _2998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_551_),
    .B(_625_),
    .C(_615_),
    .Y(_626_)
);

OAI21X1 _2999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_612_),
    .B(_578_),
    .C(_1252_),
    .Y(_627_)
);

OAI21X1 _3000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_627_),
    .B(_626_),
    .C(_1150__bF$buf1),
    .Y(_628_)
);

OAI21X1 _3001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1042_),
    .B(_1150__bF$buf0),
    .C(_628_),
    .Y(_49_)
);

OAI21X1 _3002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1396_),
    .B(_551_),
    .C(_580_),
    .Y(_629_)
);

OAI21X1 _3003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_626_),
    .B(_629_),
    .C(_1150__bF$buf4),
    .Y(_630_)
);

INVX1 _3004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_621_),
    .Y(_631_)
);

AOI22X1 _3005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(dst_reg[1]),
    .B(_1149__bF$buf1),
    .C(_531_),
    .D(_631_),
    .Y(_632_)
);

NAND2X1 _3006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_632_),
    .B(_630_),
    .Y(_50_)
);

INVX1 _3007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(load_reg),
    .Y(_633_)
);

OAI22X1 _3008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1179_),
    .B(_530_),
    .C(_578_),
    .D(_553_),
    .Y(_634_)
);

NAND2X1 _3009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_603_),
    .B(_552_),
    .Y(_635_)
);

OAI21X1 _3010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1394_),
    .B(_578_),
    .C(_635_),
    .Y(_636_)
);

NOR2X1 _3011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_636_),
    .B(_634_),
    .Y(_637_)
);

NOR2X1 _3012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1214_),
    .B(_1213_),
    .Y(_638_)
);

NAND2X1 _3013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_638_),
    .B(_609_),
    .Y(_639_)
);

INVX1 _3014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_551_),
    .Y(_640_)
);

NAND3X1 _3015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1159_),
    .B(_1178_),
    .C(_640_),
    .Y(_641_)
);

OAI21X1 _3016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1181_),
    .B(_1185_),
    .C(_1405_),
    .Y(_642_)
);

NAND3X1 _3017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_642_),
    .B(_641_),
    .C(_639_),
    .Y(_643_)
);

NOR2X1 _3018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_643_),
    .B(_620_),
    .Y(_644_)
);

AOI22X1 _3019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_633_),
    .B(_1149__bF$buf0),
    .C(_637_),
    .D(_644_),
    .Y(_51_)
);

AND2X2 _3020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf1),
    .B(res),
    .Y(_52_)
);

OAI21X1 _3021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_950_),
    .B(_1063_),
    .C(RDY_bF$buf9),
    .Y(_645_)
);

NOR2X1 _3022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .Y(_646_)
);

INVX2 _3023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_646_),
    .Y(_647_)
);

OAI21X1 _3024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[0]),
    .Y(_648_)
);

OAI21X1 _3025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_966_),
    .B(_647_),
    .C(_648_),
    .Y(_53_)
);

OAI21X1 _3026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[1]),
    .Y(_649_)
);

OAI21X1 _3027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1006_),
    .B(_647_),
    .C(_649_),
    .Y(_54_)
);

OAI21X1 _3028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[2]),
    .Y(_650_)
);

OAI21X1 _3029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1008_),
    .B(_647_),
    .C(_650_),
    .Y(_55_)
);

OAI21X1 _3030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[3]),
    .Y(_651_)
);

OAI21X1 _3031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1010_),
    .B(_647_),
    .C(_651_),
    .Y(_56_)
);

OAI21X1 _3032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[4]),
    .Y(_652_)
);

OAI21X1 _3033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_888_),
    .B(_647_),
    .C(_652_),
    .Y(_57_)
);

OAI21X1 _3034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[5]),
    .Y(_653_)
);

OAI21X1 _3035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1013_),
    .B(_647_),
    .C(_653_),
    .Y(_58_)
);

OAI21X1 _3036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[6]),
    .Y(_654_)
);

OAI21X1 _3037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1015_),
    .B(_647_),
    .C(_654_),
    .Y(_59_)
);

OAI21X1 _3038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .B(_645_),
    .C(IRHOLD[7]),
    .Y(_655_)
);

OAI21X1 _3039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .B(_647_),
    .C(_655_),
    .Y(_60_)
);

OAI21X1 _3040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1168_),
    .B(_1150__bF$buf3),
    .C(_645_),
    .Y(_61_)
);

INVX1 _3041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(bit_ins),
    .Y(_656_)
);

OAI21X1 _3042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf2),
    .B(_954_),
    .C(_1027__bF$buf0),
    .Y(_657_)
);

INVX1 _3043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_657_),
    .Y(_658_)
);

OAI21X1 _3044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_656_),
    .B(_917_),
    .C(_658_),
    .Y(_659_)
);

INVX1 _3045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_659_),
    .Y(_660_)
);

NOR2X1 _3046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(plp),
    .B(_1027__bF$buf4),
    .Y(_661_)
);

INVX1 _3047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_661_),
    .Y(_662_)
);

NOR2X1 _3048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(clv),
    .B(_662_),
    .Y(_663_)
);

AOI21X1 _3049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_308_),
    .B(_663_),
    .C(_660_),
    .Y(_664_)
);

OAI21X1 _3050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_914__bF$buf3),
    .B(_989_),
    .C(DIMUX[6]),
    .Y(_665_)
);

NAND2X1 _3051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(plp),
    .B(ADD[6]),
    .Y(_666_)
);

OAI21X1 _3052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf3),
    .B(_666_),
    .C(_665_),
    .Y(_667_)
);

AND2X2 _3053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_663_),
    .B(AV),
    .Y(_668_)
);

OAI21X1 _3054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_667_),
    .B(_668_),
    .C(_664_),
    .Y(_669_)
);

OAI21X1 _3055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1374_),
    .B(_664_),
    .C(_669_),
    .Y(_62_)
);

NOR2X1 _3056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(plp),
    .B(cld),
    .Y(_670_)
);

NAND2X1 _3057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_545_),
    .B(_670_),
    .Y(_671_)
);

OAI21X1 _3058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1027__bF$buf2),
    .B(_671_),
    .C(_657_),
    .Y(_672_)
);

NAND2X1 _3059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(D),
    .B(_672_),
    .Y(_673_)
);

INVX1 _3060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_670_),
    .Y(_674_)
);

OAI21X1 _3061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_529_),
    .B(_355_),
    .C(_674_),
    .Y(_675_)
);

MUX2X1 _3062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_675_),
    .B(DIMUX[3]),
    .S(_956_),
    .Y(_676_)
);

OAI21X1 _3063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_672_),
    .B(_676_),
    .C(_673_),
    .Y(_63_)
);

NOR2X1 _3064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(cli),
    .B(_1444_),
    .Y(_677_)
);

NAND2X1 _3065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_548_),
    .B(_677_),
    .Y(_678_)
);

AOI21X1 _3066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_658_),
    .B(_1344_),
    .C(_661_),
    .Y(_679_)
);

OAI21X1 _3067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_988_),
    .B(_679_),
    .C(_678_),
    .Y(_680_)
);

NOR2X1 _3068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_431_),
    .B(_988_),
    .Y(_681_)
);

OAI21X1 _3069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_681_),
    .B(_677_),
    .C(_956_),
    .Y(_682_)
);

OAI21X1 _3070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1008_),
    .B(_956_),
    .C(_682_),
    .Y(_683_)
);

NOR2X1 _3071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1021_),
    .B(_683_),
    .Y(_684_)
);

NAND2X1 _3072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(I),
    .B(_680_),
    .Y(_685_)
);

OAI21X1 _3073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_680_),
    .B(_684_),
    .C(_685_),
    .Y(_64_)
);

OAI21X1 _3074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1055_),
    .B(_1036_),
    .C(_1045_),
    .Y(_686_)
);

NAND2X1 _3075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1051_),
    .B(_686_),
    .Y(_687_)
);

NAND2X1 _3076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_921_),
    .B(_661_),
    .Y(_688_)
);

AOI21X1 _3077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_687_),
    .B(load_reg),
    .C(_688_),
    .Y(_689_)
);

AOI21X1 _3078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1227_),
    .B(_660_),
    .C(_689_),
    .Y(_690_)
);

AOI21X1 _3079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_662_),
    .B(_1227_),
    .C(AN),
    .Y(_691_)
);

INVX1 _3080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .Y(_692_)
);

AOI21X1 _3081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(plp),
    .B(_692_),
    .C(_1027__bF$buf1),
    .Y(_693_)
);

AOI21X1 _3082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[7]),
    .B(_1027__bF$buf0),
    .C(_693_),
    .Y(_694_)
);

AOI21X1 _3083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1227_),
    .B(_694_),
    .C(_691_),
    .Y(_695_)
);

NAND2X1 _3084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_695_),
    .B(_690_),
    .Y(_696_)
);

OAI21X1 _3085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1377_),
    .B(_690_),
    .C(_696_),
    .Y(_65_)
);

INVX1 _3086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Z),
    .Y(_697_)
);

AOI22X1 _3087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1227_),
    .B(_658_),
    .C(_689_),
    .D(_656_),
    .Y(_698_)
);

MUX2X1 _3088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[1]),
    .B(AZ),
    .S(plp),
    .Y(_699_)
);

MUX2X1 _3089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_699_),
    .B(_1006_),
    .S(_956_),
    .Y(_700_)
);

MUX2X1 _3090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_700_),
    .B(AZ),
    .S(_1227_),
    .Y(_701_)
);

MUX2X1 _3091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_701_),
    .B(_697_),
    .S(_698_),
    .Y(_66_)
);

NOR2X1 _3092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(write_back),
    .B(_1027__bF$buf4),
    .Y(_702_)
);

NOR2X1 _3093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(adc_sbc),
    .B(compare),
    .Y(_703_)
);

NAND2X1 _3094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_895_),
    .B(_703_),
    .Y(_704_)
);

INVX1 _3095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_704_),
    .Y(_705_)
);

NOR2X1 _3096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(plp),
    .B(clc),
    .Y(_706_)
);

NAND3X1 _3097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_539_),
    .B(_706_),
    .C(_705_),
    .Y(_707_)
);

OAI21X1 _3098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_895_),
    .B(_1227_),
    .C(_956_),
    .Y(_708_)
);

AOI21X1 _3099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_702_),
    .B(_707_),
    .C(_708_),
    .Y(_709_)
);

NAND2X1 _3100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(C),
    .B(_709_),
    .Y(_710_)
);

AOI21X1 _3101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(plp),
    .B(ADD[0]),
    .C(_706_),
    .Y(_711_)
);

NAND2X1 _3102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_704_),
    .Y(_712_)
);

OAI21X1 _3103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_704_),
    .B(_711_),
    .C(_712_),
    .Y(_713_)
);

MUX2X1 _3104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_713_),
    .B(DIMUX[0]),
    .S(_956_),
    .Y(_714_)
);

OAI21X1 _3105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_709_),
    .B(_714_),
    .C(_710_),
    .Y(_67_)
);

INVX1 _3106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(backwards),
    .Y(_715_)
);

NAND2X1 _3107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(DI[7]),
    .Y(_716_)
);

OAI21X1 _3108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf7),
    .B(_715_),
    .C(_716_),
    .Y(_68_)
);

OAI21X1 _3109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_935_),
    .B(_992_),
    .C(_969_),
    .Y(_717_)
);

NAND3X1 _3110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_204_),
    .B(_717_),
    .C(_1022_),
    .Y(_718_)
);

NOR2X1 _3111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_633_),
    .B(_662_),
    .Y(_719_)
);

OAI21X1 _3112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_719_),
    .B(_718_),
    .C(RDY_bF$buf6),
    .Y(_720_)
);

INVX1 _3113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf3),
    .Y(_721_)
);

NAND3X1 _3114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1051_),
    .B(_721_),
    .C(_1053_),
    .Y(_722_)
);

NAND2X1 _3115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_966_),
    .B(_1319__bF$buf2),
    .Y(_723_)
);

OAI21X1 _3116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[0]),
    .B(_1319__bF$buf1),
    .C(_723_),
    .Y(_724_)
);

NAND2X1 _3117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [0]),
    .B(_722_),
    .Y(_725_)
);

OAI21X1 _3118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_724_),
    .C(_725_),
    .Y(_69_)
);

AND2X2 _3119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(adj_bcd),
    .B(adc_bcd),
    .Y(_726_)
);

NAND2X1 _3120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(HC),
    .B(_726_),
    .Y(_727_)
);

NAND2X1 _3121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(adj_bcd),
    .B(_309_),
    .Y(_728_)
);

OAI21X1 _3122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(HC),
    .B(_728_),
    .C(_727_),
    .Y(_729_)
);

INVX1 _3123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_727_),
    .Y(_730_)
);

NOR2X1 _3124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(HC),
    .B(_728_),
    .Y(_731_)
);

OAI21X1 _3125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_731_),
    .B(_730_),
    .C(ADD[1]),
    .Y(_732_)
);

INVX1 _3126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .Y(_733_)
);

NOR2X1 _3127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf0),
    .B(_733_),
    .Y(_734_)
);

OAI21X1 _3128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[1]),
    .B(_729_),
    .C(_734_),
    .Y(_735_)
);

OAI21X1 _3129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1006_),
    .B(_1018_),
    .C(_735_),
    .Y(_736_)
);

INVX1 _3130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_736_),
    .Y(_737_)
);

NAND2X1 _3131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [1]),
    .B(_722_),
    .Y(_738_)
);

OAI21X1 _3132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_737_),
    .C(_738_),
    .Y(_70_)
);

NOR2X1 _3133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_431_),
    .B(_727_),
    .Y(_739_)
);

NOR2X1 _3134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[2]),
    .B(_730_),
    .Y(_740_)
);

OR2X2 _3135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_740_),
    .B(_739_),
    .Y(_741_)
);

OAI21X1 _3136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .B(_741_),
    .C(_1018_),
    .Y(_742_)
);

AOI21X1 _3137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .B(_741_),
    .C(_742_),
    .Y(_743_)
);

AOI21X1 _3138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[2]),
    .B(_1319__bF$buf3),
    .C(_743_),
    .Y(_744_)
);

NAND2X1 _3139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [2]),
    .B(_722_),
    .Y(_745_)
);

OAI21X1 _3140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_744_),
    .C(_745_),
    .Y(_71_)
);

NOR2X1 _3141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .B(_741_),
    .Y(_746_)
);

NOR2X1 _3142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_739_),
    .B(_746_),
    .Y(_747_)
);

OAI21X1 _3143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(HC),
    .B(_728_),
    .C(_355_),
    .Y(_748_)
);

NAND2X1 _3144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[3]),
    .B(_731_),
    .Y(_749_)
);

NAND2X1 _3145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_748_),
    .B(_749_),
    .Y(_750_)
);

AND2X2 _3146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_747_),
    .B(_750_),
    .Y(_751_)
);

NOR2X1 _3147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_750_),
    .B(_747_),
    .Y(_752_)
);

NOR2X1 _3148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_752_),
    .B(_751_),
    .Y(_753_)
);

MUX2X1 _3149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_753_),
    .B(DIMUX[3]),
    .S(_1018_),
    .Y(_754_)
);

NAND2X1 _3150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [3]),
    .B(_722_),
    .Y(_755_)
);

OAI21X1 _3151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_754_),
    .C(_755_),
    .Y(_72_)
);

OAI21X1 _3152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf1),
    .B(_1075_),
    .C(_173_),
    .Y(_756_)
);

OAI21X1 _3153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[4]),
    .B(_1018_),
    .C(_756_),
    .Y(_757_)
);

NAND2X1 _3154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [4]),
    .B(_722_),
    .Y(_758_)
);

OAI21X1 _3155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_757_),
    .C(_758_),
    .Y(_73_)
);

NAND2X1 _3156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_726_),
    .Y(_759_)
);

OAI21X1 _3157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_728_),
    .C(_759_),
    .Y(_760_)
);

OR2X2 _3158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_760_),
    .B(ADD[5]),
    .Y(_761_)
);

INVX1 _3159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_759_),
    .Y(_762_)
);

NOR2X1 _3160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_728_),
    .Y(_763_)
);

OAI21X1 _3161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_763_),
    .B(_762_),
    .C(ADD[5]),
    .Y(_764_)
);

INVX1 _3162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_764_),
    .Y(_765_)
);

NOR2X1 _3163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf2),
    .B(_765_),
    .Y(_766_)
);

AOI22X1 _3164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[5]),
    .B(_1319__bF$buf1),
    .C(_766_),
    .D(_761_),
    .Y(_767_)
);

NAND2X1 _3165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [5]),
    .B(_722_),
    .Y(_768_)
);

OAI21X1 _3166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_767_),
    .C(_768_),
    .Y(_74_)
);

INVX1 _3167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[6]),
    .Y(_769_)
);

NOR2X1 _3168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_769_),
    .B(_759_),
    .Y(_770_)
);

NOR2X1 _3169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[6]),
    .B(_762_),
    .Y(_771_)
);

NOR2X1 _3170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_770_),
    .B(_771_),
    .Y(_772_)
);

NAND2X1 _3171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_765_),
    .B(_772_),
    .Y(_773_)
);

INVX1 _3172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_773_),
    .Y(_774_)
);

NOR2X1 _3173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1319__bF$buf0),
    .B(_774_),
    .Y(_775_)
);

OAI21X1 _3174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_765_),
    .B(_772_),
    .C(_775_),
    .Y(_776_)
);

OAI21X1 _3175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1015_),
    .B(_1018_),
    .C(_776_),
    .Y(_777_)
);

INVX1 _3176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_777_),
    .Y(_778_)
);

NAND2X1 _3177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [6]),
    .B(_722_),
    .Y(_779_)
);

OAI21X1 _3178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_778_),
    .C(_779_),
    .Y(_75_)
);

OAI21X1 _3179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_769_),
    .B(_759_),
    .C(_773_),
    .Y(_780_)
);

OAI21X1 _3180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_728_),
    .C(_692_),
    .Y(_781_)
);

NAND2X1 _3181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .B(_763_),
    .Y(_782_)
);

NAND2X1 _3182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_781_),
    .B(_782_),
    .Y(_783_)
);

INVX1 _3183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_783_),
    .Y(_784_)
);

OAI21X1 _3184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_784_),
    .B(_780_),
    .C(_1018_),
    .Y(_785_)
);

AOI21X1 _3185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_780_),
    .B(_784_),
    .C(_785_),
    .Y(_786_)
);

AOI21X1 _3186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(DIMUX[7]),
    .B(_1319__bF$buf3),
    .C(_786_),
    .Y(_787_)
);

NAND2X1 _3187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[0] [7]),
    .B(_722_),
    .Y(_788_)
);

OAI21X1 _3188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_787_),
    .C(_788_),
    .Y(_76_)
);

NAND2X1 _3189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_721_),
    .B(_1047_),
    .Y(_789_)
);

OAI21X1 _3190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf2),
    .B(_687_),
    .C(\AXYS[1] [0]),
    .Y(_790_)
);

OAI21X1 _3191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .B(_789_),
    .C(_790_),
    .Y(_77_)
);

OAI21X1 _3192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf1),
    .B(_687_),
    .C(\AXYS[1] [1]),
    .Y(_791_)
);

OAI21X1 _3193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_737_),
    .B(_789_),
    .C(_791_),
    .Y(_78_)
);

OAI21X1 _3194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf0),
    .B(_687_),
    .C(\AXYS[1] [2]),
    .Y(_792_)
);

OAI21X1 _3195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_744_),
    .B(_789_),
    .C(_792_),
    .Y(_79_)
);

OAI21X1 _3196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf3),
    .B(_687_),
    .C(\AXYS[1] [3]),
    .Y(_793_)
);

OAI21X1 _3197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_754_),
    .B(_789_),
    .C(_793_),
    .Y(_80_)
);

OAI21X1 _3198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf2),
    .B(_687_),
    .C(\AXYS[1] [4]),
    .Y(_794_)
);

OAI21X1 _3199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_757_),
    .B(_789_),
    .C(_794_),
    .Y(_81_)
);

OAI21X1 _3200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf1),
    .B(_687_),
    .C(\AXYS[1] [5]),
    .Y(_795_)
);

OAI21X1 _3201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_767_),
    .B(_789_),
    .C(_795_),
    .Y(_82_)
);

OAI21X1 _3202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf0),
    .B(_687_),
    .C(\AXYS[1] [6]),
    .Y(_796_)
);

OAI21X1 _3203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_778_),
    .B(_789_),
    .C(_796_),
    .Y(_83_)
);

OAI21X1 _3204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf3),
    .B(_687_),
    .C(\AXYS[1] [7]),
    .Y(_797_)
);

OAI21X1 _3205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_787_),
    .B(_789_),
    .C(_797_),
    .Y(_84_)
);

AND2X2 _3206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1057_),
    .B(_721_),
    .Y(_798_)
);

NOR2X1 _3207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [0]),
    .B(_798_),
    .Y(_799_)
);

AOI21X1 _3208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .B(_798_),
    .C(_799_),
    .Y(_85_)
);

NOR2X1 _3209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [1]),
    .B(_798_),
    .Y(_800_)
);

AOI21X1 _3210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_737_),
    .B(_798_),
    .C(_800_),
    .Y(_86_)
);

NOR2X1 _3211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [2]),
    .B(_798_),
    .Y(_801_)
);

AOI21X1 _3212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_744_),
    .B(_798_),
    .C(_801_),
    .Y(_87_)
);

NOR2X1 _3213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [3]),
    .B(_798_),
    .Y(_802_)
);

AOI21X1 _3214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_754_),
    .B(_798_),
    .C(_802_),
    .Y(_88_)
);

NOR2X1 _3215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [4]),
    .B(_798_),
    .Y(_803_)
);

AOI21X1 _3216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_757_),
    .B(_798_),
    .C(_803_),
    .Y(_89_)
);

NOR2X1 _3217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [5]),
    .B(_798_),
    .Y(_804_)
);

AOI21X1 _3218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_767_),
    .B(_798_),
    .C(_804_),
    .Y(_90_)
);

NOR2X1 _3219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [6]),
    .B(_798_),
    .Y(_805_)
);

AOI21X1 _3220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_778_),
    .B(_798_),
    .C(_805_),
    .Y(_91_)
);

NOR2X1 _3221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\AXYS[2] [7]),
    .B(_798_),
    .Y(_806_)
);

AOI21X1 _3222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_787_),
    .B(_798_),
    .C(_806_),
    .Y(_92_)
);

NAND2X1 _3223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_721_),
    .B(_1049_),
    .Y(_807_)
);

INVX2 _3224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1049_),
    .Y(_808_)
);

OAI21X1 _3225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf2),
    .B(_808_),
    .C(\AXYS[3] [0]),
    .Y(_809_)
);

OAI21X1 _3226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .B(_807_),
    .C(_809_),
    .Y(_93_)
);

OAI21X1 _3227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf1),
    .B(_808_),
    .C(\AXYS[3] [1]),
    .Y(_810_)
);

OAI21X1 _3228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_737_),
    .B(_807_),
    .C(_810_),
    .Y(_94_)
);

OAI21X1 _3229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf0),
    .B(_808_),
    .C(\AXYS[3] [2]),
    .Y(_811_)
);

OAI21X1 _3230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_744_),
    .B(_807_),
    .C(_811_),
    .Y(_95_)
);

OAI21X1 _3231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf3),
    .B(_808_),
    .C(\AXYS[3] [3]),
    .Y(_812_)
);

OAI21X1 _3232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_754_),
    .B(_807_),
    .C(_812_),
    .Y(_96_)
);

OAI21X1 _3233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf2),
    .B(_808_),
    .C(\AXYS[3] [4]),
    .Y(_813_)
);

OAI21X1 _3234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_757_),
    .B(_807_),
    .C(_813_),
    .Y(_97_)
);

OAI21X1 _3235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf1),
    .B(_808_),
    .C(\AXYS[3] [5]),
    .Y(_814_)
);

OAI21X1 _3236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_767_),
    .B(_807_),
    .C(_814_),
    .Y(_98_)
);

OAI21X1 _3237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf0),
    .B(_808_),
    .C(\AXYS[3] [6]),
    .Y(_815_)
);

OAI21X1 _3238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_778_),
    .B(_807_),
    .C(_815_),
    .Y(_99_)
);

OAI21X1 _3239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720__bF$buf3),
    .B(_808_),
    .C(\AXYS[3] [7]),
    .Y(_816_)
);

OAI21X1 _3240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_787_),
    .B(_807_),
    .C(_816_),
    .Y(_100_)
);

OAI21X1 _3241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf0),
    .B(_1069_),
    .C(_1202_),
    .Y(_817_)
);

OAI21X1 _3242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf4),
    .B(_928_),
    .C(_1027__bF$buf3),
    .Y(_818_)
);

NOR2X1 _3243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_818_),
    .B(_817_),
    .Y(_819_)
);

OAI21X1 _3244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_902__bF$buf1),
    .B(_928_),
    .C(_1272_),
    .Y(_820_)
);

AOI21X1 _3245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_993_),
    .C(_820_),
    .Y(_821_)
);

AND2X2 _3246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_819_),
    .B(_821_),
    .Y(_822_)
);

INVX1 _3247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1030_),
    .Y(_823_)
);

OAI21X1 _3248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_935_),
    .B(_941_),
    .C(_823_),
    .Y(_824_)
);

AND2X2 _3249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1200_),
    .B(_824_),
    .Y(_825_)
);

NAND3X1 _3250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_130_),
    .B(_825_),
    .C(_822_),
    .Y(_826_)
);

OR2X2 _3251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1257_),
    .B(_818_),
    .Y(_827_)
);

NOR2X1 _3252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_817_),
    .B(_827_),
    .Y(_828_)
);

OAI21X1 _3253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .B(_1272_),
    .C(_1061_),
    .Y(_829_)
);

NOR2X1 _3254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1070_),
    .B(_829_),
    .Y(_830_)
);

AOI22X1 _3255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1303_),
    .B(_822_),
    .C(_828_),
    .D(_830_),
    .Y(_831_)
);

OAI21X1 _3256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf3),
    .B(_942_),
    .C(_974_),
    .Y(_832_)
);

NOR2X1 _3257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_950_),
    .B(_832_),
    .Y(_833_)
);

NAND3X1 _3258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_148_),
    .B(_1067_),
    .C(_833_),
    .Y(_834_)
);

OAI21X1 _3259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_834_),
    .B(_831_),
    .C(_826_),
    .Y(_835_)
);

AOI21X1 _3260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1221_),
    .B(_969_),
    .C(_1424_),
    .Y(_836_)
);

AND2X2 _3261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_836_),
    .B(_1019_),
    .Y(_837_)
);

NAND3X1 _3262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1022_),
    .B(_317_),
    .C(_837_),
    .Y(_838_)
);

OAI21X1 _3263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_952_),
    .B(_1360_),
    .C(_823_),
    .Y(_839_)
);

NOR2X1 _3264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1201_),
    .B(_1309_),
    .Y(_840_)
);

NAND3X1 _3265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_314_),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

NOR2X1 _3266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_841_),
    .B(_838_),
    .Y(_842_)
);

NAND2X1 _3267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_842_),
    .B(_835_),
    .Y(_843_)
);

OAI21X1 _3268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_977_),
    .B(_1427_),
    .C(_929_),
    .Y(_844_)
);

AND2X2 _3269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .B(_1019_),
    .Y(_845_)
);

NAND3X1 _3270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_840_),
    .B(_844_),
    .C(_845_),
    .Y(_846_)
);

NOR2X1 _3271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1021_),
    .B(_1235_),
    .Y(_847_)
);

OAI21X1 _3272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[5]),
    .B(state[4]),
    .C(_1225_),
    .Y(_848_)
);

NAND3X1 _3273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_848_),
    .B(_839_),
    .C(_847_),
    .Y(_849_)
);

OR2X2 _3274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_846_),
    .B(_849_),
    .Y(_850_)
);

OAI21X1 _3275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_931__bF$buf2),
    .B(_984_),
    .C(_210_),
    .Y(_851_)
);

NOR2X1 _3276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_975_),
    .B(_851_),
    .Y(_852_)
);

AND2X2 _3277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_836_),
    .B(_824_),
    .Y(_853_)
);

NAND3X1 _3278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_852_),
    .B(_853_),
    .C(_822_),
    .Y(_854_)
);

OAI21X1 _3279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .B(_854_),
    .C(_843_),
    .Y(_855_)
);

OAI21X1 _3280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_903__bF$buf2),
    .B(_969_),
    .C(_977_),
    .Y(_856_)
);

OAI21X1 _3281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(state[4]),
    .B(_981_),
    .C(_856_),
    .Y(_857_)
);

NOR2X1 _3282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_857_),
    .B(_1000_),
    .Y(_858_)
);

NAND2X1 _3283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_858_),
    .B(_855_),
    .Y(_859_)
);

NAND2X1 _3284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf5),
    .B(_859_),
    .Y(_860_)
);

NAND2X1 _3285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[0]),
    .B(_860_),
    .Y(_861_)
);

OAI21X1 _3286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .B(_225_),
    .C(_861_),
    .Y(_101_)
);

NAND2X1 _3287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[1]),
    .B(_860_),
    .Y(_862_)
);

OAI21X1 _3288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_231_),
    .B(_860_),
    .C(_862_),
    .Y(_102_)
);

NAND2X1 _3289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[2]),
    .B(_860_),
    .Y(_863_)
);

OAI21X1 _3290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .B(_236_),
    .C(_863_),
    .Y(_103_)
);

NAND2X1 _3291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[3]),
    .B(_860_),
    .Y(_864_)
);

OAI21X1 _3292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .B(_242_),
    .C(_864_),
    .Y(_104_)
);

NAND2X1 _3293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[4]),
    .B(_860_),
    .Y(_865_)
);

OAI21X1 _3294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .B(_249_),
    .C(_865_),
    .Y(_105_)
);

NAND2X1 _3295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[5]),
    .B(_860_),
    .Y(_866_)
);

OAI21X1 _3296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .B(_257_),
    .C(_866_),
    .Y(_106_)
);

NAND2X1 _3297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[6]),
    .B(_860_),
    .Y(_867_)
);

OAI21X1 _3298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_262_),
    .B(_860_),
    .C(_867_),
    .Y(_107_)
);

NAND2X1 _3299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABL[7]),
    .B(_860_),
    .Y(_868_)
);

OAI21X1 _3300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_267_),
    .B(_860_),
    .C(_868_),
    .Y(_108_)
);

AOI21X1 _3301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_855_),
    .B(_858_),
    .C(_886__bF$buf6),
    .Y(_869_)
);

NAND2X1 _3302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[8]),
    .B(_869_),
    .Y(_870_)
);

OAI21X1 _3303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_269_),
    .B(_869_),
    .C(_870_),
    .Y(_109_)
);

NAND2X1 _3304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[9]),
    .B(_869_),
    .Y(_871_)
);

OAI21X1 _3305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1091_),
    .B(_869_),
    .C(_871_),
    .Y(_110_)
);

NAND2X1 _3306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[10]),
    .B(_869_),
    .Y(_872_)
);

OAI21X1 _3307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1102_),
    .B(_869_),
    .C(_872_),
    .Y(_111_)
);

NAND2X1 _3308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[11]),
    .B(_869_),
    .Y(_873_)
);

OAI21X1 _3309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_448_),
    .B(_869_),
    .C(_873_),
    .Y(_112_)
);

NAND2X1 _3310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[12]),
    .B(_869_),
    .Y(_874_)
);

OAI21X1 _3311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_291_),
    .B(_869_),
    .C(_874_),
    .Y(_113_)
);

NAND2X1 _3312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[13]),
    .B(_869_),
    .Y(_875_)
);

OAI21X1 _3313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_296_),
    .B(_869_),
    .C(_875_),
    .Y(_114_)
);

NAND2X1 _3314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[14]),
    .B(_869_),
    .Y(_876_)
);

OAI21X1 _3315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1134_),
    .B(_869_),
    .C(_876_),
    .Y(_115_)
);

NAND2X1 _3316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[15]),
    .B(_869_),
    .Y(_877_)
);

OAI21X1 _3317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1144_),
    .B(_869_),
    .C(_877_),
    .Y(_116_)
);

DFFSR _3318_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_1512_[0]),
    .Q(state[0]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3319_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_1512_[1]),
    .Q(state[1]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3320_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_1512_[2]),
    .Q(state[2]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3321_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_1512_[3]),
    .Q(state[3]),
    .R(vdd),
    .S(_1__bF$buf7)
);

DFFSR _3322_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_1512_[4]),
    .Q(state[4]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3323_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_1512_[5]),
    .Q(state[5]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3324_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_2_),
    .Q(PC[0]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3325_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_3_),
    .Q(PC[1]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3326_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_4_),
    .Q(PC[2]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3327_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_5_),
    .Q(PC[3]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3328_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_6_),
    .Q(PC[4]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3329_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_7_),
    .Q(PC[5]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3330_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_8_),
    .Q(PC[6]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3331_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_9_),
    .Q(PC[7]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3332_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_10_),
    .Q(PC[8]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3333_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_11_),
    .Q(PC[9]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3334_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_12_),
    .Q(PC[10]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3335_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_13_),
    .Q(PC[11]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3336_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_14_),
    .Q(PC[12]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3337_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_15_),
    .Q(PC[13]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3338_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_16_),
    .Q(PC[14]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3339_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_17_),
    .Q(PC[15]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3340_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(NMI),
    .Q(NMI_1),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3341_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_18_),
    .Q(NMI_edge),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3342_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_19_),
    .Q(cond_code[0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3343_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_20_),
    .Q(cond_code[1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3344_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_21_),
    .Q(cond_code[2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3345_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_22_),
    .Q(plp),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3346_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_23_),
    .Q(php),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3347_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_24_),
    .Q(clc),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3348_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_25_),
    .Q(sec),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3349_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_26_),
    .Q(cld),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3350_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_27_),
    .Q(sed),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3351_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_28_),
    .Q(cli),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3352_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_29_),
    .Q(sei),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3353_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_30_),
    .Q(clv),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3354_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_31_),
    .Q(bit_ins),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3355_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_32_),
    .Q(op[0]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3356_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_33_),
    .Q(op[1]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3357_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_34_),
    .Q(op[2]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3358_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_35_),
    .Q(op[3]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3359_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_36_),
    .Q(rotate),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3360_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_37_),
    .Q(shift_right),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3361_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_38_),
    .Q(compare),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3362_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_39_),
    .Q(shift),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3363_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_40_),
    .Q(adc_bcd),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3364_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_41_),
    .Q(adc_sbc),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3365_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_42_),
    .Q(inc),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3366_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_43_),
    .Q(load_only),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3367_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_44_),
    .Q(write_back),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3368_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_45_),
    .Q(store),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3369_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_46_),
    .Q(index_y),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3370_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_47_),
    .Q(src_reg[0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3371_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_48_),
    .Q(src_reg[1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3372_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_49_),
    .Q(dst_reg[0]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3373_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_50_),
    .Q(dst_reg[1]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3374_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_51_),
    .Q(load_reg),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3375_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(DIMUX[0]),
    .Q(DIHOLD[0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3376_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(DIMUX[1]),
    .Q(DIHOLD[1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3377_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(DIMUX[2]),
    .Q(DIHOLD[2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3378_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(DIMUX[3]),
    .Q(DIHOLD[3]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3379_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(DIMUX[4]),
    .Q(DIHOLD[4]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3380_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(DIMUX[5]),
    .Q(DIHOLD[5]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3381_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(DIMUX[6]),
    .Q(DIHOLD[6]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3382_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(DIMUX[7]),
    .Q(DIHOLD[7]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3383_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_52_),
    .Q(res),
    .R(vdd),
    .S(_1__bF$buf0)
);

DFFPOSX1 _3384_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_53_),
    .Q(IRHOLD[0])
);

DFFPOSX1 _3385_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_54_),
    .Q(IRHOLD[1])
);

DFFPOSX1 _3386_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_55_),
    .Q(IRHOLD[2])
);

DFFPOSX1 _3387_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_56_),
    .Q(IRHOLD[3])
);

DFFPOSX1 _3388_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_57_),
    .Q(IRHOLD[4])
);

DFFPOSX1 _3389_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_58_),
    .Q(IRHOLD[5])
);

DFFPOSX1 _3390_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_59_),
    .Q(IRHOLD[6])
);

DFFPOSX1 _3391_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_60_),
    .Q(IRHOLD[7])
);

DFFSR _3392_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_61_),
    .Q(IRHOLD_valid),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3393_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_62_),
    .Q(V),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3394_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_63_),
    .Q(D),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3395_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_64_),
    .Q(I),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3396_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_65_),
    .Q(N),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3397_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_66_),
    .Q(Z),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3398_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_67_),
    .Q(C),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3399_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_68_),
    .Q(backwards),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3400_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_69_),
    .Q(\AXYS[0] [0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3401_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_70_),
    .Q(\AXYS[0] [1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3402_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_71_),
    .Q(\AXYS[0] [2]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3403_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_72_),
    .Q(\AXYS[0] [3]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3404_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_73_),
    .Q(\AXYS[0] [4]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3405_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_74_),
    .Q(\AXYS[0] [5]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3406_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_75_),
    .Q(\AXYS[0] [6]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3407_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_76_),
    .Q(\AXYS[0] [7]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3408_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_77_),
    .Q(\AXYS[1] [0]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3409_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_78_),
    .Q(\AXYS[1] [1]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3410_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_79_),
    .Q(\AXYS[1] [2]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3411_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_80_),
    .Q(\AXYS[1] [3]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3412_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_81_),
    .Q(\AXYS[1] [4]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3413_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_82_),
    .Q(\AXYS[1] [5]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3414_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_83_),
    .Q(\AXYS[1] [6]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3415_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_84_),
    .Q(\AXYS[1] [7]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3416_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_85_),
    .Q(\AXYS[2] [0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3417_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_86_),
    .Q(\AXYS[2] [1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3418_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_87_),
    .Q(\AXYS[2] [2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3419_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_88_),
    .Q(\AXYS[2] [3]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3420_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_89_),
    .Q(\AXYS[2] [4]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3421_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_90_),
    .Q(\AXYS[2] [5]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3422_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_91_),
    .Q(\AXYS[2] [6]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3423_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_92_),
    .Q(\AXYS[2] [7]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3424_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_0_),
    .Q(adj_bcd),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3425_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_93_),
    .Q(\AXYS[3] [0]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3426_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_94_),
    .Q(\AXYS[3] [1]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3427_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_95_),
    .Q(\AXYS[3] [2]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3428_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_96_),
    .Q(\AXYS[3] [3]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3429_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_97_),
    .Q(\AXYS[3] [4]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3430_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_98_),
    .Q(\AXYS[3] [5]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3431_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_99_),
    .Q(\AXYS[3] [6]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3432_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_100_),
    .Q(\AXYS[3] [7]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3433_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_101_),
    .Q(ABL[0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3434_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_102_),
    .Q(ABL[1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3435_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_103_),
    .Q(ABL[2]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3436_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_104_),
    .Q(ABL[3]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3437_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_105_),
    .Q(ABL[4]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3438_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_106_),
    .Q(ABL[5]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3439_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_107_),
    .Q(ABL[6]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3440_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_108_),
    .Q(ABL[7]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3441_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_109_),
    .Q(ABH[0]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3442_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_110_),
    .Q(ABH[1]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3443_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_111_),
    .Q(ABH[2]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3444_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_112_),
    .Q(ABH[3]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3445_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_113_),
    .Q(ABH[4]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3446_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_114_),
    .Q(ABH[5]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3447_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_115_),
    .Q(ABH[6]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3448_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_116_),
    .Q(ABH[7]),
    .R(_1__bF$buf9),
    .S(vdd)
);

OR2X2 _3449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[0]),
    .B(ADD[3]),
    .Y(_1698_)
);

NOR2X1 _3450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[5]),
    .B(ADD[4]),
    .Y(_1699_)
);

NOR2X1 _3451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .B(ADD[6]),
    .Y(_1700_)
);

NOR2X1 _3452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[1]),
    .B(ADD[2]),
    .Y(_1701_)
);

NAND3X1 _3453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1699_),
    .B(_1700_),
    .C(_1701_),
    .Y(_1702_)
);

NOR2X1 _3454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1698_),
    .B(_1702_),
    .Y(AZ)
);

INVX1 _3455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .Y(_1703_)
);

AND2X2 _3456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1703_),
    .B(CO),
    .Y(_1704_)
);

NOR2X1 _3457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_1703_),
    .Y(_1705_)
);

NOR2X1 _3458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1705_),
    .B(_1704_),
    .Y(_1706_)
);

INVX1 _3459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .Y(_1707_)
);

NOR2X1 _3460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.BI7 ),
    .B(_1707_),
    .Y(_1708_)
);

NAND2X1 _3461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.BI7 ),
    .B(_1707_),
    .Y(_1709_)
);

INVX1 _3462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1709_),
    .Y(_1710_)
);

OAI21X1 _3463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1708_),
    .B(_1710_),
    .C(_1706_),
    .Y(_1711_)
);

NOR2X1 _3464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1708_),
    .B(_1710_),
    .Y(_1712_)
);

OAI21X1 _3465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1704_),
    .B(_1705_),
    .C(_1712_),
    .Y(_1713_)
);

NAND2X1 _3466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1711_),
    .B(_1713_),
    .Y(AV)
);

INVX4 _3467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .Y(_1513_)
);

INVX4 _3468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf4),
    .Y(_1714_)
);

NAND2X1 _3469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CI),
    .B(alu_shift_right),
    .Y(_1715_)
);

INVX2 _3470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[1]),
    .Y(_1716_)
);

NAND2X1 _3471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_1716_),
    .Y(_1717_)
);

INVX2 _3472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .Y(_1718_)
);

AND2X2 _3473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1718_),
    .B(BI[7]),
    .Y(_1719_)
);

NAND2X1 _3474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[7]),
    .B(_1719_),
    .Y(_1720_)
);

AOI22X1 _3475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[7]),
    .B(_1716_),
    .C(_1720_),
    .D(_1717_),
    .Y(_1721_)
);

INVX2 _3476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_shift_right),
    .Y(_1722_)
);

OAI21X1 _3477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[7]),
    .B(_1719_),
    .C(_1722_),
    .Y(_1723_)
);

OAI21X1 _3478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1723_),
    .B(_1721_),
    .C(_1715_),
    .Y(_1724_)
);

INVX4 _3479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .Y(_1725_)
);

OAI21X1 _3480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[7]),
    .B(alu_op[2]),
    .C(_1725_),
    .Y(_1726_)
);

AOI21X1 _3481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[7]),
    .B(alu_op[2]),
    .C(_1726_),
    .Y(_1727_)
);

NOR2X1 _3482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .B(_1725_),
    .Y(_1728_)
);

OR2X2 _3483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1727_),
    .B(_1728_),
    .Y(_1729_)
);

OAI21X1 _3484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1727_),
    .B(_1724_),
    .C(_1729_),
    .Y(_1730_)
);

NAND2X1 _3485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.BI7 ),
    .B(_1714__bF$buf3),
    .Y(_1731_)
);

OAI21X1 _3486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf2),
    .B(_1730_),
    .C(_1731_),
    .Y(_1514_)
);

NAND2X1 _3487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_1714__bF$buf1),
    .Y(_1732_)
);

NAND2X1 _3488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_shift_right),
    .B(AI[6]),
    .Y(_1733_)
);

AND2X2 _3489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1718_),
    .B(BI[5]),
    .Y(_1734_)
);

NAND2X1 _3490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .B(_1734_),
    .Y(_1735_)
);

AOI22X1 _3491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1716_),
    .B(BI[5]),
    .C(_1735_),
    .D(_1717_),
    .Y(_1736_)
);

OAI21X1 _3492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .B(_1734_),
    .C(_1722_),
    .Y(_1737_)
);

OAI21X1 _3493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1737_),
    .B(_1736_),
    .C(_1733_),
    .Y(_1738_)
);

NAND2X1 _3494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .B(_1725_),
    .Y(_1739_)
);

INVX2 _3495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .Y(_1740_)
);

OAI21X1 _3496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .B(BI[5]),
    .C(_1740_),
    .Y(_1526_)
);

OAI21X1 _3497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[5]),
    .B(_1739_),
    .C(_1526_),
    .Y(_1527_)
);

NAND2X1 _3498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_shift_right),
    .B(AI[5]),
    .Y(_1528_)
);

AND2X2 _3499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1718_),
    .B(BI[4]),
    .Y(_1529_)
);

NAND2X1 _3500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[4]),
    .B(_1529_),
    .Y(_1530_)
);

AOI22X1 _3501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1716_),
    .B(BI[4]),
    .C(_1530_),
    .D(_1717_),
    .Y(_1531_)
);

OAI21X1 _3502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[4]),
    .B(_1529_),
    .C(_1722_),
    .Y(_1532_)
);

OAI21X1 _3503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1532_),
    .B(_1531_),
    .C(_1528_),
    .Y(_1533_)
);

OAI21X1 _3504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .B(BI[4]),
    .C(_1740_),
    .Y(_1534_)
);

OAI21X1 _3505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[4]),
    .B(_1739_),
    .C(_1534_),
    .Y(_1535_)
);

NAND2X1 _3506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1535_),
    .B(_1533_),
    .Y(_1536_)
);

INVX1 _3507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[4]),
    .Y(_1537_)
);

INVX1 _3508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[3]),
    .Y(_1538_)
);

INVX1 _3509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[3]),
    .Y(_1539_)
);

NAND2X1 _3510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[3]),
    .B(_1718_),
    .Y(_1540_)
);

OAI21X1 _3511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1539_),
    .B(_1540_),
    .C(_1717_),
    .Y(_1541_)
);

OAI21X1 _3512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[1]),
    .B(_1538_),
    .C(_1541_),
    .Y(_1542_)
);

AOI21X1 _3513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1540_),
    .B(_1539_),
    .C(alu_shift_right),
    .Y(_1543_)
);

NAND2X1 _3514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1543_),
    .B(_1542_),
    .Y(_1544_)
);

OAI21X1 _3515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1722_),
    .B(_1537_),
    .C(_1544_),
    .Y(_1545_)
);

INVX1 _3516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1728_),
    .Y(_1546_)
);

OAI21X1 _3517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .B(BI[3]),
    .C(_1740_),
    .Y(_1547_)
);

OAI21X1 _3518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[3]),
    .B(_1739_),
    .C(_1547_),
    .Y(_1548_)
);

AND2X2 _3519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1548_),
    .B(_1546_),
    .Y(_1549_)
);

OR2X2 _3520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1545_),
    .B(_1549_),
    .Y(_1550_)
);

NAND3X1 _3521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[2]),
    .B(AI[2]),
    .C(_1718_),
    .Y(_1551_)
);

AOI22X1 _3522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1716_),
    .B(BI[2]),
    .C(_1551_),
    .D(_1717_),
    .Y(_1552_)
);

INVX1 _3523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[2]),
    .Y(_1553_)
);

INVX1 _3524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[2]),
    .Y(_1554_)
);

OAI21X1 _3525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_1553_),
    .C(_1554_),
    .Y(_1555_)
);

NAND2X1 _3526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1722_),
    .B(_1555_),
    .Y(_1556_)
);

OAI22X1 _3527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1722_),
    .B(_1539_),
    .C(_1556_),
    .D(_1552_),
    .Y(_1557_)
);

NOR2X1 _3528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .B(alu_op[2]),
    .Y(_1558_)
);

AOI21X1 _3529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(_1553_),
    .C(_1740_),
    .Y(_1559_)
);

AOI21X1 _3530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1553_),
    .B(_1558_),
    .C(_1559_),
    .Y(_1560_)
);

NAND2X1 _3531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1560_),
    .B(_1557_),
    .Y(_1561_)
);

INVX1 _3532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1561_),
    .Y(_1562_)
);

NAND3X1 _3533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[1]),
    .B(AI[1]),
    .C(_1718_),
    .Y(_1563_)
);

AOI22X1 _3534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1716_),
    .B(BI[1]),
    .C(_1563_),
    .D(_1717_),
    .Y(_1564_)
);

INVX1 _3535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[1]),
    .Y(_1565_)
);

NOR2X1 _3536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_1565_),
    .Y(_1566_)
);

OAI21X1 _3537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[1]),
    .B(_1566_),
    .C(_1722_),
    .Y(_1567_)
);

OAI22X1 _3538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1722_),
    .B(_1554_),
    .C(_1564_),
    .D(_1567_),
    .Y(_1568_)
);

OAI21X1 _3539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1725_),
    .Y(_1569_)
);

AOI21X1 _3540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1569_),
    .Y(_1570_)
);

OAI21X1 _3541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1728_),
    .B(_1570_),
    .C(_1568_),
    .Y(_1571_)
);

NAND2X1 _3542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(_1718_),
    .Y(_1572_)
);

NAND2X1 _3543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[1]),
    .B(AI[0]),
    .Y(_1573_)
);

AOI22X1 _3544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(_1573_),
    .C(_1717_),
    .D(_1572_),
    .Y(_1574_)
);

INVX1 _3545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .Y(_1575_)
);

INVX1 _3546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[0]),
    .Y(_1576_)
);

OAI21X1 _3547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_1575_),
    .C(_1576_),
    .Y(_1577_)
);

NAND2X1 _3548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1722_),
    .B(_1577_),
    .Y(_1578_)
);

NAND2X1 _3549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_shift_right),
    .B(AI[1]),
    .Y(_1579_)
);

OAI21X1 _3550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1574_),
    .B(_1578_),
    .C(_1579_),
    .Y(_1580_)
);

OAI21X1 _3551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1725_),
    .Y(_1581_)
);

INVX1 _3552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1581_),
    .Y(_1582_)
);

OAI21X1 _3553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1740_),
    .B(_1575_),
    .C(_1582_),
    .Y(_1583_)
);

OAI21X1 _3554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1583_),
    .Y(_1584_)
);

OAI21X1 _3555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(_1740_),
    .C(CI),
    .Y(_1585_)
);

NOR2X1 _3556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_shift_right),
    .B(_1585_),
    .Y(_1586_)
);

MUX2X1 _3557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[1]),
    .B(_1575_),
    .S(alu_op[0]),
    .Y(_1587_)
);

NAND2X1 _3558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(_1573_),
    .Y(_1588_)
);

NAND2X1 _3559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1588_),
    .B(_1587_),
    .Y(_1589_)
);

AOI21X1 _3560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1572_),
    .B(_1576_),
    .C(alu_shift_right),
    .Y(_1590_)
);

NAND2X1 _3561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1590_),
    .B(_1589_),
    .Y(_1591_)
);

NAND3X1 _3562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1579_),
    .B(_1583_),
    .C(_1591_),
    .Y(_1592_)
);

AOI22X1 _3563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1580_),
    .B(_1584_),
    .C(_1592_),
    .D(_1586_),
    .Y(_1593_)
);

NOR2X1 _3564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1570_),
    .B(_1568_),
    .Y(_1594_)
);

OAI21X1 _3565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1594_),
    .B(_1593_),
    .C(_1571_),
    .Y(_1595_)
);

NAND2X1 _3566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(_1560_),
    .Y(_1596_)
);

INVX1 _3567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1596_),
    .Y(_1597_)
);

OAI21X1 _3568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1557_),
    .B(_1597_),
    .C(_1561_),
    .Y(_1598_)
);

INVX1 _3569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1598_),
    .Y(_1599_)
);

AND2X2 _3570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1595_),
    .B(_1599_),
    .Y(_1600_)
);

NAND2X1 _3571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1548_),
    .B(_1545_),
    .Y(_1601_)
);

OAI21X1 _3572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1545_),
    .B(_1549_),
    .C(_1601_),
    .Y(_1602_)
);

OAI21X1 _3573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1562_),
    .B(_1600_),
    .C(_1602_),
    .Y(_1603_)
);

AOI21X1 _3574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1595_),
    .B(_1599_),
    .C(_1562_),
    .Y(_1604_)
);

INVX1 _3575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1602_),
    .Y(_1605_)
);

NAND2X1 _3576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1605_),
    .B(_1604_),
    .Y(_1606_)
);

NAND2X1 _3577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1606_),
    .B(_1603_),
    .Y(_1607_)
);

INVX1 _3578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.BCD ),
    .Y(_1608_)
);

NAND2X1 _3579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1599_),
    .B(_1595_),
    .Y(_1609_)
);

AOI21X1 _3580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1581_),
    .Y(_1610_)
);

OAI21X1 _3581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1728_),
    .B(_1610_),
    .C(_1580_),
    .Y(_1611_)
);

INVX1 _3582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1586_),
    .Y(_1612_)
);

NOR2X1 _3583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1610_),
    .B(_1580_),
    .Y(_1613_)
);

OAI21X1 _3584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1612_),
    .B(_1613_),
    .C(_1611_),
    .Y(_1614_)
);

INVX1 _3585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1570_),
    .Y(_1615_)
);

OAI21X1 _3586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1615_),
    .Y(_1616_)
);

MUX2X1 _3587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1616_),
    .B(_1615_),
    .S(_1568_),
    .Y(_1617_)
);

NAND2X1 _3588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1617_),
    .B(_1614_),
    .Y(_1618_)
);

NAND3X1 _3589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1571_),
    .B(_1598_),
    .C(_1618_),
    .Y(_1619_)
);

NAND2X1 _3590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1609_),
    .B(_1619_),
    .Y(_1620_)
);

OAI21X1 _3591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1568_),
    .B(_1570_),
    .C(_1571_),
    .Y(_1621_)
);

NAND2X1 _3592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1593_),
    .B(_1621_),
    .Y(_1622_)
);

NAND2X1 _3593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1622_),
    .B(_1618_),
    .Y(_1623_)
);

AOI21X1 _3594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1620_),
    .B(_1623_),
    .C(_1608_),
    .Y(_1624_)
);

NAND2X1 _3595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1601_),
    .B(_1604_),
    .Y(_1625_)
);

AOI22X1 _3596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1550_),
    .B(_1625_),
    .C(_1607_),
    .D(_1624_),
    .Y(_1626_)
);

OAI21X1 _3597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1535_),
    .Y(_1627_)
);

INVX1 _3598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1627_),
    .Y(_1628_)
);

OAI21X1 _3599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1533_),
    .B(_1628_),
    .C(_1536_),
    .Y(_1629_)
);

OAI21X1 _3600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1629_),
    .B(_1626_),
    .C(_1536_),
    .Y(_1630_)
);

NAND2X1 _3601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1527_),
    .B(_1738_),
    .Y(_1631_)
);

OAI21X1 _3602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1527_),
    .Y(_1632_)
);

INVX1 _3603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1632_),
    .Y(_1633_)
);

OAI21X1 _3604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1738_),
    .B(_1633_),
    .C(_1631_),
    .Y(_1634_)
);

INVX1 _3605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1634_),
    .Y(_1635_)
);

AOI22X1 _3606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1738_),
    .B(_1527_),
    .C(_1630_),
    .D(_1635_),
    .Y(_1636_)
);

OAI21X1 _3607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1727_),
    .B(_1728_),
    .C(_1724_),
    .Y(_1637_)
);

OAI21X1 _3608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1724_),
    .B(_1727_),
    .C(_1637_),
    .Y(_1638_)
);

INVX1 _3609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1638_),
    .Y(_1639_)
);

NAND2X1 _3610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[7]),
    .B(alu_shift_right),
    .Y(_1640_)
);

AND2X2 _3611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1718_),
    .B(BI[6]),
    .Y(_1641_)
);

NAND2X1 _3612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[6]),
    .B(_1641_),
    .Y(_1642_)
);

AOI22X1 _3613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1716_),
    .B(BI[6]),
    .C(_1642_),
    .D(_1717_),
    .Y(_1643_)
);

OAI21X1 _3614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[6]),
    .B(_1641_),
    .C(_1722_),
    .Y(_1644_)
);

OAI21X1 _3615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1644_),
    .B(_1643_),
    .C(_1640_),
    .Y(_1645_)
);

OAI21X1 _3616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .B(BI[6]),
    .C(_1740_),
    .Y(_1646_)
);

OAI21X1 _3617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[6]),
    .B(_1739_),
    .C(_1646_),
    .Y(_1647_)
);

NAND2X1 _3618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1647_),
    .B(_1645_),
    .Y(_1648_)
);

INVX1 _3619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1648_),
    .Y(_1649_)
);

AOI22X1 _3620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1724_),
    .B(_1729_),
    .C(_1639_),
    .D(_1649_),
    .Y(_1650_)
);

OAI21X1 _3621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1647_),
    .Y(_1651_)
);

INVX1 _3622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1651_),
    .Y(_1652_)
);

OAI21X1 _3623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1645_),
    .B(_1652_),
    .C(_1648_),
    .Y(_1653_)
);

INVX1 _3624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1653_),
    .Y(_1654_)
);

NAND2X1 _3625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1654_),
    .B(_1639_),
    .Y(_1655_)
);

OAI21X1 _3626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1655_),
    .B(_1636_),
    .C(_1650_),
    .Y(_1656_)
);

NOR2X1 _3627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1722_),
    .B(_1576_),
    .Y(_1657_)
);

OR2X2 _3628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1656_),
    .B(_1657_),
    .Y(_1658_)
);

NAND2X1 _3629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1657_),
    .B(_1656_),
    .Y(_1659_)
);

OAI21X1 _3630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1653_),
    .B(_1636_),
    .C(_1648_),
    .Y(_1660_)
);

NAND2X1 _3631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1639_),
    .B(_1660_),
    .Y(_1661_)
);

NAND2X1 _3632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1602_),
    .B(_1604_),
    .Y(_1662_)
);

OAI21X1 _3633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1562_),
    .B(_1600_),
    .C(_1605_),
    .Y(_1663_)
);

NAND2X1 _3634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1662_),
    .B(_1663_),
    .Y(_1664_)
);

NOR2X1 _3635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1599_),
    .B(_1595_),
    .Y(_1665_)
);

OAI21X1 _3636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1665_),
    .B(_1600_),
    .C(_1623_),
    .Y(_1666_)
);

NAND2X1 _3637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.BCD ),
    .B(_1666_),
    .Y(_1667_)
);

OAI21X1 _3638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1545_),
    .B(_1549_),
    .C(_1625_),
    .Y(_1668_)
);

OAI21X1 _3639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1667_),
    .B(_1664_),
    .C(_1668_),
    .Y(_1669_)
);

INVX1 _3640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1629_),
    .Y(_1670_)
);

AOI22X1 _3641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1533_),
    .B(_1535_),
    .C(_1669_),
    .D(_1670_),
    .Y(_1671_)
);

OAI21X1 _3642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1634_),
    .B(_1671_),
    .C(_1631_),
    .Y(_1672_)
);

NAND2X1 _3643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1654_),
    .B(_1672_),
    .Y(_1673_)
);

NAND3X1 _3644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1638_),
    .B(_1648_),
    .C(_1673_),
    .Y(_1674_)
);

AND2X2 _3645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1661_),
    .B(_1674_),
    .Y(_1675_)
);

NAND2X1 _3646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1635_),
    .B(_1630_),
    .Y(_1676_)
);

NAND2X1 _3647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1634_),
    .B(_1671_),
    .Y(_1677_)
);

NAND2X1 _3648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1676_),
    .B(_1677_),
    .Y(_1678_)
);

NAND2X1 _3649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1653_),
    .B(_1636_),
    .Y(_1679_)
);

NAND2X1 _3650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1679_),
    .B(_1673_),
    .Y(_1680_)
);

AOI21X1 _3651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1680_),
    .B(_1678_),
    .C(_1608_),
    .Y(_1681_)
);

AOI22X1 _3652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1658_),
    .B(_1659_),
    .C(_1675_),
    .D(_1681_),
    .Y(_1682_)
);

OAI21X1 _3653_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf0),
    .B(_1682_),
    .C(_1732_),
    .Y(_1515_)
);

NAND2X1 _3654_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(HC),
    .B(_1714__bF$buf3),
    .Y(_1683_)
);

OAI21X1 _3655_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf2),
    .B(_1626_),
    .C(_1683_),
    .Y(_1516_)
);

NAND2X1 _3656_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[0]),
    .B(_1714__bF$buf1),
    .Y(_1684_)
);

AOI21X1 _3657_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1611_),
    .B(_1592_),
    .C(_1586_),
    .Y(_1685_)
);

OAI21X1 _3658_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1580_),
    .B(_1610_),
    .C(_1611_),
    .Y(_1686_)
);

OAI21X1 _3659_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1612_),
    .B(_1686_),
    .C(RDY_bF$buf3),
    .Y(_1687_)
);

OAI21X1 _3660_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1685_),
    .B(_1687_),
    .C(_1684_),
    .Y(_1517_)
);

NAND2X1 _3661_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[1]),
    .B(_1714__bF$buf0),
    .Y(_1688_)
);

OAI21X1 _3662_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf3),
    .B(_1623_),
    .C(_1688_),
    .Y(_1518_)
);

NAND2X1 _3663_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[2]),
    .B(_1714__bF$buf2),
    .Y(_1689_)
);

OAI21X1 _3664_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf1),
    .B(_1620_),
    .C(_1689_),
    .Y(_1519_)
);

NAND2X1 _3665_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[3]),
    .B(_1714__bF$buf0),
    .Y(_1690_)
);

OAI21X1 _3666_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf3),
    .B(_1664_),
    .C(_1690_),
    .Y(_1520_)
);

NAND2X1 _3667_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[4]),
    .B(_1714__bF$buf2),
    .Y(_1691_)
);

NOR2X1 _3668_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1670_),
    .B(_1669_),
    .Y(_1692_)
);

OAI21X1 _3669_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1629_),
    .B(_1626_),
    .C(RDY_bF$buf2),
    .Y(_1693_)
);

OAI21X1 _3670_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1693_),
    .B(_1692_),
    .C(_1691_),
    .Y(_1521_)
);

NAND2X1 _3671_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[5]),
    .B(_1714__bF$buf1),
    .Y(_1694_)
);

OAI21X1 _3672_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf0),
    .B(_1678_),
    .C(_1694_),
    .Y(_1522_)
);

NAND2X1 _3673_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ADD[6]),
    .B(_1714__bF$buf3),
    .Y(_1695_)
);

OAI21X1 _3674_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1714__bF$buf2),
    .B(_1680_),
    .C(_1695_),
    .Y(_1523_)
);

NAND2X1 _3675_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf1),
    .B(_1675_),
    .Y(_1696_)
);

OAI21X1 _3676_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1707_),
    .B(RDY_bF$buf0),
    .C(_1696_),
    .Y(_1524_)
);

NAND2X1 _3677_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[7]),
    .B(RDY_bF$buf9),
    .Y(_1697_)
);

OAI21X1 _3678_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(RDY_bF$buf8),
    .B(_1703_),
    .C(_1697_),
    .Y(_1525_)
);

DFFSR _3679_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_1514_),
    .Q(\u_ALU8.BI7 ),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3680_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf10),
    .D(_1515_),
    .Q(CO),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3681_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf9),
    .D(_1516_),
    .Q(HC),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3682_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf8),
    .D(_1517_),
    .Q(ADD[0]),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3683_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf7),
    .D(_1518_),
    .Q(ADD[1]),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3684_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf6),
    .D(_1519_),
    .Q(ADD[2]),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3685_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf5),
    .D(_1520_),
    .Q(ADD[3]),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3686_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_1521_),
    .Q(ADD[4]),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3687_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_1522_),
    .Q(ADD[5]),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3688_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_1523_),
    .Q(ADD[6]),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3689_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_1524_),
    .Q(AN),
    .R(_1513_),
    .S(vdd)
);

DFFSR _3690_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_1525_),
    .Q(\u_ALU8.AI7 ),
    .R(_1513_),
    .S(vdd)
);

BUFX2 _3691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[0]),
    .Y(AB[0])
);

BUFX2 _3692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[1]),
    .Y(AB[1])
);

BUFX2 _3693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[10]),
    .Y(AB[10])
);

BUFX2 _3694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[11]),
    .Y(AB[11])
);

BUFX2 _3695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[12]),
    .Y(AB[12])
);

BUFX2 _3696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[13]),
    .Y(AB[13])
);

BUFX2 _3697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[14]),
    .Y(AB[14])
);

BUFX2 _3698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[15]),
    .Y(AB[15])
);

BUFX2 _3699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[2]),
    .Y(AB[2])
);

BUFX2 _3700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[3]),
    .Y(AB[3])
);

BUFX2 _3701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[4]),
    .Y(AB[4])
);

BUFX2 _3702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[5]),
    .Y(AB[5])
);

BUFX2 _3703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[6]),
    .Y(AB[6])
);

BUFX2 _3704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[7]),
    .Y(AB[7])
);

BUFX2 _3705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[8]),
    .Y(AB[8])
);

BUFX2 _3706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1741_[9]),
    .Y(AB[9])
);

BUFX2 _3707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[0]),
    .Y(DO[0])
);

BUFX2 _3708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[1]),
    .Y(DO[1])
);

BUFX2 _3709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[2]),
    .Y(DO[2])
);

BUFX2 _3710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[3]),
    .Y(DO[3])
);

BUFX2 _3711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[4]),
    .Y(DO[4])
);

BUFX2 _3712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[5]),
    .Y(DO[5])
);

BUFX2 _3713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[6]),
    .Y(DO[6])
);

BUFX2 _3714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1742_[7]),
    .Y(DO[7])
);

BUFX2 _3715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_1743_),
    .Y(WE)
);

endmodule
