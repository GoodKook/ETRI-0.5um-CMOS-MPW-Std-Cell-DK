magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -122 -162 454 734
<< ntransistor >>
rect 71 480 81 604
rect 189 480 199 604
<< ptransistor >>
rect 43 0 53 124
rect 103 0 113 124
rect 163 0 173 124
rect 223 0 233 124
<< ndiffusion >>
rect 28 562 71 604
rect 28 550 40 562
rect 52 550 71 562
rect 28 506 71 550
rect 28 494 40 506
rect 52 494 71 506
rect 28 480 71 494
rect 81 562 124 604
rect 81 550 100 562
rect 112 550 124 562
rect 81 506 124 550
rect 81 494 100 506
rect 112 494 124 506
rect 81 480 124 494
rect 146 562 189 604
rect 146 550 158 562
rect 170 550 189 562
rect 146 506 189 550
rect 146 494 158 506
rect 170 494 189 506
rect 146 480 189 494
rect 199 562 242 604
rect 199 550 218 562
rect 230 550 242 562
rect 199 506 242 550
rect 199 494 218 506
rect 230 494 242 506
rect 199 480 242 494
<< ndcontact >>
rect 40 550 52 562
rect 40 494 52 506
rect 100 550 112 562
rect 100 494 112 506
rect 158 550 170 562
rect 158 494 170 506
rect 218 550 230 562
rect 218 494 230 506
<< psubstratepdiff >>
rect 0 110 43 124
rect 0 98 12 110
rect 24 98 43 110
rect 0 54 43 98
rect 0 42 12 54
rect 24 42 43 54
rect 0 0 43 42
rect 53 110 103 124
rect 53 98 72 110
rect 84 98 103 110
rect 53 54 103 98
rect 53 42 72 54
rect 84 42 103 54
rect 53 0 103 42
rect 113 110 163 124
rect 113 98 132 110
rect 144 98 163 110
rect 113 54 163 98
rect 113 42 132 54
rect 144 42 163 54
rect 113 0 163 42
rect 173 110 223 124
rect 173 98 192 110
rect 204 98 223 110
rect 173 54 223 98
rect 173 42 192 54
rect 204 42 223 54
rect 173 0 223 42
rect 233 110 276 124
rect 233 98 252 110
rect 264 98 276 110
rect 233 54 276 98
rect 233 42 252 54
rect 264 42 276 54
rect 233 0 276 42
<< psubstratepcontact >>
rect 12 98 24 110
rect 12 42 24 54
rect 72 98 84 110
rect 72 42 84 54
rect 132 98 144 110
rect 132 42 144 54
rect 192 98 204 110
rect 192 42 204 54
rect 252 98 264 110
rect 252 42 264 54
<< polysilicon >>
rect 71 604 81 614
rect 189 604 199 614
rect 71 456 81 480
rect 189 456 199 480
rect 43 124 53 148
rect 103 124 113 148
rect 163 124 173 148
rect 223 124 233 148
rect 43 -10 53 0
rect 103 -10 113 0
rect 163 -10 173 0
rect 223 -10 233 0
<< metal1 >>
rect 26 562 68 606
rect 26 550 40 562
rect 52 550 68 562
rect 26 506 68 550
rect 26 494 40 506
rect 52 494 68 506
rect 26 478 68 494
rect 84 562 186 606
rect 84 550 100 562
rect 112 550 158 562
rect 170 550 186 562
rect 84 506 186 550
rect 84 494 100 506
rect 112 494 158 506
rect 170 494 186 506
rect 84 478 186 494
rect 202 562 244 606
rect 202 550 218 562
rect 230 550 244 562
rect 202 506 244 550
rect 202 494 218 506
rect 230 494 244 506
rect 202 478 244 494
rect -2 418 96 462
rect 116 418 212 462
rect 2 146 126 186
rect 150 146 274 186
rect -2 110 40 126
rect -2 98 12 110
rect 24 98 40 110
rect -2 54 40 98
rect -2 42 12 54
rect 24 42 40 54
rect -2 -18 40 42
rect 56 110 100 126
rect 56 98 72 110
rect 84 98 100 110
rect 56 54 100 98
rect 56 42 72 54
rect 84 42 100 54
rect 56 -2 100 42
rect 116 110 160 126
rect 116 98 132 110
rect 144 98 160 110
rect 116 54 160 98
rect 116 42 132 54
rect 144 42 160 54
rect 116 -18 160 42
rect 176 110 220 126
rect 176 98 192 110
rect 204 98 220 110
rect 176 54 220 98
rect 176 42 192 54
rect 204 42 220 54
rect 176 -2 220 42
rect 236 110 278 126
rect 236 98 252 110
rect 264 98 278 110
rect 236 54 278 98
rect 236 42 252 54
rect 264 42 278 54
rect 236 -18 278 42
rect -2 -42 278 -18
<< metal2 >>
rect 26 478 66 606
rect 204 540 244 606
rect 204 478 334 540
rect -2 418 96 458
rect 116 418 212 458
rect 56 186 96 418
rect 172 186 212 418
rect 2 146 126 186
rect 150 146 274 186
rect 294 126 334 478
rect 58 -2 98 126
rect 178 -2 218 126
rect 238 44 334 126
rect 238 -2 278 44
<< metal3 >>
rect 26 478 66 606
rect 58 -2 98 126
rect 178 -2 218 126
use CONT  CONT_0
timestamp 1537935238
transform 1 0 106 0 1 528
box -6 -6 6 6
use CONT  CONT_1
timestamp 1537935238
transform 1 0 164 0 1 584
box -6 -6 6 6
use CONT  CONT_2
timestamp 1537935238
transform 1 0 164 0 1 528
box -6 -6 6 6
use CONT  CONT_3
timestamp 1537935238
transform 1 0 106 0 1 584
box -6 -6 6 6
use CONT  CONT_4
timestamp 1537935238
transform -1 0 138 0 -1 76
box -6 -6 6 6
use CONT  CONT_5
timestamp 1537935238
transform -1 0 138 0 -1 20
box -6 -6 6 6
use CONT  CONT_6
timestamp 1537935238
transform -1 0 18 0 -1 20
box -6 -6 6 6
use CONT  CONT_7
timestamp 1537935238
transform -1 0 18 0 -1 76
box -6 -6 6 6
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_0
timestamp 1537935238
transform -1 0 94 0 -1 458
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_1
timestamp 1537935238
transform -1 0 212 0 -1 458
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_2
timestamp 1537935238
transform 1 0 210 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_3
timestamp 1537935238
transform 1 0 150 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_4
timestamp 1537935238
transform 1 0 90 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_5
timestamp 1537935238
transform 1 0 30 0 1 146
box 0 0 36 36
use VIA1  VIA1_0
timestamp 1537935238
transform 1 0 199 0 1 166
box -8 -8 8 8
use VIA1  VIA1_1
timestamp 1537935238
transform 1 0 22 0 1 166
box -8 -8 8 8
use VIA1  VIA1_2
timestamp 1537935238
transform 1 0 46 0 1 528
box -8 -8 8 8
use VIA1  VIA1_3
timestamp 1537935238
transform 1 0 224 0 1 528
box -8 -8 8 8
use VIA1  VIA1_4
timestamp 1537935238
transform 1 0 46 0 1 584
box -8 -8 8 8
use VIA1  VIA1_5
timestamp 1537935238
transform 1 0 136 0 1 438
box -8 -8 8 8
use VIA1  VIA1_6
timestamp 1537935238
transform 1 0 224 0 1 584
box -8 -8 8 8
use VIA1  VIA1_7
timestamp 1537935238
transform 1 0 168 0 1 438
box -8 -8 8 8
use VIA1  VIA1_8
timestamp 1537935238
transform 1 0 18 0 1 438
box -8 -8 8 8
use VIA1  VIA1_9
timestamp 1537935238
transform 1 0 254 0 1 166
box -8 -8 8 8
use VIA1  VIA1_10
timestamp 1537935238
transform 1 0 78 0 1 166
box -8 -8 8 8
use VIA1  VIA1_11
timestamp 1537935238
transform 1 0 50 0 1 438
box -8 -8 8 8
use VIA1  VIA1_12
timestamp 1537935238
transform -1 0 258 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_13
timestamp 1537935238
transform -1 0 258 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_14
timestamp 1537935238
transform -1 0 198 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_15
timestamp 1537935238
transform -1 0 198 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_16
timestamp 1537935238
transform -1 0 78 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_17
timestamp 1537935238
transform -1 0 78 0 -1 20
box -8 -8 8 8
use VIA2  VIA2_0
timestamp 1537935238
transform 1 0 46 0 1 500
box -8 -8 8 8
use VIA2  VIA2_1
timestamp 1537935238
transform 1 0 46 0 1 556
box -8 -8 8 8
use VIA2  VIA2_2
timestamp 1537935238
transform -1 0 198 0 -1 48
box -8 -8 8 8
use VIA2  VIA2_3
timestamp 1537935238
transform -1 0 198 0 -1 104
box -8 -8 8 8
use VIA2  VIA2_4
timestamp 1537935238
transform -1 0 78 0 -1 48
box -8 -8 8 8
use VIA2  VIA2_5
timestamp 1537935238
transform -1 0 78 0 -1 104
box -8 -8 8 8
<< end >>
