magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect -17 39 67 79
rect -7 30 57 39
<< nwell >>
rect -7 77 57 136
<< ntransistor >>
rect 11 7 13 27
rect 16 7 18 27
rect 26 7 28 27
rect 31 7 33 27
<< ptransistor >>
rect 9 83 11 123
rect 19 83 21 123
rect 29 83 31 123
rect 39 83 41 123
<< ndiffusion >>
rect 10 7 11 27
rect 13 7 16 27
rect 18 7 19 27
rect 25 7 26 27
rect 28 7 31 27
rect 33 7 34 27
<< pdiffusion >>
rect 8 84 9 123
rect 2 83 9 84
rect 11 90 12 123
rect 18 90 19 123
rect 11 83 19 90
rect 21 84 22 123
rect 28 84 29 123
rect 21 83 29 84
rect 31 117 39 123
rect 31 83 32 117
rect 38 83 39 117
rect 41 83 42 123
<< ndcontact >>
rect 4 7 10 27
rect 19 7 25 27
rect 34 7 40 27
<< pdcontact >>
rect 2 84 8 123
rect 12 90 18 123
rect 22 84 28 123
rect 32 83 38 117
rect 42 83 48 123
<< psubstratepcontact >>
rect -3 -3 53 3
<< nsubstratencontact >>
rect -3 127 53 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 29 123 31 125
rect 39 123 41 125
rect 9 72 11 83
rect 19 72 21 83
rect 3 69 11 72
rect 16 69 21 72
rect 29 72 31 83
rect 39 72 41 83
rect 29 69 34 72
rect 39 69 44 72
rect 3 51 6 69
rect 16 64 18 69
rect 3 31 6 45
rect 3 29 13 31
rect 11 27 13 29
rect 16 27 18 58
rect 31 64 34 69
rect 31 58 32 64
rect 31 38 34 58
rect 26 36 34 38
rect 42 51 44 69
rect 26 27 28 36
rect 42 31 44 45
rect 31 29 44 31
rect 31 27 33 29
rect 11 5 13 7
rect 16 5 18 7
rect 26 5 28 7
rect 31 5 33 7
<< polycontact >>
rect 12 58 18 64
rect 2 45 8 51
rect 32 58 38 64
rect 42 45 48 51
<< metal1 >>
rect -3 133 53 134
rect -3 126 53 127
rect 12 123 18 126
rect 8 84 22 87
rect 28 120 42 123
rect 32 80 38 83
rect 22 77 38 80
rect 22 58 25 77
rect 22 27 26 51
rect 4 4 10 7
rect 34 4 40 7
rect -3 3 53 4
rect -3 -4 53 -3
<< m2contact >>
rect 1 51 8 58
rect 11 51 18 58
rect 21 51 28 58
rect 31 51 38 58
rect 41 51 48 58
<< metal2 >>
rect 3 58 7 67
rect 23 58 27 67
rect 43 58 47 67
rect 13 43 17 51
rect 33 43 37 51
<< m1p >>
rect -3 126 53 134
rect -3 -4 53 4
<< m2p >>
rect 3 59 7 67
rect 23 59 27 67
rect 43 59 47 67
rect 13 43 17 50
rect 33 43 37 50
<< labels >>
rlabel metal2 5 65 5 65 5 A
port 1 n signal input
rlabel metal2 15 44 15 44 7 B
port 2 n signal input
rlabel metal2 45 65 45 65 1 C
port 3 n signal input
rlabel metal2 35 44 35 44 5 D
port 4 n signal input
rlabel metal2 25 65 25 65 5 Y
port 5 n signal output
rlabel metal1 -3 126 53 134 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -3 -4 53 4 0 gnd
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 50 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
