magic
tech scmos
magscale 1 2
timestamp 1702310384
<< nwell >>
rect -13 154 193 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 58 14 62 54
rect 78 14 82 54
rect 98 14 102 54
rect 118 14 122 54
rect 138 14 142 54
rect 158 14 162 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
rect 58 166 62 246
rect 78 166 82 246
rect 98 166 102 246
rect 118 166 122 246
rect 138 166 142 246
rect 158 166 162 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 36 14 38 54
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
rect 76 14 78 54
rect 82 14 84 54
rect 96 14 98 54
rect 102 14 104 54
rect 116 14 118 54
rect 122 14 124 54
rect 136 14 138 54
rect 142 14 144 54
rect 156 14 158 54
rect 162 14 164 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 24 246
rect 36 166 38 246
rect 42 166 44 246
rect 56 166 58 246
rect 62 166 64 246
rect 76 166 78 246
rect 82 166 84 246
rect 96 166 98 246
rect 102 166 104 246
rect 116 166 118 246
rect 122 166 124 246
rect 136 166 138 246
rect 142 166 144 246
rect 156 166 158 246
rect 162 166 164 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
rect 64 14 76 54
rect 84 14 96 54
rect 104 14 116 54
rect 124 14 136 54
rect 144 14 156 54
rect 164 14 176 54
<< pdcontact >>
rect 4 166 16 246
rect 24 166 36 246
rect 44 166 56 246
rect 64 166 76 246
rect 84 166 96 246
rect 104 166 116 246
rect 124 166 136 246
rect 144 166 156 246
rect 164 166 176 246
<< psubstratepcontact >>
rect -6 -6 186 6
<< nsubstratencontact >>
rect -6 254 186 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 78 246 82 250
rect 98 246 102 250
rect 118 246 122 250
rect 138 246 142 250
rect 158 246 162 250
rect 18 117 22 166
rect 38 117 42 166
rect 18 108 42 117
rect 18 54 22 108
rect 38 54 42 108
rect 58 120 62 166
rect 78 120 82 166
rect 70 108 82 120
rect 58 54 62 108
rect 78 54 82 108
rect 98 120 102 166
rect 118 120 122 166
rect 110 108 122 120
rect 98 54 102 108
rect 118 54 122 108
rect 138 120 142 166
rect 158 120 162 166
rect 150 108 162 120
rect 138 54 142 108
rect 158 54 162 108
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
rect 78 10 82 14
rect 98 10 102 14
rect 118 10 122 14
rect 138 10 142 14
rect 158 10 162 14
<< polycontact >>
rect 6 105 18 117
rect 58 108 70 120
rect 98 108 110 120
rect 138 108 150 120
<< metal1 >>
rect -6 266 186 268
rect -6 252 186 254
rect 4 246 16 252
rect 44 246 56 252
rect 84 246 96 252
rect 124 246 136 252
rect 164 246 176 252
rect 24 160 36 166
rect 64 160 76 166
rect 104 160 116 166
rect 144 160 156 166
rect 24 152 46 160
rect 64 152 90 160
rect 104 152 130 160
rect 144 152 174 160
rect 3 123 17 137
rect 6 117 17 123
rect 38 116 46 152
rect 38 108 58 116
rect 82 116 90 152
rect 82 108 98 116
rect 122 116 130 152
rect 165 137 174 152
rect 163 123 177 137
rect 122 108 138 116
rect 38 68 46 108
rect 82 68 90 108
rect 122 68 130 108
rect 165 68 174 123
rect 24 60 46 68
rect 64 60 90 68
rect 104 60 130 68
rect 144 60 174 68
rect 24 54 36 60
rect 64 54 76 60
rect 104 54 116 60
rect 144 54 156 60
rect 4 8 16 14
rect 44 8 56 14
rect 84 8 96 14
rect 124 8 136 14
rect 164 8 176 14
rect -6 6 186 8
rect -6 -8 186 -6
<< m1p >>
rect -6 252 186 268
rect 3 123 17 137
rect 163 123 177 137
rect -6 -8 186 8
<< labels >>
rlabel nsubstratencontact 90 260 90 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 90 0 90 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 170 131 170 131 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
