magic
tech scmos
magscale 1 2
timestamp 1701862152
<< checkpaint >>
rect 6 142 94 159
rect 226 142 314 159
rect -14 78 94 142
rect 166 78 314 142
rect -14 61 74 78
rect 166 61 294 78
<< nwell >>
rect -13 154 313 272
rect 62 150 249 154
rect 162 136 249 150
<< ntransistor >>
rect 22 14 26 54
rect 42 14 46 54
rect 62 14 66 54
rect 82 14 86 54
rect 92 14 96 54
rect 112 14 116 54
rect 132 14 136 54
rect 152 14 156 54
rect 172 14 176 54
rect 194 14 198 54
rect 204 14 208 54
rect 214 14 218 54
rect 234 14 238 34
rect 274 14 278 34
<< ptransistor >>
rect 22 166 26 246
rect 42 166 46 246
rect 62 166 66 246
rect 82 166 86 246
rect 92 166 96 246
rect 112 166 116 246
rect 132 174 136 246
rect 152 174 156 246
rect 172 174 176 246
rect 194 150 198 246
rect 204 150 208 246
rect 214 150 218 246
rect 234 206 238 246
rect 274 206 278 246
<< ndiffusion >>
rect 20 14 22 54
rect 26 42 42 54
rect 26 14 28 42
rect 40 14 42 42
rect 46 14 48 54
rect 60 14 62 54
rect 66 46 82 54
rect 66 14 68 46
rect 80 14 82 46
rect 86 14 92 54
rect 96 50 112 54
rect 96 18 98 50
rect 110 18 112 50
rect 96 14 112 18
rect 116 52 132 54
rect 116 14 118 52
rect 130 14 132 52
rect 136 40 152 54
rect 136 18 138 40
rect 150 18 152 40
rect 136 14 152 18
rect 156 52 172 54
rect 156 14 158 52
rect 170 14 172 52
rect 176 44 194 54
rect 176 14 179 44
rect 191 14 194 44
rect 198 14 204 54
rect 208 14 214 54
rect 218 52 232 54
rect 218 14 220 52
rect 232 14 234 34
rect 238 14 240 34
rect 272 14 274 34
rect 278 14 280 34
<< pdiffusion >>
rect 20 166 22 246
rect 26 178 28 246
rect 40 178 42 246
rect 26 166 42 178
rect 46 166 48 246
rect 60 166 62 246
rect 66 176 68 246
rect 80 176 82 246
rect 66 166 82 176
rect 86 166 92 246
rect 96 166 98 246
rect 110 166 112 246
rect 116 166 118 246
rect 130 174 132 246
rect 136 186 138 246
rect 150 186 152 246
rect 136 174 152 186
rect 156 176 158 246
rect 170 176 172 246
rect 156 174 172 176
rect 176 174 179 246
rect 178 164 179 174
rect 191 164 194 246
rect 178 150 194 164
rect 198 150 204 246
rect 208 150 214 246
rect 218 150 220 246
rect 232 206 234 246
rect 238 206 240 246
rect 272 206 274 246
rect 278 206 280 246
<< ndcontact >>
rect 8 14 20 54
rect 28 14 40 42
rect 48 14 60 54
rect 68 14 80 46
rect 98 18 110 50
rect 118 14 130 52
rect 138 18 150 40
rect 158 14 170 52
rect 179 14 191 44
rect 220 14 232 52
rect 240 14 252 34
rect 260 14 272 34
rect 280 14 292 34
<< pdcontact >>
rect 8 166 20 246
rect 28 178 40 246
rect 48 166 60 246
rect 68 176 80 246
rect 98 166 110 246
rect 118 166 130 246
rect 138 186 150 246
rect 158 176 170 246
rect 179 164 191 246
rect 220 150 232 246
rect 240 206 252 246
rect 260 206 272 246
rect 280 206 292 246
<< psubstratepcontact >>
rect -6 -6 306 6
<< nsubstratencontact >>
rect -6 254 306 266
<< polysilicon >>
rect 22 246 26 250
rect 42 246 46 250
rect 62 246 66 250
rect 82 246 86 250
rect 92 246 96 250
rect 112 246 116 250
rect 132 246 136 250
rect 152 246 156 250
rect 172 246 176 250
rect 194 246 198 250
rect 204 246 208 250
rect 214 246 218 250
rect 234 246 238 250
rect 274 246 278 250
rect 22 129 26 166
rect 22 54 26 117
rect 42 91 46 166
rect 62 117 66 166
rect 42 54 46 78
rect 62 54 66 105
rect 82 91 86 166
rect 92 164 96 166
rect 112 164 116 166
rect 132 164 136 174
rect 152 172 156 174
rect 172 172 176 174
rect 92 160 116 164
rect 122 160 136 164
rect 142 168 156 172
rect 163 168 176 172
rect 82 54 86 78
rect 98 76 102 160
rect 122 91 126 160
rect 142 122 146 168
rect 163 160 168 168
rect 98 60 110 64
rect 122 62 126 78
rect 142 62 146 110
rect 160 62 165 148
rect 194 135 198 150
rect 177 131 198 135
rect 177 123 186 131
rect 204 117 208 150
rect 177 72 181 110
rect 206 104 208 117
rect 177 68 198 72
rect 92 56 116 60
rect 122 58 136 62
rect 142 58 156 62
rect 160 58 176 62
rect 92 54 96 56
rect 112 54 116 56
rect 132 54 136 58
rect 152 54 156 58
rect 172 54 176 58
rect 194 54 198 68
rect 204 54 208 104
rect 214 77 218 150
rect 234 141 238 206
rect 214 64 216 77
rect 214 54 218 64
rect 237 56 242 129
rect 234 51 242 56
rect 234 34 238 51
rect 274 34 278 206
rect 22 10 26 14
rect 42 10 46 14
rect 62 10 66 14
rect 82 10 86 14
rect 92 10 96 14
rect 112 10 116 14
rect 132 10 136 14
rect 152 10 156 14
rect 172 10 176 14
rect 194 10 198 14
rect 204 10 208 14
rect 214 10 218 14
rect 234 10 238 14
rect 274 10 278 14
<< polycontact >>
rect 22 117 34 129
rect 60 105 72 117
rect 42 78 54 91
rect 78 78 90 91
rect 134 110 146 122
rect 118 78 130 91
rect 98 64 110 76
rect 160 148 172 160
rect 174 110 186 123
rect 194 104 206 117
rect 262 164 274 176
rect 232 129 244 141
rect 216 64 228 77
<< metal1 >>
rect -6 266 306 268
rect -6 252 306 254
rect 28 246 40 252
rect 98 246 110 252
rect 138 246 150 252
rect 220 246 232 252
rect 260 246 272 252
rect 20 166 48 172
rect 68 174 80 176
rect 68 165 72 174
rect 130 176 158 180
rect 130 174 166 176
rect 178 164 179 246
rect 178 160 191 164
rect 192 146 214 152
rect 238 206 240 215
rect 238 156 244 206
rect 238 150 257 156
rect 208 141 214 146
rect 208 135 232 141
rect 72 110 134 117
rect 146 110 174 118
rect 251 117 257 150
rect 26 72 36 103
rect 194 91 206 104
rect 54 78 78 85
rect 90 84 118 91
rect 130 84 206 91
rect 26 66 98 72
rect 110 66 216 72
rect 20 48 48 54
rect 28 8 40 14
rect 98 8 110 18
rect 130 46 158 52
rect 138 8 150 18
rect 178 14 179 44
rect 251 48 257 103
rect 242 40 257 48
rect 242 34 248 40
rect 280 34 288 206
rect 220 8 228 14
rect 260 8 272 14
rect -6 6 306 8
rect -6 -8 306 -6
<< m2contact >>
rect 72 160 86 174
rect 146 148 160 162
rect 178 146 192 160
rect 250 176 264 177
rect 250 164 262 176
rect 262 164 264 176
rect 250 163 264 164
rect 22 103 36 117
rect 46 103 60 117
rect 206 103 220 117
rect 243 103 257 117
rect 266 103 280 117
rect 68 46 82 60
rect 178 44 192 58
<< metal2 >>
rect 86 166 250 172
rect 146 162 160 166
rect 46 117 54 134
rect 26 86 34 103
rect 75 60 81 160
rect 182 58 188 146
rect 266 117 274 134
rect 206 86 214 103
rect 246 86 254 103
<< m1p >>
rect -6 252 306 268
rect -6 -8 306 8
<< m2p >>
rect 46 119 54 134
rect 266 119 274 134
rect 26 86 34 101
rect 206 86 214 101
rect 246 86 254 101
<< labels >>
rlabel metal2 30 90 30 90 3 A
port 1 n signal input
rlabel metal2 210 89 210 89 3 B
port 2 n signal input
rlabel metal2 50 131 50 131 1 C
port 3 n signal input
rlabel metal2 250 88 250 88 7 YS
port 4 n signal output
rlabel metal2 270 127 270 127 5 YC
port 5 n signal output
rlabel metal1 -6 252 306 268 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -6 -8 306 8 0 gnd
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 300 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
