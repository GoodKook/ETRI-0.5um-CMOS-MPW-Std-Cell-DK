magic
tech scmos
magscale 1 2
timestamp 1702306942
<< nwell >>
rect -13 154 113 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 58 14 62 54
rect 78 14 82 54
<< ptransistor >>
rect 18 166 22 246
rect 28 166 32 246
rect 58 166 62 246
rect 68 166 72 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 45 38 54
rect 22 14 24 45
rect 36 14 38 45
rect 42 14 44 54
rect 56 14 58 54
rect 62 26 64 54
rect 76 26 78 54
rect 62 14 78 26
rect 82 14 84 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 28 246
rect 32 166 34 246
rect 56 166 58 246
rect 62 166 68 246
rect 72 166 74 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 45
rect 44 14 56 54
rect 64 26 76 54
rect 84 14 96 54
<< pdcontact >>
rect 4 166 16 246
rect 34 166 56 246
rect 74 166 86 246
<< psubstratepcontact >>
rect -7 -6 107 6
<< nsubstratencontact >>
rect -7 254 107 266
<< polysilicon >>
rect 18 246 22 250
rect 28 246 32 250
rect 58 246 62 250
rect 68 246 72 250
rect 18 164 22 166
rect 14 160 22 164
rect 28 164 32 166
rect 28 160 42 164
rect 14 117 18 160
rect 17 105 18 117
rect 14 69 18 105
rect 14 62 22 69
rect 18 54 22 62
rect 38 54 42 160
rect 58 97 62 166
rect 68 164 72 166
rect 68 160 84 164
rect 80 117 84 160
rect 80 105 83 117
rect 58 85 60 97
rect 58 54 62 85
rect 80 70 84 105
rect 78 64 84 70
rect 78 54 82 64
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
rect 78 10 82 14
<< polycontact >>
rect 5 105 17 117
rect 26 85 38 97
rect 83 105 95 117
rect 60 85 72 97
<< metal1 >>
rect -7 266 107 268
rect -7 252 107 254
rect 4 246 16 252
rect 74 246 86 252
rect 46 137 54 166
rect 3 123 17 137
rect 43 123 57 137
rect 83 123 97 137
rect 5 117 17 123
rect 23 103 37 117
rect 26 97 37 103
rect 46 78 54 123
rect 83 117 95 123
rect 63 103 77 117
rect 63 97 72 103
rect 46 71 72 78
rect 4 54 56 57
rect 66 54 72 71
rect 16 51 44 54
rect 56 14 84 20
rect 24 8 36 14
rect -7 6 107 8
rect -7 -8 107 -6
<< m1p >>
rect -7 252 107 268
rect 3 123 17 137
rect 43 123 57 137
rect 83 123 97 137
rect 23 103 37 117
rect 63 103 77 117
rect -7 -8 107 8
<< labels >>
rlabel nsubstratencontact 50 260 50 260 0 vdd
port 6 nsew power bidirectional abutment
rlabel psubstratepcontact 50 0 50 0 0 gnd
port 7 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 90 127 90 127 0 C
port 3 nsew signal input
rlabel metal1 50 130 50 130 0 Y
port 5 nsew signal output
rlabel metal1 30 106 30 106 0 B
port 2 nsew signal input
rlabel metal1 70 107 70 107 0 D
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
