magic
tech scmos
magscale 1 3
timestamp 1555589239
<< checkpaint >>
rect -60 -60 78 80
<< genericcontact >>
rect 6 7 12 13
<< metal1 >>
rect 0 0 18 20
<< pseudo_rpoly2 >>
rect 1 1 17 19
<< end >>
