magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect -7 39 37 79
rect 53 39 97 79
<< nwell >>
rect -6 77 96 136
<< ntransistor >>
rect 9 7 11 27
rect 19 7 21 27
rect 29 7 31 27
rect 39 7 41 27
rect 49 7 51 27
rect 59 7 61 27
rect 69 7 71 27
rect 79 7 81 27
<< ptransistor >>
rect 9 83 11 123
rect 19 83 21 123
rect 29 83 31 123
rect 39 83 41 123
rect 49 83 51 123
rect 59 83 61 123
rect 69 83 71 123
rect 79 83 81 123
<< ndiffusion >>
rect 8 7 9 27
rect 11 7 12 27
rect 18 7 19 27
rect 21 7 22 27
rect 28 7 29 27
rect 31 7 32 27
rect 38 7 39 27
rect 41 7 42 27
rect 48 7 49 27
rect 51 7 52 27
rect 58 7 59 27
rect 61 7 62 27
rect 68 7 69 27
rect 71 7 72 27
rect 78 7 79 27
rect 81 7 82 27
<< pdiffusion >>
rect 8 83 9 123
rect 11 83 12 123
rect 18 83 19 123
rect 21 83 22 123
rect 28 83 29 123
rect 31 83 32 123
rect 38 83 39 123
rect 41 83 42 123
rect 48 83 49 123
rect 51 83 52 123
rect 58 83 59 123
rect 61 83 62 123
rect 68 83 69 123
rect 71 83 72 123
rect 78 83 79 123
rect 81 83 82 123
<< ndcontact >>
rect 2 7 8 27
rect 12 7 18 27
rect 22 7 28 27
rect 32 7 38 27
rect 42 7 48 27
rect 52 7 58 27
rect 62 7 68 27
rect 72 7 78 27
rect 82 7 88 27
<< pdcontact >>
rect 2 83 8 123
rect 12 83 18 123
rect 22 83 28 123
rect 32 83 38 123
rect 42 83 48 123
rect 52 83 58 123
rect 62 83 68 123
rect 72 83 78 123
rect 82 83 88 123
<< psubstratepcontact >>
rect -3 -3 93 3
<< nsubstratencontact >>
rect -3 127 93 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 29 123 31 125
rect 39 123 41 125
rect 49 123 51 125
rect 59 123 61 125
rect 69 123 71 125
rect 79 123 81 125
rect 9 27 11 83
rect 19 51 21 83
rect 17 45 21 51
rect 19 27 21 45
rect 29 43 31 83
rect 39 43 41 83
rect 35 37 41 43
rect 29 27 31 37
rect 39 27 41 37
rect 49 43 51 83
rect 59 43 61 83
rect 55 37 61 43
rect 49 27 51 37
rect 59 27 61 37
rect 69 43 71 83
rect 79 43 81 83
rect 75 37 81 43
rect 69 27 71 37
rect 79 27 81 37
rect 9 5 11 7
rect 19 5 21 7
rect 29 5 31 7
rect 39 5 41 7
rect 49 5 51 7
rect 59 5 61 7
rect 69 5 71 7
rect 79 5 81 7
<< polycontact >>
rect 11 45 17 51
rect 29 37 35 43
rect 49 37 55 43
rect 69 37 75 43
<< metal1 >>
rect -3 133 93 134
rect -3 126 93 127
rect 2 123 8 126
rect 22 123 28 126
rect 42 123 48 126
rect 62 123 68 126
rect 82 123 88 126
rect 12 80 18 83
rect 32 80 38 83
rect 52 80 58 83
rect 72 80 78 83
rect 12 76 25 80
rect 32 76 45 80
rect 52 76 65 80
rect 72 76 81 80
rect 21 41 25 76
rect 21 37 29 41
rect 41 41 45 76
rect 41 37 49 41
rect 61 41 65 76
rect 61 37 69 41
rect 21 34 25 37
rect 41 34 45 37
rect 61 34 65 37
rect 78 34 81 76
rect 12 30 25 34
rect 32 30 45 34
rect 52 30 65 34
rect 72 30 81 34
rect 12 27 18 30
rect 32 27 38 30
rect 52 27 58 30
rect 72 27 78 30
rect 2 4 8 7
rect 22 4 28 7
rect 42 4 48 7
rect 62 4 68 7
rect 82 4 88 7
rect -3 3 93 4
rect -3 -4 93 -3
<< m2contact >>
rect 11 51 18 58
rect 71 51 78 58
<< metal2 >>
rect 13 58 17 67
rect 73 58 77 67
<< m1p >>
rect -3 126 93 134
rect -3 -4 93 4
<< m2p >>
rect 13 59 17 67
rect 73 59 77 67
<< labels >>
rlabel metal2 14 65 14 65 3 A
port 1 n signal input
rlabel metal2 75 65 75 65 7 Y
port 2 n signal output
rlabel metal1 -3 126 93 134 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -3 -4 93 4 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 90 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
