magic
tech scmos
magscale 1 6
timestamp 1725340883
<< checkpaint >>
rect -82 889 1054 1050
rect -124 641 1054 889
rect -124 -50 1030 641
rect -124 -86 341 -50
<< nwell >>
rect 70 760 910 910
rect 70 220 220 760
rect 760 220 910 760
rect 70 70 910 220
<< psubstratepdiff >>
rect 260 680 720 720
rect 260 300 300 680
rect 680 300 720 680
rect 260 260 720 300
<< nsubstratendiff >>
rect 90 850 890 890
rect 90 130 130 850
rect 390 390 590 590
rect 850 130 890 850
rect 90 90 890 130
<< genericcontact >>
rect 140 850 840 890
rect 90 140 130 840
rect 300 680 680 720
rect 260 300 300 680
rect 390 390 590 590
rect 680 300 720 680
rect 300 260 680 300
rect 850 140 890 840
rect 140 90 840 130
<< metal1 >>
rect 90 850 890 890
rect 90 130 130 850
rect 260 680 720 720
rect 260 300 300 680
rect 390 390 590 590
rect 680 300 720 680
rect 260 260 720 300
rect 850 130 890 850
rect 90 90 890 130
<< end >>
