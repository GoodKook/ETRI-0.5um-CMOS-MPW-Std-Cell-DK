magic
tech scmos
magscale 1 2
timestamp 1702316108
<< nwell >>
rect -14 154 113 272
<< ntransistor >>
rect 22 14 26 34
rect 64 14 68 54
rect 74 14 78 54
<< ptransistor >>
rect 22 206 26 246
rect 64 166 68 246
rect 74 166 78 246
<< ndiffusion >>
rect 20 14 22 34
rect 26 14 28 34
rect 62 14 64 54
rect 68 14 74 54
rect 78 14 80 54
<< pdiffusion >>
rect 20 206 22 246
rect 26 206 28 246
rect 62 166 64 246
rect 68 166 74 246
rect 78 166 80 246
<< ndcontact >>
rect 8 14 20 34
rect 28 14 40 34
rect 50 14 62 54
rect 80 14 92 54
<< pdcontact >>
rect 8 206 20 246
rect 28 206 40 246
rect 50 166 62 246
rect 80 166 92 246
<< psubstratepcontact >>
rect -7 -6 107 6
<< nsubstratencontact >>
rect -7 254 107 266
<< polysilicon >>
rect 22 246 26 250
rect 64 246 68 250
rect 74 246 78 250
rect 22 60 26 206
rect 64 72 68 166
rect 46 68 68 72
rect 74 117 78 166
rect 74 105 82 117
rect 22 56 68 60
rect 22 34 26 56
rect 64 54 68 56
rect 74 54 78 105
rect 22 10 26 14
rect 64 10 68 14
rect 74 10 78 14
<< polycontact >>
rect 10 105 22 117
rect 34 68 46 80
rect 82 105 94 117
<< metal1 >>
rect -7 266 107 268
rect -7 252 107 254
rect 8 246 20 252
rect 80 246 92 252
rect 3 123 17 137
rect 6 117 17 123
rect 6 105 10 117
rect 29 80 37 206
rect 46 166 50 179
rect 46 137 54 166
rect 43 123 57 137
rect 83 123 97 137
rect 46 96 54 123
rect 83 117 94 123
rect 46 87 59 96
rect 29 68 34 80
rect 29 34 40 68
rect 52 54 59 87
rect 8 8 20 14
rect 80 8 92 14
rect -7 6 107 8
rect -7 -8 107 -6
<< m1p >>
rect -7 252 107 268
rect 3 123 17 137
rect 43 123 57 137
rect 83 123 97 137
rect -7 -8 107 8
<< labels >>
rlabel nsubstratencontact 50 260 50 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 50 0 50 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 10 131 10 131 0 EN
port 2 nsew signal input
rlabel metal1 90 130 90 130 0 A
port 1 nsew signal input
rlabel metal1 51 131 51 131 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
