magic
tech scmos
magscale 1 2
timestamp 1717503367
<< metal1 >>
rect -63 2098 -3 2358
rect 2390 2342 2483 2358
rect 1153 2183 1167 2193
rect 1107 2180 1167 2183
rect 1107 2177 1163 2180
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 1817 2067 1823 2083
rect 1807 2057 1823 2067
rect 1807 2053 1820 2057
rect 2423 1838 2483 2342
rect 2390 1822 2483 1838
rect 1087 1757 1113 1763
rect 1207 1757 1233 1763
rect 1387 1743 1400 1747
rect 1387 1733 1403 1743
rect 1397 1683 1403 1733
rect 1367 1677 1403 1683
rect 1887 1677 1913 1683
rect 1867 1637 1913 1643
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 1447 1457 1473 1463
rect 200 1443 213 1447
rect 197 1433 213 1443
rect 860 1443 873 1447
rect 857 1433 873 1443
rect 1247 1443 1260 1447
rect 1247 1433 1263 1443
rect 197 1406 203 1433
rect 857 1407 863 1433
rect 1257 1407 1263 1433
rect 857 1397 873 1407
rect 860 1393 873 1397
rect 1247 1397 1263 1407
rect 1247 1393 1260 1397
rect 447 1377 473 1383
rect 1147 1377 1173 1383
rect 2423 1318 2483 1822
rect 2390 1302 2483 1318
rect 1027 1237 1073 1243
rect 467 1177 493 1183
rect 467 1157 553 1163
rect 893 1163 907 1173
rect 877 1160 907 1163
rect 873 1157 903 1160
rect 873 1147 887 1157
rect 1967 1157 2013 1163
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 1247 923 1260 927
rect 1247 913 1263 923
rect 1257 887 1263 913
rect 1247 877 1263 887
rect 1247 873 1260 877
rect 2423 798 2483 1302
rect 2390 782 2483 798
rect -63 522 30 538
rect -63 18 -3 522
rect 897 487 903 513
rect 897 306 903 413
rect 1687 337 1733 343
rect 2423 278 2483 782
rect 2390 262 2483 278
rect -63 2 30 18
rect 567 13 570 27
rect 1567 13 1570 27
rect 2207 13 2210 27
rect 2423 2 2483 262
<< m2contact >>
rect 1153 2193 1167 2207
rect 1093 2173 1107 2187
rect 2393 2093 2407 2107
rect 473 2073 487 2087
rect 1793 2053 1807 2067
rect 1073 1753 1087 1767
rect 1113 1752 1127 1766
rect 1193 1753 1207 1767
rect 1233 1753 1247 1767
rect 1373 1733 1387 1747
rect 1353 1673 1367 1687
rect 1873 1673 1887 1687
rect 1913 1673 1927 1687
rect 1853 1633 1867 1647
rect 1913 1633 1927 1647
rect 193 1553 207 1567
rect 853 1553 867 1567
rect 1253 1553 1267 1567
rect 1533 1553 1547 1567
rect 2073 1553 2087 1567
rect 1433 1453 1447 1467
rect 1473 1454 1487 1468
rect 213 1433 227 1447
rect 873 1433 887 1447
rect 1233 1433 1247 1447
rect 193 1392 207 1406
rect 873 1393 887 1407
rect 1233 1393 1247 1407
rect 433 1373 447 1387
rect 473 1373 487 1387
rect 1133 1373 1147 1387
rect 1173 1373 1187 1387
rect 1013 1233 1027 1247
rect 1073 1233 1087 1247
rect 453 1173 467 1187
rect 493 1173 507 1187
rect 893 1173 907 1187
rect 453 1152 467 1166
rect 553 1153 567 1167
rect 1953 1153 1967 1167
rect 2013 1153 2027 1167
rect 873 1133 887 1147
rect 673 1033 687 1047
rect 1013 1033 1027 1047
rect 1153 1033 1167 1047
rect 1373 1033 1387 1047
rect 1633 1033 1647 1047
rect 2393 1033 2407 1047
rect 1233 913 1247 927
rect 1233 873 1247 887
rect 893 513 907 527
rect 1693 513 1707 527
rect 2393 513 2407 527
rect 893 473 907 487
rect 893 413 907 427
rect 1673 333 1687 347
rect 1733 333 1747 347
rect 893 292 907 306
rect 553 13 567 27
rect 1553 13 1567 27
rect 2193 13 2207 27
<< metal2 >>
rect 736 2347 743 2403
rect 376 2248 383 2273
rect 76 2236 103 2243
rect 36 1988 43 2192
rect 96 2087 103 2236
rect 196 2187 203 2243
rect 436 2236 463 2243
rect 536 2236 563 2243
rect 96 1943 103 2073
rect 76 1936 103 1943
rect 196 1936 203 1993
rect 16 1607 23 1734
rect 36 1687 43 1913
rect 336 1907 343 2234
rect 356 1987 363 2173
rect 456 2167 463 2236
rect 376 1907 383 1943
rect 396 1827 403 2153
rect 556 2127 563 2236
rect 656 2147 663 2243
rect 836 2236 843 2273
rect 456 2087 463 2113
rect 467 2073 473 2087
rect 436 1728 443 1893
rect 456 1887 463 1993
rect 476 1946 483 2033
rect 536 1956 543 1993
rect 573 1960 587 1973
rect 576 1956 583 1960
rect 616 1956 623 2033
rect 636 2007 643 2053
rect 696 1967 703 2113
rect 707 1963 720 1967
rect 707 1956 723 1963
rect 756 1956 763 2013
rect 776 1967 783 2053
rect 796 2047 803 2233
rect 856 2127 863 2333
rect 896 2236 903 2293
rect 896 2027 903 2113
rect 936 2087 943 2353
rect 996 2347 1003 2403
rect 956 2227 963 2333
rect 1036 2143 1043 2293
rect 1076 2256 1083 2353
rect 1116 2307 1123 2353
rect 1116 2256 1123 2293
rect 1196 2287 1203 2403
rect 1216 2256 1243 2263
rect 1136 2220 1143 2223
rect 1133 2207 1147 2220
rect 1236 2207 1243 2256
rect 1093 2187 1107 2191
rect 1136 2167 1143 2193
rect 1153 2187 1167 2193
rect 1036 2136 1063 2143
rect 707 1953 720 1956
rect 916 1956 923 1993
rect 1036 1956 1043 2073
rect 1056 1967 1063 2136
rect 1096 1987 1103 2053
rect 1096 1956 1103 1973
rect 1136 1967 1143 2132
rect 1236 1987 1243 2193
rect 1256 2167 1263 2293
rect 1276 2256 1283 2353
rect 1296 2287 1303 2403
rect 1476 2307 1483 2403
rect 1776 2367 1783 2403
rect 1473 2260 1487 2272
rect 1476 2256 1483 2260
rect 1696 2256 1703 2313
rect 1276 2087 1283 2193
rect 1336 2127 1343 2253
rect 1816 2247 1823 2353
rect 1836 2287 1843 2403
rect 1856 2246 1863 2313
rect 1876 2236 1883 2333
rect 1256 1956 1263 1993
rect 1296 1967 1303 2093
rect 1376 2067 1383 2223
rect 1413 2207 1427 2212
rect 1416 2147 1423 2193
rect 1333 1960 1347 1973
rect 1336 1956 1343 1960
rect 1396 1967 1403 1993
rect 1436 1956 1443 2093
rect 1456 1987 1463 2013
rect 1476 1968 1483 2153
rect 1496 2027 1503 2223
rect 1516 2007 1523 2173
rect 1536 2123 1543 2213
rect 1556 2147 1563 2223
rect 1536 2116 1563 2123
rect 1536 1968 1543 2013
rect 1556 1987 1563 2116
rect 1576 1956 1583 2033
rect 1616 1956 1623 2173
rect 1676 2127 1683 2223
rect 1716 2187 1723 2223
rect 1896 2207 1903 2273
rect 2156 2243 2163 2403
rect 2156 2236 2173 2243
rect 2236 2236 2263 2243
rect 1696 1987 1703 2033
rect 1716 1983 1723 2013
rect 1736 2007 1743 2153
rect 1756 2107 1763 2193
rect 1787 2053 1793 2067
rect 1716 1976 1743 1983
rect 1736 1956 1743 1976
rect 1776 1968 1783 2013
rect 476 1787 483 1932
rect 516 1887 523 1923
rect 496 1827 503 1853
rect 536 1847 543 1893
rect 176 1716 203 1723
rect 56 1667 63 1703
rect 96 1647 103 1673
rect 136 1647 143 1683
rect 16 1327 23 1593
rect 96 1447 103 1633
rect 196 1567 203 1716
rect 296 1587 303 1723
rect 236 1543 243 1573
rect 216 1536 243 1543
rect 113 1440 127 1453
rect 216 1447 223 1536
rect 176 1440 203 1443
rect 116 1436 123 1440
rect 176 1436 207 1440
rect 193 1427 207 1436
rect 256 1436 263 1473
rect 296 1436 303 1513
rect 376 1448 383 1533
rect 436 1467 443 1714
rect 496 1587 503 1813
rect 656 1747 663 1893
rect 676 1747 683 1913
rect 716 1736 723 1833
rect 756 1748 763 1893
rect 796 1787 803 1923
rect 936 1916 963 1923
rect 976 1920 983 1923
rect 956 1863 963 1916
rect 973 1907 987 1920
rect 956 1856 983 1863
rect 936 1803 943 1853
rect 936 1796 963 1803
rect 956 1736 963 1796
rect 976 1747 983 1856
rect 1056 1736 1063 1873
rect 1076 1767 1083 1913
rect 1116 1887 1123 1923
rect 1160 1903 1173 1907
rect 1156 1893 1173 1903
rect 1116 1787 1123 1873
rect 1136 1767 1143 1793
rect 1120 1766 1143 1767
rect 1127 1756 1143 1766
rect 1127 1753 1140 1756
rect 1156 1736 1163 1893
rect 1196 1887 1203 1923
rect 1236 1867 1243 1913
rect 1176 1787 1183 1853
rect 1276 1807 1283 1923
rect 1316 1903 1323 1912
rect 1316 1896 1343 1903
rect 1336 1807 1343 1896
rect 1356 1867 1363 1923
rect 1376 1847 1383 1893
rect 1396 1887 1403 1913
rect 1193 1740 1207 1753
rect 1216 1747 1223 1793
rect 1247 1753 1253 1767
rect 1196 1736 1203 1740
rect 1273 1740 1287 1753
rect 1316 1747 1323 1773
rect 1276 1736 1283 1740
rect 1376 1747 1383 1793
rect 536 1716 563 1723
rect 556 1607 563 1716
rect 576 1667 583 1693
rect 596 1587 603 1703
rect 420 1446 440 1447
rect 420 1443 433 1446
rect 416 1436 433 1443
rect 420 1433 433 1436
rect 496 1436 503 1493
rect 516 1467 523 1533
rect 536 1447 543 1473
rect 556 1436 563 1513
rect 636 1447 643 1593
rect 676 1563 683 1693
rect 696 1667 703 1703
rect 736 1700 743 1703
rect 733 1687 747 1700
rect 656 1556 683 1563
rect 656 1487 663 1556
rect 676 1436 683 1513
rect 696 1507 703 1573
rect 716 1436 723 1473
rect 756 1436 763 1473
rect 816 1436 823 1673
rect 836 1647 843 1703
rect 856 1567 863 1673
rect 876 1627 883 1703
rect 876 1447 883 1533
rect 916 1463 923 1653
rect 936 1547 943 1692
rect 916 1456 943 1463
rect 36 1367 43 1393
rect 76 1327 83 1403
rect 16 1207 23 1253
rect 16 1047 23 1153
rect 36 1107 43 1163
rect 96 1143 103 1393
rect 136 1367 143 1403
rect 196 1347 203 1392
rect 276 1347 283 1403
rect 336 1267 343 1393
rect 356 1367 363 1403
rect 476 1400 483 1403
rect 516 1400 523 1403
rect 473 1387 487 1400
rect 513 1387 527 1400
rect 356 1206 363 1273
rect 176 1147 183 1193
rect 76 1136 103 1143
rect 76 1107 83 1136
rect 36 948 43 1093
rect 96 987 103 1033
rect 16 547 23 893
rect 96 803 103 973
rect 196 927 203 1113
rect 187 903 200 907
rect 187 896 203 903
rect 187 893 200 896
rect 96 796 123 803
rect 16 403 23 493
rect 36 447 43 793
rect 96 696 103 753
rect 116 747 123 796
rect 336 787 343 1173
rect 396 1107 403 1293
rect 416 1267 423 1373
rect 436 1347 443 1373
rect 476 1283 483 1333
rect 536 1307 543 1393
rect 576 1383 583 1403
rect 576 1380 603 1383
rect 576 1376 607 1380
rect 593 1367 607 1376
rect 696 1336 743 1343
rect 696 1303 703 1336
rect 676 1296 703 1303
rect 436 1276 483 1283
rect 436 1223 443 1276
rect 456 1228 463 1253
rect 416 1220 443 1223
rect 413 1216 443 1220
rect 413 1208 427 1216
rect 426 1200 427 1208
rect 456 1187 463 1214
rect 416 1087 423 1133
rect 396 903 403 1033
rect 416 947 423 1073
rect 376 896 403 903
rect 356 827 363 893
rect 176 708 183 773
rect 216 696 223 733
rect 256 696 263 753
rect 316 707 323 733
rect 336 696 343 773
rect 376 707 383 896
rect 436 827 443 892
rect 396 767 403 813
rect 396 696 403 753
rect 456 696 463 1152
rect 476 1047 483 1276
rect 636 1216 643 1273
rect 676 1216 683 1296
rect 696 1247 703 1273
rect 716 1227 723 1313
rect 736 1267 743 1336
rect 776 1327 783 1403
rect 836 1363 843 1403
rect 856 1387 863 1434
rect 936 1436 943 1456
rect 956 1436 963 1573
rect 976 1487 983 1673
rect 996 1467 1003 1513
rect 1016 1436 1023 1613
rect 1036 1583 1043 1703
rect 1076 1627 1083 1693
rect 1096 1627 1103 1673
rect 1136 1643 1143 1703
rect 1336 1687 1343 1703
rect 1336 1673 1353 1687
rect 1336 1647 1343 1673
rect 1136 1636 1163 1643
rect 1076 1587 1083 1613
rect 1036 1576 1063 1583
rect 1056 1507 1063 1576
rect 1116 1468 1123 1493
rect 1036 1436 1063 1443
rect 876 1363 883 1393
rect 836 1356 883 1363
rect 836 1276 873 1283
rect 776 1216 783 1253
rect 796 1247 803 1273
rect 836 1243 843 1276
rect 816 1240 843 1243
rect 813 1236 843 1240
rect 813 1227 827 1236
rect 853 1220 867 1233
rect 896 1227 903 1373
rect 916 1347 923 1403
rect 936 1287 943 1373
rect 996 1367 1003 1403
rect 1036 1367 1043 1436
rect 1136 1387 1143 1593
rect 1156 1547 1163 1636
rect 1236 1447 1243 1533
rect 1256 1507 1263 1553
rect 1176 1400 1183 1403
rect 1173 1387 1187 1400
rect 936 1228 943 1252
rect 1016 1247 1023 1293
rect 1036 1287 1043 1353
rect 1056 1347 1063 1373
rect 1076 1247 1083 1313
rect 856 1216 863 1220
rect 1116 1216 1123 1253
rect 1156 1228 1163 1273
rect 1176 1267 1183 1313
rect 1236 1247 1243 1393
rect 1256 1367 1263 1453
rect 1276 1436 1283 1593
rect 1333 1440 1347 1453
rect 1336 1436 1343 1440
rect 1256 1216 1263 1332
rect 1336 1207 1343 1333
rect 1356 1247 1363 1652
rect 1376 1627 1383 1693
rect 1396 1667 1403 1813
rect 1436 1767 1443 1893
rect 1456 1867 1463 1923
rect 1496 1827 1503 1913
rect 1536 1736 1543 1893
rect 1556 1847 1563 1923
rect 1576 1747 1583 1893
rect 1636 1867 1643 1923
rect 1816 1923 1823 2193
rect 1836 2167 1843 2203
rect 1836 1988 1843 2153
rect 2256 2107 2263 2236
rect 1876 1956 1883 2013
rect 1976 1943 1983 2053
rect 2076 2003 2083 2093
rect 2056 1996 2083 2003
rect 2056 1947 2063 1996
rect 1956 1936 1983 1943
rect 1816 1916 1843 1923
rect 1636 1743 1643 1813
rect 1713 1763 1727 1773
rect 1696 1760 1727 1763
rect 1696 1756 1723 1760
rect 1636 1736 1663 1743
rect 1696 1736 1703 1756
rect 1756 1736 1763 1912
rect 1836 1827 1843 1916
rect 1976 1843 1983 1936
rect 1976 1836 2003 1843
rect 1796 1747 1803 1793
rect 1376 1527 1383 1613
rect 1476 1468 1483 1703
rect 1516 1587 1523 1692
rect 1556 1587 1563 1703
rect 1576 1667 1583 1693
rect 1553 1567 1567 1573
rect 1547 1560 1567 1567
rect 1547 1556 1563 1560
rect 1547 1553 1560 1556
rect 1596 1527 1603 1703
rect 1433 1447 1447 1453
rect 1516 1436 1523 1473
rect 1596 1463 1603 1513
rect 1576 1456 1603 1463
rect 1576 1436 1583 1456
rect 1613 1440 1627 1453
rect 1656 1443 1663 1736
rect 1996 1736 2003 1836
rect 2016 1767 2023 1833
rect 2076 1736 2083 1793
rect 2216 1787 2223 2013
rect 2276 1943 2283 2234
rect 2316 2203 2323 2223
rect 2316 2196 2343 2203
rect 2336 1943 2343 2196
rect 2256 1936 2283 1943
rect 2296 1936 2343 1943
rect 2236 1843 2243 1934
rect 2256 1867 2263 1936
rect 2236 1836 2263 1843
rect 2256 1736 2263 1836
rect 2296 1747 2303 1936
rect 2316 1736 2323 1773
rect 2356 1768 2363 2223
rect 2376 1763 2383 2213
rect 2396 2107 2403 2333
rect 2376 1756 2403 1763
rect 2396 1736 2403 1756
rect 1736 1467 1743 1673
rect 1776 1667 1783 1703
rect 1796 1643 1803 1693
rect 1776 1636 1803 1643
rect 1616 1436 1623 1440
rect 1656 1436 1683 1443
rect 1416 1400 1423 1403
rect 1376 1327 1383 1393
rect 1413 1387 1427 1400
rect 1436 1347 1443 1393
rect 1456 1367 1463 1403
rect 1496 1307 1503 1403
rect 1596 1400 1603 1403
rect 1536 1347 1543 1393
rect 1593 1387 1607 1400
rect 1376 1247 1383 1292
rect 1616 1267 1623 1353
rect 1676 1307 1683 1436
rect 1756 1436 1763 1473
rect 1776 1447 1783 1636
rect 1816 1623 1823 1703
rect 1856 1647 1863 1703
rect 1886 1693 1887 1700
rect 1916 1700 1923 1703
rect 1873 1687 1887 1693
rect 1896 1627 1903 1693
rect 1913 1687 1927 1700
rect 1796 1616 1823 1623
rect 1796 1587 1803 1616
rect 1916 1607 1923 1633
rect 2016 1607 2023 1703
rect 1796 1467 1803 1533
rect 1816 1527 1823 1593
rect 2076 1567 2083 1593
rect 2096 1567 2103 1703
rect 2116 1587 2123 1673
rect 2136 1627 2143 1703
rect 2176 1667 2183 1693
rect 1816 1436 1823 1513
rect 1836 1467 1843 1553
rect 2016 1527 2023 1553
rect 2176 1547 2183 1653
rect 2236 1647 2243 1703
rect 1856 1436 1863 1473
rect 1976 1448 1983 1513
rect 2016 1436 2023 1473
rect 2056 1447 2063 1533
rect 2116 1436 2163 1443
rect 2196 1436 2203 1493
rect 2236 1447 2243 1573
rect 2276 1507 2283 1693
rect 2296 1643 2303 1693
rect 2296 1636 2323 1643
rect 2276 1436 2283 1493
rect 2316 1447 2323 1636
rect 2336 1627 2343 1703
rect 2356 1647 2363 1673
rect 2376 1667 2383 1703
rect 2336 1527 2343 1613
rect 2396 1567 2403 1673
rect 2416 1627 2423 1693
rect 2356 1436 2363 1473
rect 2396 1467 2403 1553
rect 2396 1436 2403 1453
rect 1636 1223 1643 1293
rect 1696 1287 1703 1353
rect 1616 1216 1643 1223
rect 1356 1196 1383 1203
rect 493 1167 507 1173
rect 516 1103 523 1183
rect 556 1180 563 1183
rect 553 1167 567 1180
rect 596 1127 603 1173
rect 736 1176 763 1183
rect 496 1096 523 1103
rect 496 987 503 1096
rect 616 1027 623 1153
rect 676 1047 683 1073
rect 716 983 723 1173
rect 736 1127 743 1176
rect 796 1147 803 1183
rect 756 1067 763 1093
rect 796 1047 803 1133
rect 696 976 723 983
rect 533 928 547 933
rect 656 916 663 973
rect 696 927 703 976
rect 716 916 723 953
rect 753 920 767 933
rect 796 927 803 973
rect 756 916 763 920
rect 816 916 823 1173
rect 836 1123 843 1183
rect 876 1163 883 1183
rect 907 1183 920 1187
rect 907 1176 923 1183
rect 907 1173 920 1176
rect 876 1156 903 1163
rect 856 1123 863 1153
rect 836 1120 863 1123
rect 836 1116 867 1120
rect 853 1107 867 1116
rect 856 947 863 1033
rect 876 1027 883 1133
rect 896 1127 903 1156
rect 1016 1163 1023 1183
rect 1016 1156 1043 1163
rect 896 1067 903 1113
rect 876 923 883 953
rect 856 916 883 923
rect 916 916 923 1153
rect 936 967 943 1033
rect 956 916 963 973
rect 976 947 983 1153
rect 1016 1047 1023 1133
rect 1036 1107 1043 1156
rect 1056 1147 1063 1172
rect 1036 928 1043 1093
rect 1076 927 1083 1033
rect 1096 987 1103 1173
rect 1136 1047 1143 1183
rect 1176 1047 1183 1183
rect 1196 1067 1203 1113
rect 1136 1036 1153 1047
rect 1140 1033 1153 1036
rect 1216 1007 1223 1173
rect 1236 1147 1243 1183
rect 1176 928 1183 953
rect 1216 916 1223 993
rect 1236 927 1243 973
rect 476 727 483 853
rect 516 787 523 883
rect 576 767 583 873
rect 596 847 603 883
rect 636 867 643 883
rect 627 856 643 867
rect 627 853 640 856
rect 656 827 663 853
rect 576 696 583 753
rect 656 727 663 773
rect 676 708 683 873
rect 776 880 783 883
rect 773 867 787 880
rect 696 747 703 813
rect 756 727 763 793
rect 816 783 823 813
rect 896 807 903 883
rect 936 827 943 883
rect 976 847 983 883
rect 1116 880 1123 883
rect 1053 867 1067 872
rect 776 776 823 783
rect 776 747 783 776
rect 136 627 143 663
rect 87 436 103 443
rect 16 396 33 403
rect 76 396 83 433
rect 96 407 103 436
rect 116 403 123 473
rect 116 396 143 403
rect 176 396 183 573
rect 236 428 243 533
rect 276 507 283 652
rect 200 363 213 367
rect 76 188 83 333
rect 156 183 163 363
rect 196 356 213 363
rect 200 353 213 356
rect 256 287 263 373
rect 276 267 283 383
rect 296 367 303 633
rect 356 627 363 663
rect 436 627 443 663
rect 616 547 623 632
rect 636 587 643 663
rect 656 483 663 653
rect 696 587 703 663
rect 876 623 883 673
rect 876 616 903 623
rect 636 480 663 483
rect 633 476 663 480
rect 633 467 647 476
rect 646 460 647 467
rect 396 376 403 413
rect 156 180 183 183
rect 156 176 187 180
rect 173 167 187 176
rect 116 67 123 123
rect 176 27 183 132
rect 416 67 423 273
rect 456 156 463 273
rect 536 267 543 413
rect 476 27 483 233
rect 513 160 527 173
rect 516 156 523 160
rect 556 127 563 373
rect 576 367 583 383
rect 576 287 583 353
rect 576 87 583 273
rect 596 247 603 453
rect 636 188 643 383
rect 656 366 663 453
rect 696 447 703 573
rect 896 527 903 616
rect 1036 547 1043 753
rect 1056 686 1063 793
rect 1076 676 1083 813
rect 1096 707 1103 873
rect 1113 867 1127 880
rect 1156 827 1163 873
rect 1196 847 1203 883
rect 1233 867 1247 873
rect 1147 756 1183 763
rect 1136 688 1143 713
rect 713 423 727 433
rect 696 420 727 423
rect 696 416 723 420
rect 696 396 703 416
rect 776 407 783 433
rect 816 396 823 473
rect 856 396 863 453
rect 896 427 903 473
rect 896 396 923 403
rect 976 396 983 533
rect 996 407 1003 513
rect 1056 427 1063 473
rect 716 267 723 363
rect 676 236 693 243
rect 547 13 553 27
rect 596 -17 603 143
rect 676 -17 683 236
rect 696 203 703 233
rect 696 196 723 203
rect 716 176 723 196
rect 736 188 743 233
rect 776 227 783 353
rect 856 247 863 333
rect 876 267 883 353
rect 896 327 903 396
rect 1076 396 1083 433
rect 1096 407 1103 672
rect 1156 423 1163 733
rect 1176 703 1183 756
rect 1176 696 1203 703
rect 1236 696 1243 793
rect 1256 723 1263 1153
rect 1276 1087 1283 1183
rect 1296 947 1303 1153
rect 1316 1107 1323 1163
rect 1336 1007 1343 1113
rect 1376 1087 1383 1196
rect 1616 1087 1623 1216
rect 1656 1196 1683 1203
rect 1716 1196 1723 1373
rect 1736 1323 1743 1403
rect 1736 1316 1763 1323
rect 1756 1247 1763 1316
rect 1776 1267 1783 1393
rect 1796 1327 1803 1403
rect 1836 1347 1843 1403
rect 1876 1347 1883 1373
rect 1896 1327 1903 1393
rect 1793 1220 1807 1233
rect 1836 1227 1843 1273
rect 1796 1216 1803 1220
rect 1676 1187 1683 1196
rect 1856 1186 1863 1253
rect 1916 1227 1923 1403
rect 1956 1216 1963 1293
rect 2016 1287 2023 1373
rect 2096 1347 2103 1392
rect 2036 1267 2043 1333
rect 2176 1327 2183 1403
rect 2196 1228 2203 1373
rect 2216 1307 2223 1403
rect 2216 1247 2223 1293
rect 1676 1163 1683 1173
rect 1676 1156 1703 1163
rect 1376 1047 1383 1073
rect 1436 967 1443 1053
rect 1296 847 1303 883
rect 1356 747 1363 953
rect 1396 916 1403 953
rect 1436 916 1443 953
rect 1476 886 1483 1073
rect 1647 1043 1660 1047
rect 1647 1033 1663 1043
rect 1496 916 1503 1033
rect 1556 927 1563 1033
rect 1616 987 1623 1013
rect 1576 916 1583 953
rect 1656 916 1663 1033
rect 1696 1007 1703 1156
rect 1776 1127 1783 1183
rect 1836 1176 1853 1183
rect 1716 1027 1723 1093
rect 1696 928 1703 953
rect 1776 928 1783 1073
rect 1816 916 1823 1113
rect 1836 967 1843 1176
rect 1856 916 1863 1033
rect 1876 987 1883 1183
rect 1916 943 1923 1173
rect 1936 1167 1943 1183
rect 2016 1180 2023 1183
rect 2013 1167 2027 1180
rect 1936 1156 1953 1167
rect 1940 1153 1953 1156
rect 2116 1147 2123 1183
rect 1956 948 1963 1013
rect 1976 967 1983 1113
rect 1996 963 2003 1133
rect 2116 1087 2123 1133
rect 2156 1047 2163 1172
rect 2256 987 2263 1393
rect 2276 1216 2283 1253
rect 2316 1243 2323 1333
rect 2336 1287 2343 1403
rect 2376 1243 2383 1392
rect 2316 1236 2343 1243
rect 1996 956 2023 963
rect 1896 936 1923 943
rect 1896 916 1903 936
rect 1256 720 1283 723
rect 1256 716 1287 720
rect 1273 707 1287 716
rect 1333 700 1347 713
rect 1336 696 1343 700
rect 1376 696 1383 873
rect 1416 727 1423 883
rect 1536 767 1543 872
rect 1616 727 1623 853
rect 1636 696 1643 753
rect 1676 696 1683 733
rect 1796 687 1803 851
rect 1976 787 1983 893
rect 1996 847 2003 903
rect 2016 787 2023 956
rect 2256 907 2263 973
rect 1136 416 1163 423
rect 1136 396 1143 416
rect 1176 396 1183 613
rect 1216 527 1223 663
rect 1296 627 1303 653
rect 1316 587 1323 663
rect 1356 660 1363 663
rect 1353 647 1367 660
rect 1316 527 1323 573
rect 1196 408 1203 453
rect 1236 396 1243 453
rect 1256 407 1263 433
rect 1376 407 1383 453
rect 1396 396 1403 653
rect 1416 547 1423 663
rect 1456 627 1463 663
rect 1456 476 1523 483
rect 1456 447 1463 476
rect 1476 407 1483 453
rect 1516 396 1523 476
rect 1536 427 1543 613
rect 1556 587 1563 663
rect 1576 627 1583 653
rect 1596 587 1603 663
rect 1556 527 1563 573
rect 1556 407 1563 513
rect 1616 396 1623 633
rect 1636 423 1643 453
rect 1656 447 1663 653
rect 1696 607 1703 663
rect 1716 543 1723 633
rect 1736 627 1743 663
rect 1707 536 1723 543
rect 1693 527 1707 533
rect 1736 487 1743 592
rect 1776 567 1783 643
rect 1836 567 1843 773
rect 2076 686 2083 773
rect 2116 676 2123 713
rect 2176 676 2183 753
rect 1636 416 1663 423
rect 1656 396 1663 416
rect 1736 408 1743 473
rect 1816 396 1823 433
rect 1916 428 1923 553
rect 1853 400 1867 413
rect 1856 396 1863 400
rect 900 306 920 307
rect 907 293 913 306
rect 956 287 963 363
rect 996 327 1003 353
rect 1016 287 1023 363
rect 856 203 863 233
rect 887 216 923 223
rect 836 196 863 203
rect 836 176 843 196
rect 696 140 703 143
rect 693 127 707 140
rect 756 87 763 143
rect 816 107 823 132
rect 856 -17 863 143
rect 916 87 923 216
rect 953 188 967 193
rect 1016 183 1023 273
rect 1056 267 1063 363
rect 1076 247 1083 313
rect 1016 176 1033 183
rect 1076 176 1083 233
rect 1096 207 1103 353
rect 1156 307 1163 363
rect 1196 247 1203 293
rect 1216 287 1223 363
rect 1316 360 1323 363
rect 1356 360 1363 363
rect 1236 267 1243 333
rect 1276 307 1283 353
rect 1313 347 1327 360
rect 1353 347 1367 360
rect 1156 176 1163 213
rect 1336 176 1343 253
rect 1376 247 1383 353
rect 1416 287 1423 363
rect 1436 176 1443 233
rect 1456 187 1463 363
rect 1476 327 1483 353
rect 1496 227 1503 353
rect 1536 327 1543 363
rect 1676 360 1683 363
rect 1496 176 1503 213
rect 1536 176 1543 313
rect 1556 187 1563 233
rect 1576 176 1583 293
rect 1596 207 1603 352
rect 1673 347 1687 360
rect 1756 347 1763 363
rect 1747 336 1763 347
rect 1747 333 1760 336
rect 1616 176 1623 213
rect 1656 187 1663 333
rect 1696 207 1703 233
rect 1716 176 1723 213
rect 1776 187 1783 293
rect 1796 247 1803 353
rect 1836 307 1843 363
rect 1956 347 1963 383
rect 1976 267 1983 413
rect 2067 383 2080 387
rect 2067 376 2083 383
rect 2067 373 2080 376
rect 2216 367 2223 713
rect 2256 696 2263 753
rect 2296 727 2303 892
rect 2316 767 2323 1033
rect 2336 947 2343 1236
rect 2356 1236 2383 1243
rect 2356 1216 2363 1236
rect 2376 903 2383 933
rect 2356 896 2383 903
rect 2356 696 2363 896
rect 2396 883 2403 1033
rect 2376 876 2403 883
rect 2376 847 2383 876
rect 2416 663 2423 693
rect 2396 656 2423 663
rect 2256 380 2263 383
rect 2253 367 2267 380
rect 2216 267 2223 353
rect 1196 107 1203 153
rect 1256 -17 1263 143
rect 1316 27 1323 143
rect 1476 140 1483 143
rect 1456 87 1463 133
rect 1473 127 1487 140
rect 1556 27 1563 113
rect 1696 27 1703 132
rect 1816 126 1823 253
rect 1756 47 1763 112
rect 1916 87 1923 163
rect 2056 67 2063 253
rect 2096 156 2103 253
rect 2316 247 2323 383
rect 2396 347 2403 513
rect 2156 156 2163 193
rect 2236 176 2243 213
rect 2316 176 2323 233
rect 2196 27 2203 153
rect 2276 -17 2283 143
rect 596 -24 623 -17
rect 676 -24 703 -17
rect 856 -24 883 -17
rect 1236 -24 1263 -17
rect 2256 -24 2283 -17
<< m3contact >>
rect 933 2353 947 2367
rect 733 2333 747 2347
rect 853 2333 867 2347
rect 373 2273 387 2287
rect 833 2273 847 2287
rect 33 2192 47 2206
rect 333 2234 347 2248
rect 373 2234 387 2248
rect 193 2173 207 2187
rect 93 2073 107 2087
rect 33 1974 47 1988
rect 193 1993 207 2007
rect 33 1913 47 1927
rect 13 1734 27 1748
rect 353 2173 367 2187
rect 493 2192 507 2206
rect 393 2153 407 2167
rect 453 2153 467 2167
rect 353 1973 367 1987
rect 333 1893 347 1907
rect 373 1893 387 1907
rect 793 2233 807 2247
rect 653 2133 667 2147
rect 453 2113 467 2127
rect 553 2113 567 2127
rect 693 2113 707 2127
rect 453 2073 467 2087
rect 633 2053 647 2067
rect 473 2033 487 2047
rect 613 2033 627 2047
rect 453 1993 467 2007
rect 433 1932 447 1946
rect 433 1893 447 1907
rect 393 1813 407 1827
rect 93 1734 107 1748
rect 533 1993 547 2007
rect 573 1973 587 1987
rect 633 1993 647 2007
rect 653 1954 667 1968
rect 773 2053 787 2067
rect 753 2013 767 2027
rect 693 1953 707 1967
rect 893 2293 907 2307
rect 853 2113 867 2127
rect 893 2113 907 2127
rect 793 2033 807 2047
rect 1073 2353 1087 2367
rect 1113 2353 1127 2367
rect 953 2333 967 2347
rect 993 2333 1007 2347
rect 1033 2293 1047 2307
rect 973 2254 987 2268
rect 953 2213 967 2227
rect 1013 2212 1027 2226
rect 1113 2293 1127 2307
rect 1273 2353 1287 2367
rect 1253 2293 1267 2307
rect 1193 2273 1207 2287
rect 1093 2212 1107 2226
rect 1173 2212 1187 2226
rect 1093 2191 1107 2205
rect 1133 2193 1147 2207
rect 1233 2193 1247 2207
rect 1153 2173 1167 2187
rect 1133 2153 1147 2167
rect 933 2073 947 2087
rect 1033 2073 1047 2087
rect 893 2013 907 2027
rect 913 1993 927 2007
rect 773 1953 787 1967
rect 813 1954 827 1968
rect 873 1954 887 1968
rect 993 1954 1007 1968
rect 1133 2132 1147 2146
rect 1093 2053 1107 2067
rect 1093 1973 1107 1987
rect 1053 1953 1067 1967
rect 1773 2353 1787 2367
rect 1813 2353 1827 2367
rect 1693 2313 1707 2327
rect 1473 2293 1487 2307
rect 1293 2273 1307 2287
rect 1473 2272 1487 2286
rect 1333 2253 1347 2267
rect 1393 2254 1407 2268
rect 1433 2254 1447 2268
rect 1513 2254 1527 2268
rect 1593 2254 1607 2268
rect 1653 2254 1667 2268
rect 1753 2254 1767 2268
rect 1313 2212 1327 2226
rect 1273 2193 1287 2207
rect 1253 2153 1267 2167
rect 1873 2333 1887 2347
rect 1853 2313 1867 2327
rect 1833 2273 1847 2287
rect 1813 2233 1827 2247
rect 1853 2232 1867 2246
rect 1893 2273 1907 2287
rect 1333 2113 1347 2127
rect 1293 2093 1307 2107
rect 1273 2073 1287 2087
rect 1253 1993 1267 2007
rect 1233 1973 1247 1987
rect 1133 1953 1147 1967
rect 1173 1954 1187 1968
rect 1213 1954 1227 1968
rect 1413 2212 1427 2226
rect 1413 2193 1427 2207
rect 1473 2153 1487 2167
rect 1413 2133 1427 2147
rect 1433 2093 1447 2107
rect 1373 2053 1387 2067
rect 1393 1993 1407 2007
rect 1333 1973 1347 1987
rect 1293 1953 1307 1967
rect 1372 1954 1386 1968
rect 1393 1953 1407 1967
rect 1453 2013 1467 2027
rect 1453 1973 1467 1987
rect 1533 2213 1547 2227
rect 1513 2173 1527 2187
rect 1493 2013 1507 2027
rect 1613 2212 1627 2226
rect 1613 2173 1627 2187
rect 1553 2133 1567 2147
rect 1533 2013 1547 2027
rect 1513 1993 1527 2007
rect 1573 2033 1587 2047
rect 1553 1973 1567 1987
rect 1473 1954 1487 1968
rect 1533 1954 1547 1968
rect 1793 2212 1807 2226
rect 1993 2232 2007 2246
rect 2393 2333 2407 2347
rect 2333 2254 2347 2268
rect 2173 2234 2187 2248
rect 1753 2193 1767 2207
rect 1813 2193 1827 2207
rect 1713 2173 1727 2187
rect 1733 2153 1747 2167
rect 1673 2113 1687 2127
rect 1693 2033 1707 2047
rect 1713 2013 1727 2027
rect 1693 1973 1707 1987
rect 1753 2093 1767 2107
rect 1773 2053 1787 2067
rect 1773 2013 1787 2027
rect 1733 1993 1747 2007
rect 1673 1954 1687 1968
rect 1773 1954 1787 1968
rect 473 1932 487 1946
rect 453 1873 467 1887
rect 553 1912 567 1926
rect 633 1912 647 1926
rect 673 1913 687 1927
rect 533 1893 547 1907
rect 653 1893 667 1907
rect 513 1873 527 1887
rect 493 1853 507 1867
rect 533 1833 547 1847
rect 493 1813 507 1827
rect 473 1773 487 1787
rect 33 1673 47 1687
rect 93 1673 107 1687
rect 53 1653 67 1667
rect 93 1633 107 1647
rect 133 1633 147 1647
rect 13 1593 27 1607
rect 53 1434 67 1448
rect 433 1714 447 1728
rect 473 1714 487 1728
rect 233 1573 247 1587
rect 293 1573 307 1587
rect 113 1453 127 1467
rect 93 1433 107 1447
rect 373 1533 387 1547
rect 293 1513 307 1527
rect 253 1473 267 1487
rect 613 1734 627 1748
rect 733 1912 747 1926
rect 753 1893 767 1907
rect 713 1833 727 1847
rect 652 1733 666 1747
rect 673 1733 687 1747
rect 893 1912 907 1926
rect 933 1853 947 1867
rect 1013 1912 1027 1926
rect 1073 1913 1087 1927
rect 973 1893 987 1907
rect 1053 1873 1067 1887
rect 793 1773 807 1787
rect 753 1734 767 1748
rect 813 1734 827 1748
rect 853 1734 867 1748
rect 973 1733 987 1747
rect 1013 1734 1027 1748
rect 1153 1912 1167 1926
rect 1173 1893 1187 1907
rect 1113 1873 1127 1887
rect 1133 1793 1147 1807
rect 1113 1773 1127 1787
rect 1113 1733 1127 1747
rect 1233 1913 1247 1927
rect 1193 1873 1207 1887
rect 1173 1853 1187 1867
rect 1233 1853 1247 1867
rect 1313 1912 1327 1926
rect 1393 1913 1407 1927
rect 1372 1893 1386 1907
rect 1353 1853 1367 1867
rect 1433 1893 1447 1907
rect 1393 1873 1407 1887
rect 1373 1833 1387 1847
rect 1393 1813 1407 1827
rect 1213 1793 1227 1807
rect 1273 1793 1287 1807
rect 1333 1793 1347 1807
rect 1373 1793 1387 1807
rect 1173 1773 1187 1787
rect 1313 1773 1327 1787
rect 1253 1753 1267 1767
rect 1273 1753 1287 1767
rect 1213 1733 1227 1747
rect 1313 1733 1327 1747
rect 1353 1734 1367 1748
rect 573 1693 587 1707
rect 573 1653 587 1667
rect 553 1593 567 1607
rect 633 1692 647 1706
rect 673 1693 687 1707
rect 633 1593 647 1607
rect 493 1573 507 1587
rect 593 1573 607 1587
rect 513 1533 527 1547
rect 493 1493 507 1507
rect 433 1453 447 1467
rect 373 1434 387 1448
rect 433 1432 447 1446
rect 553 1513 567 1527
rect 533 1473 547 1487
rect 513 1453 527 1467
rect 533 1433 547 1447
rect 612 1434 626 1448
rect 733 1673 747 1687
rect 813 1673 827 1687
rect 693 1653 707 1667
rect 693 1573 707 1587
rect 673 1513 687 1527
rect 653 1473 667 1487
rect 633 1433 647 1447
rect 693 1493 707 1507
rect 713 1473 727 1487
rect 753 1473 767 1487
rect 853 1673 867 1687
rect 833 1633 847 1647
rect 933 1692 947 1706
rect 993 1692 1007 1706
rect 913 1653 927 1667
rect 873 1613 887 1627
rect 873 1533 887 1547
rect 853 1434 867 1448
rect 973 1673 987 1687
rect 953 1573 967 1587
rect 933 1533 947 1547
rect 193 1413 207 1427
rect 33 1393 47 1407
rect 33 1353 47 1367
rect 93 1393 107 1407
rect 13 1313 27 1327
rect 73 1313 87 1327
rect 13 1253 27 1267
rect 13 1193 27 1207
rect 73 1194 87 1208
rect 13 1153 27 1167
rect 233 1392 247 1406
rect 133 1353 147 1367
rect 333 1393 347 1407
rect 193 1333 207 1347
rect 273 1333 287 1347
rect 393 1392 407 1406
rect 413 1373 427 1387
rect 533 1393 547 1407
rect 513 1373 527 1387
rect 353 1353 367 1367
rect 393 1293 407 1307
rect 353 1273 367 1287
rect 333 1253 347 1267
rect 172 1193 186 1207
rect 193 1192 207 1206
rect 352 1192 366 1206
rect 373 1194 387 1208
rect 333 1173 347 1187
rect 173 1133 187 1147
rect 193 1113 207 1127
rect 33 1093 47 1107
rect 73 1093 87 1107
rect 13 1033 27 1047
rect 93 1033 107 1047
rect 93 973 107 987
rect 33 934 47 948
rect 13 893 27 907
rect 73 892 87 906
rect 33 793 47 807
rect 193 913 207 927
rect 173 893 187 907
rect 13 533 27 547
rect 13 493 27 507
rect 93 753 107 767
rect 433 1333 447 1347
rect 473 1333 487 1347
rect 653 1392 667 1406
rect 693 1392 707 1406
rect 593 1353 607 1367
rect 533 1293 547 1307
rect 713 1313 727 1327
rect 413 1253 427 1267
rect 453 1253 467 1267
rect 453 1214 467 1228
rect 412 1194 426 1208
rect 433 1194 447 1208
rect 413 1133 427 1147
rect 393 1093 407 1107
rect 413 1073 427 1087
rect 393 1033 407 1047
rect 353 893 367 907
rect 413 933 427 947
rect 353 813 367 827
rect 173 773 187 787
rect 333 773 347 787
rect 113 733 127 747
rect 253 753 267 767
rect 213 733 227 747
rect 173 694 187 708
rect 313 733 327 747
rect 313 693 327 707
rect 433 892 447 906
rect 393 813 407 827
rect 433 813 447 827
rect 393 753 407 767
rect 373 693 387 707
rect 633 1273 647 1287
rect 533 1214 547 1228
rect 573 1214 587 1228
rect 693 1273 707 1287
rect 692 1233 706 1247
rect 893 1434 907 1448
rect 1013 1613 1027 1627
rect 993 1513 1007 1527
rect 973 1473 987 1487
rect 993 1453 1007 1467
rect 1072 1693 1086 1707
rect 1093 1673 1107 1687
rect 1173 1692 1187 1706
rect 1253 1692 1267 1706
rect 1293 1692 1307 1706
rect 1373 1693 1387 1707
rect 1353 1652 1367 1666
rect 1072 1613 1086 1627
rect 1093 1613 1107 1627
rect 1133 1593 1147 1607
rect 1073 1573 1087 1587
rect 1053 1493 1067 1507
rect 1113 1493 1127 1507
rect 1113 1454 1127 1468
rect 853 1373 867 1387
rect 893 1373 907 1387
rect 773 1313 787 1327
rect 793 1273 807 1287
rect 733 1253 747 1267
rect 773 1253 787 1267
rect 713 1213 727 1227
rect 793 1233 807 1247
rect 873 1273 887 1287
rect 813 1213 827 1227
rect 853 1233 867 1247
rect 933 1373 947 1387
rect 913 1333 927 1347
rect 1113 1433 1127 1447
rect 1073 1392 1087 1406
rect 1333 1633 1347 1647
rect 1273 1593 1287 1607
rect 1153 1533 1167 1547
rect 1233 1533 1247 1547
rect 1193 1434 1207 1448
rect 1253 1493 1267 1507
rect 1253 1453 1267 1467
rect 1213 1392 1227 1406
rect 1053 1373 1067 1387
rect 993 1353 1007 1367
rect 1033 1353 1047 1367
rect 1013 1293 1027 1307
rect 933 1273 947 1287
rect 933 1252 947 1266
rect 1053 1333 1067 1347
rect 1073 1313 1087 1327
rect 1173 1313 1187 1327
rect 1033 1273 1047 1287
rect 1153 1273 1167 1287
rect 1113 1253 1127 1267
rect 893 1213 907 1227
rect 933 1214 947 1228
rect 993 1214 1007 1228
rect 1033 1214 1047 1228
rect 1173 1253 1187 1267
rect 1333 1453 1347 1467
rect 1313 1392 1327 1406
rect 1253 1353 1267 1367
rect 1253 1332 1267 1346
rect 1333 1333 1347 1347
rect 1233 1233 1247 1247
rect 1153 1214 1167 1228
rect 1493 1913 1507 1927
rect 1453 1853 1467 1867
rect 1533 1893 1547 1907
rect 1493 1813 1507 1827
rect 1433 1753 1447 1767
rect 1453 1734 1467 1748
rect 1573 1893 1587 1907
rect 1553 1833 1567 1847
rect 1713 1912 1727 1926
rect 1753 1912 1767 1926
rect 1893 2193 1907 2207
rect 1833 2153 1847 2167
rect 2273 2234 2287 2248
rect 2073 2093 2087 2107
rect 2253 2093 2267 2107
rect 1973 2053 1987 2067
rect 1873 2013 1887 2027
rect 1833 1974 1847 1988
rect 1913 1974 1927 1988
rect 2213 2013 2227 2027
rect 1633 1853 1647 1867
rect 1633 1813 1647 1827
rect 1573 1733 1587 1747
rect 1713 1773 1727 1787
rect 2052 1933 2066 1947
rect 2073 1934 2087 1948
rect 1833 1813 1847 1827
rect 1793 1793 1807 1807
rect 1413 1692 1427 1706
rect 1393 1653 1407 1667
rect 1373 1613 1387 1627
rect 1373 1513 1387 1527
rect 1513 1692 1527 1706
rect 1573 1693 1587 1707
rect 1573 1653 1587 1667
rect 1513 1573 1527 1587
rect 1553 1573 1567 1587
rect 1593 1513 1607 1527
rect 1513 1473 1527 1487
rect 1393 1434 1407 1448
rect 1433 1433 1447 1447
rect 1473 1433 1487 1447
rect 1613 1453 1627 1467
rect 1793 1733 1807 1747
rect 1833 1734 1847 1748
rect 1933 1734 1947 1748
rect 2013 1833 2027 1847
rect 2073 1793 2087 1807
rect 2013 1753 2027 1767
rect 2033 1734 2047 1748
rect 2233 1934 2247 1948
rect 2253 1853 2267 1867
rect 2213 1773 2227 1787
rect 2113 1734 2127 1748
rect 2213 1734 2227 1748
rect 2313 1773 2327 1787
rect 2293 1733 2307 1747
rect 2373 2213 2387 2227
rect 2353 1754 2367 1768
rect 2353 1733 2367 1747
rect 1713 1692 1727 1706
rect 1733 1673 1747 1687
rect 1793 1693 1807 1707
rect 1773 1653 1787 1667
rect 1753 1473 1767 1487
rect 1733 1453 1747 1467
rect 1373 1393 1387 1407
rect 1433 1393 1447 1407
rect 1413 1373 1427 1387
rect 1453 1353 1467 1367
rect 1433 1333 1447 1347
rect 1373 1313 1387 1327
rect 1533 1393 1547 1407
rect 1633 1392 1647 1406
rect 1593 1373 1607 1387
rect 1613 1353 1627 1367
rect 1533 1333 1547 1347
rect 1373 1292 1387 1306
rect 1493 1293 1507 1307
rect 1693 1434 1707 1448
rect 1872 1693 1886 1707
rect 1893 1693 1907 1707
rect 1953 1692 1967 1706
rect 1973 1692 1987 1706
rect 1893 1613 1907 1627
rect 1813 1593 1827 1607
rect 1913 1593 1927 1607
rect 2013 1593 2027 1607
rect 2073 1593 2087 1607
rect 1793 1573 1807 1587
rect 1793 1533 1807 1547
rect 2113 1673 2127 1687
rect 2172 1693 2186 1707
rect 2193 1692 2207 1706
rect 2173 1653 2187 1667
rect 2133 1613 2147 1627
rect 2113 1573 2127 1587
rect 1833 1553 1847 1567
rect 2013 1553 2027 1567
rect 2093 1553 2107 1567
rect 1813 1513 1827 1527
rect 1793 1453 1807 1467
rect 1773 1433 1787 1447
rect 2272 1693 2286 1707
rect 2293 1693 2307 1707
rect 2233 1633 2247 1647
rect 2233 1573 2247 1587
rect 2053 1533 2067 1547
rect 2173 1533 2187 1547
rect 1973 1513 1987 1527
rect 2013 1513 2027 1527
rect 1853 1473 1867 1487
rect 1833 1453 1847 1467
rect 2013 1473 2027 1487
rect 1933 1434 1947 1448
rect 1973 1434 1987 1448
rect 2193 1493 2207 1507
rect 2053 1433 2067 1447
rect 2273 1493 2287 1507
rect 2233 1433 2247 1447
rect 2353 1673 2367 1687
rect 2413 1693 2427 1707
rect 2393 1673 2407 1687
rect 2373 1653 2387 1667
rect 2353 1633 2367 1647
rect 2333 1613 2347 1627
rect 2413 1613 2427 1627
rect 2393 1553 2407 1567
rect 2333 1513 2347 1527
rect 2353 1473 2367 1487
rect 2313 1433 2327 1447
rect 2393 1453 2407 1467
rect 1713 1373 1727 1387
rect 1693 1353 1707 1367
rect 1633 1293 1647 1307
rect 1673 1293 1687 1307
rect 1613 1253 1627 1267
rect 1352 1233 1366 1247
rect 1373 1233 1387 1247
rect 1693 1273 1707 1287
rect 1333 1193 1347 1207
rect 493 1153 507 1167
rect 593 1173 607 1187
rect 653 1172 667 1186
rect 692 1172 706 1186
rect 713 1173 727 1187
rect 613 1153 627 1167
rect 593 1113 607 1127
rect 473 1033 487 1047
rect 673 1073 687 1087
rect 613 1013 627 1027
rect 493 973 507 987
rect 653 973 667 987
rect 813 1173 827 1187
rect 793 1133 807 1147
rect 733 1113 747 1127
rect 753 1093 767 1107
rect 753 1053 767 1067
rect 793 1033 807 1047
rect 533 933 547 947
rect 493 914 507 928
rect 533 914 547 928
rect 613 914 627 928
rect 793 973 807 987
rect 713 953 727 967
rect 693 913 707 927
rect 753 933 767 947
rect 793 913 807 927
rect 853 1153 867 1167
rect 853 1093 867 1107
rect 853 1033 867 1047
rect 913 1153 927 1167
rect 973 1153 987 1167
rect 1053 1172 1067 1186
rect 1093 1173 1107 1187
rect 893 1113 907 1127
rect 893 1053 907 1067
rect 873 1013 887 1027
rect 873 953 887 967
rect 853 933 867 947
rect 933 1033 947 1047
rect 953 973 967 987
rect 933 953 947 967
rect 1013 1133 1027 1147
rect 1053 1133 1067 1147
rect 1033 1093 1047 1107
rect 973 933 987 947
rect 1073 1033 1087 1047
rect 1033 914 1047 928
rect 1213 1173 1227 1187
rect 1193 1113 1207 1127
rect 1193 1053 1207 1067
rect 1173 1033 1187 1047
rect 1253 1153 1267 1167
rect 1233 1133 1247 1147
rect 1213 993 1227 1007
rect 1093 973 1107 987
rect 1173 953 1187 967
rect 1073 913 1087 927
rect 1133 914 1147 928
rect 1173 914 1187 928
rect 1233 973 1247 987
rect 473 853 487 867
rect 573 873 587 887
rect 513 773 527 787
rect 673 873 687 887
rect 613 853 627 867
rect 653 853 667 867
rect 593 833 607 847
rect 653 813 667 827
rect 653 773 667 787
rect 573 753 587 767
rect 473 713 487 727
rect 493 694 507 708
rect 653 713 667 727
rect 733 872 747 886
rect 833 872 847 886
rect 773 853 787 867
rect 693 813 707 827
rect 813 813 827 827
rect 753 793 767 807
rect 693 733 707 747
rect 1053 872 1067 886
rect 1093 873 1107 887
rect 1053 853 1067 867
rect 973 833 987 847
rect 933 813 947 827
rect 1073 813 1087 827
rect 893 793 907 807
rect 1053 793 1067 807
rect 1033 753 1047 767
rect 773 733 787 747
rect 753 713 767 727
rect 613 694 627 708
rect 673 694 687 708
rect 773 674 787 688
rect 872 673 886 687
rect 53 652 67 666
rect 233 652 247 666
rect 273 652 287 666
rect 133 613 147 627
rect 173 573 187 587
rect 113 473 127 487
rect 33 433 47 447
rect 73 433 87 447
rect 33 394 47 408
rect 93 393 107 407
rect 233 533 247 547
rect 293 633 307 647
rect 273 493 287 507
rect 233 414 247 428
rect 253 373 267 387
rect 53 352 67 366
rect 73 333 87 347
rect 73 174 87 188
rect 213 353 227 367
rect 253 273 267 287
rect 413 652 427 666
rect 473 652 487 666
rect 553 652 567 666
rect 613 632 627 646
rect 353 613 367 627
rect 433 613 447 627
rect 653 653 667 667
rect 633 573 647 587
rect 613 533 627 547
rect 733 632 747 646
rect 893 672 907 686
rect 693 573 707 587
rect 593 453 607 467
rect 632 453 646 467
rect 653 453 667 467
rect 393 413 407 427
rect 533 413 547 427
rect 293 353 307 367
rect 413 273 427 287
rect 453 273 467 287
rect 273 253 287 267
rect 152 154 166 168
rect 173 153 187 167
rect 273 152 287 166
rect 33 132 47 146
rect 173 132 187 146
rect 113 53 127 67
rect 553 373 567 387
rect 533 253 547 267
rect 473 233 487 247
rect 413 53 427 67
rect 513 173 527 187
rect 573 353 587 367
rect 573 273 587 287
rect 553 113 567 127
rect 593 233 607 247
rect 1053 672 1067 686
rect 1153 873 1167 887
rect 1113 853 1127 867
rect 1233 853 1247 867
rect 1193 833 1207 847
rect 1153 813 1167 827
rect 1233 793 1247 807
rect 1133 753 1147 767
rect 1153 733 1167 747
rect 1133 713 1147 727
rect 1093 693 1107 707
rect 1093 672 1107 686
rect 1133 674 1147 688
rect 973 533 987 547
rect 1033 533 1047 547
rect 813 473 827 487
rect 692 433 706 447
rect 713 433 727 447
rect 773 433 787 447
rect 733 394 747 408
rect 773 393 787 407
rect 853 453 867 467
rect 993 513 1007 527
rect 1053 473 1067 487
rect 1073 433 1087 447
rect 1053 413 1067 427
rect 653 352 667 366
rect 752 352 766 366
rect 773 353 787 367
rect 713 253 727 267
rect 633 174 647 188
rect 573 73 587 87
rect 173 13 187 27
rect 473 13 487 27
rect 533 13 547 27
rect 693 233 707 247
rect 733 233 747 247
rect 833 352 847 366
rect 873 353 887 367
rect 853 333 867 347
rect 993 393 1007 407
rect 1033 394 1047 408
rect 1293 1153 1307 1167
rect 1273 1073 1287 1087
rect 1333 1113 1347 1127
rect 1313 1093 1327 1107
rect 1473 1192 1487 1206
rect 1773 1393 1787 1407
rect 1893 1393 1907 1407
rect 1873 1373 1887 1387
rect 1833 1333 1847 1347
rect 1873 1333 1887 1347
rect 1793 1313 1807 1327
rect 1893 1313 1907 1327
rect 1833 1273 1847 1287
rect 1773 1253 1787 1267
rect 1753 1233 1767 1247
rect 1793 1233 1807 1247
rect 1853 1253 1867 1267
rect 1833 1213 1847 1227
rect 1673 1173 1687 1187
rect 1892 1214 1906 1228
rect 1953 1392 1967 1406
rect 2033 1392 2047 1406
rect 2093 1392 2107 1406
rect 2013 1373 2027 1387
rect 1953 1293 1967 1307
rect 1913 1213 1927 1227
rect 2033 1333 2047 1347
rect 2093 1333 2107 1347
rect 2013 1273 2027 1287
rect 2193 1373 2207 1387
rect 2173 1313 2187 1327
rect 2033 1253 2047 1267
rect 2253 1393 2267 1407
rect 2213 1293 2227 1307
rect 2213 1233 2227 1247
rect 1993 1214 2007 1228
rect 2033 1214 2047 1228
rect 2133 1214 2147 1228
rect 2193 1214 2207 1228
rect 1373 1073 1387 1087
rect 1473 1073 1487 1087
rect 1613 1073 1627 1087
rect 1433 1053 1447 1067
rect 1333 993 1347 1007
rect 1353 953 1367 967
rect 1393 953 1407 967
rect 1433 953 1447 967
rect 1293 933 1307 947
rect 1273 914 1287 928
rect 1333 914 1347 928
rect 1293 833 1307 847
rect 1373 873 1387 887
rect 1493 1033 1507 1047
rect 1553 1033 1567 1047
rect 1613 1013 1627 1027
rect 1613 973 1627 987
rect 1573 953 1587 967
rect 1553 913 1567 927
rect 1613 914 1627 928
rect 1813 1172 1827 1186
rect 1773 1113 1787 1127
rect 1813 1113 1827 1127
rect 1713 1093 1727 1107
rect 1773 1073 1787 1087
rect 1713 1013 1727 1027
rect 1693 993 1707 1007
rect 1693 953 1707 967
rect 1693 914 1707 928
rect 1773 914 1787 928
rect 1853 1172 1867 1186
rect 1853 1033 1867 1047
rect 1833 953 1847 967
rect 1913 1173 1927 1187
rect 1873 973 1887 987
rect 2053 1172 2067 1186
rect 2153 1172 2167 1186
rect 2213 1172 2227 1186
rect 1993 1133 2007 1147
rect 2113 1133 2127 1147
rect 1973 1113 1987 1127
rect 1953 1013 1967 1027
rect 1973 953 1987 967
rect 2113 1073 2127 1087
rect 2153 1033 2167 1047
rect 2293 1392 2307 1406
rect 2313 1333 2327 1347
rect 2273 1253 2287 1267
rect 2373 1392 2387 1406
rect 2333 1273 2347 1287
rect 2313 1172 2327 1186
rect 2313 1033 2327 1047
rect 2253 973 2267 987
rect 1953 934 1967 948
rect 1973 893 1987 907
rect 1353 733 1367 747
rect 1273 693 1287 707
rect 1333 713 1347 727
rect 1473 872 1487 886
rect 1533 872 1547 886
rect 1593 872 1607 886
rect 1673 872 1687 886
rect 1713 872 1727 886
rect 1793 872 1807 886
rect 1873 872 1887 886
rect 1913 872 1927 886
rect 1613 853 1627 867
rect 1533 753 1547 767
rect 1793 851 1807 865
rect 1633 753 1647 767
rect 1413 713 1427 727
rect 1613 713 1627 727
rect 1433 694 1447 708
rect 1533 694 1547 708
rect 1673 733 1687 747
rect 1713 694 1727 708
rect 1993 833 2007 847
rect 2113 894 2127 908
rect 2253 893 2267 907
rect 2293 892 2307 906
rect 1833 773 1847 787
rect 1973 773 1987 787
rect 2013 773 2027 787
rect 2073 773 2087 787
rect 1793 673 1807 687
rect 1813 674 1827 688
rect 1173 613 1187 627
rect 1093 393 1107 407
rect 1253 652 1267 666
rect 1293 653 1307 667
rect 1293 613 1307 627
rect 1393 653 1407 667
rect 1353 633 1367 647
rect 1313 573 1327 587
rect 1213 513 1227 527
rect 1313 513 1327 527
rect 1193 453 1207 467
rect 1233 453 1247 467
rect 1373 453 1387 467
rect 1193 394 1207 408
rect 1253 433 1267 447
rect 1253 393 1267 407
rect 1293 394 1307 408
rect 1333 394 1347 408
rect 1373 393 1387 407
rect 1513 652 1527 666
rect 1453 613 1467 627
rect 1533 613 1547 627
rect 1413 533 1427 547
rect 1473 453 1487 467
rect 1453 433 1467 447
rect 1433 394 1447 408
rect 1473 393 1487 407
rect 1573 653 1587 667
rect 1573 613 1587 627
rect 1653 653 1667 667
rect 1613 633 1627 647
rect 1553 573 1567 587
rect 1593 573 1607 587
rect 1553 513 1567 527
rect 1533 413 1547 427
rect 1553 393 1567 407
rect 1633 453 1647 467
rect 1713 633 1727 647
rect 1693 593 1707 607
rect 1693 533 1707 547
rect 1733 613 1747 627
rect 1733 592 1747 606
rect 2173 753 2187 767
rect 2253 753 2267 767
rect 2113 713 2127 727
rect 1933 672 1947 686
rect 2073 672 2087 686
rect 2213 713 2227 727
rect 1773 553 1787 567
rect 1833 553 1847 567
rect 1913 553 1927 567
rect 1733 473 1747 487
rect 1653 433 1667 447
rect 1813 433 1827 447
rect 1733 394 1747 408
rect 1773 394 1787 408
rect 1853 413 1867 427
rect 1913 414 1927 428
rect 1973 413 1987 427
rect 893 313 907 327
rect 913 292 927 306
rect 993 353 1007 367
rect 993 313 1007 327
rect 953 273 967 287
rect 1013 273 1027 287
rect 873 253 887 267
rect 853 233 867 247
rect 773 213 787 227
rect 873 213 887 227
rect 733 174 747 188
rect 773 174 787 188
rect 893 174 907 188
rect 693 113 707 127
rect 813 132 827 146
rect 813 93 827 107
rect 753 73 767 87
rect 953 193 967 207
rect 953 174 967 188
rect 1092 353 1106 367
rect 1073 313 1087 327
rect 1053 253 1067 267
rect 1073 233 1087 247
rect 1033 174 1047 188
rect 1113 352 1127 366
rect 1153 293 1167 307
rect 1193 293 1207 307
rect 1273 353 1287 367
rect 1233 333 1247 347
rect 1213 273 1227 287
rect 1313 333 1327 347
rect 1373 353 1387 367
rect 1353 333 1367 347
rect 1273 293 1287 307
rect 1233 253 1247 267
rect 1333 253 1347 267
rect 1193 233 1207 247
rect 1153 213 1167 227
rect 1093 193 1107 207
rect 1213 174 1227 188
rect 1293 174 1307 188
rect 1413 273 1427 287
rect 1373 233 1387 247
rect 1433 233 1447 247
rect 1472 353 1486 367
rect 1493 353 1507 367
rect 1473 313 1487 327
rect 1593 352 1607 366
rect 1633 352 1647 366
rect 1533 313 1547 327
rect 1493 213 1507 227
rect 1453 173 1467 187
rect 1573 293 1587 307
rect 1553 233 1567 247
rect 1553 173 1567 187
rect 1793 353 1807 367
rect 1653 333 1667 347
rect 1613 213 1627 227
rect 1593 193 1607 207
rect 1773 293 1787 307
rect 1692 233 1706 247
rect 1713 213 1727 227
rect 1693 193 1707 207
rect 1653 173 1667 187
rect 1873 352 1887 366
rect 1953 333 1967 347
rect 1833 293 1847 307
rect 2053 373 2067 387
rect 2393 1172 2407 1186
rect 2333 933 2347 947
rect 2373 933 2387 947
rect 2313 753 2327 767
rect 2293 713 2307 727
rect 2373 833 2387 847
rect 2413 693 2427 707
rect 2293 652 2307 666
rect 2213 353 2227 367
rect 2253 353 2267 367
rect 1813 253 1827 267
rect 1973 253 1987 267
rect 2053 253 2067 267
rect 2093 253 2107 267
rect 2213 253 2227 267
rect 1793 233 1807 247
rect 1773 173 1787 187
rect 1193 153 1207 167
rect 1793 154 1807 168
rect 973 132 987 146
rect 1053 132 1067 146
rect 1113 132 1127 146
rect 1173 132 1187 146
rect 1193 93 1207 107
rect 913 73 927 87
rect 1353 132 1367 146
rect 1413 132 1427 146
rect 1453 133 1467 147
rect 1513 132 1527 146
rect 1593 132 1607 146
rect 1633 132 1647 146
rect 1693 132 1707 146
rect 1473 113 1487 127
rect 1553 113 1567 127
rect 1453 73 1467 87
rect 1753 112 1767 126
rect 1813 112 1827 126
rect 1913 73 1927 87
rect 2393 333 2407 347
rect 2313 233 2327 247
rect 2233 213 2247 227
rect 2153 193 2167 207
rect 2193 153 2207 167
rect 2053 53 2067 67
rect 1753 33 1767 47
rect 1313 13 1327 27
rect 1693 13 1707 27
rect 2353 132 2367 146
<< metal3 >>
rect 947 2356 1073 2364
rect 1127 2356 1273 2364
rect 1787 2356 1813 2364
rect 747 2336 853 2344
rect 967 2336 993 2344
rect 1887 2336 2393 2344
rect 1707 2316 1853 2324
rect 907 2296 1033 2304
rect 1047 2296 1113 2304
rect 1267 2296 1473 2304
rect 387 2276 833 2284
rect 1416 2276 1473 2284
rect 347 2237 373 2245
rect 976 2244 984 2254
rect 807 2236 1044 2244
rect 967 2216 1013 2224
rect 1036 2224 1044 2236
rect 1036 2216 1093 2224
rect 1196 2224 1204 2273
rect 1187 2216 1204 2224
rect 1296 2224 1304 2273
rect 1347 2256 1393 2264
rect 1416 2226 1424 2276
rect 1847 2276 1893 2284
rect 1447 2256 1513 2264
rect 1527 2256 1593 2264
rect 2347 2256 2384 2264
rect 1516 2227 1524 2254
rect 1296 2216 1313 2224
rect 1516 2216 1533 2227
rect 1520 2213 1533 2216
rect 1656 2224 1664 2254
rect 1627 2216 1664 2224
rect 1756 2207 1764 2254
rect 1813 2224 1827 2233
rect 1867 2235 1993 2243
rect 2187 2237 2273 2245
rect 2376 2227 2384 2256
rect 1807 2220 1827 2224
rect 1807 2216 1824 2220
rect 47 2196 493 2204
rect 507 2196 1093 2204
rect 1147 2196 1233 2204
rect 1287 2196 1413 2204
rect 1827 2196 1893 2204
rect 207 2176 353 2184
rect 1167 2176 1513 2184
rect 1627 2176 1713 2184
rect 407 2156 453 2164
rect 467 2156 1133 2164
rect 1267 2156 1473 2164
rect 1747 2156 1833 2164
rect 667 2136 1133 2144
rect 1427 2136 1553 2144
rect 467 2116 553 2124
rect 707 2116 853 2124
rect 907 2116 1064 2124
rect 1056 2104 1064 2116
rect 1347 2116 1673 2124
rect 1056 2096 1293 2104
rect 1307 2096 1433 2104
rect 1767 2096 2073 2104
rect 2087 2096 2253 2104
rect 107 2076 453 2084
rect 947 2076 1033 2084
rect 1047 2076 1273 2084
rect 647 2056 773 2064
rect 1107 2056 1373 2064
rect 1787 2056 1973 2064
rect 487 2036 613 2044
rect 627 2036 793 2044
rect 1587 2036 1693 2044
rect 767 2016 893 2024
rect 1467 2016 1493 2024
rect 1547 2016 1713 2024
rect 1787 2016 1873 2024
rect 1887 2016 2213 2024
rect 207 1996 453 2004
rect 547 1996 633 2004
rect 927 1996 1253 2004
rect 1267 1996 1393 2004
rect 1527 1996 1733 2004
rect 36 1927 44 1974
rect 367 1976 464 1984
rect 456 1964 464 1976
rect 587 1976 744 1984
rect 456 1956 504 1964
rect 447 1935 473 1943
rect 347 1896 373 1904
rect 387 1896 433 1904
rect 496 1904 504 1956
rect 567 1916 633 1924
rect 656 1907 664 1954
rect 696 1927 704 1953
rect 687 1916 704 1927
rect 736 1926 744 1976
rect 1036 1976 1093 1984
rect 827 1956 873 1964
rect 687 1913 700 1916
rect 496 1896 533 1904
rect 667 1896 753 1904
rect 776 1904 784 1953
rect 996 1924 1004 1954
rect 1036 1944 1044 1976
rect 1247 1976 1333 1984
rect 1567 1984 1580 1987
rect 1567 1973 1584 1984
rect 1707 1984 1720 1987
rect 1707 1973 1724 1984
rect 1847 1977 1913 1985
rect 1067 1964 1080 1967
rect 1067 1953 1084 1964
rect 1016 1936 1044 1944
rect 1016 1926 1024 1936
rect 1076 1927 1084 1953
rect 907 1916 1004 1924
rect 1136 1924 1144 1953
rect 1136 1916 1153 1924
rect 1176 1907 1184 1954
rect 1216 1944 1224 1954
rect 1293 1944 1307 1953
rect 1216 1940 1244 1944
rect 1293 1940 1324 1944
rect 1216 1936 1247 1940
rect 1296 1936 1324 1940
rect 1233 1927 1247 1936
rect 1316 1926 1324 1936
rect 1375 1907 1383 1954
rect 1396 1927 1404 1953
rect 1456 1907 1464 1973
rect 1476 1927 1484 1954
rect 1476 1916 1493 1927
rect 1480 1913 1493 1916
rect 1536 1907 1544 1954
rect 1576 1907 1584 1973
rect 1716 1964 1724 1973
rect 1716 1956 1773 1964
rect 1676 1924 1684 1954
rect 1956 1936 2052 1944
rect 1676 1916 1713 1924
rect 1956 1924 1964 1936
rect 2087 1937 2233 1945
rect 1767 1916 1964 1924
rect 776 1896 973 1904
rect 1447 1896 1464 1907
rect 1447 1893 1460 1896
rect 467 1876 513 1884
rect 1067 1876 1113 1884
rect 1207 1876 1393 1884
rect 507 1856 933 1864
rect 947 1856 1173 1864
rect 1247 1856 1353 1864
rect 1467 1856 1633 1864
rect 547 1836 713 1844
rect 1387 1836 1553 1844
rect 2253 1844 2267 1853
rect 2027 1840 2267 1844
rect 2027 1836 2264 1840
rect 407 1816 493 1824
rect 1407 1816 1493 1824
rect 1647 1816 1833 1824
rect 1147 1796 1213 1804
rect 1227 1796 1273 1804
rect 1347 1796 1373 1804
rect 1807 1796 2073 1804
rect 487 1776 793 1784
rect 1127 1784 1140 1787
rect 1127 1773 1144 1784
rect 1187 1776 1313 1784
rect 1727 1776 2213 1784
rect 1136 1764 1144 1773
rect 1136 1756 1184 1764
rect -24 1724 -16 1744
rect 27 1737 93 1745
rect 576 1736 613 1744
rect -44 1716 -16 1724
rect -44 1664 -36 1716
rect 447 1717 473 1725
rect 576 1707 584 1736
rect 640 1744 652 1747
rect 636 1733 652 1744
rect 767 1736 813 1744
rect 836 1736 853 1744
rect -24 1684 -16 1704
rect 636 1706 644 1733
rect 676 1707 684 1733
rect 836 1687 844 1736
rect 976 1704 984 1733
rect 947 1696 984 1704
rect 1016 1704 1024 1734
rect 1016 1696 1072 1704
rect 1116 1704 1124 1733
rect 1176 1706 1184 1756
rect 1267 1753 1273 1767
rect 1420 1764 1433 1767
rect 1416 1753 1433 1764
rect 1300 1744 1313 1747
rect 1227 1736 1264 1744
rect 1256 1706 1264 1736
rect 1296 1733 1313 1744
rect 1296 1706 1304 1733
rect 1356 1707 1364 1734
rect 1096 1696 1124 1704
rect 996 1687 1004 1692
rect 1096 1687 1104 1696
rect 1356 1696 1373 1707
rect 1360 1693 1373 1696
rect 1416 1706 1424 1753
rect 1456 1704 1464 1734
rect 1847 1736 1883 1744
rect 1576 1707 1584 1733
rect 1796 1707 1804 1733
rect 1875 1707 1883 1736
rect 1936 1724 1944 1734
rect 1896 1720 1944 1724
rect 1893 1716 1944 1720
rect 1893 1707 1907 1716
rect 1456 1696 1513 1704
rect 1727 1696 1793 1704
rect 1976 1706 1984 1776
rect 2227 1776 2313 1784
rect 2000 1764 2013 1767
rect 1996 1753 2013 1764
rect 2367 1764 2380 1767
rect 2367 1754 2384 1764
rect 2360 1753 2384 1754
rect -24 1676 33 1684
rect 47 1676 93 1684
rect 747 1676 813 1684
rect 836 1676 853 1687
rect 840 1673 853 1676
rect 987 1684 1004 1687
rect 987 1676 1093 1684
rect 987 1673 1000 1676
rect 1876 1684 1884 1693
rect 1967 1696 1973 1704
rect 1747 1676 1884 1684
rect 1996 1684 2004 1753
rect 2047 1736 2064 1744
rect 2056 1704 2064 1736
rect 2127 1736 2204 1744
rect 2056 1696 2172 1704
rect 2196 1706 2204 1736
rect 2216 1704 2224 1734
rect 2296 1707 2304 1733
rect 2216 1696 2272 1704
rect 2356 1687 2364 1733
rect 2376 1704 2384 1753
rect 2376 1700 2404 1704
rect 2376 1696 2407 1700
rect 2393 1687 2407 1696
rect 2427 1696 2464 1704
rect 1996 1676 2113 1684
rect -44 1656 53 1664
rect 587 1656 693 1664
rect 927 1656 1353 1664
rect 1367 1656 1393 1664
rect 1587 1656 1773 1664
rect 2187 1656 2373 1664
rect 107 1636 133 1644
rect 847 1636 1333 1644
rect 2247 1636 2353 1644
rect 887 1616 1013 1624
rect 1027 1616 1072 1624
rect 1107 1616 1373 1624
rect 1907 1616 2133 1624
rect 2347 1616 2413 1624
rect 27 1596 553 1604
rect 567 1596 633 1604
rect 1147 1596 1273 1604
rect 1287 1596 1813 1604
rect 1927 1596 2013 1604
rect 2027 1596 2073 1604
rect 247 1576 293 1584
rect 507 1576 593 1584
rect 707 1576 953 1584
rect 1087 1576 1513 1584
rect 1567 1576 1793 1584
rect 2127 1576 2233 1584
rect 1847 1556 2013 1564
rect 2107 1556 2393 1564
rect 387 1536 513 1544
rect 887 1536 933 1544
rect 1167 1536 1233 1544
rect 1247 1536 1793 1544
rect 2067 1536 2173 1544
rect 307 1516 553 1524
rect 687 1516 993 1524
rect 1387 1516 1593 1524
rect 1827 1516 1973 1524
rect 2027 1516 2333 1524
rect 507 1496 693 1504
rect 1067 1496 1113 1504
rect 1127 1496 1253 1504
rect 2207 1496 2273 1504
rect 267 1476 404 1484
rect 127 1456 184 1464
rect 36 1436 53 1444
rect 36 1407 44 1436
rect 96 1407 104 1433
rect 176 1404 184 1456
rect 376 1424 384 1434
rect 207 1416 384 1424
rect 176 1396 233 1404
rect 376 1404 384 1416
rect 396 1406 404 1476
rect 547 1476 653 1484
rect 727 1476 753 1484
rect 767 1476 973 1484
rect 1527 1476 1753 1484
rect 1867 1476 2013 1484
rect 500 1464 513 1467
rect 447 1456 484 1464
rect 347 1396 384 1404
rect 436 1387 444 1432
rect 476 1424 484 1456
rect 427 1376 444 1387
rect 456 1416 484 1424
rect 496 1453 513 1464
rect 1100 1464 1113 1467
rect 427 1373 440 1376
rect 47 1356 133 1364
rect 147 1356 353 1364
rect 367 1356 404 1364
rect 207 1336 273 1344
rect 396 1344 404 1356
rect 456 1347 464 1416
rect 496 1387 504 1453
rect 536 1407 544 1433
rect 616 1404 624 1434
rect 647 1436 704 1444
rect 696 1406 704 1436
rect 867 1437 893 1445
rect 993 1444 1007 1453
rect 1096 1454 1113 1464
rect 1096 1453 1120 1454
rect 1267 1456 1333 1464
rect 1627 1456 1733 1464
rect 1807 1456 1833 1464
rect 993 1440 1024 1444
rect 996 1436 1024 1440
rect 1016 1424 1024 1436
rect 936 1416 1024 1424
rect 616 1396 653 1404
rect 936 1387 944 1416
rect 496 1376 513 1387
rect 500 1373 513 1376
rect 867 1376 893 1384
rect 1016 1384 1024 1416
rect 1096 1404 1104 1453
rect 1127 1436 1193 1444
rect 1336 1436 1393 1444
rect 1087 1396 1104 1404
rect 1227 1396 1313 1404
rect 1336 1404 1344 1436
rect 1436 1407 1444 1433
rect 1327 1396 1373 1404
rect 1476 1404 1484 1433
rect 1476 1396 1533 1404
rect 1696 1404 1704 1434
rect 1896 1436 1933 1444
rect 1776 1407 1784 1433
rect 1896 1407 1904 1436
rect 1647 1396 1704 1404
rect 1956 1406 1964 1476
rect 2096 1476 2353 1484
rect 2040 1444 2053 1447
rect 1016 1376 1053 1384
rect 1427 1376 1593 1384
rect 1607 1376 1713 1384
rect 1727 1376 1873 1384
rect 1976 1384 1984 1434
rect 2036 1433 2053 1444
rect 2036 1406 2044 1433
rect 2096 1406 2104 1476
rect 2196 1456 2393 1464
rect 2196 1387 2204 1456
rect 2236 1407 2244 1433
rect 2236 1396 2253 1407
rect 2240 1393 2253 1396
rect 2316 1404 2324 1433
rect 2307 1396 2373 1404
rect 1976 1376 2013 1384
rect 607 1356 844 1364
rect 396 1336 433 1344
rect 456 1336 473 1347
rect 460 1333 473 1336
rect 836 1344 844 1356
rect 1007 1356 1033 1364
rect 1267 1356 1453 1364
rect 1627 1356 1693 1364
rect 836 1336 913 1344
rect 1067 1336 1253 1344
rect 1347 1336 1433 1344
rect 1547 1336 1833 1344
rect 1887 1336 2033 1344
rect 2107 1336 2313 1344
rect 27 1316 73 1324
rect 727 1316 773 1324
rect 787 1316 904 1324
rect 407 1296 533 1304
rect 896 1304 904 1316
rect 1087 1316 1173 1324
rect 1387 1316 1793 1324
rect 1907 1316 2173 1324
rect 896 1296 1013 1304
rect 1387 1296 1493 1304
rect 1647 1296 1673 1304
rect 1967 1296 2213 1304
rect 367 1276 633 1284
rect 707 1276 793 1284
rect 887 1276 933 1284
rect 1047 1276 1153 1284
rect 1707 1276 1833 1284
rect 2027 1276 2333 1284
rect 27 1256 333 1264
rect 427 1256 453 1264
rect 747 1256 773 1264
rect 947 1256 1113 1264
rect 1187 1256 1613 1264
rect 1787 1256 1853 1264
rect 2047 1256 2273 1264
rect 807 1236 853 1244
rect 1176 1236 1233 1244
rect 467 1217 533 1225
rect 587 1216 624 1224
rect 87 1196 172 1204
rect 16 1167 24 1193
rect 207 1195 352 1203
rect 387 1197 412 1205
rect 436 1184 444 1194
rect 347 1176 593 1184
rect 616 1184 624 1216
rect 695 1186 703 1233
rect 916 1216 933 1224
rect 716 1187 724 1213
rect 816 1187 824 1213
rect 616 1176 653 1184
rect 507 1156 613 1164
rect 896 1164 904 1213
rect 916 1167 924 1216
rect 1076 1216 1153 1224
rect 996 1167 1004 1214
rect 1036 1204 1044 1214
rect 1076 1204 1084 1216
rect 1176 1204 1184 1236
rect 1316 1236 1352 1244
rect 1316 1224 1324 1236
rect 1387 1236 1484 1244
rect 867 1156 904 1164
rect 987 1156 1004 1167
rect 1016 1196 1044 1204
rect 1056 1196 1084 1204
rect 1096 1200 1184 1204
rect 1093 1196 1184 1200
rect 1236 1216 1324 1224
rect 987 1153 1000 1156
rect 1016 1147 1024 1196
rect 1056 1186 1064 1196
rect 1093 1187 1107 1196
rect 1236 1187 1244 1216
rect 1227 1176 1244 1187
rect 1256 1196 1333 1204
rect 1227 1173 1240 1176
rect 1256 1167 1264 1196
rect 1476 1206 1484 1236
rect 1767 1236 1793 1244
rect 1976 1236 2024 1244
rect 1847 1216 1892 1224
rect 1916 1187 1924 1213
rect 1296 1180 1673 1184
rect 1293 1176 1673 1180
rect 1293 1167 1307 1176
rect 1827 1175 1853 1183
rect 1976 1164 1984 1236
rect 2016 1224 2024 1236
rect 2016 1216 2033 1224
rect 2056 1216 2133 1224
rect 1996 1184 2004 1214
rect 2056 1186 2064 1216
rect 2156 1216 2193 1224
rect 2156 1186 2164 1216
rect 2216 1186 2224 1233
rect 2456 1204 2464 1224
rect 2376 1196 2464 1204
rect 1996 1176 2024 1184
rect 1976 1160 2004 1164
rect 1976 1156 2007 1160
rect 1993 1147 2007 1156
rect 187 1136 413 1144
rect 436 1136 793 1144
rect 436 1124 444 1136
rect 1067 1136 1233 1144
rect 2016 1144 2024 1176
rect 2376 1184 2384 1196
rect 2327 1176 2384 1184
rect 2407 1176 2464 1184
rect 2016 1136 2113 1144
rect 207 1116 444 1124
rect 607 1116 733 1124
rect 907 1116 1193 1124
rect 1347 1116 1773 1124
rect 1827 1116 1973 1124
rect 47 1096 73 1104
rect 407 1096 753 1104
rect 867 1096 1033 1104
rect 1327 1096 1713 1104
rect 427 1076 673 1084
rect 1287 1076 1373 1084
rect 1487 1076 1613 1084
rect 1787 1076 2113 1084
rect 767 1056 893 1064
rect 1207 1056 1433 1064
rect 27 1036 93 1044
rect 407 1036 473 1044
rect 807 1036 853 1044
rect 947 1036 1073 1044
rect 1087 1036 1173 1044
rect 1187 1036 1493 1044
rect 1567 1036 1853 1044
rect 2167 1036 2313 1044
rect 627 1016 873 1024
rect 1496 1024 1504 1033
rect 1496 1016 1613 1024
rect 1727 1016 1953 1024
rect 1227 996 1333 1004
rect 1707 996 1904 1004
rect 107 976 493 984
rect 667 976 793 984
rect 967 976 1093 984
rect 1107 976 1233 984
rect 1627 976 1873 984
rect 1896 984 1904 996
rect 1896 976 2253 984
rect 727 956 784 964
rect 156 936 413 944
rect 36 907 44 934
rect 156 924 164 936
rect 547 936 753 944
rect 776 944 784 956
rect 887 956 933 964
rect 1187 956 1353 964
rect 1367 956 1393 964
rect 1447 956 1573 964
rect 1707 956 1833 964
rect 1987 964 2000 967
rect 1987 953 2004 964
rect 776 936 844 944
rect 27 896 44 907
rect 136 916 164 924
rect 27 893 40 896
rect 136 904 144 916
rect 207 920 364 924
rect 207 916 367 920
rect 353 907 367 916
rect 680 924 693 927
rect 87 896 144 904
rect 176 844 184 893
rect 496 904 504 914
rect 447 896 504 904
rect 536 884 544 914
rect 536 876 573 884
rect 616 884 624 914
rect 676 913 693 924
rect 780 924 793 927
rect 776 913 793 924
rect 676 887 684 913
rect 616 880 664 884
rect 616 876 667 880
rect 653 867 667 876
rect 776 884 784 913
rect 836 886 844 936
rect 867 936 973 944
rect 1996 944 2004 953
rect 1996 936 2333 944
rect 876 916 1033 924
rect 747 876 784 884
rect 487 856 613 864
rect 876 864 884 916
rect 1060 924 1073 927
rect 1056 913 1073 924
rect 1147 916 1173 924
rect 1196 916 1273 924
rect 1056 886 1064 913
rect 1196 904 1204 916
rect 1296 904 1304 933
rect 1096 900 1204 904
rect 1093 896 1204 900
rect 1216 896 1304 904
rect 1093 887 1107 896
rect 1216 884 1224 896
rect 1167 876 1224 884
rect 1336 884 1344 914
rect 1627 916 1693 924
rect 1336 876 1373 884
rect 1487 875 1533 883
rect 1556 884 1564 913
rect 1556 876 1593 884
rect 1687 876 1704 884
rect 787 856 884 864
rect 1067 856 1113 864
rect 1247 856 1613 864
rect 1696 864 1704 876
rect 1776 884 1784 914
rect 1956 907 1964 934
rect 2347 936 2373 944
rect 1956 896 1973 907
rect 1960 893 1973 896
rect 1727 876 1784 884
rect 1807 876 1873 884
rect 2116 884 2124 894
rect 2267 896 2293 904
rect 1927 876 2124 884
rect 1696 856 1793 864
rect 176 836 593 844
rect 1056 844 1064 853
rect 987 836 1064 844
rect 1207 836 1293 844
rect 2007 836 2373 844
rect 116 816 353 824
rect 116 804 124 816
rect 407 816 433 824
rect 667 816 693 824
rect 827 816 933 824
rect 1087 816 1153 824
rect 47 796 124 804
rect 767 796 893 804
rect 1067 796 1233 804
rect 187 776 333 784
rect 527 776 653 784
rect 1847 776 1973 784
rect 2027 776 2073 784
rect 107 756 253 764
rect 267 756 393 764
rect 436 756 573 764
rect 127 736 213 744
rect 436 744 444 756
rect 1047 756 1133 764
rect 1547 756 1633 764
rect 2187 756 2253 764
rect 2267 756 2313 764
rect 327 736 444 744
rect 707 736 773 744
rect 1167 736 1353 744
rect 1367 736 1673 744
rect 667 716 753 724
rect 1147 716 1333 724
rect 1400 724 1413 727
rect 1396 713 1413 724
rect 2127 716 2213 724
rect 2227 716 2293 724
rect -24 684 -16 704
rect 300 704 313 707
rect -24 676 4 684
rect -4 664 4 676
rect -24 624 -16 664
rect -4 656 53 664
rect 176 664 184 694
rect 296 693 313 704
rect 176 656 233 664
rect 296 664 304 693
rect 376 664 384 693
rect 476 666 484 713
rect 507 696 613 704
rect 656 696 673 704
rect 616 684 624 694
rect 596 676 624 684
rect 287 656 304 664
rect 336 656 384 664
rect 336 644 344 656
rect 427 656 473 664
rect 596 664 604 676
rect 656 667 664 696
rect 1107 696 1264 704
rect 787 676 872 684
rect 907 675 1053 683
rect 1107 677 1133 685
rect 567 656 604 664
rect 1256 666 1264 696
rect 1287 704 1300 707
rect 1287 693 1304 704
rect 1296 667 1304 693
rect 1396 667 1404 713
rect 1547 696 1584 704
rect 1436 664 1444 694
rect 1576 667 1584 696
rect 1416 656 1513 664
rect 307 636 344 644
rect 627 635 733 643
rect 1416 644 1424 656
rect 1616 647 1624 713
rect 1656 696 1713 704
rect 1656 667 1664 696
rect 2427 696 2464 704
rect 1716 676 1793 684
rect 1716 647 1724 676
rect 1807 676 1813 684
rect 1947 675 2073 683
rect 2307 656 2464 664
rect 1367 636 1424 644
rect -24 616 133 624
rect 367 616 433 624
rect 1187 616 1293 624
rect 1307 616 1453 624
rect 1467 616 1533 624
rect 1587 616 1733 624
rect 1707 596 1733 604
rect 187 576 633 584
rect 707 576 1313 584
rect 1567 576 1593 584
rect 1787 556 1833 564
rect 1847 556 1913 564
rect 27 536 233 544
rect 247 536 613 544
rect 987 536 1033 544
rect 1427 536 1693 544
rect 1007 516 1213 524
rect 1327 516 1553 524
rect 27 496 273 504
rect 16 476 113 484
rect 16 364 24 476
rect 827 476 1053 484
rect 1067 476 1733 484
rect 607 456 632 464
rect 667 456 853 464
rect 867 456 1193 464
rect 1247 456 1373 464
rect 1487 456 1633 464
rect 47 436 73 444
rect 556 436 692 444
rect 47 396 84 404
rect 16 356 53 364
rect 76 347 84 396
rect 107 396 224 404
rect 216 367 224 396
rect 236 387 244 414
rect 407 416 533 424
rect 556 387 564 436
rect 727 436 773 444
rect 1087 436 1253 444
rect 1267 436 1453 444
rect 1667 436 1813 444
rect 1236 416 1344 424
rect 236 376 253 387
rect 240 373 253 376
rect 736 384 744 394
rect 787 404 800 407
rect 980 404 993 407
rect 787 393 804 404
rect 796 384 804 393
rect 976 393 993 404
rect 1016 396 1033 404
rect 736 380 784 384
rect 736 376 787 380
rect 796 376 824 384
rect 773 367 787 376
rect 307 356 573 364
rect 667 355 752 363
rect 816 364 824 376
rect 816 356 833 364
rect 976 364 984 393
rect 1016 384 1024 396
rect 1056 384 1064 413
rect 996 380 1024 384
rect 887 356 984 364
rect 993 376 1024 380
rect 1036 376 1064 384
rect 993 367 1007 376
rect 1036 364 1044 376
rect 1096 367 1104 393
rect 1016 356 1044 364
rect 1016 344 1024 356
rect 1196 364 1204 394
rect 1127 356 1204 364
rect 1236 347 1244 416
rect 1336 408 1344 416
rect 1496 416 1533 424
rect 867 336 1024 344
rect 1256 344 1264 393
rect 1296 367 1304 394
rect 1376 367 1384 393
rect 1287 356 1304 367
rect 1287 353 1300 356
rect 1256 336 1313 344
rect 1436 344 1444 394
rect 1476 367 1484 393
rect 1496 367 1504 416
rect 1716 416 1853 424
rect 1567 396 1604 404
rect 1596 366 1604 396
rect 1716 384 1724 416
rect 1927 416 1973 424
rect 1636 376 1724 384
rect 1636 366 1644 376
rect 1367 336 1444 344
rect 1736 344 1744 394
rect 1776 367 1784 394
rect 1776 356 1793 367
rect 1780 353 1793 356
rect 2053 364 2067 373
rect 1887 360 2067 364
rect 1887 356 2064 360
rect 2227 356 2253 364
rect 1667 336 1744 344
rect 1967 336 2393 344
rect 907 316 993 324
rect 1007 316 1073 324
rect 1487 316 1533 324
rect 927 296 1153 304
rect 1207 296 1273 304
rect 1287 296 1573 304
rect 1787 296 1833 304
rect 267 276 413 284
rect 467 276 573 284
rect 967 276 1013 284
rect 1227 276 1413 284
rect 287 256 464 264
rect 456 247 464 256
rect 547 256 713 264
rect 887 256 1053 264
rect 1247 256 1333 264
rect 1827 256 1973 264
rect 2067 256 2093 264
rect 2107 256 2213 264
rect 456 236 473 247
rect 460 233 473 236
rect 607 236 693 244
rect 747 236 853 244
rect 1087 236 1193 244
rect 1387 236 1433 244
rect 1447 236 1553 244
rect 1567 236 1692 244
rect 1716 236 1793 244
rect 1716 227 1724 236
rect 1807 236 2313 244
rect 787 216 873 224
rect 1167 216 1493 224
rect 1627 216 1713 224
rect 2156 216 2233 224
rect 2156 207 2164 216
rect 967 196 1093 204
rect 1496 196 1593 204
rect 87 176 513 184
rect 647 177 733 185
rect 907 176 953 184
rect 1176 176 1213 184
rect 156 147 164 154
rect 187 155 273 163
rect 156 146 180 147
rect -24 136 33 144
rect 156 136 173 146
rect 160 133 173 136
rect 776 144 784 174
rect 776 136 813 144
rect 1036 144 1044 174
rect 1176 146 1184 176
rect 1296 164 1304 174
rect 1207 156 1304 164
rect 1456 147 1464 173
rect 987 136 1044 144
rect 1067 136 1113 144
rect 1367 136 1413 144
rect 1496 127 1504 196
rect 1707 196 2153 204
rect 1760 184 1773 187
rect 1756 173 1773 184
rect 1556 144 1564 173
rect 1527 136 1544 144
rect 1556 136 1593 144
rect 567 116 693 124
rect 1487 116 1504 127
rect 1536 127 1544 136
rect 1656 144 1664 173
rect 1647 136 1664 144
rect 1756 144 1764 173
rect 1807 156 2193 164
rect 1707 136 1764 144
rect 2367 136 2464 144
rect 1536 116 1553 127
rect 1487 113 1500 116
rect 1540 113 1553 116
rect 1767 115 1813 123
rect 827 96 1193 104
rect 587 84 600 87
rect 587 73 604 84
rect 767 76 913 84
rect 1467 76 1913 84
rect 127 56 413 64
rect 596 64 604 73
rect 427 56 564 64
rect 596 56 2053 64
rect 556 44 564 56
rect 556 36 1753 44
rect 187 16 473 24
rect 487 16 533 24
rect 1327 16 1693 24
use INVX1  _122_
timestamp 0
transform -1 0 1430 0 1 1310
box -6 -8 46 268
use NAND3X1  _123_
timestamp 0
transform -1 0 2410 0 1 1310
box -6 -8 86 268
use NOR2X1  _124_
timestamp 0
transform -1 0 1230 0 1 1310
box -6 -8 66 268
use AND2X2  _125_
timestamp 0
transform -1 0 1130 0 1 1310
box -6 -8 86 268
use INVX1  _126_
timestamp 0
transform 1 0 1690 0 -1 1830
box -6 -8 46 268
use AOI21X1  _127_
timestamp 0
transform 1 0 1650 0 1 790
box -6 -8 86 268
use NAND2X1  _128_
timestamp 0
transform -1 0 2170 0 -1 1310
box -6 -8 66 268
use INVX1  _129_
timestamp 0
transform 1 0 2190 0 -1 1310
box -6 -8 46 268
use MUX2X1  _130_
timestamp 0
transform 1 0 1870 0 -1 1310
box -6 -8 106 268
use OAI21X1  _131_
timestamp 0
transform 1 0 1990 0 -1 1310
box -6 -8 86 268
use INVX1  _132_
timestamp 0
transform -1 0 2310 0 1 1310
box -6 -8 46 268
use NAND2X1  _133_
timestamp 0
transform 1 0 1810 0 -1 1830
box -6 -8 66 268
use NAND2X1  _134_
timestamp 0
transform -1 0 1970 0 -1 1830
box -6 -8 66 268
use OAI21X1  _135_
timestamp 0
transform 1 0 2070 0 -1 1830
box -6 -8 86 268
use NAND2X1  _136_
timestamp 0
transform -1 0 2370 0 -1 2350
box -6 -8 66 268
use NAND3X1  _137_
timestamp 0
transform 1 0 1970 0 -1 1830
box -6 -8 86 268
use OAI22X1  _138_
timestamp 0
transform 1 0 2310 0 -1 1830
box -6 -8 106 268
use AOI21X1  _139_
timestamp 0
transform 1 0 2190 0 -1 1830
box -6 -8 86 268
use NAND2X1  _140_
timestamp 0
transform 1 0 1570 0 1 790
box -6 -8 66 268
use NAND2X1  _141_
timestamp 0
transform -1 0 1830 0 1 790
box -6 -8 66 268
use INVX1  _142_
timestamp 0
transform -1 0 2050 0 1 1310
box -6 -8 46 268
use INVX1  _143_
timestamp 0
transform 1 0 2090 0 1 1310
box -6 -8 46 268
use OAI21X1  _144_
timestamp 0
transform -1 0 2230 0 1 1310
box -6 -8 86 268
use NAND3X1  _145_
timestamp 0
transform -1 0 1990 0 1 1310
box -6 -8 86 268
use NAND3X1  _146_
timestamp 0
transform 1 0 1850 0 1 790
box -6 -8 86 268
use AND2X2  _147_
timestamp 0
transform 1 0 1270 0 1 1310
box -6 -8 86 268
use OAI21X1  _148_
timestamp 0
transform 1 0 1790 0 1 1310
box -6 -8 86 268
use NAND3X1  _149_
timestamp 0
transform 1 0 1570 0 1 1310
box -6 -8 86 268
use NAND2X1  _150_
timestamp 0
transform 1 0 1770 0 -1 1310
box -6 -8 66 268
use AND2X2  _151_
timestamp 0
transform 1 0 1690 0 1 1310
box -6 -8 86 268
use OAI21X1  _152_
timestamp 0
transform 1 0 1450 0 1 1310
box -6 -8 86 268
use DFFSR  _153_
timestamp 0
transform 1 0 1750 0 -1 790
box -6 -8 466 268
use DFFSR  _154_
timestamp 0
transform 1 0 1890 0 1 1830
box -6 -8 466 268
use DFFSR  _155_
timestamp 0
transform 1 0 1930 0 1 790
box -6 -8 466 268
use DFFSR  _156_
timestamp 0
transform 1 0 1290 0 -1 1310
box -6 -8 466 268
use INVX1  _157_
timestamp 0
transform -1 0 90 0 1 1310
box -6 -8 46 268
use NAND3X1  _158_
timestamp 0
transform -1 0 290 0 -1 790
box -6 -8 86 268
use NOR2X1  _159_
timestamp 0
transform 1 0 470 0 1 1310
box -6 -8 66 268
use AND2X2  _160_
timestamp 0
transform 1 0 950 0 1 1310
box -6 -8 86 268
use INVX1  _161_
timestamp 0
transform -1 0 1070 0 1 790
box -6 -8 46 268
use AOI21X1  _162_
timestamp 0
transform -1 0 1070 0 -1 1310
box -6 -8 86 268
use NAND2X1  _163_
timestamp 0
transform 1 0 30 0 1 270
box -6 -8 66 268
use INVX1  _164_
timestamp 0
transform -1 0 590 0 -1 790
box -6 -8 46 268
use MUX2X1  _165_
timestamp 0
transform -1 0 710 0 -1 790
box -6 -8 106 268
use OAI21X1  _166_
timestamp 0
transform -1 0 210 0 1 270
box -6 -8 86 268
use INVX1  _167_
timestamp 0
transform 1 0 390 0 -1 790
box -6 -8 46 268
use NAND2X1  _168_
timestamp 0
transform 1 0 1230 0 -1 1310
box -6 -8 66 268
use NAND2X1  _169_
timestamp 0
transform -1 0 870 0 1 790
box -6 -8 66 268
use OAI21X1  _170_
timestamp 0
transform -1 0 790 0 1 790
box -6 -8 86 268
use NAND2X1  _171_
timestamp 0
transform -1 0 550 0 1 790
box -6 -8 66 268
use NAND3X1  _172_
timestamp 0
transform -1 0 1190 0 -1 1310
box -6 -8 86 268
use OAI22X1  _173_
timestamp 0
transform -1 0 990 0 1 790
box -6 -8 106 268
use AOI21X1  _174_
timestamp 0
transform -1 0 670 0 1 790
box -6 -8 86 268
use NAND2X1  _175_
timestamp 0
transform -1 0 890 0 -1 1310
box -6 -8 66 268
use NAND2X1  _176_
timestamp 0
transform 1 0 750 0 -1 1310
box -6 -8 66 268
use INVX1  _177_
timestamp 0
transform -1 0 950 0 -1 1310
box -6 -8 46 268
use INVX1  _178_
timestamp 0
transform 1 0 330 0 -1 790
box -6 -8 46 268
use OAI21X1  _179_
timestamp 0
transform -1 0 510 0 -1 790
box -6 -8 86 268
use NAND3X1  _180_
timestamp 0
transform 1 0 510 0 -1 1310
box -6 -8 86 268
use NAND3X1  _181_
timestamp 0
transform -1 0 710 0 -1 1310
box -6 -8 86 268
use AND2X2  _182_
timestamp 0
transform -1 0 190 0 1 1310
box -6 -8 86 268
use OAI21X1  _183_
timestamp 0
transform 1 0 350 0 1 1310
box -6 -8 86 268
use NAND3X1  _184_
timestamp 0
transform -1 0 730 0 1 1310
box -6 -8 86 268
use NAND2X1  _185_
timestamp 0
transform -1 0 950 0 1 1310
box -6 -8 66 268
use AND2X2  _186_
timestamp 0
transform -1 0 630 0 1 1310
box -6 -8 86 268
use OAI21X1  _187_
timestamp 0
transform 1 0 230 0 1 1310
box -6 -8 86 268
use DFFSR  _188_
timestamp 0
transform 1 0 90 0 -1 270
box -6 -8 466 268
use DFFSR  _189_
timestamp 0
transform 1 0 10 0 1 790
box -6 -8 466 268
use DFFSR  _190_
timestamp 0
transform 1 0 10 0 -1 1310
box -6 -8 466 268
use DFFSR  _191_
timestamp 0
transform 1 0 110 0 -1 1830
box -6 -8 466 268
use INVX1  _192_
timestamp 0
transform 1 0 1750 0 -1 1830
box -6 -8 46 268
use NAND3X1  _193_
timestamp 0
transform -1 0 1150 0 -1 2350
box -6 -8 86 268
use NOR2X1  _194_
timestamp 0
transform -1 0 1530 0 -1 2350
box -6 -8 66 268
use AND2X2  _195_
timestamp 0
transform 1 0 1410 0 -1 1830
box -6 -8 86 268
use INVX1  _196_
timestamp 0
transform -1 0 1370 0 -1 1830
box -6 -8 46 268
use AOI21X1  _197_
timestamp 0
transform -1 0 890 0 -1 1830
box -6 -8 86 268
use NAND2X1  _198_
timestamp 0
transform 1 0 590 0 -1 1830
box -6 -8 66 268
use INVX1  _199_
timestamp 0
transform -1 0 970 0 -1 1830
box -6 -8 46 268
use MUX2X1  _200_
timestamp 0
transform 1 0 750 0 1 1310
box -6 -8 106 268
use OAI21X1  _201_
timestamp 0
transform -1 0 770 0 -1 1830
box -6 -8 86 268
use INVX1  _202_
timestamp 0
transform -1 0 1290 0 1 1830
box -6 -8 46 268
use NAND2X1  _203_
timestamp 0
transform 1 0 1510 0 -1 1830
box -6 -8 66 268
use NAND2X1  _204_
timestamp 0
transform -1 0 1590 0 1 1830
box -6 -8 66 268
use OAI21X1  _205_
timestamp 0
transform 1 0 1310 0 1 1830
box -6 -8 86 268
use NAND2X1  _206_
timestamp 0
transform -1 0 1310 0 -1 1830
box -6 -8 66 268
use NAND3X1  _207_
timestamp 0
transform 1 0 990 0 -1 1830
box -6 -8 86 268
use OAI22X1  _208_
timestamp 0
transform 1 0 1110 0 -1 1830
box -6 -8 106 268
use AOI21X1  _209_
timestamp 0
transform -1 0 1230 0 1 1830
box -6 -8 86 268
use NAND2X1  _210_
timestamp 0
transform 1 0 710 0 1 1830
box -6 -8 66 268
use NAND2X1  _211_
timestamp 0
transform 1 0 610 0 1 1830
box -6 -8 66 268
use INVX1  _212_
timestamp 0
transform -1 0 1130 0 1 1830
box -6 -8 46 268
use INVX1  _213_
timestamp 0
transform 1 0 790 0 1 1830
box -6 -8 46 268
use OAI21X1  _214_
timestamp 0
transform -1 0 950 0 1 1830
box -6 -8 86 268
use NAND3X1  _215_
timestamp 0
transform -1 0 1050 0 1 1830
box -6 -8 86 268
use NAND3X1  _216_
timestamp 0
transform -1 0 590 0 1 1830
box -6 -8 86 268
use AND2X2  _217_
timestamp 0
transform 1 0 1550 0 -1 2350
box -6 -8 86 268
use OAI21X1  _218_
timestamp 0
transform -1 0 1450 0 -1 2350
box -6 -8 86 268
use NAND3X1  _219_
timestamp 0
transform -1 0 1790 0 1 1830
box -6 -8 86 268
use NAND2X1  _220_
timestamp 0
transform -1 0 1490 0 1 1830
box -6 -8 66 268
use AND2X2  _221_
timestamp 0
transform -1 0 1690 0 1 1830
box -6 -8 86 268
use OAI21X1  _222_
timestamp 0
transform 1 0 1650 0 -1 2350
box -6 -8 86 268
use DFFSR  _223_
timestamp 0
transform 1 0 10 0 -1 2350
box -6 -8 466 268
use DFFSR  _224_
timestamp 0
transform 1 0 470 0 -1 2350
box -6 -8 466 268
use DFFSR  _225_
timestamp 0
transform 1 0 10 0 1 1830
box -6 -8 466 268
use DFFSR  _226_
timestamp 0
transform 1 0 1810 0 -1 2350
box -6 -8 466 268
use INVX1  _227_
timestamp 0
transform 1 0 950 0 -1 270
box -6 -8 46 268
use NAND3X1  _228_
timestamp 0
transform -1 0 1650 0 -1 270
box -6 -8 86 268
use NOR2X1  _229_
timestamp 0
transform 1 0 1030 0 -1 270
box -6 -8 66 268
use AND2X2  _230_
timestamp 0
transform 1 0 1110 0 -1 270
box -6 -8 86 268
use INVX1  _231_
timestamp 0
transform 1 0 1110 0 1 790
box -6 -8 46 268
use AOI21X1  _232_
timestamp 0
transform -1 0 1190 0 1 270
box -6 -8 86 268
use NAND2X1  _233_
timestamp 0
transform 1 0 810 0 1 270
box -6 -8 66 268
use INVX1  _234_
timestamp 0
transform -1 0 850 0 -1 270
box -6 -8 46 268
use MUX2X1  _235_
timestamp 0
transform 1 0 690 0 -1 270
box -6 -8 106 268
use OAI21X1  _236_
timestamp 0
transform -1 0 770 0 1 270
box -6 -8 86 268
use INVX1  _237_
timestamp 0
transform -1 0 1730 0 -1 270
box -6 -8 46 268
use NAND2X1  _238_
timestamp 0
transform -1 0 1470 0 -1 790
box -6 -8 66 268
use NAND2X1  _239_
timestamp 0
transform -1 0 1570 0 -1 790
box -6 -8 66 268
use OAI21X1  _240_
timestamp 0
transform 1 0 1670 0 -1 790
box -6 -8 86 268
use NAND2X1  _241_
timestamp 0
transform 1 0 1730 0 1 270
box -6 -8 66 268
use NAND3X1  _242_
timestamp 0
transform 1 0 1470 0 -1 270
box -6 -8 86 268
use OAI22X1  _243_
timestamp 0
transform 1 0 1590 0 1 270
box -6 -8 106 268
use AOI21X1  _244_
timestamp 0
transform 1 0 1810 0 1 270
box -6 -8 86 268
use NAND2X1  _245_
timestamp 0
transform -1 0 1450 0 1 790
box -6 -8 66 268
use NAND2X1  _246_
timestamp 0
transform -1 0 1250 0 1 270
box -6 -8 66 268
use INVX1  _247_
timestamp 0
transform -1 0 1550 0 1 270
box -6 -8 46 268
use INVX1  _248_
timestamp 0
transform -1 0 1450 0 -1 270
box -6 -8 46 268
use OAI21X1  _249_
timestamp 0
transform 1 0 1290 0 -1 270
box -6 -8 86 268
use NAND3X1  _250_
timestamp 0
transform 1 0 1290 0 1 270
box -6 -8 86 268
use NAND3X1  _251_
timestamp 0
transform 1 0 1390 0 1 270
box -6 -8 86 268
use AND2X2  _252_
timestamp 0
transform 1 0 910 0 1 270
box -6 -8 86 268
use OAI21X1  _253_
timestamp 0
transform 1 0 1010 0 1 270
box -6 -8 86 268
use NAND3X1  _254_
timestamp 0
transform 1 0 1310 0 -1 790
box -6 -8 86 268
use NAND2X1  _255_
timestamp 0
transform -1 0 1230 0 1 790
box -6 -8 66 268
use AND2X2  _256_
timestamp 0
transform -1 0 1350 0 1 790
box -6 -8 86 268
use OAI21X1  _257_
timestamp 0
transform 1 0 1190 0 -1 790
box -6 -8 86 268
use DFFSR  _258_
timestamp 0
transform 1 0 210 0 1 270
box -6 -8 466 268
use DFFSR  _259_
timestamp 0
transform 1 0 1890 0 1 270
box -6 -8 466 268
use DFFSR  _260_
timestamp 0
transform 1 0 1730 0 -1 270
box -6 -8 466 268
use DFFSR  _261_
timestamp 0
transform 1 0 710 0 -1 790
box -6 -8 466 268
use BUFX2  _262_
timestamp 0
transform 1 0 2250 0 -1 790
box -6 -8 66 268
use BUFX2  _263_
timestamp 0
transform 1 0 2350 0 -1 1310
box -6 -8 66 268
use BUFX2  _264_
timestamp 0
transform 1 0 970 0 -1 2350
box -6 -8 66 268
use BUFX2  _265_
timestamp 0
transform 1 0 1750 0 -1 2350
box -6 -8 66 268
use BUFX2  _266_
timestamp 0
transform -1 0 650 0 -1 270
box -6 -8 66 268
use BUFX2  _267_
timestamp 0
transform 1 0 2310 0 -1 270
box -6 -8 66 268
use BUFX2  _268_
timestamp 0
transform 1 0 2230 0 -1 270
box -6 -8 66 268
use BUFX2  _269_
timestamp 0
transform -1 0 910 0 -1 270
box -6 -8 66 268
use BUFX2  _270_
timestamp 0
transform 1 0 2350 0 -1 790
box -6 -8 66 268
use BUFX2  _271_
timestamp 0
transform 1 0 2270 0 -1 1310
box -6 -8 66 268
use BUFX2  _272_
timestamp 0
transform -1 0 90 0 -1 270
box -6 -8 66 268
use BUFX2  _273_
timestamp 0
transform -1 0 110 0 -1 790
box -6 -8 66 268
use BUFX2  _274_
timestamp 0
transform -1 0 190 0 -1 790
box -6 -8 66 268
use BUFX2  _275_
timestamp 0
transform -1 0 110 0 -1 1830
box -6 -8 66 268
use BUFX2  _276_
timestamp 0
transform -1 0 1230 0 -1 2350
box -6 -8 66 268
use BUFX2  _277_
timestamp 0
transform 1 0 1270 0 -1 2350
box -6 -8 66 268
use BUFX2  _278_
timestamp 0
transform 1 0 1210 0 -1 270
box -6 -8 66 268
use BUFX2  BUFX2_insert0
timestamp 0
transform -1 0 1650 0 -1 1830
box -6 -8 66 268
use BUFX2  BUFX2_insert1
timestamp 0
transform -1 0 1550 0 1 790
box -6 -8 66 268
use BUFX2  BUFX2_insert2
timestamp 0
transform -1 0 1650 0 -1 790
box -6 -8 66 268
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 1830 0 1 1830
box -6 -8 66 268
use FILL  FILL35250x4050
timestamp 0
transform 1 0 2350 0 1 270
box -6 -8 26 268
use FILL  FILL35250x27450
timestamp 0
transform 1 0 2350 0 1 1830
box -6 -8 26 268
use FILL  FILL35550x150
timestamp 0
transform -1 0 2390 0 -1 270
box -6 -8 26 268
use FILL  FILL35550x4050
timestamp 0
transform 1 0 2370 0 1 270
box -6 -8 26 268
use FILL  FILL35550x27450
timestamp 0
transform 1 0 2370 0 1 1830
box -6 -8 26 268
use FILL  FILL35550x31350
timestamp 0
transform -1 0 2390 0 -1 2350
box -6 -8 26 268
use FILL  FILL35850x150
timestamp 0
transform -1 0 2410 0 -1 270
box -6 -8 26 268
use FILL  FILL35850x4050
timestamp 0
transform 1 0 2390 0 1 270
box -6 -8 26 268
use FILL  FILL35850x11850
timestamp 0
transform 1 0 2390 0 1 790
box -6 -8 26 268
use FILL  FILL35850x27450
timestamp 0
transform 1 0 2390 0 1 1830
box -6 -8 26 268
use FILL  FILL35850x31350
timestamp 0
transform -1 0 2410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__122_
timestamp 0
transform -1 0 1370 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__123_
timestamp 0
transform -1 0 2330 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__124_
timestamp 0
transform -1 0 1150 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__125_
timestamp 0
transform -1 0 1050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__126_
timestamp 0
transform 1 0 1650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__127_
timestamp 0
transform 1 0 1630 0 1 790
box -6 -8 26 268
use FILL  FILL_0__128_
timestamp 0
transform -1 0 2090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__129_
timestamp 0
transform 1 0 2170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__130_
timestamp 0
transform 1 0 1830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__131_
timestamp 0
transform 1 0 1970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__132_
timestamp 0
transform -1 0 2250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__133_
timestamp 0
transform 1 0 1790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__134_
timestamp 0
transform -1 0 1890 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__135_
timestamp 0
transform 1 0 2050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__136_
timestamp 0
transform -1 0 2290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__138_
timestamp 0
transform 1 0 2270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__139_
timestamp 0
transform 1 0 2150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__140_
timestamp 0
transform 1 0 1550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__141_
timestamp 0
transform -1 0 1750 0 1 790
box -6 -8 26 268
use FILL  FILL_0__142_
timestamp 0
transform -1 0 2010 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__143_
timestamp 0
transform 1 0 2050 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__144_
timestamp 0
transform -1 0 2150 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__145_
timestamp 0
transform -1 0 1890 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__146_
timestamp 0
transform 1 0 1830 0 1 790
box -6 -8 26 268
use FILL  FILL_0__147_
timestamp 0
transform 1 0 1230 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__148_
timestamp 0
transform 1 0 1770 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__149_
timestamp 0
transform 1 0 1530 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__150_
timestamp 0
transform 1 0 1750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__151_
timestamp 0
transform 1 0 1650 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__152_
timestamp 0
transform 1 0 1430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__157_
timestamp 0
transform -1 0 30 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__158_
timestamp 0
transform -1 0 210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__159_
timestamp 0
transform 1 0 430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__161_
timestamp 0
transform -1 0 1010 0 1 790
box -6 -8 26 268
use FILL  FILL_0__162_
timestamp 0
transform -1 0 970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__163_
timestamp 0
transform 1 0 10 0 1 270
box -6 -8 26 268
use FILL  FILL_0__164_
timestamp 0
transform -1 0 530 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__165_
timestamp 0
transform -1 0 610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__166_
timestamp 0
transform -1 0 110 0 1 270
box -6 -8 26 268
use FILL  FILL_0__167_
timestamp 0
transform 1 0 370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__168_
timestamp 0
transform 1 0 1190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__169_
timestamp 0
transform -1 0 810 0 1 790
box -6 -8 26 268
use FILL  FILL_0__170_
timestamp 0
transform -1 0 690 0 1 790
box -6 -8 26 268
use FILL  FILL_0__171_
timestamp 0
transform -1 0 490 0 1 790
box -6 -8 26 268
use FILL  FILL_0__172_
timestamp 0
transform -1 0 1090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__173_
timestamp 0
transform -1 0 890 0 1 790
box -6 -8 26 268
use FILL  FILL_0__174_
timestamp 0
transform -1 0 570 0 1 790
box -6 -8 26 268
use FILL  FILL_0__175_
timestamp 0
transform -1 0 830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__176_
timestamp 0
transform 1 0 710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__177_
timestamp 0
transform -1 0 910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__178_
timestamp 0
transform 1 0 290 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__180_
timestamp 0
transform 1 0 470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__181_
timestamp 0
transform -1 0 610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__182_
timestamp 0
transform -1 0 110 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__183_
timestamp 0
transform 1 0 310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__184_
timestamp 0
transform -1 0 650 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__185_
timestamp 0
transform -1 0 870 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__186_
timestamp 0
transform -1 0 550 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__187_
timestamp 0
transform 1 0 190 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__192_
timestamp 0
transform 1 0 1730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__193_
timestamp 0
transform -1 0 1050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__194_
timestamp 0
transform -1 0 1470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__195_
timestamp 0
transform 1 0 1370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__196_
timestamp 0
transform -1 0 1330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__197_
timestamp 0
transform -1 0 790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__198_
timestamp 0
transform 1 0 570 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__199_
timestamp 0
transform -1 0 910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__200_
timestamp 0
transform 1 0 730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__201_
timestamp 0
transform -1 0 670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__202_
timestamp 0
transform -1 0 1250 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__203_
timestamp 0
transform 1 0 1490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__204_
timestamp 0
transform -1 0 1510 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__205_
timestamp 0
transform 1 0 1290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__206_
timestamp 0
transform -1 0 1230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__207_
timestamp 0
transform 1 0 970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__208_
timestamp 0
transform 1 0 1070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__209_
timestamp 0
transform -1 0 1150 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__210_
timestamp 0
transform 1 0 670 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__211_
timestamp 0
transform 1 0 590 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__212_
timestamp 0
transform -1 0 1070 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__213_
timestamp 0
transform 1 0 770 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__214_
timestamp 0
transform -1 0 850 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__215_
timestamp 0
transform -1 0 970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__216_
timestamp 0
transform -1 0 490 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__217_
timestamp 0
transform 1 0 1530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__218_
timestamp 0
transform -1 0 1350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__219_
timestamp 0
transform -1 0 1710 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__220_
timestamp 0
transform -1 0 1410 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__221_
timestamp 0
transform -1 0 1610 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__222_
timestamp 0
transform 1 0 1630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__227_
timestamp 0
transform 1 0 910 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__228_
timestamp 0
transform -1 0 1570 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__229_
timestamp 0
transform 1 0 990 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__230_
timestamp 0
transform 1 0 1090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__231_
timestamp 0
transform 1 0 1070 0 1 790
box -6 -8 26 268
use FILL  FILL_0__232_
timestamp 0
transform -1 0 1110 0 1 270
box -6 -8 26 268
use FILL  FILL_0__233_
timestamp 0
transform 1 0 770 0 1 270
box -6 -8 26 268
use FILL  FILL_0__234_
timestamp 0
transform -1 0 810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__235_
timestamp 0
transform 1 0 650 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__236_
timestamp 0
transform -1 0 690 0 1 270
box -6 -8 26 268
use FILL  FILL_0__237_
timestamp 0
transform -1 0 1670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__238_
timestamp 0
transform -1 0 1410 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__239_
timestamp 0
transform -1 0 1490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__240_
timestamp 0
transform 1 0 1650 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__241_
timestamp 0
transform 1 0 1690 0 1 270
box -6 -8 26 268
use FILL  FILL_0__242_
timestamp 0
transform 1 0 1450 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__243_
timestamp 0
transform 1 0 1550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__244_
timestamp 0
transform 1 0 1790 0 1 270
box -6 -8 26 268
use FILL  FILL_0__245_
timestamp 0
transform -1 0 1370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__247_
timestamp 0
transform -1 0 1490 0 1 270
box -6 -8 26 268
use FILL  FILL_0__248_
timestamp 0
transform -1 0 1390 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__249_
timestamp 0
transform 1 0 1270 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__250_
timestamp 0
transform 1 0 1250 0 1 270
box -6 -8 26 268
use FILL  FILL_0__251_
timestamp 0
transform 1 0 1370 0 1 270
box -6 -8 26 268
use FILL  FILL_0__252_
timestamp 0
transform 1 0 870 0 1 270
box -6 -8 26 268
use FILL  FILL_0__253_
timestamp 0
transform 1 0 990 0 1 270
box -6 -8 26 268
use FILL  FILL_0__254_
timestamp 0
transform 1 0 1270 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__255_
timestamp 0
transform -1 0 1170 0 1 790
box -6 -8 26 268
use FILL  FILL_0__256_
timestamp 0
transform -1 0 1250 0 1 790
box -6 -8 26 268
use FILL  FILL_0__257_
timestamp 0
transform 1 0 1170 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__262_
timestamp 0
transform 1 0 2210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__263_
timestamp 0
transform 1 0 2330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__264_
timestamp 0
transform 1 0 930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__265_
timestamp 0
transform 1 0 1730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__266_
timestamp 0
transform -1 0 570 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__267_
timestamp 0
transform 1 0 2290 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__268_
timestamp 0
transform 1 0 2190 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__270_
timestamp 0
transform 1 0 2310 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__271_
timestamp 0
transform 1 0 2230 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__272_
timestamp 0
transform -1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__273_
timestamp 0
transform -1 0 30 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__274_
timestamp 0
transform -1 0 130 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__275_
timestamp 0
transform -1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__276_
timestamp 0
transform -1 0 1170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__277_
timestamp 0
transform 1 0 1230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__278_
timestamp 0
transform 1 0 1190 0 -1 270
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform -1 0 1590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform -1 0 1470 0 1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform -1 0 1590 0 -1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 1790 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__122_
timestamp 0
transform -1 0 1390 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__124_
timestamp 0
transform -1 0 1170 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__126_
timestamp 0
transform 1 0 1670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__128_
timestamp 0
transform -1 0 2110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__130_
timestamp 0
transform 1 0 1850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__132_
timestamp 0
transform -1 0 2270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__134_
timestamp 0
transform -1 0 1910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__136_
timestamp 0
transform -1 0 2310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__138_
timestamp 0
transform 1 0 2290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__139_
timestamp 0
transform 1 0 2170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__141_
timestamp 0
transform -1 0 1770 0 1 790
box -6 -8 26 268
use FILL  FILL_1__143_
timestamp 0
transform 1 0 2070 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__145_
timestamp 0
transform -1 0 1910 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__147_
timestamp 0
transform 1 0 1250 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__149_
timestamp 0
transform 1 0 1550 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__151_
timestamp 0
transform 1 0 1670 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__157_
timestamp 0
transform -1 0 50 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__159_
timestamp 0
transform 1 0 450 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__161_
timestamp 0
transform -1 0 1030 0 1 790
box -6 -8 26 268
use FILL  FILL_1__162_
timestamp 0
transform -1 0 990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__164_
timestamp 0
transform -1 0 550 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__166_
timestamp 0
transform -1 0 130 0 1 270
box -6 -8 26 268
use FILL  FILL_1__168_
timestamp 0
transform 1 0 1210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__170_
timestamp 0
transform -1 0 710 0 1 790
box -6 -8 26 268
use FILL  FILL_1__172_
timestamp 0
transform -1 0 1110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__174_
timestamp 0
transform -1 0 590 0 1 790
box -6 -8 26 268
use FILL  FILL_1__176_
timestamp 0
transform 1 0 730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__178_
timestamp 0
transform 1 0 310 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__180_
timestamp 0
transform 1 0 490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__181_
timestamp 0
transform -1 0 630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__183_
timestamp 0
transform 1 0 330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__185_
timestamp 0
transform -1 0 890 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__187_
timestamp 0
transform 1 0 210 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__193_
timestamp 0
transform -1 0 1070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__195_
timestamp 0
transform 1 0 1390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__197_
timestamp 0
transform -1 0 810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__199_
timestamp 0
transform -1 0 930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__201_
timestamp 0
transform -1 0 690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__204_
timestamp 0
transform -1 0 1530 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__206_
timestamp 0
transform -1 0 1250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__208_
timestamp 0
transform 1 0 1090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__210_
timestamp 0
transform 1 0 690 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__212_
timestamp 0
transform -1 0 1090 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__214_
timestamp 0
transform -1 0 870 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__216_
timestamp 0
transform -1 0 510 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__218_
timestamp 0
transform -1 0 1370 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__220_
timestamp 0
transform -1 0 1430 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__227_
timestamp 0
transform 1 0 930 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__229_
timestamp 0
transform 1 0 1010 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__231_
timestamp 0
transform 1 0 1090 0 1 790
box -6 -8 26 268
use FILL  FILL_1__233_
timestamp 0
transform 1 0 790 0 1 270
box -6 -8 26 268
use FILL  FILL_1__235_
timestamp 0
transform 1 0 670 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__237_
timestamp 0
transform -1 0 1690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__239_
timestamp 0
transform -1 0 1510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__241_
timestamp 0
transform 1 0 1710 0 1 270
box -6 -8 26 268
use FILL  FILL_1__243_
timestamp 0
transform 1 0 1570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__245_
timestamp 0
transform -1 0 1390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__247_
timestamp 0
transform -1 0 1510 0 1 270
box -6 -8 26 268
use FILL  FILL_1__248_
timestamp 0
transform -1 0 1410 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__250_
timestamp 0
transform 1 0 1270 0 1 270
box -6 -8 26 268
use FILL  FILL_1__252_
timestamp 0
transform 1 0 890 0 1 270
box -6 -8 26 268
use FILL  FILL_1__254_
timestamp 0
transform 1 0 1290 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__256_
timestamp 0
transform -1 0 1270 0 1 790
box -6 -8 26 268
use FILL  FILL_1__262_
timestamp 0
transform 1 0 2230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__264_
timestamp 0
transform 1 0 950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__266_
timestamp 0
transform -1 0 590 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__268_
timestamp 0
transform 1 0 2210 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__270_
timestamp 0
transform 1 0 2330 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__271_
timestamp 0
transform 1 0 2250 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__273_
timestamp 0
transform -1 0 50 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__275_
timestamp 0
transform -1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__277_
timestamp 0
transform 1 0 1250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform -1 0 1490 0 1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform 1 0 1810 0 1 1830
box -6 -8 26 268
<< labels >>
flabel metal1 s 2423 2 2483 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 2157 2397 2163 2403 3 FreeSans 16 90 0 0 CLK
port 2 nsew
flabel metal2 s 1477 2397 1483 2403 3 FreeSans 16 90 0 0 Din[3]
port 3 nsew
flabel metal2 s 737 2397 743 2403 3 FreeSans 16 90 0 0 Din[2]
port 4 nsew
flabel metal3 s 2456 1696 2464 1704 3 FreeSans 16 0 0 0 Din[1]
port 5 nsew
flabel metal2 s 697 -23 703 -17 7 FreeSans 16 270 0 0 Din[0]
port 6 nsew
flabel metal2 s 877 -23 883 -17 7 FreeSans 16 270 0 0 Dout[15]
port 7 nsew
flabel metal2 s 2257 -23 2263 -17 7 FreeSans 16 270 0 0 Dout[14]
port 8 nsew
flabel metal3 s 2456 136 2464 144 3 FreeSans 16 0 0 0 Dout[13]
port 9 nsew
flabel metal2 s 617 -23 623 -17 7 FreeSans 16 270 0 0 Dout[12]
port 10 nsew
flabel metal2 s 1777 2397 1783 2403 3 FreeSans 16 90 0 0 Dout[11]
port 11 nsew
flabel metal2 s 997 2397 1003 2403 3 FreeSans 16 90 0 0 Dout[10]
port 12 nsew
flabel metal2 s 1297 2397 1303 2403 3 FreeSans 16 90 0 0 Dout[9]
port 13 nsew
flabel metal2 s 1197 2397 1203 2403 3 FreeSans 16 90 0 0 Dout[8]
port 14 nsew
flabel metal3 s -24 1736 -16 1744 7 FreeSans 16 0 0 0 Dout[7]
port 15 nsew
flabel metal3 s -24 656 -16 664 7 FreeSans 16 0 0 0 Dout[6]
port 16 nsew
flabel metal3 s -24 696 -16 704 7 FreeSans 16 0 0 0 Dout[5]
port 17 nsew
flabel metal3 s -24 136 -16 144 7 FreeSans 16 0 0 0 Dout[4]
port 18 nsew
flabel metal3 s 2456 1216 2464 1224 3 FreeSans 16 0 0 0 Dout[3]
port 19 nsew
flabel metal3 s 2456 696 2464 704 3 FreeSans 16 0 0 0 Dout[2]
port 20 nsew
flabel metal3 s 2456 1176 2464 1184 3 FreeSans 16 0 0 0 Dout[1]
port 21 nsew
flabel metal3 s 2456 656 2464 664 3 FreeSans 16 0 0 0 Dout[0]
port 22 nsew
flabel metal2 s 1237 -23 1243 -17 7 FreeSans 16 270 0 0 RCO
port 23 nsew
flabel metal3 s -24 1696 -16 1704 7 FreeSans 16 0 0 0 nCLR
port 24 nsew
flabel metal2 s 1837 2397 1843 2403 3 FreeSans 16 90 0 0 nLOAD
port 25 nsew
<< properties >>
string FIXED_BBOX -40 -40 2460 2400
<< end >>
