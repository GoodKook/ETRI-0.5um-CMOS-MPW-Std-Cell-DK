magic
tech scmos
magscale 1 3
timestamp 1537935238
<< checkpaint >>
rect -60 -60 330 330
<< nwell >>
rect 0 0 270 270
<< pdiffusion >>
rect 85 85 185 185
<< nsubstratendiff >>
rect 20 230 250 250
rect 20 40 40 230
rect 230 40 250 230
rect 20 20 250 40
<< metal1 >>
rect 20 230 250 250
rect 20 40 40 230
rect 85 85 185 185
rect 230 40 250 230
rect 20 20 250 40
use ntap_CDNS_7046768260514  ntap_CDNS_7046768260514_0
timestamp 1537935238
transform 1 0 226 0 1 36
box 4 4 24 194
use ntap_CDNS_7046768260514  ntap_CDNS_7046768260514_1
timestamp 1537935238
transform 0 1 36 1 0 16
box 4 4 24 194
use ntap_CDNS_7046768260514  ntap_CDNS_7046768260514_2
timestamp 1537935238
transform 0 1 36 1 0 226
box 4 4 24 194
use ntap_CDNS_7046768260514  ntap_CDNS_7046768260514_3
timestamp 1537935238
transform 1 0 16 0 1 36
box 4 4 24 194
use ptap_CDNS_7046768260515  ptap_CDNS_7046768260515_0
timestamp 1537935238
transform 1 0 81 0 1 81
box 4 4 104 104
<< end >>
