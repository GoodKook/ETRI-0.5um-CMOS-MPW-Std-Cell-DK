magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -15 -15 455 455
<< nwell >>
rect 110 110 330 330
<< pdiffusion >>
rect 195 195 245 245
<< psubstratepdiff >>
rect 45 375 395 395
rect 45 65 65 375
rect 375 65 395 375
rect 45 45 395 65
<< nsubstratendiff >>
rect 130 290 310 310
rect 130 150 150 290
rect 290 150 310 290
rect 130 130 310 150
<< metal1 >>
rect 45 375 395 395
rect 45 65 65 375
rect 130 290 310 310
rect 130 150 150 290
rect 195 195 245 245
rect 290 150 310 290
rect 130 130 310 150
rect 375 65 395 375
rect 45 45 395 65
use ntap_CDNS_7230122529117  ntap_CDNS_7230122529117_0
timestamp 1554524574
transform 1 0 286 0 1 146
box 4 4 24 144
use ntap_CDNS_7230122529117  ntap_CDNS_7230122529117_1
timestamp 1554524574
transform 0 1 146 1 0 126
box 4 4 24 144
use ntap_CDNS_7230122529117  ntap_CDNS_7230122529117_2
timestamp 1554524574
transform 0 1 146 1 0 286
box 4 4 24 144
use ntap_CDNS_7230122529117  ntap_CDNS_7230122529117_3
timestamp 1554524574
transform 1 0 126 0 1 146
box 4 4 24 144
use ptap_CDNS_7230122529118  ptap_CDNS_7230122529118_0
timestamp 1554524574
transform 0 1 71 1 0 41
box 4 4 24 294
use ptap_CDNS_7230122529118  ptap_CDNS_7230122529118_1
timestamp 1554524574
transform 1 0 41 0 1 71
box 4 4 24 294
use ptap_CDNS_7230122529118  ptap_CDNS_7230122529118_2
timestamp 1554524574
transform 0 1 71 1 0 371
box 4 4 24 294
use ptap_CDNS_7230122529118  ptap_CDNS_7230122529118_3
timestamp 1554524574
transform 1 0 371 0 1 71
box 4 4 24 294
use ptap_CDNS_7230122529119  ptap_CDNS_7230122529119_0
timestamp 1554524574
transform 1 0 191 0 1 191
box 4 4 54 54
<< end >>
