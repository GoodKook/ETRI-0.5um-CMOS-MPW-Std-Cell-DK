/* Verilog module written by vlog2Verilog (qflow) */

module fir_pe(Cin, Rdy, Vld, Xin, Xout, Yin, Yout, clk);
    input [5:0] Cin;
    input Rdy;
    output Vld;
    input [3:0] Xin;
    output [3:0] Xout;
    input [3:0] Yin;
    output [3:0] Yout;
    input clk;

wire vdd = 1'b1;
wire gnd = 1'b0;

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire [4:0] LoadCtl ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire [7:0] XinHL ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire Cin_1_bF$buf0 ;
wire Cin_1_bF$buf1 ;
wire Cin_1_bF$buf2 ;
wire Cin_1_bF$buf3 ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire LoadCtl_0_bF$buf0 ;
wire LoadCtl_0_bF$buf1 ;
wire LoadCtl_0_bF$buf2 ;
wire LoadCtl_0_bF$buf3 ;
wire LoadCtl_0_bF$buf4 ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire [3:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire [3:0] Yin0 ;
wire [3:0] Yin1 ;
wire [3:0] Yin2 ;
wire [3:0] Yin3 ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire [3:0] XinH ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire [3:0] Yout ;
wire [3:0] _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire [3:0] Xout ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire LoadCtl_4_bF$buf0 ;
wire LoadCtl_4_bF$buf1 ;
wire LoadCtl_4_bF$buf2 ;
wire LoadCtl_4_bF$buf3 ;
wire LoadCtl_4_bF$buf4 ;
wire LoadCtl_4_bF$buf5 ;
wire LoadCtl_4_bF$buf6 ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire Vld ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire [5:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire [3:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire [3:0] _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire [13:0] mul ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _135__bF$buf0 ;
wire _135__bF$buf1 ;
wire _135__bF$buf2 ;
wire _135__bF$buf3 ;
wire _135__bF$buf4 ;
wire _135__bF$buf5 ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire [15:0] rYin ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert33 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf0)
);

BUFX2 BUFX2_insert32 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf1)
);

BUFX2 BUFX2_insert31 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf2)
);

BUFX2 BUFX2_insert30 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf3)
);

BUFX2 BUFX2_insert29 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf0)
);

BUFX2 BUFX2_insert28 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf1)
);

BUFX2 BUFX2_insert27 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf2)
);

BUFX2 BUFX2_insert26 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf3)
);

BUFX2 BUFX2_insert25 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf4)
);

BUFX2 BUFX2_insert24 (
    .A(_135_),
    .Y(_135__bF$buf0)
);

BUFX2 BUFX2_insert23 (
    .A(_135_),
    .Y(_135__bF$buf1)
);

BUFX2 BUFX2_insert22 (
    .A(_135_),
    .Y(_135__bF$buf2)
);

BUFX2 BUFX2_insert21 (
    .A(_135_),
    .Y(_135__bF$buf3)
);

BUFX2 BUFX2_insert20 (
    .A(_135_),
    .Y(_135__bF$buf4)
);

BUFX2 BUFX2_insert19 (
    .A(_135_),
    .Y(_135__bF$buf5)
);

BUFX2 BUFX2_insert18 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

BUFX2 BUFX2_insert17 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert16 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert15 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert14 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert11 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert10 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert9 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert8 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert7 (
    .A(clk),
    .Y(clk_bF$buf7)
);

BUFX2 BUFX2_insert6 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf0)
);

BUFX2 BUFX2_insert5 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf1)
);

BUFX2 BUFX2_insert4 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf2)
);

BUFX2 BUFX2_insert3 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf3)
);

BUFX2 BUFX2_insert2 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf4)
);

BUFX2 BUFX2_insert1 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf5)
);

BUFX2 BUFX2_insert0 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf6)
);

NAND3X1 _1000_ (
    .A(_312_),
    .B(_309_),
    .C(_311_),
    .Y(_313_)
);

NAND3X1 _1001_ (
    .A(_308_),
    .B(_313_),
    .C(_302_),
    .Y(_314_)
);

AOI22X1 _1002_ (
    .A(XinH[0]),
    .B(Cin_1_bF$buf3),
    .C(XinH[1]),
    .D(Cin_0_bF$buf3),
    .Y(_315_)
);

OAI21X1 _1003_ (
    .A(_249_),
    .B(_315_),
    .C(_256_),
    .Y(_316_)
);

AOI22X1 _1004_ (
    .A(XinH[0]),
    .B(Cin[2]),
    .C(_311_),
    .D(_312_),
    .Y(_317_)
);

AOI21X1 _1005_ (
    .A(_305_),
    .B(_307_),
    .C(_303_),
    .Y(_318_)
);

OAI21X1 _1006_ (
    .A(_318_),
    .B(_317_),
    .C(_316_),
    .Y(_319_)
);

NAND3X1 _1007_ (
    .A(_300_),
    .B(_314_),
    .C(_319_),
    .Y(_320_)
);

AND2X2 _1008_ (
    .A(_295_),
    .B(_299_),
    .Y(_321_)
);

NAND3X1 _1009_ (
    .A(_308_),
    .B(_316_),
    .C(_313_),
    .Y(_322_)
);

OAI21X1 _1010_ (
    .A(_318_),
    .B(_317_),
    .C(_302_),
    .Y(_323_)
);

NAND3X1 _1011_ (
    .A(_322_),
    .B(_323_),
    .C(_321_),
    .Y(_324_)
);

NAND3X1 _1012_ (
    .A(_320_),
    .B(_324_),
    .C(_289_),
    .Y(_325_)
);

AOI21X1 _1013_ (
    .A(_258_),
    .B(_253_),
    .C(_247_),
    .Y(_326_)
);

OAI21X1 _1014_ (
    .A(_246_),
    .B(_326_),
    .C(_265_),
    .Y(_327_)
);

AOI21X1 _1015_ (
    .A(_323_),
    .B(_322_),
    .C(_321_),
    .Y(_328_)
);

AOI21X1 _1016_ (
    .A(_319_),
    .B(_314_),
    .C(_300_),
    .Y(_329_)
);

OAI21X1 _1017_ (
    .A(_328_),
    .B(_329_),
    .C(_327_),
    .Y(_330_)
);

NAND3X1 _1018_ (
    .A(_287_),
    .B(_330_),
    .C(_325_),
    .Y(_331_)
);

NAND3X1 _1019_ (
    .A(_320_),
    .B(_327_),
    .C(_324_),
    .Y(_332_)
);

OAI21X1 _1020_ (
    .A(_328_),
    .B(_329_),
    .C(_289_),
    .Y(_333_)
);

NAND3X1 _1021_ (
    .A(_286_),
    .B(_332_),
    .C(_333_),
    .Y(_334_)
);

NAND2X1 _1022_ (
    .A(_334_),
    .B(_331_),
    .Y(_335_)
);

XNOR2X1 _1023_ (
    .A(_335_),
    .B(_284_),
    .Y(_336_)
);

NOR2X1 _1024_ (
    .A(_282_),
    .B(_336_),
    .Y(_337_)
);

NAND3X1 _1025_ (
    .A(_334_),
    .B(_331_),
    .C(_284_),
    .Y(_338_)
);

INVX1 _1026_ (
    .A(_274_),
    .Y(_339_)
);

AOI21X1 _1027_ (
    .A(_234_),
    .B(_275_),
    .C(_339_),
    .Y(_340_)
);

AOI21X1 _1028_ (
    .A(_333_),
    .B(_332_),
    .C(_286_),
    .Y(_341_)
);

AOI21X1 _1029_ (
    .A(_325_),
    .B(_330_),
    .C(_287_),
    .Y(_342_)
);

OAI21X1 _1030_ (
    .A(_341_),
    .B(_342_),
    .C(_340_),
    .Y(_343_)
);

NAND3X1 _1031_ (
    .A(_338_),
    .B(_282_),
    .C(_343_),
    .Y(_344_)
);

NAND2X1 _1032_ (
    .A(LoadCtl_4_bF$buf6),
    .B(_344_),
    .Y(_345_)
);

OAI22X1 _1033_ (
    .A(_281_),
    .B(LoadCtl_4_bF$buf5),
    .C(_345_),
    .D(_337_),
    .Y(_26_)
);

OAI21X1 _1034_ (
    .A(_340_),
    .B(_335_),
    .C(_344_),
    .Y(_346_)
);

INVX1 _1035_ (
    .A(_332_),
    .Y(_347_)
);

AOI21X1 _1036_ (
    .A(_286_),
    .B(_333_),
    .C(_347_),
    .Y(_348_)
);

NAND2X1 _1037_ (
    .A(_297_),
    .B(_299_),
    .Y(_349_)
);

INVX1 _1038_ (
    .A(_349_),
    .Y(_350_)
);

INVX1 _1039_ (
    .A(_322_),
    .Y(_351_)
);

AOI21X1 _1040_ (
    .A(_321_),
    .B(_323_),
    .C(_351_),
    .Y(_352_)
);

NAND2X1 _1041_ (
    .A(XinHL[2]),
    .B(Cin[5]),
    .Y(_353_)
);

AND2X2 _1042_ (
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_354_)
);

OAI21X1 _1043_ (
    .A(_179_),
    .B(_214_),
    .C(_354_),
    .Y(_355_)
);

AND2X2 _1044_ (
    .A(XinHL[3]),
    .B(Cin[4]),
    .Y(_356_)
);

OAI21X1 _1045_ (
    .A(_89_),
    .B(_239_),
    .C(_356_),
    .Y(_357_)
);

NAND3X1 _1046_ (
    .A(_353_),
    .B(_355_),
    .C(_357_),
    .Y(_358_)
);

INVX1 _1047_ (
    .A(_353_),
    .Y(_359_)
);

NAND2X1 _1048_ (
    .A(_356_),
    .B(_354_),
    .Y(_360_)
);

NAND2X1 _1049_ (
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_361_)
);

OAI21X1 _1050_ (
    .A(_179_),
    .B(_214_),
    .C(_361_),
    .Y(_362_)
);

NAND3X1 _1051_ (
    .A(_362_),
    .B(_359_),
    .C(_360_),
    .Y(_363_)
);

NAND2X1 _1052_ (
    .A(_363_),
    .B(_358_),
    .Y(_364_)
);

AOI22X1 _1053_ (
    .A(_255_),
    .B(_310_),
    .C(_312_),
    .D(_309_),
    .Y(_365_)
);

NAND2X1 _1054_ (
    .A(XinH[1]),
    .B(Cin[2]),
    .Y(_366_)
);

NAND2X1 _1055_ (
    .A(XinH[3]),
    .B(Cin_1_bF$buf2),
    .Y(_367_)
);

NOR2X1 _1056_ (
    .A(_306_),
    .B(_367_),
    .Y(_368_)
);

AOI22X1 _1057_ (
    .A(XinH[2]),
    .B(Cin_1_bF$buf1),
    .C(XinH[3]),
    .D(Cin_0_bF$buf2),
    .Y(_369_)
);

OAI21X1 _1058_ (
    .A(_369_),
    .B(_368_),
    .C(_366_),
    .Y(_370_)
);

INVX1 _1059_ (
    .A(_366_),
    .Y(_371_)
);

AND2X2 _1060_ (
    .A(XinH[3]),
    .B(Cin_0_bF$buf1),
    .Y(_372_)
);

NAND2X1 _1061_ (
    .A(_310_),
    .B(_372_),
    .Y(_373_)
);

INVX1 _1062_ (
    .A(_369_),
    .Y(_374_)
);

NAND3X1 _1063_ (
    .A(_371_),
    .B(_374_),
    .C(_373_),
    .Y(_375_)
);

NAND3X1 _1064_ (
    .A(_375_),
    .B(_365_),
    .C(_370_),
    .Y(_376_)
);

AOI22X1 _1065_ (
    .A(XinH[1]),
    .B(Cin_1_bF$buf0),
    .C(XinH[2]),
    .D(Cin_0_bF$buf0),
    .Y(_377_)
);

OAI21X1 _1066_ (
    .A(_303_),
    .B(_377_),
    .C(_311_),
    .Y(_378_)
);

AOI21X1 _1067_ (
    .A(_373_),
    .B(_374_),
    .C(_371_),
    .Y(_379_)
);

OAI21X1 _1068_ (
    .A(_93_),
    .B(_151_),
    .C(_372_),
    .Y(_380_)
);

OAI21X1 _1069_ (
    .A(_95_),
    .B(_180_),
    .C(_310_),
    .Y(_381_)
);

AOI21X1 _1070_ (
    .A(_380_),
    .B(_381_),
    .C(_366_),
    .Y(_382_)
);

OAI21X1 _1071_ (
    .A(_379_),
    .B(_382_),
    .C(_378_),
    .Y(_383_)
);

NAND3X1 _1072_ (
    .A(_364_),
    .B(_376_),
    .C(_383_),
    .Y(_384_)
);

AND2X2 _1073_ (
    .A(_358_),
    .B(_363_),
    .Y(_385_)
);

NAND3X1 _1074_ (
    .A(_378_),
    .B(_375_),
    .C(_370_),
    .Y(_386_)
);

OAI21X1 _1075_ (
    .A(_379_),
    .B(_382_),
    .C(_365_),
    .Y(_387_)
);

NAND3X1 _1076_ (
    .A(_386_),
    .B(_385_),
    .C(_387_),
    .Y(_388_)
);

NAND3X1 _1077_ (
    .A(_384_),
    .B(_388_),
    .C(_352_),
    .Y(_389_)
);

AOI21X1 _1078_ (
    .A(_313_),
    .B(_308_),
    .C(_316_),
    .Y(_390_)
);

OAI21X1 _1079_ (
    .A(_300_),
    .B(_390_),
    .C(_322_),
    .Y(_391_)
);

AOI21X1 _1080_ (
    .A(_387_),
    .B(_386_),
    .C(_385_),
    .Y(_392_)
);

AOI21X1 _1081_ (
    .A(_383_),
    .B(_376_),
    .C(_364_),
    .Y(_393_)
);

OAI21X1 _1082_ (
    .A(_392_),
    .B(_393_),
    .C(_391_),
    .Y(_394_)
);

AOI21X1 _1083_ (
    .A(_389_),
    .B(_394_),
    .C(_350_),
    .Y(_395_)
);

NAND3X1 _1084_ (
    .A(_391_),
    .B(_384_),
    .C(_388_),
    .Y(_396_)
);

OAI21X1 _1085_ (
    .A(_392_),
    .B(_393_),
    .C(_352_),
    .Y(_397_)
);

AOI21X1 _1086_ (
    .A(_397_),
    .B(_396_),
    .C(_349_),
    .Y(_398_)
);

OAI21X1 _1087_ (
    .A(_398_),
    .B(_395_),
    .C(_348_),
    .Y(_399_)
);

AOI21X1 _1088_ (
    .A(_324_),
    .B(_320_),
    .C(_327_),
    .Y(_400_)
);

OAI21X1 _1089_ (
    .A(_287_),
    .B(_400_),
    .C(_332_),
    .Y(_401_)
);

NAND3X1 _1090_ (
    .A(_349_),
    .B(_396_),
    .C(_397_),
    .Y(_402_)
);

NAND3X1 _1091_ (
    .A(_350_),
    .B(_394_),
    .C(_389_),
    .Y(_403_)
);

NAND3X1 _1092_ (
    .A(_401_),
    .B(_402_),
    .C(_403_),
    .Y(_404_)
);

NAND2X1 _1093_ (
    .A(_404_),
    .B(_399_),
    .Y(_405_)
);

XOR2X1 _1094_ (
    .A(_346_),
    .B(_405_),
    .Y(_406_)
);

NAND2X1 _1095_ (
    .A(mul[7]),
    .B(_135__bF$buf5),
    .Y(_407_)
);

OAI21X1 _1096_ (
    .A(_135__bF$buf4),
    .B(_406_),
    .C(_407_),
    .Y(_27_)
);

NAND2X1 _1097_ (
    .A(mul[8]),
    .B(_135__bF$buf3),
    .Y(_408_)
);

NAND2X1 _1098_ (
    .A(_404_),
    .B(_338_),
    .Y(_409_)
);

NAND2X1 _1099_ (
    .A(_399_),
    .B(_409_),
    .Y(_410_)
);

OAI21X1 _1100_ (
    .A(_405_),
    .B(_344_),
    .C(_410_),
    .Y(_411_)
);

AOI21X1 _1101_ (
    .A(_388_),
    .B(_384_),
    .C(_391_),
    .Y(_412_)
);

OAI21X1 _1102_ (
    .A(_350_),
    .B(_412_),
    .C(_396_),
    .Y(_413_)
);

NAND2X1 _1103_ (
    .A(_360_),
    .B(_363_),
    .Y(_414_)
);

INVX1 _1104_ (
    .A(_414_),
    .Y(_415_)
);

INVX1 _1105_ (
    .A(_386_),
    .Y(_416_)
);

AOI21X1 _1106_ (
    .A(_385_),
    .B(_387_),
    .C(_416_),
    .Y(_417_)
);

INVX2 _1107_ (
    .A(Cin[5]),
    .Y(_418_)
);

NOR2X1 _1108_ (
    .A(_179_),
    .B(_418_),
    .Y(_419_)
);

AND2X2 _1109_ (
    .A(XinH[1]),
    .B(Cin[4]),
    .Y(_420_)
);

AOI22X1 _1110_ (
    .A(XinH[0]),
    .B(Cin[4]),
    .C(XinH[1]),
    .D(Cin[3]),
    .Y(_421_)
);

AOI21X1 _1111_ (
    .A(_354_),
    .B(_420_),
    .C(_421_),
    .Y(_422_)
);

XNOR2X1 _1112_ (
    .A(_422_),
    .B(_419_),
    .Y(_423_)
);

AOI21X1 _1113_ (
    .A(_371_),
    .B(_374_),
    .C(_368_),
    .Y(_424_)
);

NAND2X1 _1114_ (
    .A(XinH[2]),
    .B(Cin_1_bF$buf3),
    .Y(_425_)
);

NAND2X1 _1115_ (
    .A(XinH[3]),
    .B(Cin[2]),
    .Y(_426_)
);

NAND2X1 _1116_ (
    .A(XinH[2]),
    .B(Cin[2]),
    .Y(_427_)
);

OAI21X1 _1117_ (
    .A(_95_),
    .B(_151_),
    .C(_427_),
    .Y(_428_)
);

OAI21X1 _1118_ (
    .A(_425_),
    .B(_426_),
    .C(_428_),
    .Y(_429_)
);

NOR2X1 _1119_ (
    .A(_429_),
    .B(_424_),
    .Y(_430_)
);

OAI21X1 _1120_ (
    .A(_366_),
    .B(_369_),
    .C(_373_),
    .Y(_431_)
);

XOR2X1 _1121_ (
    .A(_367_),
    .B(_427_),
    .Y(_432_)
);

NOR2X1 _1122_ (
    .A(_431_),
    .B(_432_),
    .Y(_433_)
);

OAI21X1 _1123_ (
    .A(_433_),
    .B(_430_),
    .C(_423_),
    .Y(_434_)
);

XOR2X1 _1124_ (
    .A(_422_),
    .B(_419_),
    .Y(_435_)
);

OAI21X1 _1125_ (
    .A(_368_),
    .B(_382_),
    .C(_432_),
    .Y(_436_)
);

NAND2X1 _1126_ (
    .A(_429_),
    .B(_424_),
    .Y(_437_)
);

NAND3X1 _1127_ (
    .A(_437_),
    .B(_435_),
    .C(_436_),
    .Y(_438_)
);

NAND3X1 _1128_ (
    .A(_434_),
    .B(_438_),
    .C(_417_),
    .Y(_439_)
);

AOI21X1 _1129_ (
    .A(_370_),
    .B(_375_),
    .C(_378_),
    .Y(_440_)
);

OAI21X1 _1130_ (
    .A(_364_),
    .B(_440_),
    .C(_386_),
    .Y(_441_)
);

AOI21X1 _1131_ (
    .A(_436_),
    .B(_437_),
    .C(_435_),
    .Y(_442_)
);

NAND2X1 _1132_ (
    .A(_432_),
    .B(_424_),
    .Y(_443_)
);

OAI21X1 _1133_ (
    .A(_368_),
    .B(_382_),
    .C(_429_),
    .Y(_444_)
);

AOI21X1 _1134_ (
    .A(_444_),
    .B(_443_),
    .C(_423_),
    .Y(_445_)
);

OAI21X1 _1135_ (
    .A(_442_),
    .B(_445_),
    .C(_441_),
    .Y(_446_)
);

NAND3X1 _1136_ (
    .A(_415_),
    .B(_446_),
    .C(_439_),
    .Y(_447_)
);

NAND3X1 _1137_ (
    .A(_438_),
    .B(_434_),
    .C(_441_),
    .Y(_448_)
);

OAI21X1 _1138_ (
    .A(_442_),
    .B(_445_),
    .C(_417_),
    .Y(_449_)
);

NAND3X1 _1139_ (
    .A(_414_),
    .B(_448_),
    .C(_449_),
    .Y(_450_)
);

NAND3X1 _1140_ (
    .A(_413_),
    .B(_450_),
    .C(_447_),
    .Y(_451_)
);

INVX1 _1141_ (
    .A(_413_),
    .Y(_452_)
);

AOI21X1 _1142_ (
    .A(_449_),
    .B(_448_),
    .C(_414_),
    .Y(_453_)
);

AOI21X1 _1143_ (
    .A(_439_),
    .B(_446_),
    .C(_415_),
    .Y(_454_)
);

OAI21X1 _1144_ (
    .A(_453_),
    .B(_454_),
    .C(_452_),
    .Y(_455_)
);

NAND2X1 _1145_ (
    .A(_451_),
    .B(_455_),
    .Y(_456_)
);

XOR2X1 _1146_ (
    .A(_411_),
    .B(_456_),
    .Y(_457_)
);

OAI21X1 _1147_ (
    .A(_135__bF$buf2),
    .B(_457_),
    .C(_408_),
    .Y(_28_)
);

INVX1 _1148_ (
    .A(_451_),
    .Y(_458_)
);

AOI21X1 _1149_ (
    .A(_411_),
    .B(_455_),
    .C(_458_),
    .Y(_459_)
);

AOI22X1 _1150_ (
    .A(_354_),
    .B(_420_),
    .C(_422_),
    .D(_419_),
    .Y(_460_)
);

INVX1 _1151_ (
    .A(_460_),
    .Y(_461_)
);

OAI21X1 _1152_ (
    .A(_433_),
    .B(_423_),
    .C(_436_),
    .Y(_462_)
);

NOR2X1 _1153_ (
    .A(_89_),
    .B(_418_),
    .Y(_463_)
);

NAND2X1 _1154_ (
    .A(XinH[1]),
    .B(Cin[4]),
    .Y(_464_)
);

NAND2X1 _1155_ (
    .A(XinH[2]),
    .B(Cin[3]),
    .Y(_465_)
);

OR2X2 _1156_ (
    .A(_464_),
    .B(_465_),
    .Y(_466_)
);

OAI21X1 _1157_ (
    .A(_93_),
    .B(_239_),
    .C(_464_),
    .Y(_467_)
);

NAND3X1 _1158_ (
    .A(_463_),
    .B(_467_),
    .C(_466_),
    .Y(_468_)
);

NAND2X1 _1159_ (
    .A(XinH[1]),
    .B(Cin[3]),
    .Y(_469_)
);

NAND2X1 _1160_ (
    .A(XinH[2]),
    .B(Cin[4]),
    .Y(_470_)
);

OAI21X1 _1161_ (
    .A(_469_),
    .B(_470_),
    .C(_467_),
    .Y(_471_)
);

OAI21X1 _1162_ (
    .A(_89_),
    .B(_418_),
    .C(_471_),
    .Y(_472_)
);

NAND2X1 _1163_ (
    .A(_468_),
    .B(_472_),
    .Y(_473_)
);

OAI21X1 _1164_ (
    .A(_310_),
    .B(_426_),
    .C(_473_),
    .Y(_474_)
);

NOR2X1 _1165_ (
    .A(_426_),
    .B(_310_),
    .Y(_475_)
);

NAND3X1 _1166_ (
    .A(_468_),
    .B(_475_),
    .C(_472_),
    .Y(_476_)
);

NAND3X1 _1167_ (
    .A(_476_),
    .B(_474_),
    .C(_462_),
    .Y(_477_)
);

AOI21X1 _1168_ (
    .A(_435_),
    .B(_437_),
    .C(_430_),
    .Y(_478_)
);

AOI21X1 _1169_ (
    .A(_472_),
    .B(_468_),
    .C(_475_),
    .Y(_479_)
);

INVX1 _1170_ (
    .A(_476_),
    .Y(_480_)
);

OAI21X1 _1171_ (
    .A(_479_),
    .B(_480_),
    .C(_478_),
    .Y(_481_)
);

NAND3X1 _1172_ (
    .A(_461_),
    .B(_477_),
    .C(_481_),
    .Y(_482_)
);

NAND3X1 _1173_ (
    .A(_476_),
    .B(_474_),
    .C(_478_),
    .Y(_483_)
);

OAI21X1 _1174_ (
    .A(_479_),
    .B(_480_),
    .C(_462_),
    .Y(_484_)
);

NAND3X1 _1175_ (
    .A(_460_),
    .B(_483_),
    .C(_484_),
    .Y(_485_)
);

NAND2X1 _1176_ (
    .A(_482_),
    .B(_485_),
    .Y(_486_)
);

NAND3X1 _1177_ (
    .A(_448_),
    .B(_450_),
    .C(_486_),
    .Y(_487_)
);

AOI21X1 _1178_ (
    .A(_434_),
    .B(_438_),
    .C(_441_),
    .Y(_488_)
);

OAI21X1 _1179_ (
    .A(_415_),
    .B(_488_),
    .C(_448_),
    .Y(_489_)
);

NAND3X1 _1180_ (
    .A(_482_),
    .B(_485_),
    .C(_489_),
    .Y(_490_)
);

AND2X2 _1181_ (
    .A(_487_),
    .B(_490_),
    .Y(_491_)
);

XOR2X1 _1182_ (
    .A(_459_),
    .B(_491_),
    .Y(_492_)
);

NAND2X1 _1183_ (
    .A(mul[9]),
    .B(_135__bF$buf1),
    .Y(_493_)
);

OAI21X1 _1184_ (
    .A(_135__bF$buf0),
    .B(_492_),
    .C(_493_),
    .Y(_29_)
);

INVX1 _1185_ (
    .A(mul[10]),
    .Y(_494_)
);

NAND2X1 _1186_ (
    .A(_490_),
    .B(_487_),
    .Y(_495_)
);

NOR2X1 _1187_ (
    .A(_495_),
    .B(_456_),
    .Y(_496_)
);

NAND2X1 _1188_ (
    .A(_490_),
    .B(_451_),
    .Y(_497_)
);

NAND2X1 _1189_ (
    .A(_487_),
    .B(_497_),
    .Y(_498_)
);

INVX1 _1190_ (
    .A(_498_),
    .Y(_499_)
);

AOI21X1 _1191_ (
    .A(_411_),
    .B(_496_),
    .C(_499_),
    .Y(_500_)
);

NAND2X1 _1192_ (
    .A(_477_),
    .B(_482_),
    .Y(_501_)
);

OAI21X1 _1193_ (
    .A(_469_),
    .B(_470_),
    .C(_468_),
    .Y(_502_)
);

INVX1 _1194_ (
    .A(_502_),
    .Y(_503_)
);

OR2X2 _1195_ (
    .A(_367_),
    .B(_427_),
    .Y(_504_)
);

NOR2X1 _1196_ (
    .A(_91_),
    .B(_418_),
    .Y(_505_)
);

OAI21X1 _1197_ (
    .A(_95_),
    .B(_239_),
    .C(_470_),
    .Y(_506_)
);

NAND2X1 _1198_ (
    .A(XinH[3]),
    .B(Cin[4]),
    .Y(_507_)
);

OAI21X1 _1199_ (
    .A(_465_),
    .B(_507_),
    .C(_506_),
    .Y(_508_)
);

XOR2X1 _1200_ (
    .A(_508_),
    .B(_505_),
    .Y(_509_)
);

AOI21X1 _1201_ (
    .A(_504_),
    .B(_476_),
    .C(_509_),
    .Y(_510_)
);

NAND3X1 _1202_ (
    .A(_504_),
    .B(_476_),
    .C(_509_),
    .Y(_511_)
);

INVX1 _1203_ (
    .A(_511_),
    .Y(_512_)
);

OAI21X1 _1204_ (
    .A(_510_),
    .B(_512_),
    .C(_503_),
    .Y(_513_)
);

INVX1 _1205_ (
    .A(_510_),
    .Y(_514_)
);

NAND3X1 _1206_ (
    .A(_502_),
    .B(_511_),
    .C(_514_),
    .Y(_515_)
);

AND2X2 _1207_ (
    .A(_513_),
    .B(_515_),
    .Y(_516_)
);

NAND2X1 _1208_ (
    .A(_501_),
    .B(_516_),
    .Y(_517_)
);

OR2X2 _1209_ (
    .A(_516_),
    .B(_501_),
    .Y(_518_)
);

NAND2X1 _1210_ (
    .A(_517_),
    .B(_518_),
    .Y(_519_)
);

NAND2X1 _1211_ (
    .A(_519_),
    .B(_500_),
    .Y(_520_)
);

AND2X2 _1212_ (
    .A(_399_),
    .B(_404_),
    .Y(_521_)
);

NAND3X1 _1213_ (
    .A(_282_),
    .B(_521_),
    .C(_336_),
    .Y(_522_)
);

NAND3X1 _1214_ (
    .A(_451_),
    .B(_455_),
    .C(_491_),
    .Y(_523_)
);

AOI21X1 _1215_ (
    .A(_522_),
    .B(_410_),
    .C(_523_),
    .Y(_524_)
);

INVX1 _1216_ (
    .A(_519_),
    .Y(_525_)
);

OAI21X1 _1217_ (
    .A(_499_),
    .B(_524_),
    .C(_525_),
    .Y(_526_)
);

NAND3X1 _1218_ (
    .A(LoadCtl_4_bF$buf4),
    .B(_520_),
    .C(_526_),
    .Y(_527_)
);

OAI21X1 _1219_ (
    .A(_494_),
    .B(LoadCtl_4_bF$buf3),
    .C(_527_),
    .Y(_30_)
);

NAND2X1 _1220_ (
    .A(mul[11]),
    .B(_135__bF$buf5),
    .Y(_528_)
);

AOI21X1 _1221_ (
    .A(_502_),
    .B(_511_),
    .C(_510_),
    .Y(_529_)
);

INVX1 _1222_ (
    .A(_505_),
    .Y(_530_)
);

OAI22X1 _1223_ (
    .A(_465_),
    .B(_507_),
    .C(_530_),
    .D(_508_),
    .Y(_531_)
);

OAI21X1 _1224_ (
    .A(_93_),
    .B(_418_),
    .C(_507_),
    .Y(_532_)
);

NOR2X1 _1225_ (
    .A(_95_),
    .B(_418_),
    .Y(_533_)
);

INVX1 _1226_ (
    .A(_533_),
    .Y(_534_)
);

OR2X2 _1227_ (
    .A(_534_),
    .B(_470_),
    .Y(_535_)
);

AND2X2 _1228_ (
    .A(_535_),
    .B(_532_),
    .Y(_536_)
);

XNOR2X1 _1229_ (
    .A(_536_),
    .B(_531_),
    .Y(_537_)
);

XOR2X1 _1230_ (
    .A(_537_),
    .B(_529_),
    .Y(_538_)
);

INVX1 _1231_ (
    .A(_538_),
    .Y(_539_)
);

NAND3X1 _1232_ (
    .A(_517_),
    .B(_539_),
    .C(_526_),
    .Y(_540_)
);

OAI21X1 _1233_ (
    .A(_519_),
    .B(_500_),
    .C(_517_),
    .Y(_541_)
);

NAND2X1 _1234_ (
    .A(_538_),
    .B(_541_),
    .Y(_542_)
);

NAND3X1 _1235_ (
    .A(LoadCtl_4_bF$buf2),
    .B(_542_),
    .C(_540_),
    .Y(_543_)
);

NAND2X1 _1236_ (
    .A(_528_),
    .B(_543_),
    .Y(_31_)
);

INVX1 _1237_ (
    .A(mul[12]),
    .Y(_544_)
);

NOR2X1 _1238_ (
    .A(_529_),
    .B(_537_),
    .Y(_545_)
);

AOI21X1 _1239_ (
    .A(_529_),
    .B(_537_),
    .C(_517_),
    .Y(_546_)
);

NOR2X1 _1240_ (
    .A(_545_),
    .B(_546_),
    .Y(_547_)
);

NAND3X1 _1241_ (
    .A(_517_),
    .B(_538_),
    .C(_518_),
    .Y(_548_)
);

OAI21X1 _1242_ (
    .A(_548_),
    .B(_500_),
    .C(_547_),
    .Y(_549_)
);

NAND2X1 _1243_ (
    .A(_531_),
    .B(_536_),
    .Y(_550_)
);

OAI21X1 _1244_ (
    .A(_93_),
    .B(_214_),
    .C(_533_),
    .Y(_551_)
);

OR2X2 _1245_ (
    .A(_550_),
    .B(_551_),
    .Y(_552_)
);

INVX1 _1246_ (
    .A(_535_),
    .Y(_553_)
);

OAI21X1 _1247_ (
    .A(_534_),
    .B(_553_),
    .C(_550_),
    .Y(_554_)
);

AND2X2 _1248_ (
    .A(_552_),
    .B(_554_),
    .Y(_555_)
);

NOR2X1 _1249_ (
    .A(_555_),
    .B(_549_),
    .Y(_556_)
);

INVX1 _1250_ (
    .A(_548_),
    .Y(_557_)
);

OAI21X1 _1251_ (
    .A(_498_),
    .B(_548_),
    .C(_547_),
    .Y(_558_)
);

AOI21X1 _1252_ (
    .A(_524_),
    .B(_557_),
    .C(_558_),
    .Y(_559_)
);

INVX1 _1253_ (
    .A(_555_),
    .Y(_560_)
);

OAI21X1 _1254_ (
    .A(_560_),
    .B(_559_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_561_)
);

OAI22X1 _1255_ (
    .A(_544_),
    .B(LoadCtl_4_bF$buf0),
    .C(_556_),
    .D(_561_),
    .Y(_32_)
);

INVX1 _1256_ (
    .A(mul[13]),
    .Y(_562_)
);

AOI21X1 _1257_ (
    .A(_549_),
    .B(_555_),
    .C(_553_),
    .Y(_563_)
);

AND2X2 _1258_ (
    .A(_552_),
    .B(LoadCtl_4_bF$buf6),
    .Y(_564_)
);

AOI22X1 _1259_ (
    .A(_562_),
    .B(_135__bF$buf4),
    .C(_563_),
    .D(_564_),
    .Y(_33_)
);

NOR2X1 _1260_ (
    .A(_101_),
    .B(_133_),
    .Y(_565_)
);

INVX1 _1261_ (
    .A(_565_),
    .Y(_566_)
);

NAND2X1 _1262_ (
    .A(_101_),
    .B(_133_),
    .Y(_567_)
);

NAND2X1 _1263_ (
    .A(_567_),
    .B(_566_),
    .Y(_568_)
);

NAND2X1 _1264_ (
    .A(y[0]),
    .B(_135__bF$buf3),
    .Y(_569_)
);

OAI21X1 _1265_ (
    .A(_135__bF$buf2),
    .B(_568_),
    .C(_569_),
    .Y(_34_)
);

INVX1 _1266_ (
    .A(mul[1]),
    .Y(_570_)
);

NOR2X1 _1267_ (
    .A(_103_),
    .B(_570_),
    .Y(_571_)
);

NOR2X1 _1268_ (
    .A(rYin[1]),
    .B(mul[1]),
    .Y(_572_)
);

NOR2X1 _1269_ (
    .A(_572_),
    .B(_571_),
    .Y(_573_)
);

NAND2X1 _1270_ (
    .A(_565_),
    .B(_573_),
    .Y(_574_)
);

OAI21X1 _1271_ (
    .A(_571_),
    .B(_572_),
    .C(_566_),
    .Y(_575_)
);

NAND2X1 _1272_ (
    .A(_575_),
    .B(_574_),
    .Y(_576_)
);

NAND2X1 _1273_ (
    .A(y[1]),
    .B(_135__bF$buf1),
    .Y(_577_)
);

OAI21X1 _1274_ (
    .A(_135__bF$buf0),
    .B(_576_),
    .C(_577_),
    .Y(_35_)
);

OAI21X1 _1275_ (
    .A(_103_),
    .B(_570_),
    .C(_574_),
    .Y(_578_)
);

XOR2X1 _1276_ (
    .A(rYin[2]),
    .B(mul[2]),
    .Y(_579_)
);

XNOR2X1 _1277_ (
    .A(_578_),
    .B(_579_),
    .Y(_580_)
);

NAND2X1 _1278_ (
    .A(y[2]),
    .B(_135__bF$buf5),
    .Y(_581_)
);

OAI21X1 _1279_ (
    .A(_135__bF$buf4),
    .B(_580_),
    .C(_581_),
    .Y(_36_)
);

NOR2X1 _1280_ (
    .A(_105_),
    .B(_159_),
    .Y(_582_)
);

AOI21X1 _1281_ (
    .A(_578_),
    .B(_579_),
    .C(_582_),
    .Y(_583_)
);

NOR2X1 _1282_ (
    .A(rYin[3]),
    .B(mul[3]),
    .Y(_584_)
);

NOR2X1 _1283_ (
    .A(_107_),
    .B(_161_),
    .Y(_585_)
);

NOR2X1 _1284_ (
    .A(_584_),
    .B(_585_),
    .Y(_586_)
);

XOR2X1 _1285_ (
    .A(_583_),
    .B(_586_),
    .Y(_587_)
);

NAND2X1 _1286_ (
    .A(y[3]),
    .B(_135__bF$buf3),
    .Y(_588_)
);

OAI21X1 _1287_ (
    .A(_135__bF$buf2),
    .B(_587_),
    .C(_588_),
    .Y(_37_)
);

NAND2X1 _1288_ (
    .A(y[4]),
    .B(_135__bF$buf1),
    .Y(_589_)
);

NAND2X1 _1289_ (
    .A(_109_),
    .B(_192_),
    .Y(_590_)
);

NAND2X1 _1290_ (
    .A(rYin[4]),
    .B(mul[4]),
    .Y(_591_)
);

AND2X2 _1291_ (
    .A(_590_),
    .B(_591_),
    .Y(_592_)
);

INVX1 _1292_ (
    .A(_592_),
    .Y(_593_)
);

INVX1 _1293_ (
    .A(_585_),
    .Y(_594_)
);

OAI21X1 _1294_ (
    .A(_584_),
    .B(_583_),
    .C(_594_),
    .Y(_595_)
);

INVX1 _1295_ (
    .A(_595_),
    .Y(_596_)
);

NAND2X1 _1296_ (
    .A(_593_),
    .B(_596_),
    .Y(_597_)
);

NAND2X1 _1297_ (
    .A(_592_),
    .B(_595_),
    .Y(_598_)
);

NAND2X1 _1298_ (
    .A(_598_),
    .B(_597_),
    .Y(_599_)
);

OAI21X1 _1299_ (
    .A(_135__bF$buf0),
    .B(_599_),
    .C(_589_),
    .Y(_38_)
);

NAND2X1 _1300_ (
    .A(y[5]),
    .B(_135__bF$buf5),
    .Y(_600_)
);

OAI21X1 _1301_ (
    .A(_109_),
    .B(_192_),
    .C(_598_),
    .Y(_601_)
);

OR2X2 _1302_ (
    .A(rYin[5]),
    .B(mul[5]),
    .Y(_602_)
);

NAND2X1 _1303_ (
    .A(rYin[5]),
    .B(mul[5]),
    .Y(_603_)
);

AND2X2 _1304_ (
    .A(_602_),
    .B(_603_),
    .Y(_604_)
);

NOR2X1 _1305_ (
    .A(_604_),
    .B(_601_),
    .Y(_605_)
);

INVX1 _1306_ (
    .A(_601_),
    .Y(_606_)
);

INVX1 _1307_ (
    .A(_604_),
    .Y(_607_)
);

OAI21X1 _1308_ (
    .A(_607_),
    .B(_606_),
    .C(LoadCtl_4_bF$buf5),
    .Y(_608_)
);

OAI21X1 _1309_ (
    .A(_605_),
    .B(_608_),
    .C(_600_),
    .Y(_39_)
);

NAND2X1 _1310_ (
    .A(y[6]),
    .B(_135__bF$buf4),
    .Y(_609_)
);

OAI21X1 _1311_ (
    .A(_607_),
    .B(_606_),
    .C(_603_),
    .Y(_610_)
);

XOR2X1 _1312_ (
    .A(rYin[6]),
    .B(mul[6]),
    .Y(_611_)
);

NOR2X1 _1313_ (
    .A(_611_),
    .B(_610_),
    .Y(_612_)
);

NAND2X1 _1314_ (
    .A(_611_),
    .B(_610_),
    .Y(_613_)
);

NAND2X1 _1315_ (
    .A(LoadCtl_4_bF$buf4),
    .B(_613_),
    .Y(_614_)
);

OAI21X1 _1316_ (
    .A(_612_),
    .B(_614_),
    .C(_609_),
    .Y(_40_)
);

OAI21X1 _1317_ (
    .A(_113_),
    .B(_281_),
    .C(_613_),
    .Y(_615_)
);

NOR2X1 _1318_ (
    .A(rYin[7]),
    .B(mul[7]),
    .Y(_616_)
);

NAND2X1 _1319_ (
    .A(rYin[7]),
    .B(mul[7]),
    .Y(_617_)
);

INVX1 _1320_ (
    .A(_617_),
    .Y(_618_)
);

NOR2X1 _1321_ (
    .A(_616_),
    .B(_618_),
    .Y(_619_)
);

XNOR2X1 _1322_ (
    .A(_615_),
    .B(_619_),
    .Y(_620_)
);

NAND2X1 _1323_ (
    .A(y[7]),
    .B(_135__bF$buf3),
    .Y(_621_)
);

OAI21X1 _1324_ (
    .A(_135__bF$buf2),
    .B(_620_),
    .C(_621_),
    .Y(_41_)
);

NAND2X1 _1325_ (
    .A(y[8]),
    .B(_135__bF$buf1),
    .Y(_622_)
);

OAI21X1 _1326_ (
    .A(_591_),
    .B(_607_),
    .C(_603_),
    .Y(_623_)
);

NAND2X1 _1327_ (
    .A(rYin[6]),
    .B(mul[6]),
    .Y(_624_)
);

OAI21X1 _1328_ (
    .A(_624_),
    .B(_616_),
    .C(_617_),
    .Y(_625_)
);

AND2X2 _1329_ (
    .A(_619_),
    .B(_611_),
    .Y(_626_)
);

AOI21X1 _1330_ (
    .A(_623_),
    .B(_626_),
    .C(_625_),
    .Y(_627_)
);

NOR2X1 _1331_ (
    .A(_607_),
    .B(_593_),
    .Y(_628_)
);

NAND3X1 _1332_ (
    .A(_628_),
    .B(_626_),
    .C(_595_),
    .Y(_629_)
);

NAND2X1 _1333_ (
    .A(_627_),
    .B(_629_),
    .Y(_630_)
);

OR2X2 _1334_ (
    .A(rYin[8]),
    .B(mul[8]),
    .Y(_631_)
);

NAND2X1 _1335_ (
    .A(rYin[8]),
    .B(mul[8]),
    .Y(_632_)
);

AND2X2 _1336_ (
    .A(_631_),
    .B(_632_),
    .Y(_633_)
);

NOR2X1 _1337_ (
    .A(_633_),
    .B(_630_),
    .Y(_634_)
);

INVX1 _1338_ (
    .A(_630_),
    .Y(_635_)
);

INVX1 _1339_ (
    .A(_633_),
    .Y(_636_)
);

OAI21X1 _1340_ (
    .A(_636_),
    .B(_635_),
    .C(LoadCtl_4_bF$buf3),
    .Y(_637_)
);

OAI21X1 _1341_ (
    .A(_634_),
    .B(_637_),
    .C(_622_),
    .Y(_42_)
);

OAI21X1 _1342_ (
    .A(_636_),
    .B(_635_),
    .C(_632_),
    .Y(_638_)
);

NOR2X1 _1343_ (
    .A(rYin[9]),
    .B(mul[9]),
    .Y(_639_)
);

NAND2X1 _1344_ (
    .A(rYin[9]),
    .B(mul[9]),
    .Y(_640_)
);

INVX1 _1345_ (
    .A(_640_),
    .Y(_641_)
);

NOR2X1 _1346_ (
    .A(_639_),
    .B(_641_),
    .Y(_642_)
);

INVX1 _1347_ (
    .A(_642_),
    .Y(_643_)
);

XOR2X1 _1348_ (
    .A(_638_),
    .B(_643_),
    .Y(_644_)
);

NAND2X1 _1349_ (
    .A(y[9]),
    .B(_135__bF$buf0),
    .Y(_645_)
);

OAI21X1 _1350_ (
    .A(_135__bF$buf5),
    .B(_644_),
    .C(_645_),
    .Y(_43_)
);

NAND2X1 _1351_ (
    .A(y[10]),
    .B(_135__bF$buf4),
    .Y(_646_)
);

NOR2X1 _1352_ (
    .A(_643_),
    .B(_636_),
    .Y(_647_)
);

OAI21X1 _1353_ (
    .A(_632_),
    .B(_639_),
    .C(_640_),
    .Y(_648_)
);

AOI21X1 _1354_ (
    .A(_630_),
    .B(_647_),
    .C(_648_),
    .Y(_649_)
);

NOR2X1 _1355_ (
    .A(rYin[10]),
    .B(mul[10]),
    .Y(_650_)
);

NOR2X1 _1356_ (
    .A(_121_),
    .B(_494_),
    .Y(_651_)
);

NOR2X1 _1357_ (
    .A(_650_),
    .B(_651_),
    .Y(_652_)
);

INVX1 _1358_ (
    .A(_652_),
    .Y(_653_)
);

AND2X2 _1359_ (
    .A(_649_),
    .B(_653_),
    .Y(_654_)
);

OAI21X1 _1360_ (
    .A(_653_),
    .B(_649_),
    .C(LoadCtl_4_bF$buf2),
    .Y(_655_)
);

OAI21X1 _1361_ (
    .A(_655_),
    .B(_654_),
    .C(_646_),
    .Y(_44_)
);

NOR2X1 _1362_ (
    .A(_653_),
    .B(_649_),
    .Y(_656_)
);

NOR2X1 _1363_ (
    .A(_651_),
    .B(_656_),
    .Y(_657_)
);

NOR2X1 _1364_ (
    .A(rYin[11]),
    .B(mul[11]),
    .Y(_658_)
);

NAND2X1 _1365_ (
    .A(rYin[11]),
    .B(mul[11]),
    .Y(_659_)
);

INVX1 _1366_ (
    .A(_659_),
    .Y(_660_)
);

NOR2X1 _1367_ (
    .A(_658_),
    .B(_660_),
    .Y(_661_)
);

XOR2X1 _1368_ (
    .A(_657_),
    .B(_661_),
    .Y(_662_)
);

NAND2X1 _1369_ (
    .A(y[11]),
    .B(_135__bF$buf3),
    .Y(_663_)
);

OAI21X1 _1370_ (
    .A(_135__bF$buf2),
    .B(_662_),
    .C(_663_),
    .Y(_45_)
);

NAND2X1 _1371_ (
    .A(y[12]),
    .B(_135__bF$buf1),
    .Y(_664_)
);

AOI21X1 _1372_ (
    .A(_661_),
    .B(_651_),
    .C(_660_),
    .Y(_665_)
);

NAND2X1 _1373_ (
    .A(_661_),
    .B(_652_),
    .Y(_666_)
);

OAI21X1 _1374_ (
    .A(_666_),
    .B(_649_),
    .C(_665_),
    .Y(_667_)
);

NAND2X1 _1375_ (
    .A(_125_),
    .B(_544_),
    .Y(_668_)
);

NOR2X1 _1376_ (
    .A(_125_),
    .B(_544_),
    .Y(_669_)
);

INVX1 _1377_ (
    .A(_669_),
    .Y(_670_)
);

AND2X2 _1378_ (
    .A(_670_),
    .B(_668_),
    .Y(_671_)
);

NOR2X1 _1379_ (
    .A(_671_),
    .B(_667_),
    .Y(_672_)
);

INVX1 _1380_ (
    .A(_667_),
    .Y(_673_)
);

INVX1 _1381_ (
    .A(_671_),
    .Y(_674_)
);

OAI21X1 _1382_ (
    .A(_674_),
    .B(_673_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_675_)
);

OAI21X1 _1383_ (
    .A(_672_),
    .B(_675_),
    .C(_664_),
    .Y(_46_)
);

OAI21X1 _1384_ (
    .A(_674_),
    .B(_673_),
    .C(_670_),
    .Y(_676_)
);

NOR2X1 _1385_ (
    .A(rYin[13]),
    .B(mul[13]),
    .Y(_677_)
);

NOR2X1 _1386_ (
    .A(_127_),
    .B(_562_),
    .Y(_678_)
);

NOR2X1 _1387_ (
    .A(_677_),
    .B(_678_),
    .Y(_679_)
);

INVX1 _1388_ (
    .A(_679_),
    .Y(_680_)
);

OR2X2 _1389_ (
    .A(_676_),
    .B(_680_),
    .Y(_681_)
);

AOI21X1 _1390_ (
    .A(_676_),
    .B(_680_),
    .C(_135__bF$buf0),
    .Y(_682_)
);

AOI22X1 _1391_ (
    .A(_78_),
    .B(_135__bF$buf5),
    .C(_681_),
    .D(_682_),
    .Y(_47_)
);

AOI21X1 _1392_ (
    .A(_679_),
    .B(_669_),
    .C(_678_),
    .Y(_683_)
);

INVX1 _1393_ (
    .A(_683_),
    .Y(_684_)
);

NOR2X1 _1394_ (
    .A(_680_),
    .B(_674_),
    .Y(_685_)
);

AOI21X1 _1395_ (
    .A(_667_),
    .B(_685_),
    .C(_684_),
    .Y(_686_)
);

INVX1 _1396_ (
    .A(_686_),
    .Y(_687_)
);

NOR2X1 _1397_ (
    .A(rYin[14]),
    .B(_687_),
    .Y(_688_)
);

OAI21X1 _1398_ (
    .A(_129_),
    .B(_686_),
    .C(LoadCtl_4_bF$buf0),
    .Y(_689_)
);

OAI22X1 _1399_ (
    .A(_82_),
    .B(LoadCtl_4_bF$buf6),
    .C(_689_),
    .D(_688_),
    .Y(_48_)
);

NAND2X1 _1400_ (
    .A(y[15]),
    .B(_135__bF$buf4),
    .Y(_690_)
);

NAND3X1 _1401_ (
    .A(rYin[14]),
    .B(rYin[15]),
    .C(_687_),
    .Y(_691_)
);

OAI21X1 _1402_ (
    .A(_129_),
    .B(_686_),
    .C(_131_),
    .Y(_692_)
);

NAND2X1 _1403_ (
    .A(_692_),
    .B(_691_),
    .Y(_693_)
);

OAI21X1 _1404_ (
    .A(_135__bF$buf3),
    .B(_693_),
    .C(_690_),
    .Y(_49_)
);

INVX1 _1405_ (
    .A(Yin[0]),
    .Y(_694_)
);

NAND3X1 _1406_ (
    .A(LoadCtl[3]),
    .B(_71_),
    .C(_72_),
    .Y(_695_)
);

NAND2X1 _1407_ (
    .A(Yin3[0]),
    .B(_695_),
    .Y(_696_)
);

OAI21X1 _1408_ (
    .A(_694_),
    .B(_695_),
    .C(_696_),
    .Y(_50_)
);

INVX1 _1409_ (
    .A(Yin[1]),
    .Y(_697_)
);

NAND2X1 _1410_ (
    .A(Yin3[1]),
    .B(_695_),
    .Y(_698_)
);

OAI21X1 _1411_ (
    .A(_697_),
    .B(_695_),
    .C(_698_),
    .Y(_51_)
);

INVX1 _1412_ (
    .A(Yin[2]),
    .Y(_699_)
);

NAND2X1 _1413_ (
    .A(Yin3[2]),
    .B(_695_),
    .Y(_700_)
);

OAI21X1 _1414_ (
    .A(_699_),
    .B(_695_),
    .C(_700_),
    .Y(_52_)
);

INVX1 _1415_ (
    .A(Yin[3]),
    .Y(_701_)
);

NAND2X1 _1416_ (
    .A(Yin3[3]),
    .B(_695_),
    .Y(_702_)
);

OAI21X1 _1417_ (
    .A(_701_),
    .B(_695_),
    .C(_702_),
    .Y(_53_)
);

NOR2X1 _1418_ (
    .A(_71_),
    .B(_77_),
    .Y(_703_)
);

NOR2X1 _1419_ (
    .A(Yin2[0]),
    .B(_703_),
    .Y(_704_)
);

AOI21X1 _1420_ (
    .A(_694_),
    .B(_703_),
    .C(_704_),
    .Y(_54_)
);

NOR2X1 _1421_ (
    .A(Yin2[1]),
    .B(_703_),
    .Y(_705_)
);

AOI21X1 _1422_ (
    .A(_697_),
    .B(_703_),
    .C(_705_),
    .Y(_55_)
);

NOR2X1 _1423_ (
    .A(Yin2[2]),
    .B(_703_),
    .Y(_706_)
);

AOI21X1 _1424_ (
    .A(_699_),
    .B(_703_),
    .C(_706_),
    .Y(_56_)
);

NOR2X1 _1425_ (
    .A(Yin2[3]),
    .B(_703_),
    .Y(_707_)
);

AOI21X1 _1426_ (
    .A(_701_),
    .B(_703_),
    .C(_707_),
    .Y(_57_)
);

INVX1 _1427_ (
    .A(_75_),
    .Y(_708_)
);

OAI21X1 _1428_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_74_),
    .C(Yin1[0]),
    .Y(_709_)
);

OAI21X1 _1429_ (
    .A(_694_),
    .B(_708_),
    .C(_709_),
    .Y(_58_)
);

OAI21X1 _1430_ (
    .A(LoadCtl_0_bF$buf3),
    .B(_74_),
    .C(Yin1[1]),
    .Y(_710_)
);

OAI21X1 _1431_ (
    .A(_697_),
    .B(_708_),
    .C(_710_),
    .Y(_59_)
);

OAI21X1 _1432_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_74_),
    .C(Yin1[2]),
    .Y(_711_)
);

OAI21X1 _1433_ (
    .A(_699_),
    .B(_708_),
    .C(_711_),
    .Y(_60_)
);

OAI21X1 _1434_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_74_),
    .C(Yin1[3]),
    .Y(_712_)
);

OAI21X1 _1435_ (
    .A(_701_),
    .B(_708_),
    .C(_712_),
    .Y(_61_)
);

NOR2X1 _1436_ (
    .A(LoadCtl_0_bF$buf0),
    .B(Yin0[0]),
    .Y(_713_)
);

AOI21X1 _1437_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_694_),
    .C(_713_),
    .Y(_62_)
);

NOR2X1 _1438_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Yin0[1]),
    .Y(_714_)
);

AOI21X1 _1439_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_697_),
    .C(_714_),
    .Y(_63_)
);

NOR2X1 _1440_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Yin0[2]),
    .Y(_715_)
);

AOI21X1 _1441_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_699_),
    .C(_715_),
    .Y(_64_)
);

NOR2X1 _1442_ (
    .A(LoadCtl_0_bF$buf4),
    .B(Yin0[3]),
    .Y(_716_)
);

AOI21X1 _1443_ (
    .A(LoadCtl_0_bF$buf3),
    .B(_701_),
    .C(_716_),
    .Y(_65_)
);

NAND2X1 _1444_ (
    .A(LoadCtl_0_bF$buf2),
    .B(Xin[0]),
    .Y(_717_)
);

OAI21X1 _1445_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_213_),
    .C(_717_),
    .Y(_66_)
);

NAND2X1 _1446_ (
    .A(LoadCtl_0_bF$buf0),
    .B(Xin[1]),
    .Y(_718_)
);

OAI21X1 _1447_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_150_),
    .C(_718_),
    .Y(_67_)
);

NAND2X1 _1448_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Xin[2]),
    .Y(_719_)
);

OAI21X1 _1449_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_177_),
    .C(_719_),
    .Y(_68_)
);

NAND2X1 _1450_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Xin[3]),
    .Y(_720_)
);

OAI21X1 _1451_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_179_),
    .C(_720_),
    .Y(_69_)
);

DFFPOSX1 _1452_ (
    .CLK(clk_bF$buf7),
    .D(_0_),
    .Q(XinH[0])
);

DFFPOSX1 _1453_ (
    .CLK(clk_bF$buf6),
    .D(_1_),
    .Q(XinH[1])
);

DFFPOSX1 _1454_ (
    .CLK(clk_bF$buf5),
    .D(_2_),
    .Q(XinH[2])
);

DFFPOSX1 _1455_ (
    .CLK(clk_bF$buf4),
    .D(_3_),
    .Q(XinH[3])
);

DFFPOSX1 _1456_ (
    .CLK(clk_bF$buf3),
    .D(_4_),
    .Q(rYin[0])
);

DFFPOSX1 _1457_ (
    .CLK(clk_bF$buf2),
    .D(_5_),
    .Q(rYin[1])
);

DFFPOSX1 _1458_ (
    .CLK(clk_bF$buf1),
    .D(_6_),
    .Q(rYin[2])
);

DFFPOSX1 _1459_ (
    .CLK(clk_bF$buf0),
    .D(_7_),
    .Q(rYin[3])
);

DFFPOSX1 _1460_ (
    .CLK(clk_bF$buf7),
    .D(_8_),
    .Q(rYin[4])
);

DFFPOSX1 _1461_ (
    .CLK(clk_bF$buf6),
    .D(_9_),
    .Q(rYin[5])
);

DFFPOSX1 _1462_ (
    .CLK(clk_bF$buf5),
    .D(_10_),
    .Q(rYin[6])
);

DFFPOSX1 _1463_ (
    .CLK(clk_bF$buf4),
    .D(_11_),
    .Q(rYin[7])
);

DFFPOSX1 _1464_ (
    .CLK(clk_bF$buf3),
    .D(_12_),
    .Q(rYin[8])
);

DFFPOSX1 _1465_ (
    .CLK(clk_bF$buf2),
    .D(_13_),
    .Q(rYin[9])
);

DFFPOSX1 _1466_ (
    .CLK(clk_bF$buf1),
    .D(_14_),
    .Q(rYin[10])
);

DFFPOSX1 _1467_ (
    .CLK(clk_bF$buf0),
    .D(_15_),
    .Q(rYin[11])
);

DFFPOSX1 _1468_ (
    .CLK(clk_bF$buf7),
    .D(_16_),
    .Q(rYin[12])
);

DFFPOSX1 _1469_ (
    .CLK(clk_bF$buf6),
    .D(_17_),
    .Q(rYin[13])
);

DFFPOSX1 _1470_ (
    .CLK(clk_bF$buf5),
    .D(_18_),
    .Q(rYin[14])
);

DFFPOSX1 _1471_ (
    .CLK(clk_bF$buf4),
    .D(_19_),
    .Q(rYin[15])
);

DFFPOSX1 _1472_ (
    .CLK(clk_bF$buf3),
    .D(_20_),
    .Q(mul[0])
);

DFFPOSX1 _1473_ (
    .CLK(clk_bF$buf2),
    .D(_21_),
    .Q(mul[1])
);

DFFPOSX1 _1474_ (
    .CLK(clk_bF$buf1),
    .D(_22_),
    .Q(mul[2])
);

DFFPOSX1 _1475_ (
    .CLK(clk_bF$buf0),
    .D(_23_),
    .Q(mul[3])
);

DFFPOSX1 _1476_ (
    .CLK(clk_bF$buf7),
    .D(_24_),
    .Q(mul[4])
);

DFFPOSX1 _1477_ (
    .CLK(clk_bF$buf6),
    .D(_25_),
    .Q(mul[5])
);

DFFPOSX1 _1478_ (
    .CLK(clk_bF$buf5),
    .D(_26_),
    .Q(mul[6])
);

DFFPOSX1 _1479_ (
    .CLK(clk_bF$buf4),
    .D(_27_),
    .Q(mul[7])
);

DFFPOSX1 _1480_ (
    .CLK(clk_bF$buf3),
    .D(_28_),
    .Q(mul[8])
);

DFFPOSX1 _1481_ (
    .CLK(clk_bF$buf2),
    .D(_29_),
    .Q(mul[9])
);

DFFPOSX1 _1482_ (
    .CLK(clk_bF$buf1),
    .D(_30_),
    .Q(mul[10])
);

DFFPOSX1 _1483_ (
    .CLK(clk_bF$buf0),
    .D(_31_),
    .Q(mul[11])
);

DFFPOSX1 _1484_ (
    .CLK(clk_bF$buf7),
    .D(_32_),
    .Q(mul[12])
);

DFFPOSX1 _1485_ (
    .CLK(clk_bF$buf6),
    .D(_33_),
    .Q(mul[13])
);

DFFPOSX1 _1486_ (
    .CLK(clk_bF$buf5),
    .D(_34_),
    .Q(y[0])
);

DFFPOSX1 _1487_ (
    .CLK(clk_bF$buf4),
    .D(_35_),
    .Q(y[1])
);

DFFPOSX1 _1488_ (
    .CLK(clk_bF$buf3),
    .D(_36_),
    .Q(y[2])
);

DFFPOSX1 _1489_ (
    .CLK(clk_bF$buf2),
    .D(_37_),
    .Q(y[3])
);

DFFPOSX1 _1490_ (
    .CLK(clk_bF$buf1),
    .D(_38_),
    .Q(y[4])
);

DFFPOSX1 _1491_ (
    .CLK(clk_bF$buf0),
    .D(_39_),
    .Q(y[5])
);

DFFPOSX1 _1492_ (
    .CLK(clk_bF$buf7),
    .D(_40_),
    .Q(y[6])
);

DFFPOSX1 _1493_ (
    .CLK(clk_bF$buf6),
    .D(_41_),
    .Q(y[7])
);

DFFPOSX1 _1494_ (
    .CLK(clk_bF$buf5),
    .D(_42_),
    .Q(y[8])
);

DFFPOSX1 _1495_ (
    .CLK(clk_bF$buf4),
    .D(_43_),
    .Q(y[9])
);

DFFPOSX1 _1496_ (
    .CLK(clk_bF$buf3),
    .D(_44_),
    .Q(y[10])
);

DFFPOSX1 _1497_ (
    .CLK(clk_bF$buf2),
    .D(_45_),
    .Q(y[11])
);

DFFPOSX1 _1498_ (
    .CLK(clk_bF$buf1),
    .D(_46_),
    .Q(y[12])
);

DFFPOSX1 _1499_ (
    .CLK(clk_bF$buf0),
    .D(_47_),
    .Q(y[13])
);

DFFPOSX1 _1500_ (
    .CLK(clk_bF$buf7),
    .D(_48_),
    .Q(y[14])
);

DFFPOSX1 _1501_ (
    .CLK(clk_bF$buf6),
    .D(_49_),
    .Q(y[15])
);

DFFPOSX1 _1502_ (
    .CLK(clk_bF$buf5),
    .D(_50_),
    .Q(Yin3[0])
);

DFFPOSX1 _1503_ (
    .CLK(clk_bF$buf4),
    .D(_51_),
    .Q(Yin3[1])
);

DFFPOSX1 _1504_ (
    .CLK(clk_bF$buf3),
    .D(_52_),
    .Q(Yin3[2])
);

DFFPOSX1 _1505_ (
    .CLK(clk_bF$buf2),
    .D(_53_),
    .Q(Yin3[3])
);

DFFPOSX1 _1506_ (
    .CLK(clk_bF$buf1),
    .D(_54_),
    .Q(Yin2[0])
);

DFFPOSX1 _1507_ (
    .CLK(clk_bF$buf0),
    .D(_55_),
    .Q(Yin2[1])
);

DFFPOSX1 _1508_ (
    .CLK(clk_bF$buf7),
    .D(_56_),
    .Q(Yin2[2])
);

DFFPOSX1 _1509_ (
    .CLK(clk_bF$buf6),
    .D(_57_),
    .Q(Yin2[3])
);

DFFPOSX1 _1510_ (
    .CLK(clk_bF$buf5),
    .D(_58_),
    .Q(Yin1[0])
);

DFFPOSX1 _1511_ (
    .CLK(clk_bF$buf4),
    .D(_59_),
    .Q(Yin1[1])
);

DFFPOSX1 _1512_ (
    .CLK(clk_bF$buf3),
    .D(_60_),
    .Q(Yin1[2])
);

DFFPOSX1 _1513_ (
    .CLK(clk_bF$buf2),
    .D(_61_),
    .Q(Yin1[3])
);

DFFPOSX1 _1514_ (
    .CLK(clk_bF$buf1),
    .D(_62_),
    .Q(Yin0[0])
);

DFFPOSX1 _1515_ (
    .CLK(clk_bF$buf0),
    .D(_63_),
    .Q(Yin0[1])
);

DFFPOSX1 _1516_ (
    .CLK(clk_bF$buf7),
    .D(_64_),
    .Q(Yin0[2])
);

DFFPOSX1 _1517_ (
    .CLK(clk_bF$buf6),
    .D(_65_),
    .Q(Yin0[3])
);

DFFPOSX1 _1518_ (
    .CLK(clk_bF$buf5),
    .D(_66_),
    .Q(XinHL[0])
);

DFFPOSX1 _1519_ (
    .CLK(clk_bF$buf4),
    .D(_67_),
    .Q(XinHL[1])
);

DFFPOSX1 _1520_ (
    .CLK(clk_bF$buf3),
    .D(_68_),
    .Q(XinHL[2])
);

DFFPOSX1 _1521_ (
    .CLK(clk_bF$buf2),
    .D(_69_),
    .Q(XinHL[3])
);

DFFPOSX1 _1522_ (
    .CLK(clk_bF$buf1),
    .D(Rdy),
    .Q(LoadCtl[0])
);

DFFPOSX1 _1523_ (
    .CLK(clk_bF$buf0),
    .D(LoadCtl_0_bF$buf4),
    .Q(LoadCtl[1])
);

DFFPOSX1 _1524_ (
    .CLK(clk_bF$buf7),
    .D(LoadCtl[1]),
    .Q(LoadCtl[2])
);

DFFPOSX1 _1525_ (
    .CLK(clk_bF$buf6),
    .D(LoadCtl[2]),
    .Q(LoadCtl[3])
);

DFFPOSX1 _1526_ (
    .CLK(clk_bF$buf5),
    .D(LoadCtl[3]),
    .Q(LoadCtl[4])
);

BUFX2 _1527_ (
    .A(LoadCtl_4_bF$buf5),
    .Y(Vld)
);

BUFX2 _1528_ (
    .A(_721_[0]),
    .Y(Xout[0])
);

BUFX2 _1529_ (
    .A(_721_[1]),
    .Y(Xout[1])
);

BUFX2 _1530_ (
    .A(_721_[2]),
    .Y(Xout[2])
);

BUFX2 _1531_ (
    .A(_721_[3]),
    .Y(Xout[3])
);

BUFX2 _1532_ (
    .A(_722_[0]),
    .Y(Yout[0])
);

BUFX2 _1533_ (
    .A(_722_[1]),
    .Y(Yout[1])
);

BUFX2 _1534_ (
    .A(_722_[2]),
    .Y(Yout[2])
);

BUFX2 _1535_ (
    .A(_722_[3]),
    .Y(Yout[3])
);

NOR2X1 _723_ (
    .A(LoadCtl[2]),
    .B(y[12]),
    .Y(_70_)
);

INVX2 _724_ (
    .A(LoadCtl[2]),
    .Y(_71_)
);

NOR2X1 _725_ (
    .A(LoadCtl[1]),
    .B(LoadCtl_0_bF$buf3),
    .Y(_72_)
);

OAI21X1 _726_ (
    .A(_71_),
    .B(y[8]),
    .C(_72_),
    .Y(_73_)
);

INVX2 _727_ (
    .A(LoadCtl[1]),
    .Y(_74_)
);

NOR2X1 _728_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_74_),
    .Y(_75_)
);

AOI22X1 _729_ (
    .A(LoadCtl_0_bF$buf1),
    .B(y[0]),
    .C(_75_),
    .D(y[4]),
    .Y(_76_)
);

OAI21X1 _730_ (
    .A(_70_),
    .B(_73_),
    .C(_76_),
    .Y(_722_[0])
);

INVX1 _731_ (
    .A(_72_),
    .Y(_77_)
);

INVX1 _732_ (
    .A(y[13]),
    .Y(_78_)
);

NAND2X1 _733_ (
    .A(_71_),
    .B(_78_),
    .Y(_79_)
);

OAI21X1 _734_ (
    .A(_71_),
    .B(y[9]),
    .C(_79_),
    .Y(_80_)
);

AOI22X1 _735_ (
    .A(LoadCtl_0_bF$buf0),
    .B(y[1]),
    .C(_75_),
    .D(y[5]),
    .Y(_81_)
);

OAI21X1 _736_ (
    .A(_77_),
    .B(_80_),
    .C(_81_),
    .Y(_722_[1])
);

INVX1 _737_ (
    .A(y[14]),
    .Y(_82_)
);

NAND2X1 _738_ (
    .A(_71_),
    .B(_82_),
    .Y(_83_)
);

OAI21X1 _739_ (
    .A(_71_),
    .B(y[10]),
    .C(_83_),
    .Y(_84_)
);

AOI22X1 _740_ (
    .A(LoadCtl_0_bF$buf4),
    .B(y[2]),
    .C(_75_),
    .D(y[6]),
    .Y(_85_)
);

OAI21X1 _741_ (
    .A(_77_),
    .B(_84_),
    .C(_85_),
    .Y(_722_[2])
);

NOR2X1 _742_ (
    .A(LoadCtl[2]),
    .B(y[15]),
    .Y(_86_)
);

OAI21X1 _743_ (
    .A(_71_),
    .B(y[11]),
    .C(_72_),
    .Y(_87_)
);

AOI22X1 _744_ (
    .A(LoadCtl_0_bF$buf3),
    .B(y[3]),
    .C(_75_),
    .D(y[7]),
    .Y(_88_)
);

OAI21X1 _745_ (
    .A(_86_),
    .B(_87_),
    .C(_88_),
    .Y(_722_[3])
);

INVX2 _746_ (
    .A(XinH[0]),
    .Y(_89_)
);

NAND2X1 _747_ (
    .A(LoadCtl_0_bF$buf2),
    .B(XinHL[0]),
    .Y(_90_)
);

OAI21X1 _748_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_89_),
    .C(_90_),
    .Y(_721_[0])
);

INVX1 _749_ (
    .A(XinH[1]),
    .Y(_91_)
);

NAND2X1 _750_ (
    .A(LoadCtl_0_bF$buf0),
    .B(XinHL[1]),
    .Y(_92_)
);

OAI21X1 _751_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_91_),
    .C(_92_),
    .Y(_721_[1])
);

INVX2 _752_ (
    .A(XinH[2]),
    .Y(_93_)
);

NAND2X1 _753_ (
    .A(LoadCtl_0_bF$buf3),
    .B(XinHL[2]),
    .Y(_94_)
);

OAI21X1 _754_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_93_),
    .C(_94_),
    .Y(_721_[2])
);

INVX2 _755_ (
    .A(XinH[3]),
    .Y(_95_)
);

NAND2X1 _756_ (
    .A(LoadCtl_0_bF$buf1),
    .B(XinHL[3]),
    .Y(_96_)
);

OAI21X1 _757_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_95_),
    .C(_96_),
    .Y(_721_[3])
);

NAND2X1 _758_ (
    .A(Xin[0]),
    .B(_75_),
    .Y(_97_)
);

OAI21X1 _759_ (
    .A(_89_),
    .B(_75_),
    .C(_97_),
    .Y(_0_)
);

NAND2X1 _760_ (
    .A(Xin[1]),
    .B(_75_),
    .Y(_98_)
);

OAI21X1 _761_ (
    .A(_91_),
    .B(_75_),
    .C(_98_),
    .Y(_1_)
);

NAND2X1 _762_ (
    .A(Xin[2]),
    .B(_75_),
    .Y(_99_)
);

OAI21X1 _763_ (
    .A(_93_),
    .B(_75_),
    .C(_99_),
    .Y(_2_)
);

NAND2X1 _764_ (
    .A(Xin[3]),
    .B(_75_),
    .Y(_100_)
);

OAI21X1 _765_ (
    .A(_95_),
    .B(_75_),
    .C(_100_),
    .Y(_3_)
);

INVX1 _766_ (
    .A(rYin[0]),
    .Y(_101_)
);

NAND2X1 _767_ (
    .A(Yin0[0]),
    .B(LoadCtl_4_bF$buf4),
    .Y(_102_)
);

OAI21X1 _768_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_101_),
    .C(_102_),
    .Y(_4_)
);

INVX1 _769_ (
    .A(rYin[1]),
    .Y(_103_)
);

NAND2X1 _770_ (
    .A(LoadCtl_4_bF$buf2),
    .B(Yin0[1]),
    .Y(_104_)
);

OAI21X1 _771_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_103_),
    .C(_104_),
    .Y(_5_)
);

INVX1 _772_ (
    .A(rYin[2]),
    .Y(_105_)
);

NAND2X1 _773_ (
    .A(LoadCtl_4_bF$buf0),
    .B(Yin0[2]),
    .Y(_106_)
);

OAI21X1 _774_ (
    .A(LoadCtl_4_bF$buf6),
    .B(_105_),
    .C(_106_),
    .Y(_6_)
);

INVX1 _775_ (
    .A(rYin[3]),
    .Y(_107_)
);

NAND2X1 _776_ (
    .A(LoadCtl_4_bF$buf5),
    .B(Yin0[3]),
    .Y(_108_)
);

OAI21X1 _777_ (
    .A(LoadCtl_4_bF$buf4),
    .B(_107_),
    .C(_108_),
    .Y(_7_)
);

INVX1 _778_ (
    .A(rYin[4]),
    .Y(_109_)
);

NAND2X1 _779_ (
    .A(LoadCtl_4_bF$buf3),
    .B(Yin1[0]),
    .Y(_110_)
);

OAI21X1 _780_ (
    .A(LoadCtl_4_bF$buf2),
    .B(_109_),
    .C(_110_),
    .Y(_8_)
);

INVX1 _781_ (
    .A(rYin[5]),
    .Y(_111_)
);

NAND2X1 _782_ (
    .A(LoadCtl_4_bF$buf1),
    .B(Yin1[1]),
    .Y(_112_)
);

OAI21X1 _783_ (
    .A(LoadCtl_4_bF$buf0),
    .B(_111_),
    .C(_112_),
    .Y(_9_)
);

INVX1 _784_ (
    .A(rYin[6]),
    .Y(_113_)
);

NAND2X1 _785_ (
    .A(LoadCtl_4_bF$buf6),
    .B(Yin1[2]),
    .Y(_114_)
);

OAI21X1 _786_ (
    .A(LoadCtl_4_bF$buf5),
    .B(_113_),
    .C(_114_),
    .Y(_10_)
);

INVX1 _787_ (
    .A(rYin[7]),
    .Y(_115_)
);

NAND2X1 _788_ (
    .A(LoadCtl_4_bF$buf4),
    .B(Yin1[3]),
    .Y(_116_)
);

OAI21X1 _789_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_115_),
    .C(_116_),
    .Y(_11_)
);

INVX1 _790_ (
    .A(rYin[8]),
    .Y(_117_)
);

NAND2X1 _791_ (
    .A(LoadCtl_4_bF$buf2),
    .B(Yin2[0]),
    .Y(_118_)
);

OAI21X1 _792_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_117_),
    .C(_118_),
    .Y(_12_)
);

INVX1 _793_ (
    .A(rYin[9]),
    .Y(_119_)
);

NAND2X1 _794_ (
    .A(LoadCtl_4_bF$buf0),
    .B(Yin2[1]),
    .Y(_120_)
);

OAI21X1 _795_ (
    .A(LoadCtl_4_bF$buf6),
    .B(_119_),
    .C(_120_),
    .Y(_13_)
);

INVX1 _796_ (
    .A(rYin[10]),
    .Y(_121_)
);

NAND2X1 _797_ (
    .A(LoadCtl_4_bF$buf5),
    .B(Yin2[2]),
    .Y(_122_)
);

OAI21X1 _798_ (
    .A(LoadCtl_4_bF$buf4),
    .B(_121_),
    .C(_122_),
    .Y(_14_)
);

INVX1 _799_ (
    .A(rYin[11]),
    .Y(_123_)
);

NAND2X1 _800_ (
    .A(LoadCtl_4_bF$buf3),
    .B(Yin2[3]),
    .Y(_124_)
);

OAI21X1 _801_ (
    .A(LoadCtl_4_bF$buf2),
    .B(_123_),
    .C(_124_),
    .Y(_15_)
);

INVX1 _802_ (
    .A(rYin[12]),
    .Y(_125_)
);

NAND2X1 _803_ (
    .A(LoadCtl_4_bF$buf1),
    .B(Yin3[0]),
    .Y(_126_)
);

OAI21X1 _804_ (
    .A(LoadCtl_4_bF$buf0),
    .B(_125_),
    .C(_126_),
    .Y(_16_)
);

INVX1 _805_ (
    .A(rYin[13]),
    .Y(_127_)
);

NAND2X1 _806_ (
    .A(LoadCtl_4_bF$buf6),
    .B(Yin3[1]),
    .Y(_128_)
);

OAI21X1 _807_ (
    .A(LoadCtl_4_bF$buf5),
    .B(_127_),
    .C(_128_),
    .Y(_17_)
);

INVX1 _808_ (
    .A(rYin[14]),
    .Y(_129_)
);

NAND2X1 _809_ (
    .A(LoadCtl_4_bF$buf4),
    .B(Yin3[2]),
    .Y(_130_)
);

OAI21X1 _810_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_129_),
    .C(_130_),
    .Y(_18_)
);

INVX1 _811_ (
    .A(rYin[15]),
    .Y(_131_)
);

NAND2X1 _812_ (
    .A(LoadCtl_4_bF$buf2),
    .B(Yin3[3]),
    .Y(_132_)
);

OAI21X1 _813_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_131_),
    .C(_132_),
    .Y(_19_)
);

INVX1 _814_ (
    .A(mul[0]),
    .Y(_133_)
);

NAND3X1 _815_ (
    .A(XinHL[0]),
    .B(Cin_0_bF$buf3),
    .C(LoadCtl_4_bF$buf0),
    .Y(_134_)
);

OAI21X1 _816_ (
    .A(_133_),
    .B(LoadCtl_4_bF$buf6),
    .C(_134_),
    .Y(_20_)
);

INVX8 _817_ (
    .A(LoadCtl_4_bF$buf5),
    .Y(_135_)
);

NAND2X1 _818_ (
    .A(XinHL[0]),
    .B(Cin_1_bF$buf2),
    .Y(_136_)
);

NAND2X1 _819_ (
    .A(XinHL[1]),
    .B(Cin_0_bF$buf2),
    .Y(_137_)
);

XNOR2X1 _820_ (
    .A(_136_),
    .B(_137_),
    .Y(_138_)
);

NAND2X1 _821_ (
    .A(mul[1]),
    .B(_135__bF$buf2),
    .Y(_139_)
);

OAI21X1 _822_ (
    .A(_135__bF$buf1),
    .B(_138_),
    .C(_139_),
    .Y(_21_)
);

NOR2X1 _823_ (
    .A(_136_),
    .B(_137_),
    .Y(_140_)
);

NAND2X1 _824_ (
    .A(XinHL[0]),
    .B(Cin[2]),
    .Y(_141_)
);

NAND2X1 _825_ (
    .A(XinHL[2]),
    .B(Cin_1_bF$buf1),
    .Y(_142_)
);

NOR2X1 _826_ (
    .A(_137_),
    .B(_142_),
    .Y(_143_)
);

AOI22X1 _827_ (
    .A(XinHL[1]),
    .B(Cin_1_bF$buf0),
    .C(XinHL[2]),
    .D(Cin_0_bF$buf1),
    .Y(_144_)
);

OAI21X1 _828_ (
    .A(_144_),
    .B(_143_),
    .C(_141_),
    .Y(_145_)
);

INVX1 _829_ (
    .A(_141_),
    .Y(_146_)
);

AND2X2 _830_ (
    .A(XinHL[1]),
    .B(Cin_0_bF$buf0),
    .Y(_147_)
);

AND2X2 _831_ (
    .A(XinHL[2]),
    .B(Cin_1_bF$buf3),
    .Y(_148_)
);

NAND2X1 _832_ (
    .A(_147_),
    .B(_148_),
    .Y(_149_)
);

INVX1 _833_ (
    .A(XinHL[1]),
    .Y(_150_)
);

INVX1 _834_ (
    .A(Cin_1_bF$buf2),
    .Y(_151_)
);

NAND2X1 _835_ (
    .A(XinHL[2]),
    .B(Cin_0_bF$buf3),
    .Y(_152_)
);

OAI21X1 _836_ (
    .A(_150_),
    .B(_151_),
    .C(_152_),
    .Y(_153_)
);

NAND3X1 _837_ (
    .A(_153_),
    .B(_146_),
    .C(_149_),
    .Y(_154_)
);

NAND3X1 _838_ (
    .A(_140_),
    .B(_154_),
    .C(_145_),
    .Y(_155_)
);

INVX1 _839_ (
    .A(_155_),
    .Y(_156_)
);

AOI21X1 _840_ (
    .A(_145_),
    .B(_154_),
    .C(_140_),
    .Y(_157_)
);

OAI21X1 _841_ (
    .A(_157_),
    .B(_156_),
    .C(LoadCtl_4_bF$buf4),
    .Y(_158_)
);

INVX1 _842_ (
    .A(mul[2]),
    .Y(_159_)
);

NAND2X1 _843_ (
    .A(_159_),
    .B(_135__bF$buf0),
    .Y(_160_)
);

AND2X2 _844_ (
    .A(_158_),
    .B(_160_),
    .Y(_22_)
);

INVX1 _845_ (
    .A(mul[3]),
    .Y(_161_)
);

NAND2X1 _846_ (
    .A(XinHL[0]),
    .B(Cin[3]),
    .Y(_162_)
);

AOI21X1 _847_ (
    .A(_146_),
    .B(_153_),
    .C(_143_),
    .Y(_163_)
);

NAND2X1 _848_ (
    .A(XinHL[1]),
    .B(Cin[2]),
    .Y(_164_)
);

NAND2X1 _849_ (
    .A(XinHL[3]),
    .B(Cin_0_bF$buf2),
    .Y(_165_)
);

NOR2X1 _850_ (
    .A(_142_),
    .B(_165_),
    .Y(_166_)
);

AOI22X1 _851_ (
    .A(XinHL[2]),
    .B(Cin_1_bF$buf1),
    .C(XinHL[3]),
    .D(Cin_0_bF$buf1),
    .Y(_167_)
);

OAI21X1 _852_ (
    .A(_167_),
    .B(_166_),
    .C(_164_),
    .Y(_168_)
);

INVX1 _853_ (
    .A(_164_),
    .Y(_169_)
);

AND2X2 _854_ (
    .A(XinHL[3]),
    .B(Cin_0_bF$buf0),
    .Y(_170_)
);

NAND2X1 _855_ (
    .A(_148_),
    .B(_170_),
    .Y(_171_)
);

INVX1 _856_ (
    .A(_167_),
    .Y(_172_)
);

NAND3X1 _857_ (
    .A(_169_),
    .B(_172_),
    .C(_171_),
    .Y(_173_)
);

NAND3X1 _858_ (
    .A(_173_),
    .B(_168_),
    .C(_163_),
    .Y(_174_)
);

OAI21X1 _859_ (
    .A(_141_),
    .B(_144_),
    .C(_149_),
    .Y(_175_)
);

AOI21X1 _860_ (
    .A(_171_),
    .B(_172_),
    .C(_169_),
    .Y(_176_)
);

INVX2 _861_ (
    .A(XinHL[2]),
    .Y(_177_)
);

OAI21X1 _862_ (
    .A(_177_),
    .B(_151_),
    .C(_170_),
    .Y(_178_)
);

INVX2 _863_ (
    .A(XinHL[3]),
    .Y(_179_)
);

INVX1 _864_ (
    .A(Cin_0_bF$buf3),
    .Y(_180_)
);

OAI21X1 _865_ (
    .A(_179_),
    .B(_180_),
    .C(_148_),
    .Y(_181_)
);

AOI21X1 _866_ (
    .A(_178_),
    .B(_181_),
    .C(_164_),
    .Y(_182_)
);

OAI21X1 _867_ (
    .A(_176_),
    .B(_182_),
    .C(_175_),
    .Y(_183_)
);

NAND3X1 _868_ (
    .A(_162_),
    .B(_174_),
    .C(_183_),
    .Y(_184_)
);

INVX1 _869_ (
    .A(_162_),
    .Y(_185_)
);

NAND3X1 _870_ (
    .A(_175_),
    .B(_173_),
    .C(_168_),
    .Y(_186_)
);

OAI21X1 _871_ (
    .A(_176_),
    .B(_182_),
    .C(_163_),
    .Y(_187_)
);

NAND3X1 _872_ (
    .A(_185_),
    .B(_186_),
    .C(_187_),
    .Y(_188_)
);

AOI21X1 _873_ (
    .A(_184_),
    .B(_188_),
    .C(_156_),
    .Y(_189_)
);

NAND3X1 _874_ (
    .A(_156_),
    .B(_184_),
    .C(_188_),
    .Y(_190_)
);

NAND2X1 _875_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_190_),
    .Y(_191_)
);

OAI22X1 _876_ (
    .A(_161_),
    .B(LoadCtl_4_bF$buf2),
    .C(_189_),
    .D(_191_),
    .Y(_23_)
);

INVX1 _877_ (
    .A(mul[4]),
    .Y(_192_)
);

INVX1 _878_ (
    .A(_190_),
    .Y(_193_)
);

AOI21X1 _879_ (
    .A(_168_),
    .B(_173_),
    .C(_175_),
    .Y(_194_)
);

OAI21X1 _880_ (
    .A(_162_),
    .B(_194_),
    .C(_186_),
    .Y(_195_)
);

OAI21X1 _881_ (
    .A(_164_),
    .B(_167_),
    .C(_171_),
    .Y(_196_)
);

AND2X2 _882_ (
    .A(XinH[0]),
    .B(Cin_1_bF$buf0),
    .Y(_197_)
);

NAND2X1 _883_ (
    .A(_170_),
    .B(_197_),
    .Y(_198_)
);

AOI22X1 _884_ (
    .A(XinH[0]),
    .B(Cin_0_bF$buf2),
    .C(XinHL[3]),
    .D(Cin_1_bF$buf3),
    .Y(_199_)
);

INVX1 _885_ (
    .A(_199_),
    .Y(_200_)
);

NAND2X1 _886_ (
    .A(XinHL[2]),
    .B(Cin[2]),
    .Y(_201_)
);

INVX1 _887_ (
    .A(_201_),
    .Y(_202_)
);

NAND3X1 _888_ (
    .A(_202_),
    .B(_200_),
    .C(_198_),
    .Y(_203_)
);

NAND2X1 _889_ (
    .A(XinH[0]),
    .B(Cin_1_bF$buf2),
    .Y(_204_)
);

NOR2X1 _890_ (
    .A(_165_),
    .B(_204_),
    .Y(_205_)
);

OAI21X1 _891_ (
    .A(_199_),
    .B(_205_),
    .C(_201_),
    .Y(_206_)
);

AOI21X1 _892_ (
    .A(_206_),
    .B(_203_),
    .C(_196_),
    .Y(_207_)
);

AOI21X1 _893_ (
    .A(_169_),
    .B(_172_),
    .C(_166_),
    .Y(_208_)
);

NAND3X1 _894_ (
    .A(_201_),
    .B(_200_),
    .C(_198_),
    .Y(_209_)
);

OAI21X1 _895_ (
    .A(_199_),
    .B(_205_),
    .C(_202_),
    .Y(_210_)
);

AOI21X1 _896_ (
    .A(_210_),
    .B(_209_),
    .C(_208_),
    .Y(_211_)
);

NAND2X1 _897_ (
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_212_)
);

INVX1 _898_ (
    .A(XinHL[0]),
    .Y(_213_)
);

INVX2 _899_ (
    .A(Cin[4]),
    .Y(_214_)
);

NAND2X1 _900_ (
    .A(XinHL[1]),
    .B(Cin[3]),
    .Y(_215_)
);

OAI21X1 _901_ (
    .A(_213_),
    .B(_214_),
    .C(_215_),
    .Y(_216_)
);

OAI21X1 _902_ (
    .A(_162_),
    .B(_212_),
    .C(_216_),
    .Y(_217_)
);

OAI21X1 _903_ (
    .A(_207_),
    .B(_211_),
    .C(_217_),
    .Y(_218_)
);

NAND3X1 _904_ (
    .A(_209_),
    .B(_210_),
    .C(_208_),
    .Y(_219_)
);

NAND3X1 _905_ (
    .A(_196_),
    .B(_203_),
    .C(_206_),
    .Y(_220_)
);

INVX1 _906_ (
    .A(_217_),
    .Y(_221_)
);

NAND3X1 _907_ (
    .A(_221_),
    .B(_220_),
    .C(_219_),
    .Y(_222_)
);

NAND3X1 _908_ (
    .A(_222_),
    .B(_195_),
    .C(_218_),
    .Y(_223_)
);

INVX1 _909_ (
    .A(_186_),
    .Y(_224_)
);

AOI21X1 _910_ (
    .A(_185_),
    .B(_187_),
    .C(_224_),
    .Y(_225_)
);

AOI21X1 _911_ (
    .A(_219_),
    .B(_220_),
    .C(_221_),
    .Y(_226_)
);

INVX1 _912_ (
    .A(_222_),
    .Y(_227_)
);

OAI21X1 _913_ (
    .A(_226_),
    .B(_227_),
    .C(_225_),
    .Y(_228_)
);

AOI21X1 _914_ (
    .A(_223_),
    .B(_228_),
    .C(_193_),
    .Y(_229_)
);

NAND3X1 _915_ (
    .A(_223_),
    .B(_228_),
    .C(_193_),
    .Y(_230_)
);

NAND2X1 _916_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_230_),
    .Y(_231_)
);

OAI22X1 _917_ (
    .A(_192_),
    .B(LoadCtl_4_bF$buf0),
    .C(_229_),
    .D(_231_),
    .Y(_24_)
);

AND2X2 _918_ (
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_232_)
);

NAND2X1 _919_ (
    .A(_232_),
    .B(_185_),
    .Y(_233_)
);

INVX1 _920_ (
    .A(_233_),
    .Y(_234_)
);

AOI21X1 _921_ (
    .A(_219_),
    .B(_221_),
    .C(_211_),
    .Y(_235_)
);

NAND2X1 _922_ (
    .A(XinHL[0]),
    .B(Cin[5]),
    .Y(_236_)
);

AND2X2 _923_ (
    .A(XinHL[2]),
    .B(Cin[3]),
    .Y(_237_)
);

OAI21X1 _924_ (
    .A(_150_),
    .B(_214_),
    .C(_237_),
    .Y(_238_)
);

INVX2 _925_ (
    .A(Cin[3]),
    .Y(_239_)
);

OAI21X1 _926_ (
    .A(_177_),
    .B(_239_),
    .C(_232_),
    .Y(_240_)
);

NAND3X1 _927_ (
    .A(_236_),
    .B(_238_),
    .C(_240_),
    .Y(_241_)
);

INVX1 _928_ (
    .A(_236_),
    .Y(_242_)
);

NAND2X1 _929_ (
    .A(_232_),
    .B(_237_),
    .Y(_243_)
);

OAI21X1 _930_ (
    .A(_177_),
    .B(_239_),
    .C(_212_),
    .Y(_244_)
);

NAND3X1 _931_ (
    .A(_244_),
    .B(_242_),
    .C(_243_),
    .Y(_245_)
);

NAND2X1 _932_ (
    .A(_245_),
    .B(_241_),
    .Y(_246_)
);

OAI22X1 _933_ (
    .A(_165_),
    .B(_204_),
    .C(_201_),
    .D(_199_),
    .Y(_247_)
);

INVX1 _934_ (
    .A(_247_),
    .Y(_248_)
);

NAND2X1 _935_ (
    .A(XinHL[3]),
    .B(Cin[2]),
    .Y(_249_)
);

NAND3X1 _936_ (
    .A(XinH[1]),
    .B(Cin_0_bF$buf1),
    .C(_204_),
    .Y(_250_)
);

NAND2X1 _937_ (
    .A(XinH[1]),
    .B(Cin_0_bF$buf0),
    .Y(_251_)
);

NAND3X1 _938_ (
    .A(XinH[0]),
    .B(Cin_1_bF$buf1),
    .C(_251_),
    .Y(_252_)
);

NAND3X1 _939_ (
    .A(_249_),
    .B(_250_),
    .C(_252_),
    .Y(_253_)
);

INVX1 _940_ (
    .A(_249_),
    .Y(_254_)
);

AND2X2 _941_ (
    .A(XinH[1]),
    .B(Cin_0_bF$buf3),
    .Y(_255_)
);

NAND2X1 _942_ (
    .A(_197_),
    .B(_255_),
    .Y(_256_)
);

OAI21X1 _943_ (
    .A(_91_),
    .B(_180_),
    .C(_204_),
    .Y(_257_)
);

NAND3X1 _944_ (
    .A(_254_),
    .B(_257_),
    .C(_256_),
    .Y(_258_)
);

NAND3X1 _945_ (
    .A(_253_),
    .B(_258_),
    .C(_248_),
    .Y(_259_)
);

AOI21X1 _946_ (
    .A(_256_),
    .B(_257_),
    .C(_254_),
    .Y(_260_)
);

AOI21X1 _947_ (
    .A(_250_),
    .B(_252_),
    .C(_249_),
    .Y(_261_)
);

OAI21X1 _948_ (
    .A(_261_),
    .B(_260_),
    .C(_247_),
    .Y(_262_)
);

NAND3X1 _949_ (
    .A(_246_),
    .B(_259_),
    .C(_262_),
    .Y(_263_)
);

AND2X2 _950_ (
    .A(_241_),
    .B(_245_),
    .Y(_264_)
);

NAND3X1 _951_ (
    .A(_247_),
    .B(_253_),
    .C(_258_),
    .Y(_265_)
);

OAI21X1 _952_ (
    .A(_261_),
    .B(_260_),
    .C(_248_),
    .Y(_266_)
);

NAND3X1 _953_ (
    .A(_265_),
    .B(_264_),
    .C(_266_),
    .Y(_267_)
);

NAND3X1 _954_ (
    .A(_263_),
    .B(_267_),
    .C(_235_),
    .Y(_268_)
);

OAI21X1 _955_ (
    .A(_217_),
    .B(_207_),
    .C(_220_),
    .Y(_269_)
);

AOI21X1 _956_ (
    .A(_266_),
    .B(_265_),
    .C(_264_),
    .Y(_270_)
);

AOI21X1 _957_ (
    .A(_262_),
    .B(_259_),
    .C(_246_),
    .Y(_271_)
);

OAI21X1 _958_ (
    .A(_270_),
    .B(_271_),
    .C(_269_),
    .Y(_272_)
);

NAND3X1 _959_ (
    .A(_234_),
    .B(_268_),
    .C(_272_),
    .Y(_273_)
);

NAND3X1 _960_ (
    .A(_263_),
    .B(_267_),
    .C(_269_),
    .Y(_274_)
);

OAI21X1 _961_ (
    .A(_270_),
    .B(_271_),
    .C(_235_),
    .Y(_275_)
);

NAND3X1 _962_ (
    .A(_233_),
    .B(_274_),
    .C(_275_),
    .Y(_276_)
);

NAND2X1 _963_ (
    .A(_273_),
    .B(_276_),
    .Y(_277_)
);

NAND2X1 _964_ (
    .A(_223_),
    .B(_230_),
    .Y(_278_)
);

XNOR2X1 _965_ (
    .A(_278_),
    .B(_277_),
    .Y(_279_)
);

NAND2X1 _966_ (
    .A(mul[5]),
    .B(_135__bF$buf5),
    .Y(_280_)
);

OAI21X1 _967_ (
    .A(_135__bF$buf4),
    .B(_279_),
    .C(_280_),
    .Y(_25_)
);

INVX1 _968_ (
    .A(mul[6]),
    .Y(_281_)
);

AOI22X1 _969_ (
    .A(_273_),
    .B(_276_),
    .C(_230_),
    .D(_223_),
    .Y(_282_)
);

AOI21X1 _970_ (
    .A(_263_),
    .B(_267_),
    .C(_269_),
    .Y(_283_)
);

OAI21X1 _971_ (
    .A(_233_),
    .B(_283_),
    .C(_274_),
    .Y(_284_)
);

NAND2X1 _972_ (
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_285_)
);

OAI21X1 _973_ (
    .A(_215_),
    .B(_285_),
    .C(_245_),
    .Y(_286_)
);

INVX1 _974_ (
    .A(_286_),
    .Y(_287_)
);

INVX1 _975_ (
    .A(_265_),
    .Y(_288_)
);

AOI21X1 _976_ (
    .A(_264_),
    .B(_266_),
    .C(_288_),
    .Y(_289_)
);

NAND2X1 _977_ (
    .A(XinHL[1]),
    .B(Cin[5]),
    .Y(_290_)
);

AND2X2 _978_ (
    .A(XinHL[3]),
    .B(Cin[3]),
    .Y(_291_)
);

OAI21X1 _979_ (
    .A(_177_),
    .B(_214_),
    .C(_291_),
    .Y(_292_)
);

AND2X2 _980_ (
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_293_)
);

OAI21X1 _981_ (
    .A(_179_),
    .B(_239_),
    .C(_293_),
    .Y(_294_)
);

NAND3X1 _982_ (
    .A(_290_),
    .B(_292_),
    .C(_294_),
    .Y(_295_)
);

INVX1 _983_ (
    .A(_290_),
    .Y(_296_)
);

NAND2X1 _984_ (
    .A(_293_),
    .B(_291_),
    .Y(_297_)
);

OAI21X1 _985_ (
    .A(_179_),
    .B(_239_),
    .C(_285_),
    .Y(_298_)
);

NAND3X1 _986_ (
    .A(_298_),
    .B(_296_),
    .C(_297_),
    .Y(_299_)
);

NAND2X1 _987_ (
    .A(_299_),
    .B(_295_),
    .Y(_300_)
);

NOR2X1 _988_ (
    .A(_204_),
    .B(_251_),
    .Y(_301_)
);

AOI21X1 _989_ (
    .A(_254_),
    .B(_257_),
    .C(_301_),
    .Y(_302_)
);

NAND2X1 _990_ (
    .A(XinH[0]),
    .B(Cin[2]),
    .Y(_303_)
);

NAND2X1 _991_ (
    .A(XinH[1]),
    .B(Cin_1_bF$buf0),
    .Y(_304_)
);

NAND3X1 _992_ (
    .A(XinH[2]),
    .B(Cin_0_bF$buf2),
    .C(_304_),
    .Y(_305_)
);

NAND2X1 _993_ (
    .A(XinH[2]),
    .B(Cin_0_bF$buf1),
    .Y(_306_)
);

NAND3X1 _994_ (
    .A(XinH[1]),
    .B(Cin_1_bF$buf3),
    .C(_306_),
    .Y(_307_)
);

NAND3X1 _995_ (
    .A(_303_),
    .B(_305_),
    .C(_307_),
    .Y(_308_)
);

INVX1 _996_ (
    .A(_303_),
    .Y(_309_)
);

AND2X2 _997_ (
    .A(XinH[2]),
    .B(Cin_1_bF$buf2),
    .Y(_310_)
);

NAND2X1 _998_ (
    .A(_255_),
    .B(_310_),
    .Y(_311_)
);

OAI21X1 _999_ (
    .A(_93_),
    .B(_180_),
    .C(_304_),
    .Y(_312_)
);

endmodule
