magic
tech scmos
magscale 1 6
timestamp 1709081121
<< checkpaint >>
rect 46 4691 482 5132
rect 45 4081 482 4691
rect 47 3959 482 4081
rect 39 2121 482 3959
rect 50 -120 475 1680
<< nwell >>
rect 0 4201 362 4571
rect 0 2241 362 3839
<< psubstratepdiff >>
rect 27 4680 335 5012
rect 27 0 335 1560
<< nsubstratendiff >>
rect 27 4220 335 4552
rect 27 2260 335 3820
<< genericcontact >>
rect 49 4926 61 4938
rect 113 4926 125 4938
rect 197 4926 209 4938
rect 261 4926 273 4938
rect 49 4862 61 4874
rect 113 4862 125 4874
rect 197 4862 209 4874
rect 261 4862 273 4874
rect 49 4798 61 4810
rect 113 4798 125 4810
rect 197 4798 209 4810
rect 261 4798 273 4810
rect 49 4734 61 4746
rect 113 4734 125 4746
rect 197 4734 209 4746
rect 261 4734 273 4746
rect 49 4450 61 4462
rect 113 4450 125 4462
rect 197 4450 209 4462
rect 261 4450 273 4462
rect 49 4386 61 4398
rect 113 4386 125 4398
rect 197 4386 209 4398
rect 261 4386 273 4398
rect 49 4322 61 4334
rect 113 4322 125 4334
rect 197 4322 209 4334
rect 261 4322 273 4334
rect 49 4258 61 4270
rect 113 4258 125 4270
rect 197 4258 209 4270
rect 261 4258 273 4270
rect 49 3766 61 3778
rect 113 3766 125 3778
rect 197 3766 209 3778
rect 261 3766 273 3778
rect 49 3702 61 3714
rect 113 3702 125 3714
rect 197 3702 209 3714
rect 261 3702 273 3714
rect 49 3638 61 3650
rect 113 3638 125 3650
rect 197 3638 209 3650
rect 261 3638 273 3650
rect 49 3574 61 3586
rect 113 3574 125 3586
rect 197 3574 209 3586
rect 261 3574 273 3586
rect 49 3510 61 3522
rect 113 3510 125 3522
rect 197 3510 209 3522
rect 261 3510 273 3522
rect 49 3446 61 3458
rect 113 3446 125 3458
rect 197 3446 209 3458
rect 261 3446 273 3458
rect 49 3382 61 3394
rect 113 3382 125 3394
rect 197 3382 209 3394
rect 261 3382 273 3394
rect 49 3318 61 3330
rect 113 3318 125 3330
rect 197 3318 209 3330
rect 261 3318 273 3330
rect 49 3254 61 3266
rect 113 3254 125 3266
rect 197 3254 209 3266
rect 261 3254 273 3266
rect 49 3190 61 3202
rect 113 3190 125 3202
rect 197 3190 209 3202
rect 261 3190 273 3202
rect 49 3126 61 3138
rect 113 3126 125 3138
rect 197 3126 209 3138
rect 261 3126 273 3138
rect 49 3062 61 3074
rect 113 3062 125 3074
rect 197 3062 209 3074
rect 261 3062 273 3074
rect 49 2998 61 3010
rect 113 2998 125 3010
rect 197 2998 209 3010
rect 261 2998 273 3010
rect 49 2934 61 2946
rect 113 2934 125 2946
rect 197 2934 209 2946
rect 261 2934 273 2946
rect 49 2870 61 2882
rect 113 2870 125 2882
rect 197 2870 209 2882
rect 261 2870 273 2882
rect 49 2806 61 2818
rect 113 2806 125 2818
rect 197 2806 209 2818
rect 261 2806 273 2818
rect 49 2742 61 2754
rect 113 2742 125 2754
rect 197 2742 209 2754
rect 261 2742 273 2754
rect 49 2678 61 2690
rect 113 2678 125 2690
rect 197 2678 209 2690
rect 261 2678 273 2690
rect 49 2614 61 2626
rect 113 2614 125 2626
rect 197 2614 209 2626
rect 261 2614 273 2626
rect 49 2550 61 2562
rect 113 2550 125 2562
rect 197 2550 209 2562
rect 261 2550 273 2562
rect 49 2486 61 2498
rect 113 2486 125 2498
rect 197 2486 209 2498
rect 261 2486 273 2498
rect 49 2422 61 2434
rect 113 2422 125 2434
rect 197 2422 209 2434
rect 261 2422 273 2434
rect 49 2358 61 2370
rect 113 2358 125 2370
rect 197 2358 209 2370
rect 261 2358 273 2370
rect 49 2294 61 2306
rect 113 2294 125 2306
rect 197 2294 209 2306
rect 261 2294 273 2306
rect 55 1488 67 1500
rect 119 1488 131 1500
rect 203 1488 215 1500
rect 267 1488 279 1500
rect 55 1424 67 1436
rect 119 1424 131 1436
rect 203 1424 215 1436
rect 267 1424 279 1436
rect 55 1360 67 1372
rect 119 1360 131 1372
rect 203 1360 215 1372
rect 267 1360 279 1372
rect 55 1296 67 1308
rect 119 1296 131 1308
rect 203 1296 215 1308
rect 267 1296 279 1308
rect 55 1232 67 1244
rect 119 1232 131 1244
rect 203 1232 215 1244
rect 267 1232 279 1244
rect 55 1168 67 1180
rect 119 1168 131 1180
rect 203 1168 215 1180
rect 267 1168 279 1180
rect 55 1104 67 1116
rect 119 1104 131 1116
rect 203 1104 215 1116
rect 267 1104 279 1116
rect 55 1040 67 1052
rect 119 1040 131 1052
rect 203 1040 215 1052
rect 267 1040 279 1052
rect 55 976 67 988
rect 119 976 131 988
rect 203 976 215 988
rect 267 976 279 988
rect 55 912 67 924
rect 119 912 131 924
rect 203 912 215 924
rect 267 912 279 924
rect 55 848 67 860
rect 119 848 131 860
rect 203 848 215 860
rect 267 848 279 860
rect 55 784 67 796
rect 119 784 131 796
rect 203 784 215 796
rect 267 784 279 796
rect 55 720 67 732
rect 119 720 131 732
rect 203 720 215 732
rect 267 720 279 732
rect 55 656 67 668
rect 119 656 131 668
rect 203 656 215 668
rect 267 656 279 668
rect 55 592 67 604
rect 119 592 131 604
rect 203 592 215 604
rect 267 592 279 604
rect 55 528 67 540
rect 119 528 131 540
rect 203 528 215 540
rect 267 528 279 540
rect 55 464 67 476
rect 119 464 131 476
rect 203 464 215 476
rect 267 464 279 476
rect 55 400 67 412
rect 119 400 131 412
rect 203 400 215 412
rect 267 400 279 412
rect 55 336 67 348
rect 119 336 131 348
rect 203 336 215 348
rect 267 336 279 348
rect 55 272 67 284
rect 119 272 131 284
rect 203 272 215 284
rect 267 272 279 284
rect 55 208 67 220
rect 119 208 131 220
rect 203 208 215 220
rect 267 208 279 220
rect 55 144 67 156
rect 119 144 131 156
rect 203 144 215 156
rect 267 144 279 156
rect 55 80 67 92
rect 119 80 131 92
rect 203 80 215 92
rect 267 80 279 92
rect 55 16 67 28
rect 119 16 131 28
rect 203 16 215 28
rect 267 16 279 28
<< metal1 >>
rect 31 4680 331 5012
rect 31 4220 331 4552
rect 31 2260 331 3820
rect 31 0 331 1560
<< metal2 >>
rect 31 4680 331 5012
rect 31 4220 331 4552
rect 31 2260 331 3820
rect 31 0 331 1560
<< gv1 >>
rect 79 4892 95 4908
rect 143 4892 159 4908
rect 227 4892 243 4908
rect 291 4892 307 4908
rect 79 4828 95 4844
rect 143 4828 159 4844
rect 227 4828 243 4844
rect 291 4828 307 4844
rect 79 4764 95 4780
rect 143 4764 159 4780
rect 227 4764 243 4780
rect 291 4764 307 4780
rect 79 4416 95 4432
rect 143 4416 159 4432
rect 227 4416 243 4432
rect 291 4416 307 4432
rect 79 4352 95 4368
rect 143 4352 159 4368
rect 227 4352 243 4368
rect 291 4352 307 4368
rect 79 4288 95 4304
rect 143 4288 159 4304
rect 227 4288 243 4304
rect 291 4288 307 4304
rect 79 3732 95 3748
rect 143 3732 159 3748
rect 227 3732 243 3748
rect 291 3732 307 3748
rect 79 3668 95 3684
rect 143 3668 159 3684
rect 227 3668 243 3684
rect 291 3668 307 3684
rect 79 3604 95 3620
rect 143 3604 159 3620
rect 227 3604 243 3620
rect 291 3604 307 3620
rect 79 3540 95 3556
rect 143 3540 159 3556
rect 227 3540 243 3556
rect 291 3540 307 3556
rect 79 3476 95 3492
rect 143 3476 159 3492
rect 227 3476 243 3492
rect 291 3476 307 3492
rect 79 3412 95 3428
rect 143 3412 159 3428
rect 227 3412 243 3428
rect 291 3412 307 3428
rect 79 3348 95 3364
rect 143 3348 159 3364
rect 227 3348 243 3364
rect 291 3348 307 3364
rect 79 3284 95 3300
rect 143 3284 159 3300
rect 227 3284 243 3300
rect 291 3284 307 3300
rect 79 3220 95 3236
rect 143 3220 159 3236
rect 227 3220 243 3236
rect 291 3220 307 3236
rect 79 3156 95 3172
rect 143 3156 159 3172
rect 227 3156 243 3172
rect 291 3156 307 3172
rect 79 3092 95 3108
rect 143 3092 159 3108
rect 227 3092 243 3108
rect 291 3092 307 3108
rect 79 3028 95 3044
rect 143 3028 159 3044
rect 227 3028 243 3044
rect 291 3028 307 3044
rect 79 2964 95 2980
rect 143 2964 159 2980
rect 227 2964 243 2980
rect 291 2964 307 2980
rect 79 2900 95 2916
rect 143 2900 159 2916
rect 227 2900 243 2916
rect 291 2900 307 2916
rect 79 2836 95 2852
rect 143 2836 159 2852
rect 227 2836 243 2852
rect 291 2836 307 2852
rect 79 2772 95 2788
rect 143 2772 159 2788
rect 227 2772 243 2788
rect 291 2772 307 2788
rect 79 2708 95 2724
rect 143 2708 159 2724
rect 227 2708 243 2724
rect 291 2708 307 2724
rect 79 2644 95 2660
rect 143 2644 159 2660
rect 227 2644 243 2660
rect 291 2644 307 2660
rect 79 2580 95 2596
rect 143 2580 159 2596
rect 227 2580 243 2596
rect 291 2580 307 2596
rect 79 2516 95 2532
rect 143 2516 159 2532
rect 227 2516 243 2532
rect 291 2516 307 2532
rect 79 2452 95 2468
rect 143 2452 159 2468
rect 227 2452 243 2468
rect 291 2452 307 2468
rect 79 2388 95 2404
rect 143 2388 159 2404
rect 227 2388 243 2404
rect 291 2388 307 2404
rect 79 2324 95 2340
rect 143 2324 159 2340
rect 227 2324 243 2340
rect 291 2324 307 2340
rect 85 1454 101 1470
rect 149 1454 165 1470
rect 233 1454 249 1470
rect 297 1454 313 1470
rect 85 1390 101 1406
rect 149 1390 165 1406
rect 233 1390 249 1406
rect 297 1390 313 1406
rect 85 1326 101 1342
rect 149 1326 165 1342
rect 233 1326 249 1342
rect 297 1326 313 1342
rect 85 1262 101 1278
rect 149 1262 165 1278
rect 233 1262 249 1278
rect 297 1262 313 1278
rect 85 1198 101 1214
rect 149 1198 165 1214
rect 233 1198 249 1214
rect 297 1198 313 1214
rect 85 1134 101 1150
rect 149 1134 165 1150
rect 233 1134 249 1150
rect 297 1134 313 1150
rect 85 1070 101 1086
rect 149 1070 165 1086
rect 233 1070 249 1086
rect 297 1070 313 1086
rect 85 1006 101 1022
rect 149 1006 165 1022
rect 233 1006 249 1022
rect 297 1006 313 1022
rect 85 942 101 958
rect 149 942 165 958
rect 233 942 249 958
rect 297 942 313 958
rect 85 878 101 894
rect 149 878 165 894
rect 233 878 249 894
rect 297 878 313 894
rect 85 814 101 830
rect 149 814 165 830
rect 233 814 249 830
rect 297 814 313 830
rect 85 750 101 766
rect 149 750 165 766
rect 233 750 249 766
rect 297 750 313 766
rect 85 686 101 702
rect 149 686 165 702
rect 233 686 249 702
rect 297 686 313 702
rect 85 622 101 638
rect 149 622 165 638
rect 233 622 249 638
rect 297 622 313 638
rect 85 558 101 574
rect 149 558 165 574
rect 233 558 249 574
rect 297 558 313 574
rect 85 494 101 510
rect 149 494 165 510
rect 233 494 249 510
rect 297 494 313 510
rect 85 430 101 446
rect 149 430 165 446
rect 233 430 249 446
rect 297 430 313 446
rect 85 366 101 382
rect 149 366 165 382
rect 233 366 249 382
rect 297 366 313 382
rect 85 302 101 318
rect 149 302 165 318
rect 233 302 249 318
rect 297 302 313 318
rect 85 238 101 254
rect 149 238 165 254
rect 233 238 249 254
rect 297 238 313 254
rect 85 174 101 190
rect 149 174 165 190
rect 233 174 249 190
rect 297 174 313 190
rect 85 110 101 126
rect 149 110 165 126
rect 233 110 249 126
rect 297 110 313 126
rect 85 46 101 62
rect 149 46 165 62
rect 233 46 249 62
rect 297 46 313 62
<< metal3 >>
rect 7 4680 355 5012
rect 7 4220 355 4552
rect 7 2260 355 3820
rect 7 0 355 1560
<< gv2 >>
rect 47 4924 63 4940
rect 111 4924 127 4940
rect 195 4924 211 4940
rect 259 4924 275 4940
rect 47 4860 63 4876
rect 111 4860 127 4876
rect 195 4860 211 4876
rect 259 4860 275 4876
rect 47 4796 63 4812
rect 111 4796 127 4812
rect 195 4796 211 4812
rect 259 4796 275 4812
rect 47 4732 63 4748
rect 111 4732 127 4748
rect 195 4732 211 4748
rect 259 4732 275 4748
rect 47 4448 63 4464
rect 111 4448 127 4464
rect 195 4448 211 4464
rect 259 4448 275 4464
rect 47 4384 63 4400
rect 111 4384 127 4400
rect 195 4384 211 4400
rect 259 4384 275 4400
rect 47 4320 63 4336
rect 111 4320 127 4336
rect 195 4320 211 4336
rect 259 4320 275 4336
rect 47 4256 63 4272
rect 111 4256 127 4272
rect 195 4256 211 4272
rect 259 4256 275 4272
rect 47 3764 63 3780
rect 111 3764 127 3780
rect 195 3764 211 3780
rect 259 3764 275 3780
rect 47 3700 63 3716
rect 111 3700 127 3716
rect 195 3700 211 3716
rect 259 3700 275 3716
rect 47 3636 63 3652
rect 111 3636 127 3652
rect 195 3636 211 3652
rect 259 3636 275 3652
rect 47 3572 63 3588
rect 111 3572 127 3588
rect 195 3572 211 3588
rect 259 3572 275 3588
rect 47 3508 63 3524
rect 111 3508 127 3524
rect 195 3508 211 3524
rect 259 3508 275 3524
rect 47 3444 63 3460
rect 111 3444 127 3460
rect 195 3444 211 3460
rect 259 3444 275 3460
rect 47 3380 63 3396
rect 111 3380 127 3396
rect 195 3380 211 3396
rect 259 3380 275 3396
rect 47 3316 63 3332
rect 111 3316 127 3332
rect 195 3316 211 3332
rect 259 3316 275 3332
rect 47 3252 63 3268
rect 111 3252 127 3268
rect 195 3252 211 3268
rect 259 3252 275 3268
rect 47 3188 63 3204
rect 111 3188 127 3204
rect 195 3188 211 3204
rect 259 3188 275 3204
rect 47 3124 63 3140
rect 111 3124 127 3140
rect 195 3124 211 3140
rect 259 3124 275 3140
rect 47 3060 63 3076
rect 111 3060 127 3076
rect 195 3060 211 3076
rect 259 3060 275 3076
rect 47 2996 63 3012
rect 111 2996 127 3012
rect 195 2996 211 3012
rect 259 2996 275 3012
rect 47 2932 63 2948
rect 111 2932 127 2948
rect 195 2932 211 2948
rect 259 2932 275 2948
rect 47 2868 63 2884
rect 111 2868 127 2884
rect 195 2868 211 2884
rect 259 2868 275 2884
rect 47 2804 63 2820
rect 111 2804 127 2820
rect 195 2804 211 2820
rect 259 2804 275 2820
rect 47 2740 63 2756
rect 111 2740 127 2756
rect 195 2740 211 2756
rect 259 2740 275 2756
rect 47 2676 63 2692
rect 111 2676 127 2692
rect 195 2676 211 2692
rect 259 2676 275 2692
rect 47 2612 63 2628
rect 111 2612 127 2628
rect 195 2612 211 2628
rect 259 2612 275 2628
rect 47 2548 63 2564
rect 111 2548 127 2564
rect 195 2548 211 2564
rect 259 2548 275 2564
rect 47 2484 63 2500
rect 111 2484 127 2500
rect 195 2484 211 2500
rect 259 2484 275 2500
rect 47 2420 63 2436
rect 111 2420 127 2436
rect 195 2420 211 2436
rect 259 2420 275 2436
rect 47 2356 63 2372
rect 111 2356 127 2372
rect 195 2356 211 2372
rect 259 2356 275 2372
rect 47 2292 63 2308
rect 111 2292 127 2308
rect 195 2292 211 2308
rect 259 2292 275 2308
rect 53 1486 69 1502
rect 117 1486 133 1502
rect 201 1486 217 1502
rect 265 1486 281 1502
rect 53 1422 69 1438
rect 117 1422 133 1438
rect 201 1422 217 1438
rect 265 1422 281 1438
rect 53 1358 69 1374
rect 117 1358 133 1374
rect 201 1358 217 1374
rect 265 1358 281 1374
rect 53 1294 69 1310
rect 117 1294 133 1310
rect 201 1294 217 1310
rect 265 1294 281 1310
rect 53 1230 69 1246
rect 117 1230 133 1246
rect 201 1230 217 1246
rect 265 1230 281 1246
rect 53 1166 69 1182
rect 117 1166 133 1182
rect 201 1166 217 1182
rect 265 1166 281 1182
rect 53 1102 69 1118
rect 117 1102 133 1118
rect 201 1102 217 1118
rect 265 1102 281 1118
rect 53 1038 69 1054
rect 117 1038 133 1054
rect 201 1038 217 1054
rect 265 1038 281 1054
rect 53 974 69 990
rect 117 974 133 990
rect 201 974 217 990
rect 265 974 281 990
rect 53 910 69 926
rect 117 910 133 926
rect 201 910 217 926
rect 265 910 281 926
rect 53 846 69 862
rect 117 846 133 862
rect 201 846 217 862
rect 265 846 281 862
rect 53 782 69 798
rect 117 782 133 798
rect 201 782 217 798
rect 265 782 281 798
rect 53 718 69 734
rect 117 718 133 734
rect 201 718 217 734
rect 265 718 281 734
rect 53 654 69 670
rect 117 654 133 670
rect 201 654 217 670
rect 265 654 281 670
rect 53 590 69 606
rect 117 590 133 606
rect 201 590 217 606
rect 265 590 281 606
rect 53 526 69 542
rect 117 526 133 542
rect 201 526 217 542
rect 265 526 281 542
rect 53 462 69 478
rect 117 462 133 478
rect 201 462 217 478
rect 265 462 281 478
rect 53 398 69 414
rect 117 398 133 414
rect 201 398 217 414
rect 265 398 281 414
rect 53 334 69 350
rect 117 334 133 350
rect 201 334 217 350
rect 265 334 281 350
rect 53 270 69 286
rect 117 270 133 286
rect 201 270 217 286
rect 265 270 281 286
rect 53 206 69 222
rect 117 206 133 222
rect 201 206 217 222
rect 265 206 281 222
rect 53 142 69 158
rect 117 142 133 158
rect 201 142 217 158
rect 265 142 281 158
rect 53 78 69 94
rect 117 78 133 94
rect 201 78 217 94
rect 265 78 281 94
rect 53 14 69 30
rect 117 14 133 30
rect 201 14 217 30
rect 265 14 281 30
<< end >>
