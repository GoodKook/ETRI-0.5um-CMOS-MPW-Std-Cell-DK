magic
tech scmos
magscale 1 6
timestamp 1569139307
<< checkpaint >>
rect -120 -120 5180 5180
<< metal1 >>
rect 0 2260 1560 5030
rect 2260 4220 3820 5030
rect 4220 4552 4552 5030
rect 4680 4991 4991 5036
tri 4991 4991 5036 5036 sw
rect 4680 4817 5036 4991
tri 4680 4680 4817 4817 ne
rect 4817 4680 5036 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5030 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5030 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5030 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5030 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5030 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5030 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5030 1560
<< metal2 >>
rect 0 2260 1560 5030
rect 2260 4220 3820 5030
rect 4220 4552 4552 5031
rect 4680 4991 4991 5036
tri 4991 4991 5036 5036 sw
rect 4680 4817 5036 4991
tri 4680 4680 4817 4817 ne
rect 4817 4680 5036 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5030 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5030 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5030 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5030 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5030 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5030 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5030 1560
<< metal3 >>
rect 0 2260 1560 5060
rect 2260 4220 3820 5060
rect 4220 4552 4552 5060
rect 4680 5012 5012 5060
tri 5012 5012 5060 5060 sw
rect 4680 4817 5060 5012
tri 4680 4680 4817 4817 ne
rect 4817 4680 5060 4817
tri 4552 4552 4641 4641 sw
rect 4220 4483 5060 4552
tri 4220 4249 4454 4483 ne
rect 4454 4249 5060 4483
tri 3820 4220 3849 4249 sw
tri 4454 4220 4483 4249 ne
rect 4483 4220 5060 4249
rect 2260 3820 3849 4220
tri 3849 3820 4249 4220 sw
rect 2260 3381 5060 3820
tri 2260 2952 2689 3381 ne
rect 2689 2952 5060 3381
tri 1560 2260 2252 2952 sw
tri 2689 2260 3381 2952 ne
rect 3381 2260 5060 2952
rect 0 1752 2252 2260
tri 0 0 1752 1752 ne
rect 1752 1560 2252 1752
tri 2252 1560 2952 2260 sw
rect 1752 0 5060 1560
use VIA1  VIA1_0
timestamp 1569139307
transform 1 0 4744 0 1 136
box -8 -8 8 8
use VIA1  VIA1_1
timestamp 1569139307
transform 1 0 4872 0 1 264
box -8 -8 8 8
use VIA1  VIA1_2
timestamp 1569139307
transform 1 0 4808 0 1 328
box -8 -8 8 8
use VIA1  VIA1_3
timestamp 1569139307
transform 1 0 4680 0 1 328
box -8 -8 8 8
use VIA1  VIA1_4
timestamp 1569139307
transform 1 0 4680 0 1 72
box -8 -8 8 8
use VIA1  VIA1_5
timestamp 1569139307
transform 1 0 4744 0 1 264
box -8 -8 8 8
use VIA1  VIA1_6
timestamp 1569139307
transform 1 0 4744 0 1 328
box -8 -8 8 8
use VIA1  VIA1_7
timestamp 1569139307
transform 1 0 4872 0 1 72
box -8 -8 8 8
use VIA1  VIA1_8
timestamp 1569139307
transform 1 0 4680 0 1 200
box -8 -8 8 8
use VIA1  VIA1_9
timestamp 1569139307
transform 1 0 4808 0 1 72
box -8 -8 8 8
use VIA1  VIA1_10
timestamp 1569139307
transform 1 0 4872 0 1 136
box -8 -8 8 8
use VIA1  VIA1_11
timestamp 1569139307
transform 1 0 4680 0 1 136
box -8 -8 8 8
use VIA1  VIA1_12
timestamp 1569139307
transform 1 0 4808 0 1 264
box -8 -8 8 8
use VIA1  VIA1_13
timestamp 1569139307
transform 1 0 4744 0 1 72
box -8 -8 8 8
use VIA1  VIA1_14
timestamp 1569139307
transform 1 0 4680 0 1 264
box -8 -8 8 8
use VIA1  VIA1_15
timestamp 1569139307
transform 1 0 4808 0 1 136
box -8 -8 8 8
use VIA1  VIA1_16
timestamp 1569139307
transform 1 0 4808 0 1 200
box -8 -8 8 8
use VIA1  VIA1_17
timestamp 1569139307
transform 1 0 4872 0 1 328
box -8 -8 8 8
use VIA1  VIA1_18
timestamp 1569139307
transform 1 0 4744 0 1 200
box -8 -8 8 8
use VIA1  VIA1_19
timestamp 1569139307
transform 1 0 4872 0 1 200
box -8 -8 8 8
use VIA1  VIA1_20
timestamp 1569139307
transform 1 0 4552 0 1 72
box -8 -8 8 8
use VIA1  VIA1_21
timestamp 1569139307
transform 1 0 4488 0 1 200
box -8 -8 8 8
use VIA1  VIA1_22
timestamp 1569139307
transform 1 0 4616 0 1 264
box -8 -8 8 8
use VIA1  VIA1_23
timestamp 1569139307
transform 1 0 4552 0 1 264
box -8 -8 8 8
use VIA1  VIA1_24
timestamp 1569139307
transform 1 0 4616 0 1 200
box -8 -8 8 8
use VIA1  VIA1_25
timestamp 1569139307
transform 1 0 4488 0 1 264
box -8 -8 8 8
use VIA1  VIA1_26
timestamp 1569139307
transform 1 0 4424 0 1 136
box -8 -8 8 8
use VIA1  VIA1_27
timestamp 1569139307
transform 1 0 4616 0 1 328
box -8 -8 8 8
use VIA1  VIA1_28
timestamp 1569139307
transform 1 0 4552 0 1 136
box -8 -8 8 8
use VIA1  VIA1_29
timestamp 1569139307
transform 1 0 4488 0 1 328
box -8 -8 8 8
use VIA1  VIA1_30
timestamp 1569139307
transform 1 0 4424 0 1 328
box -8 -8 8 8
use VIA1  VIA1_31
timestamp 1569139307
transform 1 0 4424 0 1 264
box -8 -8 8 8
use VIA1  VIA1_32
timestamp 1569139307
transform 1 0 4552 0 1 328
box -8 -8 8 8
use VIA1  VIA1_33
timestamp 1569139307
transform 1 0 4616 0 1 72
box -8 -8 8 8
use VIA1  VIA1_34
timestamp 1569139307
transform 1 0 4424 0 1 200
box -8 -8 8 8
use VIA1  VIA1_35
timestamp 1569139307
transform 1 0 4424 0 1 72
box -8 -8 8 8
use VIA1  VIA1_36
timestamp 1569139307
transform 1 0 4552 0 1 200
box -8 -8 8 8
use VIA1  VIA1_37
timestamp 1569139307
transform 1 0 4488 0 1 136
box -8 -8 8 8
use VIA1  VIA1_38
timestamp 1569139307
transform 1 0 4488 0 1 72
box -8 -8 8 8
use VIA1  VIA1_39
timestamp 1569139307
transform 1 0 4616 0 1 136
box -8 -8 8 8
use VIA1  VIA1_40
timestamp 1569139307
transform 1 0 4616 0 1 584
box -8 -8 8 8
use VIA1  VIA1_41
timestamp 1569139307
transform 1 0 4424 0 1 584
box -8 -8 8 8
use VIA1  VIA1_42
timestamp 1569139307
transform 1 0 4424 0 1 456
box -8 -8 8 8
use VIA1  VIA1_43
timestamp 1569139307
transform 1 0 4552 0 1 584
box -8 -8 8 8
use VIA1  VIA1_44
timestamp 1569139307
transform 1 0 4488 0 1 392
box -8 -8 8 8
use VIA1  VIA1_45
timestamp 1569139307
transform 1 0 4488 0 1 520
box -8 -8 8 8
use VIA1  VIA1_46
timestamp 1569139307
transform 1 0 4552 0 1 392
box -8 -8 8 8
use VIA1  VIA1_47
timestamp 1569139307
transform 1 0 4424 0 1 392
box -8 -8 8 8
use VIA1  VIA1_48
timestamp 1569139307
transform 1 0 4552 0 1 520
box -8 -8 8 8
use VIA1  VIA1_49
timestamp 1569139307
transform 1 0 4616 0 1 392
box -8 -8 8 8
use VIA1  VIA1_50
timestamp 1569139307
transform 1 0 4552 0 1 456
box -8 -8 8 8
use VIA1  VIA1_51
timestamp 1569139307
transform 1 0 4616 0 1 520
box -8 -8 8 8
use VIA1  VIA1_52
timestamp 1569139307
transform 1 0 4616 0 1 456
box -8 -8 8 8
use VIA1  VIA1_53
timestamp 1569139307
transform 1 0 4488 0 1 584
box -8 -8 8 8
use VIA1  VIA1_54
timestamp 1569139307
transform 1 0 4488 0 1 456
box -8 -8 8 8
use VIA1  VIA1_55
timestamp 1569139307
transform 1 0 4424 0 1 520
box -8 -8 8 8
use VIA1  VIA1_56
timestamp 1569139307
transform 1 0 4872 0 1 520
box -8 -8 8 8
use VIA1  VIA1_57
timestamp 1569139307
transform 1 0 4680 0 1 520
box -8 -8 8 8
use VIA1  VIA1_58
timestamp 1569139307
transform 1 0 4808 0 1 392
box -8 -8 8 8
use VIA1  VIA1_59
timestamp 1569139307
transform 1 0 4872 0 1 584
box -8 -8 8 8
use VIA1  VIA1_60
timestamp 1569139307
transform 1 0 4808 0 1 584
box -8 -8 8 8
use VIA1  VIA1_61
timestamp 1569139307
transform 1 0 4744 0 1 456
box -8 -8 8 8
use VIA1  VIA1_62
timestamp 1569139307
transform 1 0 4744 0 1 520
box -8 -8 8 8
use VIA1  VIA1_63
timestamp 1569139307
transform 1 0 4808 0 1 456
box -8 -8 8 8
use VIA1  VIA1_64
timestamp 1569139307
transform 1 0 4680 0 1 584
box -8 -8 8 8
use VIA1  VIA1_65
timestamp 1569139307
transform 1 0 4872 0 1 392
box -8 -8 8 8
use VIA1  VIA1_66
timestamp 1569139307
transform 1 0 4808 0 1 520
box -8 -8 8 8
use VIA1  VIA1_67
timestamp 1569139307
transform 1 0 4744 0 1 392
box -8 -8 8 8
use VIA1  VIA1_68
timestamp 1569139307
transform 1 0 4872 0 1 456
box -8 -8 8 8
use VIA1  VIA1_69
timestamp 1569139307
transform 1 0 4680 0 1 456
box -8 -8 8 8
use VIA1  VIA1_70
timestamp 1569139307
transform 1 0 4680 0 1 392
box -8 -8 8 8
use VIA1  VIA1_71
timestamp 1569139307
transform 1 0 4744 0 1 584
box -8 -8 8 8
use VIA1  VIA1_72
timestamp 1569139307
transform 1 0 4232 0 1 264
box -8 -8 8 8
use VIA1  VIA1_73
timestamp 1569139307
transform 1 0 4168 0 1 72
box -8 -8 8 8
use VIA1  VIA1_74
timestamp 1569139307
transform 1 0 4168 0 1 200
box -8 -8 8 8
use VIA1  VIA1_75
timestamp 1569139307
transform 1 0 4296 0 1 200
box -8 -8 8 8
use VIA1  VIA1_76
timestamp 1569139307
transform 1 0 4296 0 1 264
box -8 -8 8 8
use VIA1  VIA1_77
timestamp 1569139307
transform 1 0 4296 0 1 72
box -8 -8 8 8
use VIA1  VIA1_78
timestamp 1569139307
transform 1 0 4232 0 1 136
box -8 -8 8 8
use VIA1  VIA1_79
timestamp 1569139307
transform 1 0 4104 0 1 328
box -8 -8 8 8
use VIA1  VIA1_80
timestamp 1569139307
transform 1 0 4168 0 1 136
box -8 -8 8 8
use VIA1  VIA1_81
timestamp 1569139307
transform 1 0 4168 0 1 264
box -8 -8 8 8
use VIA1  VIA1_82
timestamp 1569139307
transform 1 0 4232 0 1 328
box -8 -8 8 8
use VIA1  VIA1_83
timestamp 1569139307
transform 1 0 4104 0 1 200
box -8 -8 8 8
use VIA1  VIA1_84
timestamp 1569139307
transform 1 0 4104 0 1 72
box -8 -8 8 8
use VIA1  VIA1_85
timestamp 1569139307
transform 1 0 4104 0 1 264
box -8 -8 8 8
use VIA1  VIA1_86
timestamp 1569139307
transform 1 0 4232 0 1 72
box -8 -8 8 8
use VIA1  VIA1_87
timestamp 1569139307
transform 1 0 4232 0 1 200
box -8 -8 8 8
use VIA1  VIA1_88
timestamp 1569139307
transform 1 0 4104 0 1 136
box -8 -8 8 8
use VIA1  VIA1_89
timestamp 1569139307
transform 1 0 4296 0 1 136
box -8 -8 8 8
use VIA1  VIA1_90
timestamp 1569139307
transform 1 0 4296 0 1 328
box -8 -8 8 8
use VIA1  VIA1_91
timestamp 1569139307
transform 1 0 4168 0 1 328
box -8 -8 8 8
use VIA1  VIA1_92
timestamp 1569139307
transform 1 0 3784 0 1 328
box -8 -8 8 8
use VIA1  VIA1_93
timestamp 1569139307
transform 1 0 3848 0 1 328
box -8 -8 8 8
use VIA1  VIA1_94
timestamp 1569139307
transform 1 0 3912 0 1 72
box -8 -8 8 8
use VIA1  VIA1_95
timestamp 1569139307
transform 1 0 4040 0 1 136
box -8 -8 8 8
use VIA1  VIA1_96
timestamp 1569139307
transform 1 0 4040 0 1 200
box -8 -8 8 8
use VIA1  VIA1_97
timestamp 1569139307
transform 1 0 3912 0 1 264
box -8 -8 8 8
use VIA1  VIA1_98
timestamp 1569139307
transform 1 0 3848 0 1 72
box -8 -8 8 8
use VIA1  VIA1_99
timestamp 1569139307
transform 1 0 3976 0 1 72
box -8 -8 8 8
use VIA1  VIA1_100
timestamp 1569139307
transform 1 0 3784 0 1 136
box -8 -8 8 8
use VIA1  VIA1_101
timestamp 1569139307
transform 1 0 3912 0 1 328
box -8 -8 8 8
use VIA1  VIA1_102
timestamp 1569139307
transform 1 0 4040 0 1 264
box -8 -8 8 8
use VIA1  VIA1_103
timestamp 1569139307
transform 1 0 3976 0 1 264
box -8 -8 8 8
use VIA1  VIA1_104
timestamp 1569139307
transform 1 0 4040 0 1 72
box -8 -8 8 8
use VIA1  VIA1_105
timestamp 1569139307
transform 1 0 3848 0 1 136
box -8 -8 8 8
use VIA1  VIA1_106
timestamp 1569139307
transform 1 0 3848 0 1 200
box -8 -8 8 8
use VIA1  VIA1_107
timestamp 1569139307
transform 1 0 3912 0 1 136
box -8 -8 8 8
use VIA1  VIA1_108
timestamp 1569139307
transform 1 0 4040 0 1 328
box -8 -8 8 8
use VIA1  VIA1_109
timestamp 1569139307
transform 1 0 3976 0 1 328
box -8 -8 8 8
use VIA1  VIA1_110
timestamp 1569139307
transform 1 0 3912 0 1 200
box -8 -8 8 8
use VIA1  VIA1_111
timestamp 1569139307
transform 1 0 3784 0 1 200
box -8 -8 8 8
use VIA1  VIA1_112
timestamp 1569139307
transform 1 0 3848 0 1 264
box -8 -8 8 8
use VIA1  VIA1_113
timestamp 1569139307
transform 1 0 3784 0 1 264
box -8 -8 8 8
use VIA1  VIA1_114
timestamp 1569139307
transform 1 0 3784 0 1 72
box -8 -8 8 8
use VIA1  VIA1_115
timestamp 1569139307
transform 1 0 3976 0 1 200
box -8 -8 8 8
use VIA1  VIA1_116
timestamp 1569139307
transform 1 0 3976 0 1 136
box -8 -8 8 8
use VIA1  VIA1_117
timestamp 1569139307
transform 1 0 3784 0 1 584
box -8 -8 8 8
use VIA1  VIA1_118
timestamp 1569139307
transform 1 0 3912 0 1 584
box -8 -8 8 8
use VIA1  VIA1_119
timestamp 1569139307
transform 1 0 3976 0 1 520
box -8 -8 8 8
use VIA1  VIA1_120
timestamp 1569139307
transform 1 0 3848 0 1 456
box -8 -8 8 8
use VIA1  VIA1_121
timestamp 1569139307
transform 1 0 4040 0 1 392
box -8 -8 8 8
use VIA1  VIA1_122
timestamp 1569139307
transform 1 0 3912 0 1 520
box -8 -8 8 8
use VIA1  VIA1_123
timestamp 1569139307
transform 1 0 4040 0 1 520
box -8 -8 8 8
use VIA1  VIA1_124
timestamp 1569139307
transform 1 0 3976 0 1 392
box -8 -8 8 8
use VIA1  VIA1_125
timestamp 1569139307
transform 1 0 3976 0 1 584
box -8 -8 8 8
use VIA1  VIA1_126
timestamp 1569139307
transform 1 0 3912 0 1 456
box -8 -8 8 8
use VIA1  VIA1_127
timestamp 1569139307
transform 1 0 3976 0 1 456
box -8 -8 8 8
use VIA1  VIA1_128
timestamp 1569139307
transform 1 0 3848 0 1 520
box -8 -8 8 8
use VIA1  VIA1_129
timestamp 1569139307
transform 1 0 3784 0 1 520
box -8 -8 8 8
use VIA1  VIA1_130
timestamp 1569139307
transform 1 0 4040 0 1 584
box -8 -8 8 8
use VIA1  VIA1_131
timestamp 1569139307
transform 1 0 3912 0 1 392
box -8 -8 8 8
use VIA1  VIA1_132
timestamp 1569139307
transform 1 0 3784 0 1 392
box -8 -8 8 8
use VIA1  VIA1_133
timestamp 1569139307
transform 1 0 3848 0 1 584
box -8 -8 8 8
use VIA1  VIA1_134
timestamp 1569139307
transform 1 0 4040 0 1 456
box -8 -8 8 8
use VIA1  VIA1_135
timestamp 1569139307
transform 1 0 3848 0 1 392
box -8 -8 8 8
use VIA1  VIA1_136
timestamp 1569139307
transform 1 0 3784 0 1 456
box -8 -8 8 8
use VIA1  VIA1_137
timestamp 1569139307
transform 1 0 4104 0 1 392
box -8 -8 8 8
use VIA1  VIA1_138
timestamp 1569139307
transform 1 0 4296 0 1 584
box -8 -8 8 8
use VIA1  VIA1_139
timestamp 1569139307
transform 1 0 4168 0 1 584
box -8 -8 8 8
use VIA1  VIA1_140
timestamp 1569139307
transform 1 0 4168 0 1 520
box -8 -8 8 8
use VIA1  VIA1_141
timestamp 1569139307
transform 1 0 4104 0 1 456
box -8 -8 8 8
use VIA1  VIA1_142
timestamp 1569139307
transform 1 0 4104 0 1 520
box -8 -8 8 8
use VIA1  VIA1_143
timestamp 1569139307
transform 1 0 4232 0 1 392
box -8 -8 8 8
use VIA1  VIA1_144
timestamp 1569139307
transform 1 0 4232 0 1 456
box -8 -8 8 8
use VIA1  VIA1_145
timestamp 1569139307
transform 1 0 4232 0 1 520
box -8 -8 8 8
use VIA1  VIA1_146
timestamp 1569139307
transform 1 0 4168 0 1 456
box -8 -8 8 8
use VIA1  VIA1_147
timestamp 1569139307
transform 1 0 4168 0 1 392
box -8 -8 8 8
use VIA1  VIA1_148
timestamp 1569139307
transform 1 0 4232 0 1 584
box -8 -8 8 8
use VIA1  VIA1_149
timestamp 1569139307
transform 1 0 4104 0 1 584
box -8 -8 8 8
use VIA1  VIA1_150
timestamp 1569139307
transform 1 0 4296 0 1 392
box -8 -8 8 8
use VIA1  VIA1_151
timestamp 1569139307
transform 1 0 4296 0 1 456
box -8 -8 8 8
use VIA1  VIA1_152
timestamp 1569139307
transform 1 0 4296 0 1 520
box -8 -8 8 8
use VIA1  VIA1_153
timestamp 1569139307
transform 1 0 4232 0 1 712
box -8 -8 8 8
use VIA1  VIA1_154
timestamp 1569139307
transform 1 0 4104 0 1 712
box -8 -8 8 8
use VIA1  VIA1_155
timestamp 1569139307
transform 1 0 4232 0 1 840
box -8 -8 8 8
use VIA1  VIA1_156
timestamp 1569139307
transform 1 0 4168 0 1 840
box -8 -8 8 8
use VIA1  VIA1_157
timestamp 1569139307
transform 1 0 4168 0 1 712
box -8 -8 8 8
use VIA1  VIA1_158
timestamp 1569139307
transform 1 0 4168 0 1 904
box -8 -8 8 8
use VIA1  VIA1_159
timestamp 1569139307
transform 1 0 4168 0 1 776
box -8 -8 8 8
use VIA1  VIA1_160
timestamp 1569139307
transform 1 0 4232 0 1 776
box -8 -8 8 8
use VIA1  VIA1_161
timestamp 1569139307
transform 1 0 4104 0 1 776
box -8 -8 8 8
use VIA1  VIA1_162
timestamp 1569139307
transform 1 0 4296 0 1 840
box -8 -8 8 8
use VIA1  VIA1_163
timestamp 1569139307
transform 1 0 4296 0 1 776
box -8 -8 8 8
use VIA1  VIA1_164
timestamp 1569139307
transform 1 0 4232 0 1 904
box -8 -8 8 8
use VIA1  VIA1_165
timestamp 1569139307
transform 1 0 4296 0 1 712
box -8 -8 8 8
use VIA1  VIA1_166
timestamp 1569139307
transform 1 0 4104 0 1 840
box -8 -8 8 8
use VIA1  VIA1_167
timestamp 1569139307
transform 1 0 4296 0 1 904
box -8 -8 8 8
use VIA1  VIA1_168
timestamp 1569139307
transform 1 0 4104 0 1 904
box -8 -8 8 8
use VIA1  VIA1_169
timestamp 1569139307
transform 1 0 3976 0 1 840
box -8 -8 8 8
use VIA1  VIA1_170
timestamp 1569139307
transform 1 0 3976 0 1 904
box -8 -8 8 8
use VIA1  VIA1_171
timestamp 1569139307
transform 1 0 3912 0 1 776
box -8 -8 8 8
use VIA1  VIA1_172
timestamp 1569139307
transform 1 0 4040 0 1 904
box -8 -8 8 8
use VIA1  VIA1_173
timestamp 1569139307
transform 1 0 3848 0 1 776
box -8 -8 8 8
use VIA1  VIA1_174
timestamp 1569139307
transform 1 0 3848 0 1 904
box -8 -8 8 8
use VIA1  VIA1_175
timestamp 1569139307
transform 1 0 3784 0 1 840
box -8 -8 8 8
use VIA1  VIA1_176
timestamp 1569139307
transform 1 0 3784 0 1 712
box -8 -8 8 8
use VIA1  VIA1_177
timestamp 1569139307
transform 1 0 3912 0 1 904
box -8 -8 8 8
use VIA1  VIA1_178
timestamp 1569139307
transform 1 0 3848 0 1 840
box -8 -8 8 8
use VIA1  VIA1_179
timestamp 1569139307
transform 1 0 4040 0 1 712
box -8 -8 8 8
use VIA1  VIA1_180
timestamp 1569139307
transform 1 0 3784 0 1 776
box -8 -8 8 8
use VIA1  VIA1_181
timestamp 1569139307
transform 1 0 3912 0 1 840
box -8 -8 8 8
use VIA1  VIA1_182
timestamp 1569139307
transform 1 0 3976 0 1 712
box -8 -8 8 8
use VIA1  VIA1_183
timestamp 1569139307
transform 1 0 3912 0 1 712
box -8 -8 8 8
use VIA1  VIA1_184
timestamp 1569139307
transform 1 0 3976 0 1 776
box -8 -8 8 8
use VIA1  VIA1_185
timestamp 1569139307
transform 1 0 4040 0 1 840
box -8 -8 8 8
use VIA1  VIA1_186
timestamp 1569139307
transform 1 0 3784 0 1 904
box -8 -8 8 8
use VIA1  VIA1_187
timestamp 1569139307
transform 1 0 4040 0 1 776
box -8 -8 8 8
use VIA1  VIA1_188
timestamp 1569139307
transform 1 0 3848 0 1 712
box -8 -8 8 8
use VIA1  VIA1_189
timestamp 1569139307
transform 1 0 3848 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_190
timestamp 1569139307
transform 1 0 4040 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_191
timestamp 1569139307
transform 1 0 3848 0 1 968
box -8 -8 8 8
use VIA1  VIA1_192
timestamp 1569139307
transform 1 0 3784 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_193
timestamp 1569139307
transform 1 0 4040 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_194
timestamp 1569139307
transform 1 0 4040 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_195
timestamp 1569139307
transform 1 0 3848 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_196
timestamp 1569139307
transform 1 0 3976 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_197
timestamp 1569139307
transform 1 0 3848 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_198
timestamp 1569139307
transform 1 0 3976 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_199
timestamp 1569139307
transform 1 0 3784 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_200
timestamp 1569139307
transform 1 0 3976 0 1 968
box -8 -8 8 8
use VIA1  VIA1_201
timestamp 1569139307
transform 1 0 3912 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_202
timestamp 1569139307
transform 1 0 3784 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_203
timestamp 1569139307
transform 1 0 3912 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_204
timestamp 1569139307
transform 1 0 3784 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_205
timestamp 1569139307
transform 1 0 3912 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_206
timestamp 1569139307
transform 1 0 4040 0 1 968
box -8 -8 8 8
use VIA1  VIA1_207
timestamp 1569139307
transform 1 0 3976 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_208
timestamp 1569139307
transform 1 0 3912 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_209
timestamp 1569139307
transform 1 0 3784 0 1 968
box -8 -8 8 8
use VIA1  VIA1_210
timestamp 1569139307
transform 1 0 3848 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_211
timestamp 1569139307
transform 1 0 4040 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_212
timestamp 1569139307
transform 1 0 3976 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_213
timestamp 1569139307
transform 1 0 3912 0 1 968
box -8 -8 8 8
use VIA1  VIA1_214
timestamp 1569139307
transform 1 0 4104 0 1 968
box -8 -8 8 8
use VIA1  VIA1_215
timestamp 1569139307
transform 1 0 4104 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_216
timestamp 1569139307
transform 1 0 4296 0 1 968
box -8 -8 8 8
use VIA1  VIA1_217
timestamp 1569139307
transform 1 0 4104 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_218
timestamp 1569139307
transform 1 0 4104 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_219
timestamp 1569139307
transform 1 0 4104 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_220
timestamp 1569139307
transform 1 0 4296 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_221
timestamp 1569139307
transform 1 0 4296 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_222
timestamp 1569139307
transform 1 0 4168 0 1 968
box -8 -8 8 8
use VIA1  VIA1_223
timestamp 1569139307
transform 1 0 4296 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_224
timestamp 1569139307
transform 1 0 4168 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_225
timestamp 1569139307
transform 1 0 4168 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_226
timestamp 1569139307
transform 1 0 4168 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_227
timestamp 1569139307
transform 1 0 4168 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_228
timestamp 1569139307
transform 1 0 4296 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_229
timestamp 1569139307
transform 1 0 4232 0 1 968
box -8 -8 8 8
use VIA1  VIA1_230
timestamp 1569139307
transform 1 0 4232 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_231
timestamp 1569139307
transform 1 0 4232 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_232
timestamp 1569139307
transform 1 0 4232 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_233
timestamp 1569139307
transform 1 0 4232 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_234
timestamp 1569139307
transform 1 0 4680 0 1 776
box -8 -8 8 8
use VIA1  VIA1_235
timestamp 1569139307
transform 1 0 4744 0 1 712
box -8 -8 8 8
use VIA1  VIA1_236
timestamp 1569139307
transform 1 0 4808 0 1 840
box -8 -8 8 8
use VIA1  VIA1_237
timestamp 1569139307
transform 1 0 4808 0 1 904
box -8 -8 8 8
use VIA1  VIA1_238
timestamp 1569139307
transform 1 0 4808 0 1 712
box -8 -8 8 8
use VIA1  VIA1_239
timestamp 1569139307
transform 1 0 4744 0 1 776
box -8 -8 8 8
use VIA1  VIA1_240
timestamp 1569139307
transform 1 0 4872 0 1 712
box -8 -8 8 8
use VIA1  VIA1_241
timestamp 1569139307
transform 1 0 4680 0 1 904
box -8 -8 8 8
use VIA1  VIA1_242
timestamp 1569139307
transform 1 0 4744 0 1 840
box -8 -8 8 8
use VIA1  VIA1_243
timestamp 1569139307
transform 1 0 4744 0 1 904
box -8 -8 8 8
use VIA1  VIA1_244
timestamp 1569139307
transform 1 0 4872 0 1 776
box -8 -8 8 8
use VIA1  VIA1_245
timestamp 1569139307
transform 1 0 4808 0 1 776
box -8 -8 8 8
use VIA1  VIA1_246
timestamp 1569139307
transform 1 0 4680 0 1 712
box -8 -8 8 8
use VIA1  VIA1_247
timestamp 1569139307
transform 1 0 4872 0 1 840
box -8 -8 8 8
use VIA1  VIA1_248
timestamp 1569139307
transform 1 0 4872 0 1 904
box -8 -8 8 8
use VIA1  VIA1_249
timestamp 1569139307
transform 1 0 4680 0 1 840
box -8 -8 8 8
use VIA1  VIA1_250
timestamp 1569139307
transform 1 0 4616 0 1 776
box -8 -8 8 8
use VIA1  VIA1_251
timestamp 1569139307
transform 1 0 4488 0 1 840
box -8 -8 8 8
use VIA1  VIA1_252
timestamp 1569139307
transform 1 0 4552 0 1 904
box -8 -8 8 8
use VIA1  VIA1_253
timestamp 1569139307
transform 1 0 4424 0 1 776
box -8 -8 8 8
use VIA1  VIA1_254
timestamp 1569139307
transform 1 0 4424 0 1 840
box -8 -8 8 8
use VIA1  VIA1_255
timestamp 1569139307
transform 1 0 4424 0 1 712
box -8 -8 8 8
use VIA1  VIA1_256
timestamp 1569139307
transform 1 0 4488 0 1 904
box -8 -8 8 8
use VIA1  VIA1_257
timestamp 1569139307
transform 1 0 4616 0 1 840
box -8 -8 8 8
use VIA1  VIA1_258
timestamp 1569139307
transform 1 0 4616 0 1 712
box -8 -8 8 8
use VIA1  VIA1_259
timestamp 1569139307
transform 1 0 4552 0 1 712
box -8 -8 8 8
use VIA1  VIA1_260
timestamp 1569139307
transform 1 0 4616 0 1 904
box -8 -8 8 8
use VIA1  VIA1_261
timestamp 1569139307
transform 1 0 4488 0 1 776
box -8 -8 8 8
use VIA1  VIA1_262
timestamp 1569139307
transform 1 0 4552 0 1 776
box -8 -8 8 8
use VIA1  VIA1_263
timestamp 1569139307
transform 1 0 4424 0 1 904
box -8 -8 8 8
use VIA1  VIA1_264
timestamp 1569139307
transform 1 0 4552 0 1 840
box -8 -8 8 8
use VIA1  VIA1_265
timestamp 1569139307
transform 1 0 4488 0 1 712
box -8 -8 8 8
use VIA1  VIA1_266
timestamp 1569139307
transform 1 0 4488 0 1 968
box -8 -8 8 8
use VIA1  VIA1_267
timestamp 1569139307
transform 1 0 4488 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_268
timestamp 1569139307
transform 1 0 4488 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_269
timestamp 1569139307
transform 1 0 4552 0 1 968
box -8 -8 8 8
use VIA1  VIA1_270
timestamp 1569139307
transform 1 0 4424 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_271
timestamp 1569139307
transform 1 0 4424 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_272
timestamp 1569139307
transform 1 0 4616 0 1 968
box -8 -8 8 8
use VIA1  VIA1_273
timestamp 1569139307
transform 1 0 4424 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_274
timestamp 1569139307
transform 1 0 4488 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_275
timestamp 1569139307
transform 1 0 4616 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_276
timestamp 1569139307
transform 1 0 4488 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_277
timestamp 1569139307
transform 1 0 4424 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_278
timestamp 1569139307
transform 1 0 4616 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_279
timestamp 1569139307
transform 1 0 4552 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_280
timestamp 1569139307
transform 1 0 4552 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_281
timestamp 1569139307
transform 1 0 4552 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_282
timestamp 1569139307
transform 1 0 4424 0 1 968
box -8 -8 8 8
use VIA1  VIA1_283
timestamp 1569139307
transform 1 0 4552 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_284
timestamp 1569139307
transform 1 0 4616 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_285
timestamp 1569139307
transform 1 0 4616 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_286
timestamp 1569139307
transform 1 0 4680 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_287
timestamp 1569139307
transform 1 0 4680 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_288
timestamp 1569139307
transform 1 0 4680 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_289
timestamp 1569139307
transform 1 0 4680 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_290
timestamp 1569139307
transform 1 0 4744 0 1 968
box -8 -8 8 8
use VIA1  VIA1_291
timestamp 1569139307
transform 1 0 4744 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_292
timestamp 1569139307
transform 1 0 4744 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_293
timestamp 1569139307
transform 1 0 4744 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_294
timestamp 1569139307
transform 1 0 4744 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_295
timestamp 1569139307
transform 1 0 4808 0 1 968
box -8 -8 8 8
use VIA1  VIA1_296
timestamp 1569139307
transform 1 0 4808 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_297
timestamp 1569139307
transform 1 0 4808 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_298
timestamp 1569139307
transform 1 0 4808 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_299
timestamp 1569139307
transform 1 0 4808 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_300
timestamp 1569139307
transform 1 0 4872 0 1 968
box -8 -8 8 8
use VIA1  VIA1_301
timestamp 1569139307
transform 1 0 4872 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_302
timestamp 1569139307
transform 1 0 4872 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_303
timestamp 1569139307
transform 1 0 4872 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_304
timestamp 1569139307
transform 1 0 4872 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_305
timestamp 1569139307
transform 1 0 4680 0 1 968
box -8 -8 8 8
use VIA1  VIA1_306
timestamp 1569139307
transform 1 0 3976 0 1 648
box -8 -8 8 8
use VIA1  VIA1_307
timestamp 1569139307
transform 1 0 3784 0 1 648
box -8 -8 8 8
use VIA1  VIA1_308
timestamp 1569139307
transform 1 0 4424 0 1 648
box -8 -8 8 8
use VIA1  VIA1_309
timestamp 1569139307
transform 1 0 4616 0 1 648
box -8 -8 8 8
use VIA1  VIA1_310
timestamp 1569139307
transform 1 0 4360 0 1 776
box -8 -8 8 8
use VIA1  VIA1_311
timestamp 1569139307
transform 1 0 3848 0 1 648
box -8 -8 8 8
use VIA1  VIA1_312
timestamp 1569139307
transform 1 0 4488 0 1 648
box -8 -8 8 8
use VIA1  VIA1_313
timestamp 1569139307
transform 1 0 4104 0 1 648
box -8 -8 8 8
use VIA1  VIA1_314
timestamp 1569139307
transform 1 0 4744 0 1 648
box -8 -8 8 8
use VIA1  VIA1_315
timestamp 1569139307
transform 1 0 4360 0 1 72
box -8 -8 8 8
use VIA1  VIA1_316
timestamp 1569139307
transform 1 0 3912 0 1 648
box -8 -8 8 8
use VIA1  VIA1_317
timestamp 1569139307
transform 1 0 4552 0 1 648
box -8 -8 8 8
use VIA1  VIA1_318
timestamp 1569139307
transform 1 0 4232 0 1 648
box -8 -8 8 8
use VIA1  VIA1_319
timestamp 1569139307
transform 1 0 4872 0 1 648
box -8 -8 8 8
use VIA1  VIA1_320
timestamp 1569139307
transform 1 0 4360 0 1 840
box -8 -8 8 8
use VIA1  VIA1_321
timestamp 1569139307
transform 1 0 4040 0 1 648
box -8 -8 8 8
use VIA1  VIA1_322
timestamp 1569139307
transform 1 0 4680 0 1 648
box -8 -8 8 8
use VIA1  VIA1_323
timestamp 1569139307
transform 1 0 4360 0 1 904
box -8 -8 8 8
use VIA1  VIA1_324
timestamp 1569139307
transform 1 0 4296 0 1 648
box -8 -8 8 8
use VIA1  VIA1_325
timestamp 1569139307
transform 1 0 4360 0 1 968
box -8 -8 8 8
use VIA1  VIA1_326
timestamp 1569139307
transform 1 0 4360 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_327
timestamp 1569139307
transform 1 0 4360 0 1 136
box -8 -8 8 8
use VIA1  VIA1_328
timestamp 1569139307
transform 1 0 4360 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_329
timestamp 1569139307
transform 1 0 4360 0 1 200
box -8 -8 8 8
use VIA1  VIA1_330
timestamp 1569139307
transform 1 0 4360 0 1 264
box -8 -8 8 8
use VIA1  VIA1_331
timestamp 1569139307
transform 1 0 4360 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_332
timestamp 1569139307
transform 1 0 4360 0 1 328
box -8 -8 8 8
use VIA1  VIA1_333
timestamp 1569139307
transform 1 0 4360 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_334
timestamp 1569139307
transform 1 0 4360 0 1 392
box -8 -8 8 8
use VIA1  VIA1_335
timestamp 1569139307
transform 1 0 4360 0 1 456
box -8 -8 8 8
use VIA1  VIA1_336
timestamp 1569139307
transform 1 0 4168 0 1 648
box -8 -8 8 8
use VIA1  VIA1_337
timestamp 1569139307
transform 1 0 4360 0 1 520
box -8 -8 8 8
use VIA1  VIA1_338
timestamp 1569139307
transform 1 0 4360 0 1 584
box -8 -8 8 8
use VIA1  VIA1_339
timestamp 1569139307
transform 1 0 4808 0 1 648
box -8 -8 8 8
use VIA1  VIA1_340
timestamp 1569139307
transform 1 0 4360 0 1 648
box -8 -8 8 8
use VIA1  VIA1_341
timestamp 1569139307
transform 1 0 4360 0 1 712
box -8 -8 8 8
use VIA1  VIA1_342
timestamp 1569139307
transform 1 0 3592 0 1 328
box -8 -8 8 8
use VIA1  VIA1_343
timestamp 1569139307
transform 1 0 3656 0 1 200
box -8 -8 8 8
use VIA1  VIA1_344
timestamp 1569139307
transform 1 0 3592 0 1 200
box -8 -8 8 8
use VIA1  VIA1_345
timestamp 1569139307
transform 1 0 3592 0 1 72
box -8 -8 8 8
use VIA1  VIA1_346
timestamp 1569139307
transform 1 0 3464 0 1 200
box -8 -8 8 8
use VIA1  VIA1_347
timestamp 1569139307
transform 1 0 3592 0 1 136
box -8 -8 8 8
use VIA1  VIA1_348
timestamp 1569139307
transform 1 0 3656 0 1 136
box -8 -8 8 8
use VIA1  VIA1_349
timestamp 1569139307
transform 1 0 3720 0 1 200
box -8 -8 8 8
use VIA1  VIA1_350
timestamp 1569139307
transform 1 0 3656 0 1 328
box -8 -8 8 8
use VIA1  VIA1_351
timestamp 1569139307
transform 1 0 3720 0 1 72
box -8 -8 8 8
use VIA1  VIA1_352
timestamp 1569139307
transform 1 0 3720 0 1 136
box -8 -8 8 8
use VIA1  VIA1_353
timestamp 1569139307
transform 1 0 3656 0 1 264
box -8 -8 8 8
use VIA1  VIA1_354
timestamp 1569139307
transform 1 0 3592 0 1 264
box -8 -8 8 8
use VIA1  VIA1_355
timestamp 1569139307
transform 1 0 3528 0 1 72
box -8 -8 8 8
use VIA1  VIA1_356
timestamp 1569139307
transform 1 0 3528 0 1 264
box -8 -8 8 8
use VIA1  VIA1_357
timestamp 1569139307
transform 1 0 3464 0 1 136
box -8 -8 8 8
use VIA1  VIA1_358
timestamp 1569139307
transform 1 0 3720 0 1 264
box -8 -8 8 8
use VIA1  VIA1_359
timestamp 1569139307
transform 1 0 3528 0 1 200
box -8 -8 8 8
use VIA1  VIA1_360
timestamp 1569139307
transform 1 0 3464 0 1 72
box -8 -8 8 8
use VIA1  VIA1_361
timestamp 1569139307
transform 1 0 3464 0 1 264
box -8 -8 8 8
use VIA1  VIA1_362
timestamp 1569139307
transform 1 0 3528 0 1 136
box -8 -8 8 8
use VIA1  VIA1_363
timestamp 1569139307
transform 1 0 3656 0 1 72
box -8 -8 8 8
use VIA1  VIA1_364
timestamp 1569139307
transform 1 0 3720 0 1 328
box -8 -8 8 8
use VIA1  VIA1_365
timestamp 1569139307
transform 1 0 3464 0 1 328
box -8 -8 8 8
use VIA1  VIA1_366
timestamp 1569139307
transform 1 0 3528 0 1 328
box -8 -8 8 8
use VIA1  VIA1_367
timestamp 1569139307
transform 1 0 3400 0 1 264
box -8 -8 8 8
use VIA1  VIA1_368
timestamp 1569139307
transform 1 0 3336 0 1 328
box -8 -8 8 8
use VIA1  VIA1_369
timestamp 1569139307
transform 1 0 3336 0 1 72
box -8 -8 8 8
use VIA1  VIA1_370
timestamp 1569139307
transform 1 0 3272 0 1 200
box -8 -8 8 8
use VIA1  VIA1_371
timestamp 1569139307
transform 1 0 3400 0 1 136
box -8 -8 8 8
use VIA1  VIA1_372
timestamp 1569139307
transform 1 0 3400 0 1 328
box -8 -8 8 8
use VIA1  VIA1_373
timestamp 1569139307
transform 1 0 3144 0 1 136
box -8 -8 8 8
use VIA1  VIA1_374
timestamp 1569139307
transform 1 0 3144 0 1 200
box -8 -8 8 8
use VIA1  VIA1_375
timestamp 1569139307
transform 1 0 3272 0 1 328
box -8 -8 8 8
use VIA1  VIA1_376
timestamp 1569139307
transform 1 0 3336 0 1 200
box -8 -8 8 8
use VIA1  VIA1_377
timestamp 1569139307
transform 1 0 3144 0 1 264
box -8 -8 8 8
use VIA1  VIA1_378
timestamp 1569139307
transform 1 0 3144 0 1 328
box -8 -8 8 8
use VIA1  VIA1_379
timestamp 1569139307
transform 1 0 3144 0 1 72
box -8 -8 8 8
use VIA1  VIA1_380
timestamp 1569139307
transform 1 0 3272 0 1 72
box -8 -8 8 8
use VIA1  VIA1_381
timestamp 1569139307
transform 1 0 3272 0 1 264
box -8 -8 8 8
use VIA1  VIA1_382
timestamp 1569139307
transform 1 0 3400 0 1 72
box -8 -8 8 8
use VIA1  VIA1_383
timestamp 1569139307
transform 1 0 3208 0 1 136
box -8 -8 8 8
use VIA1  VIA1_384
timestamp 1569139307
transform 1 0 3336 0 1 136
box -8 -8 8 8
use VIA1  VIA1_385
timestamp 1569139307
transform 1 0 3208 0 1 200
box -8 -8 8 8
use VIA1  VIA1_386
timestamp 1569139307
transform 1 0 3208 0 1 264
box -8 -8 8 8
use VIA1  VIA1_387
timestamp 1569139307
transform 1 0 3336 0 1 264
box -8 -8 8 8
use VIA1  VIA1_388
timestamp 1569139307
transform 1 0 3400 0 1 200
box -8 -8 8 8
use VIA1  VIA1_389
timestamp 1569139307
transform 1 0 3208 0 1 72
box -8 -8 8 8
use VIA1  VIA1_390
timestamp 1569139307
transform 1 0 3208 0 1 328
box -8 -8 8 8
use VIA1  VIA1_391
timestamp 1569139307
transform 1 0 3272 0 1 136
box -8 -8 8 8
use VIA1  VIA1_392
timestamp 1569139307
transform 1 0 3336 0 1 584
box -8 -8 8 8
use VIA1  VIA1_393
timestamp 1569139307
transform 1 0 3272 0 1 584
box -8 -8 8 8
use VIA1  VIA1_394
timestamp 1569139307
transform 1 0 3272 0 1 392
box -8 -8 8 8
use VIA1  VIA1_395
timestamp 1569139307
transform 1 0 3208 0 1 392
box -8 -8 8 8
use VIA1  VIA1_396
timestamp 1569139307
transform 1 0 3272 0 1 520
box -8 -8 8 8
use VIA1  VIA1_397
timestamp 1569139307
transform 1 0 3336 0 1 456
box -8 -8 8 8
use VIA1  VIA1_398
timestamp 1569139307
transform 1 0 3144 0 1 392
box -8 -8 8 8
use VIA1  VIA1_399
timestamp 1569139307
transform 1 0 3208 0 1 456
box -8 -8 8 8
use VIA1  VIA1_400
timestamp 1569139307
transform 1 0 3208 0 1 520
box -8 -8 8 8
use VIA1  VIA1_401
timestamp 1569139307
transform 1 0 3400 0 1 584
box -8 -8 8 8
use VIA1  VIA1_402
timestamp 1569139307
transform 1 0 3208 0 1 584
box -8 -8 8 8
use VIA1  VIA1_403
timestamp 1569139307
transform 1 0 3272 0 1 456
box -8 -8 8 8
use VIA1  VIA1_404
timestamp 1569139307
transform 1 0 3400 0 1 456
box -8 -8 8 8
use VIA1  VIA1_405
timestamp 1569139307
transform 1 0 3144 0 1 456
box -8 -8 8 8
use VIA1  VIA1_406
timestamp 1569139307
transform 1 0 3144 0 1 520
box -8 -8 8 8
use VIA1  VIA1_407
timestamp 1569139307
transform 1 0 3336 0 1 392
box -8 -8 8 8
use VIA1  VIA1_408
timestamp 1569139307
transform 1 0 3400 0 1 392
box -8 -8 8 8
use VIA1  VIA1_409
timestamp 1569139307
transform 1 0 3336 0 1 520
box -8 -8 8 8
use VIA1  VIA1_410
timestamp 1569139307
transform 1 0 3400 0 1 520
box -8 -8 8 8
use VIA1  VIA1_411
timestamp 1569139307
transform 1 0 3144 0 1 584
box -8 -8 8 8
use VIA1  VIA1_412
timestamp 1569139307
transform 1 0 3656 0 1 392
box -8 -8 8 8
use VIA1  VIA1_413
timestamp 1569139307
transform 1 0 3720 0 1 456
box -8 -8 8 8
use VIA1  VIA1_414
timestamp 1569139307
transform 1 0 3656 0 1 584
box -8 -8 8 8
use VIA1  VIA1_415
timestamp 1569139307
transform 1 0 3656 0 1 520
box -8 -8 8 8
use VIA1  VIA1_416
timestamp 1569139307
transform 1 0 3656 0 1 456
box -8 -8 8 8
use VIA1  VIA1_417
timestamp 1569139307
transform 1 0 3464 0 1 456
box -8 -8 8 8
use VIA1  VIA1_418
timestamp 1569139307
transform 1 0 3464 0 1 584
box -8 -8 8 8
use VIA1  VIA1_419
timestamp 1569139307
transform 1 0 3528 0 1 392
box -8 -8 8 8
use VIA1  VIA1_420
timestamp 1569139307
transform 1 0 3592 0 1 392
box -8 -8 8 8
use VIA1  VIA1_421
timestamp 1569139307
transform 1 0 3528 0 1 584
box -8 -8 8 8
use VIA1  VIA1_422
timestamp 1569139307
transform 1 0 3464 0 1 392
box -8 -8 8 8
use VIA1  VIA1_423
timestamp 1569139307
transform 1 0 3592 0 1 456
box -8 -8 8 8
use VIA1  VIA1_424
timestamp 1569139307
transform 1 0 3528 0 1 456
box -8 -8 8 8
use VIA1  VIA1_425
timestamp 1569139307
transform 1 0 3528 0 1 520
box -8 -8 8 8
use VIA1  VIA1_426
timestamp 1569139307
transform 1 0 3592 0 1 520
box -8 -8 8 8
use VIA1  VIA1_427
timestamp 1569139307
transform 1 0 3720 0 1 584
box -8 -8 8 8
use VIA1  VIA1_428
timestamp 1569139307
transform 1 0 3720 0 1 392
box -8 -8 8 8
use VIA1  VIA1_429
timestamp 1569139307
transform 1 0 3592 0 1 584
box -8 -8 8 8
use VIA1  VIA1_430
timestamp 1569139307
transform 1 0 3464 0 1 520
box -8 -8 8 8
use VIA1  VIA1_431
timestamp 1569139307
transform 1 0 3720 0 1 520
box -8 -8 8 8
use VIA1  VIA1_432
timestamp 1569139307
transform 1 0 2824 0 1 264
box -8 -8 8 8
use VIA1  VIA1_433
timestamp 1569139307
transform 1 0 3016 0 1 328
box -8 -8 8 8
use VIA1  VIA1_434
timestamp 1569139307
transform 1 0 2888 0 1 72
box -8 -8 8 8
use VIA1  VIA1_435
timestamp 1569139307
transform 1 0 3080 0 1 200
box -8 -8 8 8
use VIA1  VIA1_436
timestamp 1569139307
transform 1 0 3016 0 1 72
box -8 -8 8 8
use VIA1  VIA1_437
timestamp 1569139307
transform 1 0 3016 0 1 200
box -8 -8 8 8
use VIA1  VIA1_438
timestamp 1569139307
transform 1 0 3080 0 1 136
box -8 -8 8 8
use VIA1  VIA1_439
timestamp 1569139307
transform 1 0 2888 0 1 200
box -8 -8 8 8
use VIA1  VIA1_440
timestamp 1569139307
transform 1 0 2952 0 1 200
box -8 -8 8 8
use VIA1  VIA1_441
timestamp 1569139307
transform 1 0 2888 0 1 136
box -8 -8 8 8
use VIA1  VIA1_442
timestamp 1569139307
transform 1 0 2824 0 1 328
box -8 -8 8 8
use VIA1  VIA1_443
timestamp 1569139307
transform 1 0 2888 0 1 264
box -8 -8 8 8
use VIA1  VIA1_444
timestamp 1569139307
transform 1 0 2952 0 1 264
box -8 -8 8 8
use VIA1  VIA1_445
timestamp 1569139307
transform 1 0 2952 0 1 328
box -8 -8 8 8
use VIA1  VIA1_446
timestamp 1569139307
transform 1 0 2888 0 1 328
box -8 -8 8 8
use VIA1  VIA1_447
timestamp 1569139307
transform 1 0 2824 0 1 136
box -8 -8 8 8
use VIA1  VIA1_448
timestamp 1569139307
transform 1 0 2824 0 1 200
box -8 -8 8 8
use VIA1  VIA1_449
timestamp 1569139307
transform 1 0 3080 0 1 328
box -8 -8 8 8
use VIA1  VIA1_450
timestamp 1569139307
transform 1 0 2824 0 1 72
box -8 -8 8 8
use VIA1  VIA1_451
timestamp 1569139307
transform 1 0 3016 0 1 136
box -8 -8 8 8
use VIA1  VIA1_452
timestamp 1569139307
transform 1 0 2952 0 1 72
box -8 -8 8 8
use VIA1  VIA1_453
timestamp 1569139307
transform 1 0 3080 0 1 264
box -8 -8 8 8
use VIA1  VIA1_454
timestamp 1569139307
transform 1 0 3080 0 1 72
box -8 -8 8 8
use VIA1  VIA1_455
timestamp 1569139307
transform 1 0 3016 0 1 264
box -8 -8 8 8
use VIA1  VIA1_456
timestamp 1569139307
transform 1 0 2952 0 1 136
box -8 -8 8 8
use VIA1  VIA1_457
timestamp 1569139307
transform 1 0 2760 0 1 328
box -8 -8 8 8
use VIA1  VIA1_458
timestamp 1569139307
transform 1 0 2632 0 1 264
box -8 -8 8 8
use VIA1  VIA1_459
timestamp 1569139307
transform 1 0 2568 0 1 200
box -8 -8 8 8
use VIA1  VIA1_460
timestamp 1569139307
transform 1 0 2568 0 1 72
box -8 -8 8 8
use VIA1  VIA1_461
timestamp 1569139307
transform 1 0 2632 0 1 136
box -8 -8 8 8
use VIA1  VIA1_462
timestamp 1569139307
transform 1 0 2760 0 1 200
box -8 -8 8 8
use VIA1  VIA1_463
timestamp 1569139307
transform 1 0 2696 0 1 200
box -8 -8 8 8
use VIA1  VIA1_464
timestamp 1569139307
transform 1 0 2696 0 1 72
box -8 -8 8 8
use VIA1  VIA1_465
timestamp 1569139307
transform 1 0 2696 0 1 328
box -8 -8 8 8
use VIA1  VIA1_466
timestamp 1569139307
transform 1 0 2760 0 1 264
box -8 -8 8 8
use VIA1  VIA1_467
timestamp 1569139307
transform 1 0 2696 0 1 264
box -8 -8 8 8
use VIA1  VIA1_468
timestamp 1569139307
transform 1 0 2760 0 1 136
box -8 -8 8 8
use VIA1  VIA1_469
timestamp 1569139307
transform 1 0 2632 0 1 328
box -8 -8 8 8
use VIA1  VIA1_470
timestamp 1569139307
transform 1 0 2568 0 1 264
box -8 -8 8 8
use VIA1  VIA1_471
timestamp 1569139307
transform 1 0 2696 0 1 136
box -8 -8 8 8
use VIA1  VIA1_472
timestamp 1569139307
transform 1 0 2632 0 1 72
box -8 -8 8 8
use VIA1  VIA1_473
timestamp 1569139307
transform 1 0 2632 0 1 200
box -8 -8 8 8
use VIA1  VIA1_474
timestamp 1569139307
transform 1 0 2760 0 1 72
box -8 -8 8 8
use VIA1  VIA1_475
timestamp 1569139307
transform 1 0 2568 0 1 328
box -8 -8 8 8
use VIA1  VIA1_476
timestamp 1569139307
transform 1 0 2568 0 1 136
box -8 -8 8 8
use VIA1  VIA1_477
timestamp 1569139307
transform 1 0 2696 0 1 456
box -8 -8 8 8
use VIA1  VIA1_478
timestamp 1569139307
transform 1 0 2760 0 1 392
box -8 -8 8 8
use VIA1  VIA1_479
timestamp 1569139307
transform 1 0 2568 0 1 392
box -8 -8 8 8
use VIA1  VIA1_480
timestamp 1569139307
transform 1 0 2568 0 1 456
box -8 -8 8 8
use VIA1  VIA1_481
timestamp 1569139307
transform 1 0 2632 0 1 584
box -8 -8 8 8
use VIA1  VIA1_482
timestamp 1569139307
transform 1 0 2568 0 1 520
box -8 -8 8 8
use VIA1  VIA1_483
timestamp 1569139307
transform 1 0 2568 0 1 584
box -8 -8 8 8
use VIA1  VIA1_484
timestamp 1569139307
transform 1 0 2696 0 1 520
box -8 -8 8 8
use VIA1  VIA1_485
timestamp 1569139307
transform 1 0 2632 0 1 392
box -8 -8 8 8
use VIA1  VIA1_486
timestamp 1569139307
transform 1 0 2696 0 1 584
box -8 -8 8 8
use VIA1  VIA1_487
timestamp 1569139307
transform 1 0 2760 0 1 456
box -8 -8 8 8
use VIA1  VIA1_488
timestamp 1569139307
transform 1 0 2632 0 1 456
box -8 -8 8 8
use VIA1  VIA1_489
timestamp 1569139307
transform 1 0 2760 0 1 584
box -8 -8 8 8
use VIA1  VIA1_490
timestamp 1569139307
transform 1 0 2696 0 1 392
box -8 -8 8 8
use VIA1  VIA1_491
timestamp 1569139307
transform 1 0 2760 0 1 520
box -8 -8 8 8
use VIA1  VIA1_492
timestamp 1569139307
transform 1 0 2632 0 1 520
box -8 -8 8 8
use VIA1  VIA1_493
timestamp 1569139307
transform 1 0 2888 0 1 584
box -8 -8 8 8
use VIA1  VIA1_494
timestamp 1569139307
transform 1 0 2824 0 1 392
box -8 -8 8 8
use VIA1  VIA1_495
timestamp 1569139307
transform 1 0 3016 0 1 392
box -8 -8 8 8
use VIA1  VIA1_496
timestamp 1569139307
transform 1 0 3016 0 1 456
box -8 -8 8 8
use VIA1  VIA1_497
timestamp 1569139307
transform 1 0 2824 0 1 456
box -8 -8 8 8
use VIA1  VIA1_498
timestamp 1569139307
transform 1 0 2952 0 1 392
box -8 -8 8 8
use VIA1  VIA1_499
timestamp 1569139307
transform 1 0 2952 0 1 456
box -8 -8 8 8
use VIA1  VIA1_500
timestamp 1569139307
transform 1 0 2824 0 1 520
box -8 -8 8 8
use VIA1  VIA1_501
timestamp 1569139307
transform 1 0 3016 0 1 520
box -8 -8 8 8
use VIA1  VIA1_502
timestamp 1569139307
transform 1 0 2952 0 1 520
box -8 -8 8 8
use VIA1  VIA1_503
timestamp 1569139307
transform 1 0 3080 0 1 456
box -8 -8 8 8
use VIA1  VIA1_504
timestamp 1569139307
transform 1 0 2952 0 1 584
box -8 -8 8 8
use VIA1  VIA1_505
timestamp 1569139307
transform 1 0 3016 0 1 584
box -8 -8 8 8
use VIA1  VIA1_506
timestamp 1569139307
transform 1 0 3080 0 1 520
box -8 -8 8 8
use VIA1  VIA1_507
timestamp 1569139307
transform 1 0 3080 0 1 584
box -8 -8 8 8
use VIA1  VIA1_508
timestamp 1569139307
transform 1 0 3080 0 1 392
box -8 -8 8 8
use VIA1  VIA1_509
timestamp 1569139307
transform 1 0 2888 0 1 392
box -8 -8 8 8
use VIA1  VIA1_510
timestamp 1569139307
transform 1 0 2824 0 1 584
box -8 -8 8 8
use VIA1  VIA1_511
timestamp 1569139307
transform 1 0 2888 0 1 456
box -8 -8 8 8
use VIA1  VIA1_512
timestamp 1569139307
transform 1 0 2888 0 1 520
box -8 -8 8 8
use VIA1  VIA1_513
timestamp 1569139307
transform 1 0 2888 0 1 712
box -8 -8 8 8
use VIA1  VIA1_514
timestamp 1569139307
transform 1 0 2888 0 1 776
box -8 -8 8 8
use VIA1  VIA1_515
timestamp 1569139307
transform 1 0 3016 0 1 840
box -8 -8 8 8
use VIA1  VIA1_516
timestamp 1569139307
transform 1 0 2952 0 1 840
box -8 -8 8 8
use VIA1  VIA1_517
timestamp 1569139307
transform 1 0 3080 0 1 840
box -8 -8 8 8
use VIA1  VIA1_518
timestamp 1569139307
transform 1 0 3080 0 1 712
box -8 -8 8 8
use VIA1  VIA1_519
timestamp 1569139307
transform 1 0 3080 0 1 904
box -8 -8 8 8
use VIA1  VIA1_520
timestamp 1569139307
transform 1 0 3080 0 1 776
box -8 -8 8 8
use VIA1  VIA1_521
timestamp 1569139307
transform 1 0 2952 0 1 904
box -8 -8 8 8
use VIA1  VIA1_522
timestamp 1569139307
transform 1 0 2824 0 1 840
box -8 -8 8 8
use VIA1  VIA1_523
timestamp 1569139307
transform 1 0 2824 0 1 776
box -8 -8 8 8
use VIA1  VIA1_524
timestamp 1569139307
transform 1 0 2824 0 1 904
box -8 -8 8 8
use VIA1  VIA1_525
timestamp 1569139307
transform 1 0 2952 0 1 776
box -8 -8 8 8
use VIA1  VIA1_526
timestamp 1569139307
transform 1 0 3016 0 1 776
box -8 -8 8 8
use VIA1  VIA1_527
timestamp 1569139307
transform 1 0 3016 0 1 904
box -8 -8 8 8
use VIA1  VIA1_528
timestamp 1569139307
transform 1 0 3016 0 1 712
box -8 -8 8 8
use VIA1  VIA1_529
timestamp 1569139307
transform 1 0 2888 0 1 840
box -8 -8 8 8
use VIA1  VIA1_530
timestamp 1569139307
transform 1 0 2824 0 1 712
box -8 -8 8 8
use VIA1  VIA1_531
timestamp 1569139307
transform 1 0 2888 0 1 904
box -8 -8 8 8
use VIA1  VIA1_532
timestamp 1569139307
transform 1 0 2952 0 1 712
box -8 -8 8 8
use VIA1  VIA1_533
timestamp 1569139307
transform 1 0 2568 0 1 840
box -8 -8 8 8
use VIA1  VIA1_534
timestamp 1569139307
transform 1 0 2696 0 1 776
box -8 -8 8 8
use VIA1  VIA1_535
timestamp 1569139307
transform 1 0 2632 0 1 840
box -8 -8 8 8
use VIA1  VIA1_536
timestamp 1569139307
transform 1 0 2760 0 1 904
box -8 -8 8 8
use VIA1  VIA1_537
timestamp 1569139307
transform 1 0 2760 0 1 776
box -8 -8 8 8
use VIA1  VIA1_538
timestamp 1569139307
transform 1 0 2696 0 1 904
box -8 -8 8 8
use VIA1  VIA1_539
timestamp 1569139307
transform 1 0 2632 0 1 904
box -8 -8 8 8
use VIA1  VIA1_540
timestamp 1569139307
transform 1 0 2568 0 1 712
box -8 -8 8 8
use VIA1  VIA1_541
timestamp 1569139307
transform 1 0 2696 0 1 840
box -8 -8 8 8
use VIA1  VIA1_542
timestamp 1569139307
transform 1 0 2568 0 1 776
box -8 -8 8 8
use VIA1  VIA1_543
timestamp 1569139307
transform 1 0 2632 0 1 712
box -8 -8 8 8
use VIA1  VIA1_544
timestamp 1569139307
transform 1 0 2760 0 1 840
box -8 -8 8 8
use VIA1  VIA1_545
timestamp 1569139307
transform 1 0 2632 0 1 776
box -8 -8 8 8
use VIA1  VIA1_546
timestamp 1569139307
transform 1 0 2696 0 1 712
box -8 -8 8 8
use VIA1  VIA1_547
timestamp 1569139307
transform 1 0 2568 0 1 904
box -8 -8 8 8
use VIA1  VIA1_548
timestamp 1569139307
transform 1 0 2760 0 1 712
box -8 -8 8 8
use VIA1  VIA1_549
timestamp 1569139307
transform 1 0 2760 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_550
timestamp 1569139307
transform 1 0 2632 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_551
timestamp 1569139307
transform 1 0 2760 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_552
timestamp 1569139307
transform 1 0 2760 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_553
timestamp 1569139307
transform 1 0 2696 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_554
timestamp 1569139307
transform 1 0 2696 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_555
timestamp 1569139307
transform 1 0 2568 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_556
timestamp 1569139307
transform 1 0 2632 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_557
timestamp 1569139307
transform 1 0 2632 0 1 968
box -8 -8 8 8
use VIA1  VIA1_558
timestamp 1569139307
transform 1 0 2760 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_559
timestamp 1569139307
transform 1 0 2568 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_560
timestamp 1569139307
transform 1 0 2696 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_561
timestamp 1569139307
transform 1 0 2568 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_562
timestamp 1569139307
transform 1 0 2696 0 1 968
box -8 -8 8 8
use VIA1  VIA1_563
timestamp 1569139307
transform 1 0 2568 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_564
timestamp 1569139307
transform 1 0 2632 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_565
timestamp 1569139307
transform 1 0 2696 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_566
timestamp 1569139307
transform 1 0 2568 0 1 968
box -8 -8 8 8
use VIA1  VIA1_567
timestamp 1569139307
transform 1 0 2760 0 1 968
box -8 -8 8 8
use VIA1  VIA1_568
timestamp 1569139307
transform 1 0 2632 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_569
timestamp 1569139307
transform 1 0 3080 0 1 968
box -8 -8 8 8
use VIA1  VIA1_570
timestamp 1569139307
transform 1 0 2824 0 1 968
box -8 -8 8 8
use VIA1  VIA1_571
timestamp 1569139307
transform 1 0 3080 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_572
timestamp 1569139307
transform 1 0 2824 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_573
timestamp 1569139307
transform 1 0 2824 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_574
timestamp 1569139307
transform 1 0 3080 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_575
timestamp 1569139307
transform 1 0 2824 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_576
timestamp 1569139307
transform 1 0 2824 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_577
timestamp 1569139307
transform 1 0 3080 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_578
timestamp 1569139307
transform 1 0 3080 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_579
timestamp 1569139307
transform 1 0 2888 0 1 968
box -8 -8 8 8
use VIA1  VIA1_580
timestamp 1569139307
transform 1 0 2888 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_581
timestamp 1569139307
transform 1 0 2888 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_582
timestamp 1569139307
transform 1 0 2888 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_583
timestamp 1569139307
transform 1 0 2888 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_584
timestamp 1569139307
transform 1 0 2952 0 1 968
box -8 -8 8 8
use VIA1  VIA1_585
timestamp 1569139307
transform 1 0 2952 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_586
timestamp 1569139307
transform 1 0 2952 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_587
timestamp 1569139307
transform 1 0 2952 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_588
timestamp 1569139307
transform 1 0 2952 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_589
timestamp 1569139307
transform 1 0 3016 0 1 968
box -8 -8 8 8
use VIA1  VIA1_590
timestamp 1569139307
transform 1 0 3016 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_591
timestamp 1569139307
transform 1 0 3016 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_592
timestamp 1569139307
transform 1 0 3016 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_593
timestamp 1569139307
transform 1 0 3016 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_594
timestamp 1569139307
transform 1 0 3656 0 1 840
box -8 -8 8 8
use VIA1  VIA1_595
timestamp 1569139307
transform 1 0 3592 0 1 840
box -8 -8 8 8
use VIA1  VIA1_596
timestamp 1569139307
transform 1 0 3592 0 1 904
box -8 -8 8 8
use VIA1  VIA1_597
timestamp 1569139307
transform 1 0 3720 0 1 712
box -8 -8 8 8
use VIA1  VIA1_598
timestamp 1569139307
transform 1 0 3528 0 1 776
box -8 -8 8 8
use VIA1  VIA1_599
timestamp 1569139307
transform 1 0 3720 0 1 776
box -8 -8 8 8
use VIA1  VIA1_600
timestamp 1569139307
transform 1 0 3464 0 1 840
box -8 -8 8 8
use VIA1  VIA1_601
timestamp 1569139307
transform 1 0 3464 0 1 904
box -8 -8 8 8
use VIA1  VIA1_602
timestamp 1569139307
transform 1 0 3720 0 1 840
box -8 -8 8 8
use VIA1  VIA1_603
timestamp 1569139307
transform 1 0 3656 0 1 904
box -8 -8 8 8
use VIA1  VIA1_604
timestamp 1569139307
transform 1 0 3720 0 1 904
box -8 -8 8 8
use VIA1  VIA1_605
timestamp 1569139307
transform 1 0 3656 0 1 712
box -8 -8 8 8
use VIA1  VIA1_606
timestamp 1569139307
transform 1 0 3592 0 1 712
box -8 -8 8 8
use VIA1  VIA1_607
timestamp 1569139307
transform 1 0 3464 0 1 776
box -8 -8 8 8
use VIA1  VIA1_608
timestamp 1569139307
transform 1 0 3528 0 1 840
box -8 -8 8 8
use VIA1  VIA1_609
timestamp 1569139307
transform 1 0 3528 0 1 904
box -8 -8 8 8
use VIA1  VIA1_610
timestamp 1569139307
transform 1 0 3656 0 1 776
box -8 -8 8 8
use VIA1  VIA1_611
timestamp 1569139307
transform 1 0 3464 0 1 712
box -8 -8 8 8
use VIA1  VIA1_612
timestamp 1569139307
transform 1 0 3528 0 1 712
box -8 -8 8 8
use VIA1  VIA1_613
timestamp 1569139307
transform 1 0 3592 0 1 776
box -8 -8 8 8
use VIA1  VIA1_614
timestamp 1569139307
transform 1 0 3272 0 1 840
box -8 -8 8 8
use VIA1  VIA1_615
timestamp 1569139307
transform 1 0 3336 0 1 712
box -8 -8 8 8
use VIA1  VIA1_616
timestamp 1569139307
transform 1 0 3400 0 1 904
box -8 -8 8 8
use VIA1  VIA1_617
timestamp 1569139307
transform 1 0 3400 0 1 840
box -8 -8 8 8
use VIA1  VIA1_618
timestamp 1569139307
transform 1 0 3336 0 1 904
box -8 -8 8 8
use VIA1  VIA1_619
timestamp 1569139307
transform 1 0 3208 0 1 904
box -8 -8 8 8
use VIA1  VIA1_620
timestamp 1569139307
transform 1 0 3144 0 1 712
box -8 -8 8 8
use VIA1  VIA1_621
timestamp 1569139307
transform 1 0 3144 0 1 776
box -8 -8 8 8
use VIA1  VIA1_622
timestamp 1569139307
transform 1 0 3272 0 1 712
box -8 -8 8 8
use VIA1  VIA1_623
timestamp 1569139307
transform 1 0 3400 0 1 712
box -8 -8 8 8
use VIA1  VIA1_624
timestamp 1569139307
transform 1 0 3144 0 1 840
box -8 -8 8 8
use VIA1  VIA1_625
timestamp 1569139307
transform 1 0 3208 0 1 712
box -8 -8 8 8
use VIA1  VIA1_626
timestamp 1569139307
transform 1 0 3144 0 1 904
box -8 -8 8 8
use VIA1  VIA1_627
timestamp 1569139307
transform 1 0 3208 0 1 776
box -8 -8 8 8
use VIA1  VIA1_628
timestamp 1569139307
transform 1 0 3272 0 1 776
box -8 -8 8 8
use VIA1  VIA1_629
timestamp 1569139307
transform 1 0 3208 0 1 840
box -8 -8 8 8
use VIA1  VIA1_630
timestamp 1569139307
transform 1 0 3400 0 1 776
box -8 -8 8 8
use VIA1  VIA1_631
timestamp 1569139307
transform 1 0 3336 0 1 840
box -8 -8 8 8
use VIA1  VIA1_632
timestamp 1569139307
transform 1 0 3272 0 1 904
box -8 -8 8 8
use VIA1  VIA1_633
timestamp 1569139307
transform 1 0 3336 0 1 776
box -8 -8 8 8
use VIA1  VIA1_634
timestamp 1569139307
transform 1 0 3400 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_635
timestamp 1569139307
transform 1 0 3400 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_636
timestamp 1569139307
transform 1 0 3400 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_637
timestamp 1569139307
transform 1 0 3208 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_638
timestamp 1569139307
transform 1 0 3208 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_639
timestamp 1569139307
transform 1 0 3208 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_640
timestamp 1569139307
transform 1 0 3272 0 1 968
box -8 -8 8 8
use VIA1  VIA1_641
timestamp 1569139307
transform 1 0 3336 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_642
timestamp 1569139307
transform 1 0 3272 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_643
timestamp 1569139307
transform 1 0 3144 0 1 968
box -8 -8 8 8
use VIA1  VIA1_644
timestamp 1569139307
transform 1 0 3144 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_645
timestamp 1569139307
transform 1 0 3144 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_646
timestamp 1569139307
transform 1 0 3144 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_647
timestamp 1569139307
transform 1 0 3272 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_648
timestamp 1569139307
transform 1 0 3208 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_649
timestamp 1569139307
transform 1 0 3144 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_650
timestamp 1569139307
transform 1 0 3272 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_651
timestamp 1569139307
transform 1 0 3336 0 1 968
box -8 -8 8 8
use VIA1  VIA1_652
timestamp 1569139307
transform 1 0 3336 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_653
timestamp 1569139307
transform 1 0 3336 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_654
timestamp 1569139307
transform 1 0 3272 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_655
timestamp 1569139307
transform 1 0 3400 0 1 968
box -8 -8 8 8
use VIA1  VIA1_656
timestamp 1569139307
transform 1 0 3336 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_657
timestamp 1569139307
transform 1 0 3208 0 1 968
box -8 -8 8 8
use VIA1  VIA1_658
timestamp 1569139307
transform 1 0 3400 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_659
timestamp 1569139307
transform 1 0 3464 0 1 968
box -8 -8 8 8
use VIA1  VIA1_660
timestamp 1569139307
transform 1 0 3464 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_661
timestamp 1569139307
transform 1 0 3464 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_662
timestamp 1569139307
transform 1 0 3464 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_663
timestamp 1569139307
transform 1 0 3464 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_664
timestamp 1569139307
transform 1 0 3528 0 1 968
box -8 -8 8 8
use VIA1  VIA1_665
timestamp 1569139307
transform 1 0 3528 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_666
timestamp 1569139307
transform 1 0 3528 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_667
timestamp 1569139307
transform 1 0 3528 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_668
timestamp 1569139307
transform 1 0 3528 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_669
timestamp 1569139307
transform 1 0 3592 0 1 968
box -8 -8 8 8
use VIA1  VIA1_670
timestamp 1569139307
transform 1 0 3592 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_671
timestamp 1569139307
transform 1 0 3592 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_672
timestamp 1569139307
transform 1 0 3592 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_673
timestamp 1569139307
transform 1 0 3592 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_674
timestamp 1569139307
transform 1 0 3656 0 1 968
box -8 -8 8 8
use VIA1  VIA1_675
timestamp 1569139307
transform 1 0 3656 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_676
timestamp 1569139307
transform 1 0 3656 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_677
timestamp 1569139307
transform 1 0 3656 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_678
timestamp 1569139307
transform 1 0 3656 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_679
timestamp 1569139307
transform 1 0 3720 0 1 968
box -8 -8 8 8
use VIA1  VIA1_680
timestamp 1569139307
transform 1 0 3720 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_681
timestamp 1569139307
transform 1 0 3720 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_682
timestamp 1569139307
transform 1 0 3720 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_683
timestamp 1569139307
transform 1 0 3720 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_684
timestamp 1569139307
transform 1 0 3080 0 1 648
box -8 -8 8 8
use VIA1  VIA1_685
timestamp 1569139307
transform 1 0 3720 0 1 648
box -8 -8 8 8
use VIA1  VIA1_686
timestamp 1569139307
transform 1 0 3144 0 1 648
box -8 -8 8 8
use VIA1  VIA1_687
timestamp 1569139307
transform 1 0 2568 0 1 648
box -8 -8 8 8
use VIA1  VIA1_688
timestamp 1569139307
transform 1 0 3208 0 1 648
box -8 -8 8 8
use VIA1  VIA1_689
timestamp 1569139307
transform 1 0 2632 0 1 648
box -8 -8 8 8
use VIA1  VIA1_690
timestamp 1569139307
transform 1 0 3272 0 1 648
box -8 -8 8 8
use VIA1  VIA1_691
timestamp 1569139307
transform 1 0 2888 0 1 648
box -8 -8 8 8
use VIA1  VIA1_692
timestamp 1569139307
transform 1 0 3528 0 1 648
box -8 -8 8 8
use VIA1  VIA1_693
timestamp 1569139307
transform 1 0 2696 0 1 648
box -8 -8 8 8
use VIA1  VIA1_694
timestamp 1569139307
transform 1 0 3336 0 1 648
box -8 -8 8 8
use VIA1  VIA1_695
timestamp 1569139307
transform 1 0 2760 0 1 648
box -8 -8 8 8
use VIA1  VIA1_696
timestamp 1569139307
transform 1 0 3400 0 1 648
box -8 -8 8 8
use VIA1  VIA1_697
timestamp 1569139307
transform 1 0 2952 0 1 648
box -8 -8 8 8
use VIA1  VIA1_698
timestamp 1569139307
transform 1 0 3592 0 1 648
box -8 -8 8 8
use VIA1  VIA1_699
timestamp 1569139307
transform 1 0 3016 0 1 648
box -8 -8 8 8
use VIA1  VIA1_700
timestamp 1569139307
transform 1 0 3656 0 1 648
box -8 -8 8 8
use VIA1  VIA1_701
timestamp 1569139307
transform 1 0 2824 0 1 648
box -8 -8 8 8
use VIA1  VIA1_702
timestamp 1569139307
transform 1 0 3464 0 1 648
box -8 -8 8 8
use VIA1  VIA1_703
timestamp 1569139307
transform 1 0 3144 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_704
timestamp 1569139307
transform 1 0 3208 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_705
timestamp 1569139307
transform 1 0 3400 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_706
timestamp 1569139307
transform 1 0 3592 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_707
timestamp 1569139307
transform 1 0 3144 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_708
timestamp 1569139307
transform 1 0 3400 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_709
timestamp 1569139307
transform 1 0 3656 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_710
timestamp 1569139307
transform 1 0 3592 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_711
timestamp 1569139307
transform 1 0 3720 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_712
timestamp 1569139307
transform 1 0 3400 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_713
timestamp 1569139307
transform 1 0 3208 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_714
timestamp 1569139307
transform 1 0 3272 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_715
timestamp 1569139307
transform 1 0 3400 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_716
timestamp 1569139307
transform 1 0 3656 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_717
timestamp 1569139307
transform 1 0 3144 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_718
timestamp 1569139307
transform 1 0 3144 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_719
timestamp 1569139307
transform 1 0 3336 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_720
timestamp 1569139307
transform 1 0 3336 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_721
timestamp 1569139307
transform 1 0 3464 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_722
timestamp 1569139307
transform 1 0 3656 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_723
timestamp 1569139307
transform 1 0 3592 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_724
timestamp 1569139307
transform 1 0 3464 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_725
timestamp 1569139307
transform 1 0 3720 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_726
timestamp 1569139307
transform 1 0 3272 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_727
timestamp 1569139307
transform 1 0 3464 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_728
timestamp 1569139307
transform 1 0 3464 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_729
timestamp 1569139307
transform 1 0 3208 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_730
timestamp 1569139307
transform 1 0 3528 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_731
timestamp 1569139307
transform 1 0 3592 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_732
timestamp 1569139307
transform 1 0 3528 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_733
timestamp 1569139307
transform 1 0 3272 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_734
timestamp 1569139307
transform 1 0 3528 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_735
timestamp 1569139307
transform 1 0 3528 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_736
timestamp 1569139307
transform 1 0 3720 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_737
timestamp 1569139307
transform 1 0 3272 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_738
timestamp 1569139307
transform 1 0 3336 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_739
timestamp 1569139307
transform 1 0 3656 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_740
timestamp 1569139307
transform 1 0 3720 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_741
timestamp 1569139307
transform 1 0 3336 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_742
timestamp 1569139307
transform 1 0 3208 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_743
timestamp 1569139307
transform 1 0 2824 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_744
timestamp 1569139307
transform 1 0 3016 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_745
timestamp 1569139307
transform 1 0 2888 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_746
timestamp 1569139307
transform 1 0 2952 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_747
timestamp 1569139307
transform 1 0 2952 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_748
timestamp 1569139307
transform 1 0 2952 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_749
timestamp 1569139307
transform 1 0 3016 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_750
timestamp 1569139307
transform 1 0 2888 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_751
timestamp 1569139307
transform 1 0 3080 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_752
timestamp 1569139307
transform 1 0 3080 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_753
timestamp 1569139307
transform 1 0 3016 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_754
timestamp 1569139307
transform 1 0 2824 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_755
timestamp 1569139307
transform 1 0 2824 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_756
timestamp 1569139307
transform 1 0 2824 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_757
timestamp 1569139307
transform 1 0 2888 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_758
timestamp 1569139307
transform 1 0 3016 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_759
timestamp 1569139307
transform 1 0 2888 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_760
timestamp 1569139307
transform 1 0 2888 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_761
timestamp 1569139307
transform 1 0 3080 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_762
timestamp 1569139307
transform 1 0 3080 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_763
timestamp 1569139307
transform 1 0 2952 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_764
timestamp 1569139307
transform 1 0 2824 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_765
timestamp 1569139307
transform 1 0 2696 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_766
timestamp 1569139307
transform 1 0 2760 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_767
timestamp 1569139307
transform 1 0 2760 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_768
timestamp 1569139307
transform 1 0 2632 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_769
timestamp 1569139307
transform 1 0 2760 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_770
timestamp 1569139307
transform 1 0 2568 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_771
timestamp 1569139307
transform 1 0 2568 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_772
timestamp 1569139307
transform 1 0 2632 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_773
timestamp 1569139307
transform 1 0 2632 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_774
timestamp 1569139307
transform 1 0 2568 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_775
timestamp 1569139307
transform 1 0 2696 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_776
timestamp 1569139307
transform 1 0 2696 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_777
timestamp 1569139307
transform 1 0 2696 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_778
timestamp 1569139307
transform 1 0 2632 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_779
timestamp 1569139307
transform 1 0 2568 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_780
timestamp 1569139307
transform 1 0 2696 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_781
timestamp 1569139307
transform 1 0 2760 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_782
timestamp 1569139307
transform 1 0 2760 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_783
timestamp 1569139307
transform 1 0 2568 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_784
timestamp 1569139307
transform 1 0 2632 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_785
timestamp 1569139307
transform 1 0 2568 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_786
timestamp 1569139307
transform 1 0 2632 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_787
timestamp 1569139307
transform 1 0 2632 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_788
timestamp 1569139307
transform 1 0 2632 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_789
timestamp 1569139307
transform 1 0 2632 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_790
timestamp 1569139307
transform 1 0 2568 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_791
timestamp 1569139307
transform 1 0 2568 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_792
timestamp 1569139307
transform 1 0 2696 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_793
timestamp 1569139307
transform 1 0 2696 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_794
timestamp 1569139307
transform 1 0 2696 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_795
timestamp 1569139307
transform 1 0 2760 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_796
timestamp 1569139307
transform 1 0 2760 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_797
timestamp 1569139307
transform 1 0 2568 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_798
timestamp 1569139307
transform 1 0 2568 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_799
timestamp 1569139307
transform 1 0 2824 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_800
timestamp 1569139307
transform 1 0 3400 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_801
timestamp 1569139307
transform 1 0 3720 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_802
timestamp 1569139307
transform 1 0 3464 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_803
timestamp 1569139307
transform 1 0 3528 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_804
timestamp 1569139307
transform 1 0 3272 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_805
timestamp 1569139307
transform 1 0 3592 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_806
timestamp 1569139307
transform 1 0 3656 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_807
timestamp 1569139307
transform 1 0 3336 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_808
timestamp 1569139307
transform 1 0 3592 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_809
timestamp 1569139307
transform 1 0 3336 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_810
timestamp 1569139307
transform 1 0 3656 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_811
timestamp 1569139307
transform 1 0 3400 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_812
timestamp 1569139307
transform 1 0 3720 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_813
timestamp 1569139307
transform 1 0 3464 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_814
timestamp 1569139307
transform 1 0 3464 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_815
timestamp 1569139307
transform 1 0 3528 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_816
timestamp 1569139307
transform 1 0 3592 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_817
timestamp 1569139307
transform 1 0 3528 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_818
timestamp 1569139307
transform 1 0 3400 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_819
timestamp 1569139307
transform 1 0 3656 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_820
timestamp 1569139307
transform 1 0 3720 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_821
timestamp 1569139307
transform 1 0 4744 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_822
timestamp 1569139307
transform 1 0 4680 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_823
timestamp 1569139307
transform 1 0 4680 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_824
timestamp 1569139307
transform 1 0 4872 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_825
timestamp 1569139307
transform 1 0 4552 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_826
timestamp 1569139307
transform 1 0 4424 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_827
timestamp 1569139307
transform 1 0 4616 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_828
timestamp 1569139307
transform 1 0 4488 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_829
timestamp 1569139307
transform 1 0 4424 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_830
timestamp 1569139307
transform 1 0 4744 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_831
timestamp 1569139307
transform 1 0 4744 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_832
timestamp 1569139307
transform 1 0 4680 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_833
timestamp 1569139307
transform 1 0 4808 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_834
timestamp 1569139307
transform 1 0 4488 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_835
timestamp 1569139307
transform 1 0 4808 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_836
timestamp 1569139307
transform 1 0 4424 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_837
timestamp 1569139307
transform 1 0 4808 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_838
timestamp 1569139307
transform 1 0 4552 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_839
timestamp 1569139307
transform 1 0 4616 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_840
timestamp 1569139307
transform 1 0 4616 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_841
timestamp 1569139307
transform 1 0 4552 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_842
timestamp 1569139307
transform 1 0 4680 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_843
timestamp 1569139307
transform 1 0 4744 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_844
timestamp 1569139307
transform 1 0 4616 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_845
timestamp 1569139307
transform 1 0 4488 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_846
timestamp 1569139307
transform 1 0 4808 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_847
timestamp 1569139307
transform 1 0 4552 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_848
timestamp 1569139307
transform 1 0 4872 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_849
timestamp 1569139307
transform 1 0 4488 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_850
timestamp 1569139307
transform 1 0 4872 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_851
timestamp 1569139307
transform 1 0 4424 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_852
timestamp 1569139307
transform 1 0 4872 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_853
timestamp 1569139307
transform 1 0 3848 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_854
timestamp 1569139307
transform 1 0 4040 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_855
timestamp 1569139307
transform 1 0 4040 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_856
timestamp 1569139307
transform 1 0 4232 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_857
timestamp 1569139307
transform 1 0 4040 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_858
timestamp 1569139307
transform 1 0 4232 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_859
timestamp 1569139307
transform 1 0 4232 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_860
timestamp 1569139307
transform 1 0 3848 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_861
timestamp 1569139307
transform 1 0 3848 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_862
timestamp 1569139307
transform 1 0 4232 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_863
timestamp 1569139307
transform 1 0 4104 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_864
timestamp 1569139307
transform 1 0 4104 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_865
timestamp 1569139307
transform 1 0 4104 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_866
timestamp 1569139307
transform 1 0 4168 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_867
timestamp 1569139307
transform 1 0 4168 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_868
timestamp 1569139307
transform 1 0 4168 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_869
timestamp 1569139307
transform 1 0 3912 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_870
timestamp 1569139307
transform 1 0 3976 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_871
timestamp 1569139307
transform 1 0 4040 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_872
timestamp 1569139307
transform 1 0 4104 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_873
timestamp 1569139307
transform 1 0 4168 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_874
timestamp 1569139307
transform 1 0 4296 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_875
timestamp 1569139307
transform 1 0 4296 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_876
timestamp 1569139307
transform 1 0 4296 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_877
timestamp 1569139307
transform 1 0 4296 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_878
timestamp 1569139307
transform 1 0 3976 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_879
timestamp 1569139307
transform 1 0 3976 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_880
timestamp 1569139307
transform 1 0 3912 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_881
timestamp 1569139307
transform 1 0 3784 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_882
timestamp 1569139307
transform 1 0 3848 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_883
timestamp 1569139307
transform 1 0 3912 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_884
timestamp 1569139307
transform 1 0 3784 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_885
timestamp 1569139307
transform 1 0 3784 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_886
timestamp 1569139307
transform 1 0 3784 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_887
timestamp 1569139307
transform 1 0 3912 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_888
timestamp 1569139307
transform 1 0 3976 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_889
timestamp 1569139307
transform 1 0 4168 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_890
timestamp 1569139307
transform 1 0 3912 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_891
timestamp 1569139307
transform 1 0 4296 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_892
timestamp 1569139307
transform 1 0 4232 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_893
timestamp 1569139307
transform 1 0 3976 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_894
timestamp 1569139307
transform 1 0 3784 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_895
timestamp 1569139307
transform 1 0 4296 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_896
timestamp 1569139307
transform 1 0 4040 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_897
timestamp 1569139307
transform 1 0 3848 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_898
timestamp 1569139307
transform 1 0 4040 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_899
timestamp 1569139307
transform 1 0 4104 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_900
timestamp 1569139307
transform 1 0 3912 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_901
timestamp 1569139307
transform 1 0 3848 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_902
timestamp 1569139307
transform 1 0 4168 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_903
timestamp 1569139307
transform 1 0 3976 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_904
timestamp 1569139307
transform 1 0 4232 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_905
timestamp 1569139307
transform 1 0 4040 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_906
timestamp 1569139307
transform 1 0 3784 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_907
timestamp 1569139307
transform 1 0 4296 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_908
timestamp 1569139307
transform 1 0 4104 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_909
timestamp 1569139307
transform 1 0 3848 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_910
timestamp 1569139307
transform 1 0 4232 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_911
timestamp 1569139307
transform 1 0 3784 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_912
timestamp 1569139307
transform 1 0 4168 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_913
timestamp 1569139307
transform 1 0 3912 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_914
timestamp 1569139307
transform 1 0 3976 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_915
timestamp 1569139307
transform 1 0 4104 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_916
timestamp 1569139307
transform 1 0 4680 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_917
timestamp 1569139307
transform 1 0 4488 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_918
timestamp 1569139307
transform 1 0 4744 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_919
timestamp 1569139307
transform 1 0 4552 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_920
timestamp 1569139307
transform 1 0 4808 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_921
timestamp 1569139307
transform 1 0 4616 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_922
timestamp 1569139307
transform 1 0 4552 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_923
timestamp 1569139307
transform 1 0 4872 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_924
timestamp 1569139307
transform 1 0 4680 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_925
timestamp 1569139307
transform 1 0 4424 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_926
timestamp 1569139307
transform 1 0 4744 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_927
timestamp 1569139307
transform 1 0 4488 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_928
timestamp 1569139307
transform 1 0 4808 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_929
timestamp 1569139307
transform 1 0 4552 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_930
timestamp 1569139307
transform 1 0 4872 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_931
timestamp 1569139307
transform 1 0 4616 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_932
timestamp 1569139307
transform 1 0 4680 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_933
timestamp 1569139307
transform 1 0 4424 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_934
timestamp 1569139307
transform 1 0 4424 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_935
timestamp 1569139307
transform 1 0 4872 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_936
timestamp 1569139307
transform 1 0 4616 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_937
timestamp 1569139307
transform 1 0 4744 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_938
timestamp 1569139307
transform 1 0 4488 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_939
timestamp 1569139307
transform 1 0 4808 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_940
timestamp 1569139307
transform 1 0 4360 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_941
timestamp 1569139307
transform 1 0 4360 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_942
timestamp 1569139307
transform 1 0 4360 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_943
timestamp 1569139307
transform 1 0 4360 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_944
timestamp 1569139307
transform 1 0 4360 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_945
timestamp 1569139307
transform 1 0 4360 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_946
timestamp 1569139307
transform 1 0 4360 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_947
timestamp 1569139307
transform 1 0 2376 0 1 72
box -8 -8 8 8
use VIA1  VIA1_948
timestamp 1569139307
transform 1 0 2312 0 1 72
box -8 -8 8 8
use VIA1  VIA1_949
timestamp 1569139307
transform 1 0 2440 0 1 72
box -8 -8 8 8
use VIA1  VIA1_950
timestamp 1569139307
transform 1 0 2248 0 1 328
box -8 -8 8 8
use VIA1  VIA1_951
timestamp 1569139307
transform 1 0 2312 0 1 136
box -8 -8 8 8
use VIA1  VIA1_952
timestamp 1569139307
transform 1 0 2248 0 1 264
box -8 -8 8 8
use VIA1  VIA1_953
timestamp 1569139307
transform 1 0 2312 0 1 200
box -8 -8 8 8
use VIA1  VIA1_954
timestamp 1569139307
transform 1 0 2376 0 1 136
box -8 -8 8 8
use VIA1  VIA1_955
timestamp 1569139307
transform 1 0 2312 0 1 264
box -8 -8 8 8
use VIA1  VIA1_956
timestamp 1569139307
transform 1 0 2440 0 1 136
box -8 -8 8 8
use VIA1  VIA1_957
timestamp 1569139307
transform 1 0 2376 0 1 200
box -8 -8 8 8
use VIA1  VIA1_958
timestamp 1569139307
transform 1 0 2440 0 1 200
box -8 -8 8 8
use VIA1  VIA1_959
timestamp 1569139307
transform 1 0 2248 0 1 200
box -8 -8 8 8
use VIA1  VIA1_960
timestamp 1569139307
transform 1 0 2312 0 1 328
box -8 -8 8 8
use VIA1  VIA1_961
timestamp 1569139307
transform 1 0 2248 0 1 136
box -8 -8 8 8
use VIA1  VIA1_962
timestamp 1569139307
transform 1 0 2376 0 1 328
box -8 -8 8 8
use VIA1  VIA1_963
timestamp 1569139307
transform 1 0 2440 0 1 328
box -8 -8 8 8
use VIA1  VIA1_964
timestamp 1569139307
transform 1 0 2376 0 1 264
box -8 -8 8 8
use VIA1  VIA1_965
timestamp 1569139307
transform 1 0 2440 0 1 264
box -8 -8 8 8
use VIA1  VIA1_966
timestamp 1569139307
transform 1 0 2248 0 1 72
box -8 -8 8 8
use VIA1  VIA1_967
timestamp 1569139307
transform 1 0 2184 0 1 328
box -8 -8 8 8
use VIA1  VIA1_968
timestamp 1569139307
transform 1 0 2056 0 1 136
box -8 -8 8 8
use VIA1  VIA1_969
timestamp 1569139307
transform 1 0 1928 0 1 136
box -8 -8 8 8
use VIA1  VIA1_970
timestamp 1569139307
transform 1 0 2120 0 1 136
box -8 -8 8 8
use VIA1  VIA1_971
timestamp 1569139307
transform 1 0 2120 0 1 200
box -8 -8 8 8
use VIA1  VIA1_972
timestamp 1569139307
transform 1 0 2120 0 1 264
box -8 -8 8 8
use VIA1  VIA1_973
timestamp 1569139307
transform 1 0 1928 0 1 200
box -8 -8 8 8
use VIA1  VIA1_974
timestamp 1569139307
transform 1 0 2120 0 1 328
box -8 -8 8 8
use VIA1  VIA1_975
timestamp 1569139307
transform 1 0 1928 0 1 264
box -8 -8 8 8
use VIA1  VIA1_976
timestamp 1569139307
transform 1 0 1992 0 1 72
box -8 -8 8 8
use VIA1  VIA1_977
timestamp 1569139307
transform 1 0 2120 0 1 72
box -8 -8 8 8
use VIA1  VIA1_978
timestamp 1569139307
transform 1 0 1928 0 1 328
box -8 -8 8 8
use VIA1  VIA1_979
timestamp 1569139307
transform 1 0 1992 0 1 136
box -8 -8 8 8
use VIA1  VIA1_980
timestamp 1569139307
transform 1 0 1992 0 1 200
box -8 -8 8 8
use VIA1  VIA1_981
timestamp 1569139307
transform 1 0 2184 0 1 136
box -8 -8 8 8
use VIA1  VIA1_982
timestamp 1569139307
transform 1 0 1992 0 1 264
box -8 -8 8 8
use VIA1  VIA1_983
timestamp 1569139307
transform 1 0 2184 0 1 200
box -8 -8 8 8
use VIA1  VIA1_984
timestamp 1569139307
transform 1 0 1992 0 1 328
box -8 -8 8 8
use VIA1  VIA1_985
timestamp 1569139307
transform 1 0 1928 0 1 72
box -8 -8 8 8
use VIA1  VIA1_986
timestamp 1569139307
transform 1 0 2056 0 1 72
box -8 -8 8 8
use VIA1  VIA1_987
timestamp 1569139307
transform 1 0 2056 0 1 264
box -8 -8 8 8
use VIA1  VIA1_988
timestamp 1569139307
transform 1 0 2184 0 1 72
box -8 -8 8 8
use VIA1  VIA1_989
timestamp 1569139307
transform 1 0 2056 0 1 200
box -8 -8 8 8
use VIA1  VIA1_990
timestamp 1569139307
transform 1 0 2056 0 1 328
box -8 -8 8 8
use VIA1  VIA1_991
timestamp 1569139307
transform 1 0 2184 0 1 264
box -8 -8 8 8
use VIA1  VIA1_992
timestamp 1569139307
transform 1 0 1928 0 1 584
box -8 -8 8 8
use VIA1  VIA1_993
timestamp 1569139307
transform 1 0 2120 0 1 392
box -8 -8 8 8
use VIA1  VIA1_994
timestamp 1569139307
transform 1 0 2184 0 1 584
box -8 -8 8 8
use VIA1  VIA1_995
timestamp 1569139307
transform 1 0 2120 0 1 456
box -8 -8 8 8
use VIA1  VIA1_996
timestamp 1569139307
transform 1 0 2120 0 1 520
box -8 -8 8 8
use VIA1  VIA1_997
timestamp 1569139307
transform 1 0 1928 0 1 520
box -8 -8 8 8
use VIA1  VIA1_998
timestamp 1569139307
transform 1 0 2120 0 1 584
box -8 -8 8 8
use VIA1  VIA1_999
timestamp 1569139307
transform 1 0 2056 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1000
timestamp 1569139307
transform 1 0 1928 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1001
timestamp 1569139307
transform 1 0 2056 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1002
timestamp 1569139307
transform 1 0 1992 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1003
timestamp 1569139307
transform 1 0 1992 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1004
timestamp 1569139307
transform 1 0 1992 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1005
timestamp 1569139307
transform 1 0 1928 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1006
timestamp 1569139307
transform 1 0 2184 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1007
timestamp 1569139307
transform 1 0 1992 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1008
timestamp 1569139307
transform 1 0 2184 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1009
timestamp 1569139307
transform 1 0 2056 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1010
timestamp 1569139307
transform 1 0 2056 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1011
timestamp 1569139307
transform 1 0 2184 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1012
timestamp 1569139307
transform 1 0 2376 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1013
timestamp 1569139307
transform 1 0 2440 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1014
timestamp 1569139307
transform 1 0 2376 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1015
timestamp 1569139307
transform 1 0 2376 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1016
timestamp 1569139307
transform 1 0 2376 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1017
timestamp 1569139307
transform 1 0 2312 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1018
timestamp 1569139307
transform 1 0 2312 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1019
timestamp 1569139307
transform 1 0 2312 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1020
timestamp 1569139307
transform 1 0 2312 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1021
timestamp 1569139307
transform 1 0 2440 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1022
timestamp 1569139307
transform 1 0 2440 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1023
timestamp 1569139307
transform 1 0 2248 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1024
timestamp 1569139307
transform 1 0 2248 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1025
timestamp 1569139307
transform 1 0 2248 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1026
timestamp 1569139307
transform 1 0 2248 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1027
timestamp 1569139307
transform 1 0 2440 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1028
timestamp 1569139307
transform 1 0 1864 0 1 328
box -8 -8 8 8
use VIA1  VIA1_1029
timestamp 1569139307
transform 1 0 1864 0 1 136
box -8 -8 8 8
use VIA1  VIA1_1030
timestamp 1569139307
transform 1 0 1736 0 1 264
box -8 -8 8 8
use VIA1  VIA1_1031
timestamp 1569139307
transform 1 0 1736 0 1 72
box -8 -8 8 8
use VIA1  VIA1_1032
timestamp 1569139307
transform 1 0 1864 0 1 72
box -8 -8 8 8
use VIA1  VIA1_1033
timestamp 1569139307
transform 1 0 1800 0 1 72
box -8 -8 8 8
use VIA1  VIA1_1034
timestamp 1569139307
transform 1 0 1672 0 1 136
box -8 -8 8 8
use VIA1  VIA1_1035
timestamp 1569139307
transform 1 0 1672 0 1 200
box -8 -8 8 8
use VIA1  VIA1_1036
timestamp 1569139307
transform 1 0 1672 0 1 264
box -8 -8 8 8
use VIA1  VIA1_1037
timestamp 1569139307
transform 1 0 1672 0 1 328
box -8 -8 8 8
use VIA1  VIA1_1038
timestamp 1569139307
transform 1 0 1736 0 1 328
box -8 -8 8 8
use VIA1  VIA1_1039
timestamp 1569139307
transform 1 0 1800 0 1 136
box -8 -8 8 8
use VIA1  VIA1_1040
timestamp 1569139307
transform 1 0 1800 0 1 200
box -8 -8 8 8
use VIA1  VIA1_1041
timestamp 1569139307
transform 1 0 1864 0 1 264
box -8 -8 8 8
use VIA1  VIA1_1042
timestamp 1569139307
transform 1 0 1608 0 1 200
box -8 -8 8 8
use VIA1  VIA1_1043
timestamp 1569139307
transform 1 0 1608 0 1 264
box -8 -8 8 8
use VIA1  VIA1_1044
timestamp 1569139307
transform 1 0 1608 0 1 328
box -8 -8 8 8
use VIA1  VIA1_1045
timestamp 1569139307
transform 1 0 1736 0 1 136
box -8 -8 8 8
use VIA1  VIA1_1046
timestamp 1569139307
transform 1 0 1864 0 1 200
box -8 -8 8 8
use VIA1  VIA1_1047
timestamp 1569139307
transform 1 0 1800 0 1 264
box -8 -8 8 8
use VIA1  VIA1_1048
timestamp 1569139307
transform 1 0 1800 0 1 328
box -8 -8 8 8
use VIA1  VIA1_1049
timestamp 1569139307
transform 1 0 1736 0 1 200
box -8 -8 8 8
use VIA1  VIA1_1050
timestamp 1569139307
transform 1 0 1544 0 1 264
box -8 -8 8 8
use VIA1  VIA1_1051
timestamp 1569139307
transform 1 0 1544 0 1 328
box -8 -8 8 8
use VIA1  VIA1_1052
timestamp 1569139307
transform 1 0 1480 0 1 328
box -8 -8 8 8
use VIA1  VIA1_1053
timestamp 1569139307
transform 1 0 1544 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1054
timestamp 1569139307
transform 1 0 1544 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1055
timestamp 1569139307
transform 1 0 1544 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1056
timestamp 1569139307
transform 1 0 1544 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1057
timestamp 1569139307
transform 1 0 1288 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1058
timestamp 1569139307
transform 1 0 1416 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1059
timestamp 1569139307
transform 1 0 1416 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1060
timestamp 1569139307
transform 1 0 1416 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1061
timestamp 1569139307
transform 1 0 1416 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1062
timestamp 1569139307
transform 1 0 1480 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1063
timestamp 1569139307
transform 1 0 1480 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1064
timestamp 1569139307
transform 1 0 1480 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1065
timestamp 1569139307
transform 1 0 1352 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1066
timestamp 1569139307
transform 1 0 1352 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1067
timestamp 1569139307
transform 1 0 1352 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1068
timestamp 1569139307
transform 1 0 1480 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1069
timestamp 1569139307
transform 1 0 1288 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1070
timestamp 1569139307
transform 1 0 1736 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1071
timestamp 1569139307
transform 1 0 1608 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1072
timestamp 1569139307
transform 1 0 1608 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1073
timestamp 1569139307
transform 1 0 1608 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1074
timestamp 1569139307
transform 1 0 1608 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1075
timestamp 1569139307
transform 1 0 1800 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1076
timestamp 1569139307
transform 1 0 1736 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1077
timestamp 1569139307
transform 1 0 1800 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1078
timestamp 1569139307
transform 1 0 1736 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1079
timestamp 1569139307
transform 1 0 1736 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1080
timestamp 1569139307
transform 1 0 1672 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1081
timestamp 1569139307
transform 1 0 1672 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1082
timestamp 1569139307
transform 1 0 1672 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1083
timestamp 1569139307
transform 1 0 1672 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1084
timestamp 1569139307
transform 1 0 1864 0 1 392
box -8 -8 8 8
use VIA1  VIA1_1085
timestamp 1569139307
transform 1 0 1864 0 1 456
box -8 -8 8 8
use VIA1  VIA1_1086
timestamp 1569139307
transform 1 0 1864 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1087
timestamp 1569139307
transform 1 0 1800 0 1 520
box -8 -8 8 8
use VIA1  VIA1_1088
timestamp 1569139307
transform 1 0 1864 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1089
timestamp 1569139307
transform 1 0 1800 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1090
timestamp 1569139307
transform 1 0 1736 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1091
timestamp 1569139307
transform 1 0 1800 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1092
timestamp 1569139307
transform 1 0 1736 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1093
timestamp 1569139307
transform 1 0 1864 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1094
timestamp 1569139307
transform 1 0 1672 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1095
timestamp 1569139307
transform 1 0 1864 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1096
timestamp 1569139307
transform 1 0 1672 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1097
timestamp 1569139307
transform 1 0 1736 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1098
timestamp 1569139307
transform 1 0 1864 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1099
timestamp 1569139307
transform 1 0 1864 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1100
timestamp 1569139307
transform 1 0 1608 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1101
timestamp 1569139307
transform 1 0 1800 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1102
timestamp 1569139307
transform 1 0 1672 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1103
timestamp 1569139307
transform 1 0 1736 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1104
timestamp 1569139307
transform 1 0 1608 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1105
timestamp 1569139307
transform 1 0 1608 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1106
timestamp 1569139307
transform 1 0 1800 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1107
timestamp 1569139307
transform 1 0 1800 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1108
timestamp 1569139307
transform 1 0 1672 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1109
timestamp 1569139307
transform 1 0 1608 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1110
timestamp 1569139307
transform 1 0 1544 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1111
timestamp 1569139307
transform 1 0 1416 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1112
timestamp 1569139307
transform 1 0 1480 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1113
timestamp 1569139307
transform 1 0 1544 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1114
timestamp 1569139307
transform 1 0 1288 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1115
timestamp 1569139307
transform 1 0 1416 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1116
timestamp 1569139307
transform 1 0 1544 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1117
timestamp 1569139307
transform 1 0 1416 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1118
timestamp 1569139307
transform 1 0 1480 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1119
timestamp 1569139307
transform 1 0 1352 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1120
timestamp 1569139307
transform 1 0 1352 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1121
timestamp 1569139307
transform 1 0 1288 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1122
timestamp 1569139307
transform 1 0 1480 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1123
timestamp 1569139307
transform 1 0 1352 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1124
timestamp 1569139307
transform 1 0 1544 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1125
timestamp 1569139307
transform 1 0 1352 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1126
timestamp 1569139307
transform 1 0 1480 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1127
timestamp 1569139307
transform 1 0 1288 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1128
timestamp 1569139307
transform 1 0 1288 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1129
timestamp 1569139307
transform 1 0 1416 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1130
timestamp 1569139307
transform 1 0 1352 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1131
timestamp 1569139307
transform 1 0 1544 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1132
timestamp 1569139307
transform 1 0 1544 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1133
timestamp 1569139307
transform 1 0 1416 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1134
timestamp 1569139307
transform 1 0 1288 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1135
timestamp 1569139307
transform 1 0 1480 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1136
timestamp 1569139307
transform 1 0 1288 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1137
timestamp 1569139307
transform 1 0 1288 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1138
timestamp 1569139307
transform 1 0 1416 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1139
timestamp 1569139307
transform 1 0 1480 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1140
timestamp 1569139307
transform 1 0 1416 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1141
timestamp 1569139307
transform 1 0 1544 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1142
timestamp 1569139307
transform 1 0 1288 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1143
timestamp 1569139307
transform 1 0 1416 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1144
timestamp 1569139307
transform 1 0 1480 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1145
timestamp 1569139307
transform 1 0 1544 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1146
timestamp 1569139307
transform 1 0 1288 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1147
timestamp 1569139307
transform 1 0 1352 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1148
timestamp 1569139307
transform 1 0 1416 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1149
timestamp 1569139307
transform 1 0 1352 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1150
timestamp 1569139307
transform 1 0 1352 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1151
timestamp 1569139307
transform 1 0 1480 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1152
timestamp 1569139307
transform 1 0 1480 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1153
timestamp 1569139307
transform 1 0 1544 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1154
timestamp 1569139307
transform 1 0 1352 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1155
timestamp 1569139307
transform 1 0 1672 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1156
timestamp 1569139307
transform 1 0 1672 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1157
timestamp 1569139307
transform 1 0 1736 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1158
timestamp 1569139307
transform 1 0 1736 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1159
timestamp 1569139307
transform 1 0 1736 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1160
timestamp 1569139307
transform 1 0 1736 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1161
timestamp 1569139307
transform 1 0 1736 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1162
timestamp 1569139307
transform 1 0 1800 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1163
timestamp 1569139307
transform 1 0 1800 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1164
timestamp 1569139307
transform 1 0 1800 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1165
timestamp 1569139307
transform 1 0 1800 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1166
timestamp 1569139307
transform 1 0 1800 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1167
timestamp 1569139307
transform 1 0 1672 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1168
timestamp 1569139307
transform 1 0 1608 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1169
timestamp 1569139307
transform 1 0 1864 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1170
timestamp 1569139307
transform 1 0 1864 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1171
timestamp 1569139307
transform 1 0 1608 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1172
timestamp 1569139307
transform 1 0 1864 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1173
timestamp 1569139307
transform 1 0 1672 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1174
timestamp 1569139307
transform 1 0 1608 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1175
timestamp 1569139307
transform 1 0 1864 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1176
timestamp 1569139307
transform 1 0 1864 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1177
timestamp 1569139307
transform 1 0 1608 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1178
timestamp 1569139307
transform 1 0 1672 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1179
timestamp 1569139307
transform 1 0 1608 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1180
timestamp 1569139307
transform 1 0 2248 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1181
timestamp 1569139307
transform 1 0 2376 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1182
timestamp 1569139307
transform 1 0 2440 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1183
timestamp 1569139307
transform 1 0 2376 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1184
timestamp 1569139307
transform 1 0 2440 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1185
timestamp 1569139307
transform 1 0 2376 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1186
timestamp 1569139307
transform 1 0 2312 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1187
timestamp 1569139307
transform 1 0 2312 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1188
timestamp 1569139307
transform 1 0 2376 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1189
timestamp 1569139307
transform 1 0 2248 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1190
timestamp 1569139307
transform 1 0 2312 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1191
timestamp 1569139307
transform 1 0 2312 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1192
timestamp 1569139307
transform 1 0 2248 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1193
timestamp 1569139307
transform 1 0 2248 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1194
timestamp 1569139307
transform 1 0 2440 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1195
timestamp 1569139307
transform 1 0 2440 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1196
timestamp 1569139307
transform 1 0 1992 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1197
timestamp 1569139307
transform 1 0 1992 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1198
timestamp 1569139307
transform 1 0 2056 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1199
timestamp 1569139307
transform 1 0 2120 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1200
timestamp 1569139307
transform 1 0 2184 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1201
timestamp 1569139307
transform 1 0 2184 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1202
timestamp 1569139307
transform 1 0 1992 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1203
timestamp 1569139307
transform 1 0 1992 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1204
timestamp 1569139307
transform 1 0 1928 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1205
timestamp 1569139307
transform 1 0 1928 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1206
timestamp 1569139307
transform 1 0 2120 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1207
timestamp 1569139307
transform 1 0 2056 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1208
timestamp 1569139307
transform 1 0 2056 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1209
timestamp 1569139307
transform 1 0 2056 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1210
timestamp 1569139307
transform 1 0 1928 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1211
timestamp 1569139307
transform 1 0 1928 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1212
timestamp 1569139307
transform 1 0 2120 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1213
timestamp 1569139307
transform 1 0 2120 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1214
timestamp 1569139307
transform 1 0 2184 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1215
timestamp 1569139307
transform 1 0 2184 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1216
timestamp 1569139307
transform 1 0 1928 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1217
timestamp 1569139307
transform 1 0 2120 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1218
timestamp 1569139307
transform 1 0 1928 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1219
timestamp 1569139307
transform 1 0 2120 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1220
timestamp 1569139307
transform 1 0 2120 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1221
timestamp 1569139307
transform 1 0 2120 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1222
timestamp 1569139307
transform 1 0 2120 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1223
timestamp 1569139307
transform 1 0 2184 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1224
timestamp 1569139307
transform 1 0 2184 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1225
timestamp 1569139307
transform 1 0 2184 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1226
timestamp 1569139307
transform 1 0 1992 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1227
timestamp 1569139307
transform 1 0 1992 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1228
timestamp 1569139307
transform 1 0 1992 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1229
timestamp 1569139307
transform 1 0 1992 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1230
timestamp 1569139307
transform 1 0 1992 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1231
timestamp 1569139307
transform 1 0 2056 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1232
timestamp 1569139307
transform 1 0 2056 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1233
timestamp 1569139307
transform 1 0 2056 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1234
timestamp 1569139307
transform 1 0 2056 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1235
timestamp 1569139307
transform 1 0 2056 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1236
timestamp 1569139307
transform 1 0 2184 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1237
timestamp 1569139307
transform 1 0 2184 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1238
timestamp 1569139307
transform 1 0 1928 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1239
timestamp 1569139307
transform 1 0 1928 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1240
timestamp 1569139307
transform 1 0 1928 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1241
timestamp 1569139307
transform 1 0 2376 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1242
timestamp 1569139307
transform 1 0 2376 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1243
timestamp 1569139307
transform 1 0 2376 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1244
timestamp 1569139307
transform 1 0 2376 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1245
timestamp 1569139307
transform 1 0 2376 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1246
timestamp 1569139307
transform 1 0 2440 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1247
timestamp 1569139307
transform 1 0 2440 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1248
timestamp 1569139307
transform 1 0 2440 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1249
timestamp 1569139307
transform 1 0 2440 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1250
timestamp 1569139307
transform 1 0 2440 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1251
timestamp 1569139307
transform 1 0 2248 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1252
timestamp 1569139307
transform 1 0 2312 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1253
timestamp 1569139307
transform 1 0 2312 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1254
timestamp 1569139307
transform 1 0 2312 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1255
timestamp 1569139307
transform 1 0 2312 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1256
timestamp 1569139307
transform 1 0 2312 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1257
timestamp 1569139307
transform 1 0 2248 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1258
timestamp 1569139307
transform 1 0 2248 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1259
timestamp 1569139307
transform 1 0 2248 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1260
timestamp 1569139307
transform 1 0 2248 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1261
timestamp 1569139307
transform 1 0 1672 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1262
timestamp 1569139307
transform 1 0 2312 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1263
timestamp 1569139307
transform 1 0 1352 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1264
timestamp 1569139307
transform 1 0 1992 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1265
timestamp 1569139307
transform 1 0 1416 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1266
timestamp 1569139307
transform 1 0 2056 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1267
timestamp 1569139307
transform 1 0 1480 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1268
timestamp 1569139307
transform 1 0 2120 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1269
timestamp 1569139307
transform 1 0 1544 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1270
timestamp 1569139307
transform 1 0 2184 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1271
timestamp 1569139307
transform 1 0 1608 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1272
timestamp 1569139307
transform 1 0 2248 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1273
timestamp 1569139307
transform 1 0 1736 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1274
timestamp 1569139307
transform 1 0 2376 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1275
timestamp 1569139307
transform 1 0 1800 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1276
timestamp 1569139307
transform 1 0 2440 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1277
timestamp 1569139307
transform 1 0 1864 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1278
timestamp 1569139307
transform 1 0 1288 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1279
timestamp 1569139307
transform 1 0 1928 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1280
timestamp 1569139307
transform 1 0 1224 0 1 584
box -8 -8 8 8
use VIA1  VIA1_1281
timestamp 1569139307
transform 1 0 584 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1282
timestamp 1569139307
transform 1 0 968 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1283
timestamp 1569139307
transform 1 0 968 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1284
timestamp 1569139307
transform 1 0 1160 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1285
timestamp 1569139307
transform 1 0 1224 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1286
timestamp 1569139307
transform 1 0 1224 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1287
timestamp 1569139307
transform 1 0 1032 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1288
timestamp 1569139307
transform 1 0 1096 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1289
timestamp 1569139307
transform 1 0 1096 0 1 776
box -8 -8 8 8
use VIA1  VIA1_1290
timestamp 1569139307
transform 1 0 1032 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1291
timestamp 1569139307
transform 1 0 1032 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1292
timestamp 1569139307
transform 1 0 1096 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1293
timestamp 1569139307
transform 1 0 1096 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1294
timestamp 1569139307
transform 1 0 1224 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1295
timestamp 1569139307
transform 1 0 1160 0 1 712
box -8 -8 8 8
use VIA1  VIA1_1296
timestamp 1569139307
transform 1 0 1224 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1297
timestamp 1569139307
transform 1 0 1160 0 1 840
box -8 -8 8 8
use VIA1  VIA1_1298
timestamp 1569139307
transform 1 0 1160 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1299
timestamp 1569139307
transform 1 0 904 0 1 904
box -8 -8 8 8
use VIA1  VIA1_1300
timestamp 1569139307
transform 1 0 904 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1301
timestamp 1569139307
transform 1 0 904 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1302
timestamp 1569139307
transform 1 0 904 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1303
timestamp 1569139307
transform 1 0 904 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1304
timestamp 1569139307
transform 1 0 904 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1305
timestamp 1569139307
transform 1 0 840 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1306
timestamp 1569139307
transform 1 0 840 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1307
timestamp 1569139307
transform 1 0 840 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1308
timestamp 1569139307
transform 1 0 840 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1309
timestamp 1569139307
transform 1 0 840 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1310
timestamp 1569139307
transform 1 0 712 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1311
timestamp 1569139307
transform 1 0 712 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1312
timestamp 1569139307
transform 1 0 712 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1313
timestamp 1569139307
transform 1 0 776 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1314
timestamp 1569139307
transform 1 0 776 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1315
timestamp 1569139307
transform 1 0 776 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1316
timestamp 1569139307
transform 1 0 776 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1317
timestamp 1569139307
transform 1 0 1032 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1318
timestamp 1569139307
transform 1 0 1032 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1319
timestamp 1569139307
transform 1 0 1032 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1320
timestamp 1569139307
transform 1 0 1096 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1321
timestamp 1569139307
transform 1 0 1096 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1322
timestamp 1569139307
transform 1 0 1096 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1323
timestamp 1569139307
transform 1 0 1096 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1324
timestamp 1569139307
transform 1 0 1096 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1325
timestamp 1569139307
transform 1 0 1160 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1326
timestamp 1569139307
transform 1 0 1160 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1327
timestamp 1569139307
transform 1 0 1160 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1328
timestamp 1569139307
transform 1 0 1160 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1329
timestamp 1569139307
transform 1 0 1160 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1330
timestamp 1569139307
transform 1 0 968 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1331
timestamp 1569139307
transform 1 0 968 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1332
timestamp 1569139307
transform 1 0 968 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1333
timestamp 1569139307
transform 1 0 968 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1334
timestamp 1569139307
transform 1 0 968 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1335
timestamp 1569139307
transform 1 0 1224 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1336
timestamp 1569139307
transform 1 0 1224 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1337
timestamp 1569139307
transform 1 0 1224 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_1338
timestamp 1569139307
transform 1 0 1224 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1339
timestamp 1569139307
transform 1 0 1224 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1340
timestamp 1569139307
transform 1 0 1032 0 1 968
box -8 -8 8 8
use VIA1  VIA1_1341
timestamp 1569139307
transform 1 0 1032 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_1342
timestamp 1569139307
transform 1 0 648 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_1343
timestamp 1569139307
transform 1 0 648 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_1344
timestamp 1569139307
transform 1 0 1160 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1345
timestamp 1569139307
transform 1 0 1224 0 1 648
box -8 -8 8 8
use VIA1  VIA1_1346
timestamp 1569139307
transform 1 0 1160 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1347
timestamp 1569139307
transform 1 0 1096 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1348
timestamp 1569139307
transform 1 0 1160 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1349
timestamp 1569139307
transform 1 0 1096 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1350
timestamp 1569139307
transform 1 0 1032 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1351
timestamp 1569139307
transform 1 0 968 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1352
timestamp 1569139307
transform 1 0 1160 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1353
timestamp 1569139307
transform 1 0 1160 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1354
timestamp 1569139307
transform 1 0 1096 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1355
timestamp 1569139307
transform 1 0 968 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1356
timestamp 1569139307
transform 1 0 1096 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1357
timestamp 1569139307
transform 1 0 1096 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1358
timestamp 1569139307
transform 1 0 1032 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1359
timestamp 1569139307
transform 1 0 968 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1360
timestamp 1569139307
transform 1 0 1224 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1361
timestamp 1569139307
transform 1 0 1032 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1362
timestamp 1569139307
transform 1 0 968 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1363
timestamp 1569139307
transform 1 0 1224 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1364
timestamp 1569139307
transform 1 0 968 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1365
timestamp 1569139307
transform 1 0 1224 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1366
timestamp 1569139307
transform 1 0 1032 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1367
timestamp 1569139307
transform 1 0 1224 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1368
timestamp 1569139307
transform 1 0 1224 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1369
timestamp 1569139307
transform 1 0 1160 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1370
timestamp 1569139307
transform 1 0 1032 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1371
timestamp 1569139307
transform 1 0 776 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1372
timestamp 1569139307
transform 1 0 840 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1373
timestamp 1569139307
transform 1 0 904 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1374
timestamp 1569139307
transform 1 0 840 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1375
timestamp 1569139307
transform 1 0 712 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1376
timestamp 1569139307
transform 1 0 904 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1377
timestamp 1569139307
transform 1 0 776 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1378
timestamp 1569139307
transform 1 0 712 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1379
timestamp 1569139307
transform 1 0 904 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1380
timestamp 1569139307
transform 1 0 712 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1381
timestamp 1569139307
transform 1 0 840 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1382
timestamp 1569139307
transform 1 0 904 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1383
timestamp 1569139307
transform 1 0 712 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1384
timestamp 1569139307
transform 1 0 840 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1385
timestamp 1569139307
transform 1 0 904 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1386
timestamp 1569139307
transform 1 0 712 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1387
timestamp 1569139307
transform 1 0 840 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1388
timestamp 1569139307
transform 1 0 776 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1389
timestamp 1569139307
transform 1 0 776 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1390
timestamp 1569139307
transform 1 0 776 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1391
timestamp 1569139307
transform 1 0 776 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1392
timestamp 1569139307
transform 1 0 904 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1393
timestamp 1569139307
transform 1 0 776 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1394
timestamp 1569139307
transform 1 0 840 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1395
timestamp 1569139307
transform 1 0 904 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1396
timestamp 1569139307
transform 1 0 776 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1397
timestamp 1569139307
transform 1 0 840 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1398
timestamp 1569139307
transform 1 0 712 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1399
timestamp 1569139307
transform 1 0 840 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1400
timestamp 1569139307
transform 1 0 776 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1401
timestamp 1569139307
transform 1 0 712 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1402
timestamp 1569139307
transform 1 0 904 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1403
timestamp 1569139307
transform 1 0 840 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1404
timestamp 1569139307
transform 1 0 712 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1405
timestamp 1569139307
transform 1 0 904 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1406
timestamp 1569139307
transform 1 0 712 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1407
timestamp 1569139307
transform 1 0 840 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1408
timestamp 1569139307
transform 1 0 712 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1409
timestamp 1569139307
transform 1 0 776 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1410
timestamp 1569139307
transform 1 0 904 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1411
timestamp 1569139307
transform 1 0 1224 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1412
timestamp 1569139307
transform 1 0 1096 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1413
timestamp 1569139307
transform 1 0 1096 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1414
timestamp 1569139307
transform 1 0 1224 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1415
timestamp 1569139307
transform 1 0 1096 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1416
timestamp 1569139307
transform 1 0 1096 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1417
timestamp 1569139307
transform 1 0 1224 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1418
timestamp 1569139307
transform 1 0 1224 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1419
timestamp 1569139307
transform 1 0 1096 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1420
timestamp 1569139307
transform 1 0 1032 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1421
timestamp 1569139307
transform 1 0 1160 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1422
timestamp 1569139307
transform 1 0 968 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1423
timestamp 1569139307
transform 1 0 1032 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1424
timestamp 1569139307
transform 1 0 1160 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1425
timestamp 1569139307
transform 1 0 968 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1426
timestamp 1569139307
transform 1 0 1160 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1427
timestamp 1569139307
transform 1 0 1032 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1428
timestamp 1569139307
transform 1 0 1160 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1429
timestamp 1569139307
transform 1 0 968 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1430
timestamp 1569139307
transform 1 0 1160 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1431
timestamp 1569139307
transform 1 0 968 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1432
timestamp 1569139307
transform 1 0 1224 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1433
timestamp 1569139307
transform 1 0 968 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1434
timestamp 1569139307
transform 1 0 1032 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1435
timestamp 1569139307
transform 1 0 1032 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1436
timestamp 1569139307
transform 1 0 392 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1437
timestamp 1569139307
transform 1 0 584 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1438
timestamp 1569139307
transform 1 0 520 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1439
timestamp 1569139307
transform 1 0 520 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1440
timestamp 1569139307
transform 1 0 392 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1441
timestamp 1569139307
transform 1 0 456 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1442
timestamp 1569139307
transform 1 0 584 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1443
timestamp 1569139307
transform 1 0 520 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1444
timestamp 1569139307
transform 1 0 456 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1445
timestamp 1569139307
transform 1 0 520 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1446
timestamp 1569139307
transform 1 0 456 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1447
timestamp 1569139307
transform 1 0 584 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1448
timestamp 1569139307
transform 1 0 584 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1449
timestamp 1569139307
transform 1 0 584 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1450
timestamp 1569139307
transform 1 0 392 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1451
timestamp 1569139307
transform 1 0 456 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1452
timestamp 1569139307
transform 1 0 520 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1453
timestamp 1569139307
transform 1 0 328 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1454
timestamp 1569139307
transform 1 0 264 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1455
timestamp 1569139307
transform 1 0 328 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1456
timestamp 1569139307
transform 1 0 328 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1457
timestamp 1569139307
transform 1 0 200 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1458
timestamp 1569139307
transform 1 0 136 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1459
timestamp 1569139307
transform 1 0 264 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1460
timestamp 1569139307
transform 1 0 200 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1461
timestamp 1569139307
transform 1 0 72 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1462
timestamp 1569139307
transform 1 0 72 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1463
timestamp 1569139307
transform 1 0 200 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1464
timestamp 1569139307
transform 1 0 136 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1465
timestamp 1569139307
transform 1 0 328 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1466
timestamp 1569139307
transform 1 0 72 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1467
timestamp 1569139307
transform 1 0 200 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1468
timestamp 1569139307
transform 1 0 328 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1469
timestamp 1569139307
transform 1 0 264 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1470
timestamp 1569139307
transform 1 0 136 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1471
timestamp 1569139307
transform 1 0 264 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1472
timestamp 1569139307
transform 1 0 328 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1473
timestamp 1569139307
transform 1 0 328 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1474
timestamp 1569139307
transform 1 0 264 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1475
timestamp 1569139307
transform 1 0 136 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1476
timestamp 1569139307
transform 1 0 264 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1477
timestamp 1569139307
transform 1 0 200 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1478
timestamp 1569139307
transform 1 0 456 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1479
timestamp 1569139307
transform 1 0 584 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1480
timestamp 1569139307
transform 1 0 456 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1481
timestamp 1569139307
transform 1 0 456 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1482
timestamp 1569139307
transform 1 0 456 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1483
timestamp 1569139307
transform 1 0 584 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1484
timestamp 1569139307
transform 1 0 456 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1485
timestamp 1569139307
transform 1 0 392 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1486
timestamp 1569139307
transform 1 0 392 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1487
timestamp 1569139307
transform 1 0 520 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1488
timestamp 1569139307
transform 1 0 584 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1489
timestamp 1569139307
transform 1 0 520 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1490
timestamp 1569139307
transform 1 0 520 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1491
timestamp 1569139307
transform 1 0 392 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1492
timestamp 1569139307
transform 1 0 520 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1493
timestamp 1569139307
transform 1 0 520 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1494
timestamp 1569139307
transform 1 0 392 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1495
timestamp 1569139307
transform 1 0 584 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1496
timestamp 1569139307
transform 1 0 584 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1497
timestamp 1569139307
transform 1 0 392 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1498
timestamp 1569139307
transform 1 0 392 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1499
timestamp 1569139307
transform 1 0 392 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1500
timestamp 1569139307
transform 1 0 456 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1501
timestamp 1569139307
transform 1 0 520 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1502
timestamp 1569139307
transform 1 0 456 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1503
timestamp 1569139307
transform 1 0 520 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1504
timestamp 1569139307
transform 1 0 456 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1505
timestamp 1569139307
transform 1 0 456 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1506
timestamp 1569139307
transform 1 0 392 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1507
timestamp 1569139307
transform 1 0 584 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1508
timestamp 1569139307
transform 1 0 520 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1509
timestamp 1569139307
transform 1 0 584 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1510
timestamp 1569139307
transform 1 0 520 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1511
timestamp 1569139307
transform 1 0 584 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1512
timestamp 1569139307
transform 1 0 456 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1513
timestamp 1569139307
transform 1 0 392 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1514
timestamp 1569139307
transform 1 0 520 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1515
timestamp 1569139307
transform 1 0 584 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1516
timestamp 1569139307
transform 1 0 392 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1517
timestamp 1569139307
transform 1 0 584 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1518
timestamp 1569139307
transform 1 0 200 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1519
timestamp 1569139307
transform 1 0 200 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1520
timestamp 1569139307
transform 1 0 328 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1521
timestamp 1569139307
transform 1 0 72 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1522
timestamp 1569139307
transform 1 0 136 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1523
timestamp 1569139307
transform 1 0 72 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1524
timestamp 1569139307
transform 1 0 264 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1525
timestamp 1569139307
transform 1 0 200 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1526
timestamp 1569139307
transform 1 0 136 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1527
timestamp 1569139307
transform 1 0 328 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1528
timestamp 1569139307
transform 1 0 328 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1529
timestamp 1569139307
transform 1 0 136 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1530
timestamp 1569139307
transform 1 0 72 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1531
timestamp 1569139307
transform 1 0 136 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1532
timestamp 1569139307
transform 1 0 72 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1533
timestamp 1569139307
transform 1 0 328 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1534
timestamp 1569139307
transform 1 0 264 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1535
timestamp 1569139307
transform 1 0 264 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1536
timestamp 1569139307
transform 1 0 200 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1537
timestamp 1569139307
transform 1 0 72 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1538
timestamp 1569139307
transform 1 0 328 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1539
timestamp 1569139307
transform 1 0 200 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1540
timestamp 1569139307
transform 1 0 264 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1541
timestamp 1569139307
transform 1 0 264 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1542
timestamp 1569139307
transform 1 0 136 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1543
timestamp 1569139307
transform 1 0 136 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1544
timestamp 1569139307
transform 1 0 200 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1545
timestamp 1569139307
transform 1 0 264 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1546
timestamp 1569139307
transform 1 0 72 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1547
timestamp 1569139307
transform 1 0 136 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1548
timestamp 1569139307
transform 1 0 328 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1549
timestamp 1569139307
transform 1 0 264 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1550
timestamp 1569139307
transform 1 0 200 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1551
timestamp 1569139307
transform 1 0 328 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1552
timestamp 1569139307
transform 1 0 72 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1553
timestamp 1569139307
transform 1 0 328 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1554
timestamp 1569139307
transform 1 0 200 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1555
timestamp 1569139307
transform 1 0 136 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1556
timestamp 1569139307
transform 1 0 264 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1557
timestamp 1569139307
transform 1 0 328 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1558
timestamp 1569139307
transform 1 0 264 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1559
timestamp 1569139307
transform 1 0 72 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1560
timestamp 1569139307
transform 1 0 72 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1561
timestamp 1569139307
transform 1 0 136 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1562
timestamp 1569139307
transform 1 0 200 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1563
timestamp 1569139307
transform 1 0 392 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1564
timestamp 1569139307
transform 1 0 456 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1565
timestamp 1569139307
transform 1 0 456 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1566
timestamp 1569139307
transform 1 0 584 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1567
timestamp 1569139307
transform 1 0 456 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1568
timestamp 1569139307
transform 1 0 584 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1569
timestamp 1569139307
transform 1 0 520 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1570
timestamp 1569139307
transform 1 0 456 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1571
timestamp 1569139307
transform 1 0 584 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1572
timestamp 1569139307
transform 1 0 392 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1573
timestamp 1569139307
transform 1 0 584 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1574
timestamp 1569139307
transform 1 0 392 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1575
timestamp 1569139307
transform 1 0 520 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1576
timestamp 1569139307
transform 1 0 392 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1577
timestamp 1569139307
transform 1 0 520 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1578
timestamp 1569139307
transform 1 0 520 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1579
timestamp 1569139307
transform 1 0 968 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1580
timestamp 1569139307
transform 1 0 1096 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1581
timestamp 1569139307
transform 1 0 1096 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1582
timestamp 1569139307
transform 1 0 1096 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1583
timestamp 1569139307
transform 1 0 968 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1584
timestamp 1569139307
transform 1 0 1160 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1585
timestamp 1569139307
transform 1 0 1160 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1586
timestamp 1569139307
transform 1 0 1224 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1587
timestamp 1569139307
transform 1 0 1160 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1588
timestamp 1569139307
transform 1 0 1032 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1589
timestamp 1569139307
transform 1 0 968 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1590
timestamp 1569139307
transform 1 0 1096 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1591
timestamp 1569139307
transform 1 0 1032 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1592
timestamp 1569139307
transform 1 0 1160 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1593
timestamp 1569139307
transform 1 0 1032 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1594
timestamp 1569139307
transform 1 0 968 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1595
timestamp 1569139307
transform 1 0 1224 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1596
timestamp 1569139307
transform 1 0 1096 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1597
timestamp 1569139307
transform 1 0 1032 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1598
timestamp 1569139307
transform 1 0 1224 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1599
timestamp 1569139307
transform 1 0 1160 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1600
timestamp 1569139307
transform 1 0 1224 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1601
timestamp 1569139307
transform 1 0 1224 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1602
timestamp 1569139307
transform 1 0 968 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1603
timestamp 1569139307
transform 1 0 1032 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1604
timestamp 1569139307
transform 1 0 840 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1605
timestamp 1569139307
transform 1 0 776 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1606
timestamp 1569139307
transform 1 0 840 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1607
timestamp 1569139307
transform 1 0 776 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1608
timestamp 1569139307
transform 1 0 712 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1609
timestamp 1569139307
transform 1 0 712 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1610
timestamp 1569139307
transform 1 0 840 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1611
timestamp 1569139307
transform 1 0 712 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1612
timestamp 1569139307
transform 1 0 712 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1613
timestamp 1569139307
transform 1 0 904 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1614
timestamp 1569139307
transform 1 0 776 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1615
timestamp 1569139307
transform 1 0 712 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1616
timestamp 1569139307
transform 1 0 776 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1617
timestamp 1569139307
transform 1 0 904 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1618
timestamp 1569139307
transform 1 0 776 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1619
timestamp 1569139307
transform 1 0 840 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1620
timestamp 1569139307
transform 1 0 904 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1621
timestamp 1569139307
transform 1 0 904 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1622
timestamp 1569139307
transform 1 0 840 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1623
timestamp 1569139307
transform 1 0 904 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1624
timestamp 1569139307
transform 1 0 904 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1625
timestamp 1569139307
transform 1 0 776 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1626
timestamp 1569139307
transform 1 0 840 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1627
timestamp 1569139307
transform 1 0 840 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1628
timestamp 1569139307
transform 1 0 840 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1629
timestamp 1569139307
transform 1 0 776 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1630
timestamp 1569139307
transform 1 0 712 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1631
timestamp 1569139307
transform 1 0 904 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1632
timestamp 1569139307
transform 1 0 840 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1633
timestamp 1569139307
transform 1 0 776 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1634
timestamp 1569139307
transform 1 0 904 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1635
timestamp 1569139307
transform 1 0 712 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1636
timestamp 1569139307
transform 1 0 904 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1637
timestamp 1569139307
transform 1 0 712 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1638
timestamp 1569139307
transform 1 0 712 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1639
timestamp 1569139307
transform 1 0 776 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1640
timestamp 1569139307
transform 1 0 1224 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1641
timestamp 1569139307
transform 1 0 968 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1642
timestamp 1569139307
transform 1 0 1160 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1643
timestamp 1569139307
transform 1 0 1032 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1644
timestamp 1569139307
transform 1 0 1224 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1645
timestamp 1569139307
transform 1 0 968 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1646
timestamp 1569139307
transform 1 0 1096 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1647
timestamp 1569139307
transform 1 0 1032 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1648
timestamp 1569139307
transform 1 0 1096 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1649
timestamp 1569139307
transform 1 0 1032 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1650
timestamp 1569139307
transform 1 0 1032 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1651
timestamp 1569139307
transform 1 0 1096 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1652
timestamp 1569139307
transform 1 0 1096 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1653
timestamp 1569139307
transform 1 0 1160 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1654
timestamp 1569139307
transform 1 0 1160 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1655
timestamp 1569139307
transform 1 0 1160 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1656
timestamp 1569139307
transform 1 0 1224 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1657
timestamp 1569139307
transform 1 0 968 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1658
timestamp 1569139307
transform 1 0 1224 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1659
timestamp 1569139307
transform 1 0 968 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1660
timestamp 1569139307
transform 1 0 648 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1661
timestamp 1569139307
transform 1 0 648 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1662
timestamp 1569139307
transform 1 0 648 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1663
timestamp 1569139307
transform 1 0 648 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1664
timestamp 1569139307
transform 1 0 648 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1665
timestamp 1569139307
transform 1 0 648 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1666
timestamp 1569139307
transform 1 0 648 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1667
timestamp 1569139307
transform 1 0 648 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1668
timestamp 1569139307
transform 1 0 648 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1669
timestamp 1569139307
transform 1 0 648 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1670
timestamp 1569139307
transform 1 0 648 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1671
timestamp 1569139307
transform 1 0 648 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1672
timestamp 1569139307
transform 1 0 648 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1673
timestamp 1569139307
transform 1 0 648 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1674
timestamp 1569139307
transform 1 0 648 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1675
timestamp 1569139307
transform 1 0 648 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1676
timestamp 1569139307
transform 1 0 648 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1677
timestamp 1569139307
transform 1 0 648 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1678
timestamp 1569139307
transform 1 0 648 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1679
timestamp 1569139307
transform 1 0 2248 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1680
timestamp 1569139307
transform 1 0 2376 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1681
timestamp 1569139307
transform 1 0 2376 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1682
timestamp 1569139307
transform 1 0 2312 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1683
timestamp 1569139307
transform 1 0 2248 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1684
timestamp 1569139307
transform 1 0 2440 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1685
timestamp 1569139307
transform 1 0 2248 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1686
timestamp 1569139307
transform 1 0 2312 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1687
timestamp 1569139307
transform 1 0 2248 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1688
timestamp 1569139307
transform 1 0 2440 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1689
timestamp 1569139307
transform 1 0 2312 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1690
timestamp 1569139307
transform 1 0 2376 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1691
timestamp 1569139307
transform 1 0 2440 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1692
timestamp 1569139307
transform 1 0 2312 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1693
timestamp 1569139307
transform 1 0 2376 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1694
timestamp 1569139307
transform 1 0 2440 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1695
timestamp 1569139307
transform 1 0 2376 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1696
timestamp 1569139307
transform 1 0 2248 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1697
timestamp 1569139307
transform 1 0 2312 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1698
timestamp 1569139307
transform 1 0 2440 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1699
timestamp 1569139307
transform 1 0 2056 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1700
timestamp 1569139307
transform 1 0 1928 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1701
timestamp 1569139307
transform 1 0 2056 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1702
timestamp 1569139307
transform 1 0 2056 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1703
timestamp 1569139307
transform 1 0 2056 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1704
timestamp 1569139307
transform 1 0 1928 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1705
timestamp 1569139307
transform 1 0 2120 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1706
timestamp 1569139307
transform 1 0 2120 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1707
timestamp 1569139307
transform 1 0 2184 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1708
timestamp 1569139307
transform 1 0 2120 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1709
timestamp 1569139307
transform 1 0 1992 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1710
timestamp 1569139307
transform 1 0 2120 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1711
timestamp 1569139307
transform 1 0 2120 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1712
timestamp 1569139307
transform 1 0 2184 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1713
timestamp 1569139307
transform 1 0 2184 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1714
timestamp 1569139307
transform 1 0 2056 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1715
timestamp 1569139307
transform 1 0 2184 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1716
timestamp 1569139307
transform 1 0 2184 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1717
timestamp 1569139307
transform 1 0 1928 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1718
timestamp 1569139307
transform 1 0 1992 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1719
timestamp 1569139307
transform 1 0 1992 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1720
timestamp 1569139307
transform 1 0 1928 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1721
timestamp 1569139307
transform 1 0 1928 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1722
timestamp 1569139307
transform 1 0 1992 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1723
timestamp 1569139307
transform 1 0 1992 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1724
timestamp 1569139307
transform 1 0 2056 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1725
timestamp 1569139307
transform 1 0 2184 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1726
timestamp 1569139307
transform 1 0 2056 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1727
timestamp 1569139307
transform 1 0 2056 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1728
timestamp 1569139307
transform 1 0 1928 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1729
timestamp 1569139307
transform 1 0 2056 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1730
timestamp 1569139307
transform 1 0 2056 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1731
timestamp 1569139307
transform 1 0 2184 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1732
timestamp 1569139307
transform 1 0 2184 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1733
timestamp 1569139307
transform 1 0 2184 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1734
timestamp 1569139307
transform 1 0 2184 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1735
timestamp 1569139307
transform 1 0 2120 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1736
timestamp 1569139307
transform 1 0 1992 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1737
timestamp 1569139307
transform 1 0 2120 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1738
timestamp 1569139307
transform 1 0 2120 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1739
timestamp 1569139307
transform 1 0 1928 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1740
timestamp 1569139307
transform 1 0 2120 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1741
timestamp 1569139307
transform 1 0 2120 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1742
timestamp 1569139307
transform 1 0 1928 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1743
timestamp 1569139307
transform 1 0 1928 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1744
timestamp 1569139307
transform 1 0 1928 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1745
timestamp 1569139307
transform 1 0 1992 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1746
timestamp 1569139307
transform 1 0 1992 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1747
timestamp 1569139307
transform 1 0 1992 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1748
timestamp 1569139307
transform 1 0 1992 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1749
timestamp 1569139307
transform 1 0 2376 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1750
timestamp 1569139307
transform 1 0 2440 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1751
timestamp 1569139307
transform 1 0 2440 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1752
timestamp 1569139307
transform 1 0 2376 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1753
timestamp 1569139307
transform 1 0 2440 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1754
timestamp 1569139307
transform 1 0 2440 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1755
timestamp 1569139307
transform 1 0 2440 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1756
timestamp 1569139307
transform 1 0 2312 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1757
timestamp 1569139307
transform 1 0 2248 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1758
timestamp 1569139307
transform 1 0 2248 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1759
timestamp 1569139307
transform 1 0 2312 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1760
timestamp 1569139307
transform 1 0 2248 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1761
timestamp 1569139307
transform 1 0 2248 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1762
timestamp 1569139307
transform 1 0 2312 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1763
timestamp 1569139307
transform 1 0 2248 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1764
timestamp 1569139307
transform 1 0 2312 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1765
timestamp 1569139307
transform 1 0 2312 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1766
timestamp 1569139307
transform 1 0 2376 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1767
timestamp 1569139307
transform 1 0 2376 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1768
timestamp 1569139307
transform 1 0 2376 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1769
timestamp 1569139307
transform 1 0 1672 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1770
timestamp 1569139307
transform 1 0 1672 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1771
timestamp 1569139307
transform 1 0 1608 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1772
timestamp 1569139307
transform 1 0 1608 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1773
timestamp 1569139307
transform 1 0 1800 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1774
timestamp 1569139307
transform 1 0 1800 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1775
timestamp 1569139307
transform 1 0 1672 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1776
timestamp 1569139307
transform 1 0 1672 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1777
timestamp 1569139307
transform 1 0 1672 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1778
timestamp 1569139307
transform 1 0 1736 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1779
timestamp 1569139307
transform 1 0 1864 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1780
timestamp 1569139307
transform 1 0 1736 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1781
timestamp 1569139307
transform 1 0 1736 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1782
timestamp 1569139307
transform 1 0 1800 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1783
timestamp 1569139307
transform 1 0 1800 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1784
timestamp 1569139307
transform 1 0 1800 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1785
timestamp 1569139307
transform 1 0 1736 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1786
timestamp 1569139307
transform 1 0 1736 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1787
timestamp 1569139307
transform 1 0 1864 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1788
timestamp 1569139307
transform 1 0 1864 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1789
timestamp 1569139307
transform 1 0 1864 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1790
timestamp 1569139307
transform 1 0 1864 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1791
timestamp 1569139307
transform 1 0 1608 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1792
timestamp 1569139307
transform 1 0 1608 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1793
timestamp 1569139307
transform 1 0 1608 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1794
timestamp 1569139307
transform 1 0 1544 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1795
timestamp 1569139307
transform 1 0 1544 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1796
timestamp 1569139307
transform 1 0 1288 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1797
timestamp 1569139307
transform 1 0 1288 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1798
timestamp 1569139307
transform 1 0 1288 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1799
timestamp 1569139307
transform 1 0 1288 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1800
timestamp 1569139307
transform 1 0 1288 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1801
timestamp 1569139307
transform 1 0 1480 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1802
timestamp 1569139307
transform 1 0 1416 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1803
timestamp 1569139307
transform 1 0 1416 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1804
timestamp 1569139307
transform 1 0 1480 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1805
timestamp 1569139307
transform 1 0 1352 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1806
timestamp 1569139307
transform 1 0 1352 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1807
timestamp 1569139307
transform 1 0 1352 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1808
timestamp 1569139307
transform 1 0 1416 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1809
timestamp 1569139307
transform 1 0 1416 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1810
timestamp 1569139307
transform 1 0 1416 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1811
timestamp 1569139307
transform 1 0 1480 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1812
timestamp 1569139307
transform 1 0 1480 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1813
timestamp 1569139307
transform 1 0 1480 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1814
timestamp 1569139307
transform 1 0 1544 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_1815
timestamp 1569139307
transform 1 0 1544 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_1816
timestamp 1569139307
transform 1 0 1544 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_1817
timestamp 1569139307
transform 1 0 1352 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_1818
timestamp 1569139307
transform 1 0 1352 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_1819
timestamp 1569139307
transform 1 0 1544 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1820
timestamp 1569139307
transform 1 0 1352 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1821
timestamp 1569139307
transform 1 0 1352 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1822
timestamp 1569139307
transform 1 0 1352 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1823
timestamp 1569139307
transform 1 0 1352 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1824
timestamp 1569139307
transform 1 0 1352 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1825
timestamp 1569139307
transform 1 0 1544 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1826
timestamp 1569139307
transform 1 0 1544 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1827
timestamp 1569139307
transform 1 0 1544 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1828
timestamp 1569139307
transform 1 0 1416 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1829
timestamp 1569139307
transform 1 0 1416 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1830
timestamp 1569139307
transform 1 0 1288 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1831
timestamp 1569139307
transform 1 0 1416 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1832
timestamp 1569139307
transform 1 0 1416 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1833
timestamp 1569139307
transform 1 0 1416 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1834
timestamp 1569139307
transform 1 0 1288 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1835
timestamp 1569139307
transform 1 0 1288 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1836
timestamp 1569139307
transform 1 0 1480 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1837
timestamp 1569139307
transform 1 0 1480 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1838
timestamp 1569139307
transform 1 0 1480 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1839
timestamp 1569139307
transform 1 0 1480 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1840
timestamp 1569139307
transform 1 0 1480 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1841
timestamp 1569139307
transform 1 0 1288 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1842
timestamp 1569139307
transform 1 0 1288 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1843
timestamp 1569139307
transform 1 0 1544 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1844
timestamp 1569139307
transform 1 0 1800 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1845
timestamp 1569139307
transform 1 0 1800 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1846
timestamp 1569139307
transform 1 0 1608 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1847
timestamp 1569139307
transform 1 0 1608 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1848
timestamp 1569139307
transform 1 0 1608 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1849
timestamp 1569139307
transform 1 0 1608 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1850
timestamp 1569139307
transform 1 0 1608 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1851
timestamp 1569139307
transform 1 0 1800 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1852
timestamp 1569139307
transform 1 0 1800 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1853
timestamp 1569139307
transform 1 0 1864 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1854
timestamp 1569139307
transform 1 0 1864 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1855
timestamp 1569139307
transform 1 0 1864 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1856
timestamp 1569139307
transform 1 0 1672 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1857
timestamp 1569139307
transform 1 0 1672 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1858
timestamp 1569139307
transform 1 0 1672 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1859
timestamp 1569139307
transform 1 0 1672 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1860
timestamp 1569139307
transform 1 0 1672 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1861
timestamp 1569139307
transform 1 0 1864 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1862
timestamp 1569139307
transform 1 0 1736 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1863
timestamp 1569139307
transform 1 0 1736 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_1864
timestamp 1569139307
transform 1 0 1736 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_1865
timestamp 1569139307
transform 1 0 1736 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1866
timestamp 1569139307
transform 1 0 1736 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_1867
timestamp 1569139307
transform 1 0 1864 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_1868
timestamp 1569139307
transform 1 0 1800 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_1869
timestamp 1569139307
transform 1 0 1800 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1870
timestamp 1569139307
transform 1 0 1608 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1871
timestamp 1569139307
transform 1 0 1864 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1872
timestamp 1569139307
transform 1 0 1608 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1873
timestamp 1569139307
transform 1 0 1800 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1874
timestamp 1569139307
transform 1 0 1672 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1875
timestamp 1569139307
transform 1 0 1864 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1876
timestamp 1569139307
transform 1 0 1672 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1877
timestamp 1569139307
transform 1 0 1864 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1878
timestamp 1569139307
transform 1 0 1672 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1879
timestamp 1569139307
transform 1 0 1864 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1880
timestamp 1569139307
transform 1 0 1672 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1881
timestamp 1569139307
transform 1 0 1672 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1882
timestamp 1569139307
transform 1 0 1736 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1883
timestamp 1569139307
transform 1 0 1800 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1884
timestamp 1569139307
transform 1 0 1736 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1885
timestamp 1569139307
transform 1 0 1736 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1886
timestamp 1569139307
transform 1 0 1608 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1887
timestamp 1569139307
transform 1 0 1736 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1888
timestamp 1569139307
transform 1 0 1608 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1889
timestamp 1569139307
transform 1 0 1736 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1890
timestamp 1569139307
transform 1 0 1608 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1891
timestamp 1569139307
transform 1 0 1864 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1892
timestamp 1569139307
transform 1 0 1800 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1893
timestamp 1569139307
transform 1 0 1800 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1894
timestamp 1569139307
transform 1 0 1352 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1895
timestamp 1569139307
transform 1 0 1480 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1896
timestamp 1569139307
transform 1 0 1480 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1897
timestamp 1569139307
transform 1 0 1544 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1898
timestamp 1569139307
transform 1 0 1544 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1899
timestamp 1569139307
transform 1 0 1416 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1900
timestamp 1569139307
transform 1 0 1288 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1901
timestamp 1569139307
transform 1 0 1544 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1902
timestamp 1569139307
transform 1 0 1416 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1903
timestamp 1569139307
transform 1 0 1544 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1904
timestamp 1569139307
transform 1 0 1288 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1905
timestamp 1569139307
transform 1 0 1544 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1906
timestamp 1569139307
transform 1 0 1480 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1907
timestamp 1569139307
transform 1 0 1288 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1908
timestamp 1569139307
transform 1 0 1480 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1909
timestamp 1569139307
transform 1 0 1288 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1910
timestamp 1569139307
transform 1 0 1352 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1911
timestamp 1569139307
transform 1 0 1352 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1912
timestamp 1569139307
transform 1 0 1352 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1913
timestamp 1569139307
transform 1 0 1288 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1914
timestamp 1569139307
transform 1 0 1352 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1915
timestamp 1569139307
transform 1 0 1416 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1916
timestamp 1569139307
transform 1 0 1416 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1917
timestamp 1569139307
transform 1 0 1416 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1918
timestamp 1569139307
transform 1 0 1480 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1919
timestamp 1569139307
transform 1 0 1352 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1920
timestamp 1569139307
transform 1 0 1288 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1921
timestamp 1569139307
transform 1 0 1544 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1922
timestamp 1569139307
transform 1 0 1352 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1923
timestamp 1569139307
transform 1 0 1288 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1924
timestamp 1569139307
transform 1 0 1416 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1925
timestamp 1569139307
transform 1 0 1416 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1926
timestamp 1569139307
transform 1 0 1480 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1927
timestamp 1569139307
transform 1 0 1480 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1928
timestamp 1569139307
transform 1 0 1480 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1929
timestamp 1569139307
transform 1 0 1352 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1930
timestamp 1569139307
transform 1 0 1480 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1931
timestamp 1569139307
transform 1 0 1544 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1932
timestamp 1569139307
transform 1 0 1416 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1933
timestamp 1569139307
transform 1 0 1544 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1934
timestamp 1569139307
transform 1 0 1288 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1935
timestamp 1569139307
transform 1 0 1544 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1936
timestamp 1569139307
transform 1 0 1416 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1937
timestamp 1569139307
transform 1 0 1288 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1938
timestamp 1569139307
transform 1 0 1352 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1939
timestamp 1569139307
transform 1 0 1608 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1940
timestamp 1569139307
transform 1 0 1864 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1941
timestamp 1569139307
transform 1 0 1608 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1942
timestamp 1569139307
transform 1 0 1672 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1943
timestamp 1569139307
transform 1 0 1672 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1944
timestamp 1569139307
transform 1 0 1672 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1945
timestamp 1569139307
transform 1 0 1736 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1946
timestamp 1569139307
transform 1 0 1736 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1947
timestamp 1569139307
transform 1 0 1800 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1948
timestamp 1569139307
transform 1 0 1736 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1949
timestamp 1569139307
transform 1 0 1800 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1950
timestamp 1569139307
transform 1 0 1864 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1951
timestamp 1569139307
transform 1 0 1800 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1952
timestamp 1569139307
transform 1 0 1608 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1953
timestamp 1569139307
transform 1 0 1800 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1954
timestamp 1569139307
transform 1 0 1864 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_1955
timestamp 1569139307
transform 1 0 1608 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1956
timestamp 1569139307
transform 1 0 1864 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_1957
timestamp 1569139307
transform 1 0 1672 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1958
timestamp 1569139307
transform 1 0 1736 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_1959
timestamp 1569139307
transform 1 0 2376 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1960
timestamp 1569139307
transform 1 0 2376 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1961
timestamp 1569139307
transform 1 0 2248 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1962
timestamp 1569139307
transform 1 0 2440 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1963
timestamp 1569139307
transform 1 0 2440 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1964
timestamp 1569139307
transform 1 0 2312 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1965
timestamp 1569139307
transform 1 0 2376 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1966
timestamp 1569139307
transform 1 0 2248 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1967
timestamp 1569139307
transform 1 0 2248 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1968
timestamp 1569139307
transform 1 0 2312 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1969
timestamp 1569139307
transform 1 0 2312 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1970
timestamp 1569139307
transform 1 0 2248 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1971
timestamp 1569139307
transform 1 0 2248 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1972
timestamp 1569139307
transform 1 0 2312 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1973
timestamp 1569139307
transform 1 0 1992 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1974
timestamp 1569139307
transform 1 0 1992 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1975
timestamp 1569139307
transform 1 0 1928 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1976
timestamp 1569139307
transform 1 0 2056 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1977
timestamp 1569139307
transform 1 0 2056 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1978
timestamp 1569139307
transform 1 0 1992 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1979
timestamp 1569139307
transform 1 0 2120 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1980
timestamp 1569139307
transform 1 0 2120 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1981
timestamp 1569139307
transform 1 0 2056 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1982
timestamp 1569139307
transform 1 0 2184 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1983
timestamp 1569139307
transform 1 0 2184 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1984
timestamp 1569139307
transform 1 0 2120 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1985
timestamp 1569139307
transform 1 0 2056 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1986
timestamp 1569139307
transform 1 0 2056 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1987
timestamp 1569139307
transform 1 0 2120 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1988
timestamp 1569139307
transform 1 0 2120 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1989
timestamp 1569139307
transform 1 0 2184 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1990
timestamp 1569139307
transform 1 0 1928 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1991
timestamp 1569139307
transform 1 0 2184 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1992
timestamp 1569139307
transform 1 0 1992 0 1 2184
box -8 -8 8 8
use VIA1  VIA1_1993
timestamp 1569139307
transform 1 0 2184 0 1 2056
box -8 -8 8 8
use VIA1  VIA1_1994
timestamp 1569139307
transform 1 0 1928 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_1995
timestamp 1569139307
transform 1 0 1928 0 1 1992
box -8 -8 8 8
use VIA1  VIA1_1996
timestamp 1569139307
transform 1 0 1928 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1997
timestamp 1569139307
transform 1 0 1992 0 1 2120
box -8 -8 8 8
use VIA1  VIA1_1998
timestamp 1569139307
transform 1 0 2056 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_1999
timestamp 1569139307
transform 1 0 1928 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_2000
timestamp 1569139307
transform 1 0 1928 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_2001
timestamp 1569139307
transform 1 0 1992 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_2002
timestamp 1569139307
transform 1 0 1992 0 1 2440
box -8 -8 8 8
use VIA1  VIA1_2003
timestamp 1569139307
transform 1 0 2184 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_2004
timestamp 1569139307
transform 1 0 1928 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_2005
timestamp 1569139307
transform 1 0 2056 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_2006
timestamp 1569139307
transform 1 0 1992 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_2007
timestamp 1569139307
transform 1 0 2120 0 1 2248
box -8 -8 8 8
use VIA1  VIA1_2008
timestamp 1569139307
transform 1 0 2056 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_2009
timestamp 1569139307
transform 1 0 2120 0 1 2312
box -8 -8 8 8
use VIA1  VIA1_2010
timestamp 1569139307
transform 1 0 1928 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_2011
timestamp 1569139307
transform 1 0 1992 0 1 2376
box -8 -8 8 8
use VIA1  VIA1_2012
timestamp 1569139307
transform 1 0 1864 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2013
timestamp 1569139307
transform 1 0 1672 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2014
timestamp 1569139307
transform 1 0 1672 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2015
timestamp 1569139307
transform 1 0 1608 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2016
timestamp 1569139307
transform 1 0 1736 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2017
timestamp 1569139307
transform 1 0 1608 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2018
timestamp 1569139307
transform 1 0 1800 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2019
timestamp 1569139307
transform 1 0 1672 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2020
timestamp 1569139307
transform 1 0 1800 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2021
timestamp 1569139307
transform 1 0 1672 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2022
timestamp 1569139307
transform 1 0 1736 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2023
timestamp 1569139307
transform 1 0 1608 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2024
timestamp 1569139307
transform 1 0 1608 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2025
timestamp 1569139307
transform 1 0 1480 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2026
timestamp 1569139307
transform 1 0 1416 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2027
timestamp 1569139307
transform 1 0 1352 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2028
timestamp 1569139307
transform 1 0 1416 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2029
timestamp 1569139307
transform 1 0 1416 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2030
timestamp 1569139307
transform 1 0 1416 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2031
timestamp 1569139307
transform 1 0 1352 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2032
timestamp 1569139307
transform 1 0 1352 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2033
timestamp 1569139307
transform 1 0 1288 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2034
timestamp 1569139307
transform 1 0 1544 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2035
timestamp 1569139307
transform 1 0 1288 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2036
timestamp 1569139307
transform 1 0 1544 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2037
timestamp 1569139307
transform 1 0 1288 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2038
timestamp 1569139307
transform 1 0 1352 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2039
timestamp 1569139307
transform 1 0 1480 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2040
timestamp 1569139307
transform 1 0 1544 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2041
timestamp 1569139307
transform 1 0 1480 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2042
timestamp 1569139307
transform 1 0 1544 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2043
timestamp 1569139307
transform 1 0 1480 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2044
timestamp 1569139307
transform 1 0 1288 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2045
timestamp 1569139307
transform 1 0 1288 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2046
timestamp 1569139307
transform 1 0 1288 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2047
timestamp 1569139307
transform 1 0 1288 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2048
timestamp 1569139307
transform 1 0 1544 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2049
timestamp 1569139307
transform 1 0 1544 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2050
timestamp 1569139307
transform 1 0 1416 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2051
timestamp 1569139307
transform 1 0 1288 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2052
timestamp 1569139307
transform 1 0 1416 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2053
timestamp 1569139307
transform 1 0 1352 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2054
timestamp 1569139307
transform 1 0 1352 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2055
timestamp 1569139307
transform 1 0 1416 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2056
timestamp 1569139307
transform 1 0 1480 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2057
timestamp 1569139307
transform 1 0 1288 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2058
timestamp 1569139307
transform 1 0 1416 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2059
timestamp 1569139307
transform 1 0 1480 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2060
timestamp 1569139307
transform 1 0 1352 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2061
timestamp 1569139307
transform 1 0 1480 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2062
timestamp 1569139307
transform 1 0 1352 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2063
timestamp 1569139307
transform 1 0 1416 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2064
timestamp 1569139307
transform 1 0 1352 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2065
timestamp 1569139307
transform 1 0 1480 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2066
timestamp 1569139307
transform 1 0 1480 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2067
timestamp 1569139307
transform 1 0 1608 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2068
timestamp 1569139307
transform 1 0 1480 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2069
timestamp 1569139307
transform 1 0 1480 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2070
timestamp 1569139307
transform 1 0 1480 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2071
timestamp 1569139307
transform 1 0 1352 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2072
timestamp 1569139307
transform 1 0 1288 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2073
timestamp 1569139307
transform 1 0 1480 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2074
timestamp 1569139307
transform 1 0 1480 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2075
timestamp 1569139307
transform 1 0 1352 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2076
timestamp 1569139307
transform 1 0 1416 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2077
timestamp 1569139307
transform 1 0 1480 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2078
timestamp 1569139307
transform 1 0 1288 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2079
timestamp 1569139307
transform 1 0 1288 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2080
timestamp 1569139307
transform 1 0 1416 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2081
timestamp 1569139307
transform 1 0 1480 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2082
timestamp 1569139307
transform 1 0 1480 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2083
timestamp 1569139307
transform 1 0 1352 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2084
timestamp 1569139307
transform 1 0 1352 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2085
timestamp 1569139307
transform 1 0 1352 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2086
timestamp 1569139307
transform 1 0 1288 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2087
timestamp 1569139307
transform 1 0 1288 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2088
timestamp 1569139307
transform 1 0 1352 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2089
timestamp 1569139307
transform 1 0 1352 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2090
timestamp 1569139307
transform 1 0 1288 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2091
timestamp 1569139307
transform 1 0 1416 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2092
timestamp 1569139307
transform 1 0 1352 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2093
timestamp 1569139307
transform 1 0 1416 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2094
timestamp 1569139307
transform 1 0 1480 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2095
timestamp 1569139307
transform 1 0 1288 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2096
timestamp 1569139307
transform 1 0 1416 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2097
timestamp 1569139307
transform 1 0 1416 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2098
timestamp 1569139307
transform 1 0 1352 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2099
timestamp 1569139307
transform 1 0 1288 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2100
timestamp 1569139307
transform 1 0 1352 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2101
timestamp 1569139307
transform 1 0 1416 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2102
timestamp 1569139307
transform 1 0 1480 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2103
timestamp 1569139307
transform 1 0 1288 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2104
timestamp 1569139307
transform 1 0 1416 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2105
timestamp 1569139307
transform 1 0 1416 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2106
timestamp 1569139307
transform 1 0 1288 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2107
timestamp 1569139307
transform 1 0 1416 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2108
timestamp 1569139307
transform 1 0 2440 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2109
timestamp 1569139307
transform 1 0 2440 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2110
timestamp 1569139307
transform 1 0 2440 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2111
timestamp 1569139307
transform 1 0 2376 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2112
timestamp 1569139307
transform 1 0 2376 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2113
timestamp 1569139307
transform 1 0 2440 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2114
timestamp 1569139307
transform 1 0 2376 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2115
timestamp 1569139307
transform 1 0 2312 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2116
timestamp 1569139307
transform 1 0 2376 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2117
timestamp 1569139307
transform 1 0 2440 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2118
timestamp 1569139307
transform 1 0 2376 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2119
timestamp 1569139307
transform 1 0 2376 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2120
timestamp 1569139307
transform 1 0 2376 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2121
timestamp 1569139307
transform 1 0 2312 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2122
timestamp 1569139307
transform 1 0 2312 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2123
timestamp 1569139307
transform 1 0 2312 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2124
timestamp 1569139307
transform 1 0 2312 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2125
timestamp 1569139307
transform 1 0 2312 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2126
timestamp 1569139307
transform 1 0 2440 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2127
timestamp 1569139307
transform 1 0 2440 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2128
timestamp 1569139307
transform 1 0 2440 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2129
timestamp 1569139307
transform 1 0 1096 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2130
timestamp 1569139307
transform 1 0 1160 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2131
timestamp 1569139307
transform 1 0 968 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2132
timestamp 1569139307
transform 1 0 1096 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2133
timestamp 1569139307
transform 1 0 1032 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2134
timestamp 1569139307
transform 1 0 968 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2135
timestamp 1569139307
transform 1 0 1160 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2136
timestamp 1569139307
transform 1 0 1224 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2137
timestamp 1569139307
transform 1 0 1032 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2138
timestamp 1569139307
transform 1 0 1160 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2139
timestamp 1569139307
transform 1 0 1224 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2140
timestamp 1569139307
transform 1 0 1160 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2141
timestamp 1569139307
transform 1 0 968 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2142
timestamp 1569139307
transform 1 0 1096 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2143
timestamp 1569139307
transform 1 0 1032 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2144
timestamp 1569139307
transform 1 0 1096 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2145
timestamp 1569139307
transform 1 0 1032 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2146
timestamp 1569139307
transform 1 0 1224 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2147
timestamp 1569139307
transform 1 0 1224 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2148
timestamp 1569139307
transform 1 0 968 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2149
timestamp 1569139307
transform 1 0 904 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2150
timestamp 1569139307
transform 1 0 904 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2151
timestamp 1569139307
transform 1 0 840 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2152
timestamp 1569139307
transform 1 0 776 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2153
timestamp 1569139307
transform 1 0 840 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2154
timestamp 1569139307
transform 1 0 712 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2155
timestamp 1569139307
transform 1 0 904 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2156
timestamp 1569139307
transform 1 0 712 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2157
timestamp 1569139307
transform 1 0 776 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2158
timestamp 1569139307
transform 1 0 712 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2159
timestamp 1569139307
transform 1 0 776 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2160
timestamp 1569139307
transform 1 0 776 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2161
timestamp 1569139307
transform 1 0 840 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2162
timestamp 1569139307
transform 1 0 904 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2163
timestamp 1569139307
transform 1 0 712 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2164
timestamp 1569139307
transform 1 0 840 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2165
timestamp 1569139307
transform 1 0 840 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2166
timestamp 1569139307
transform 1 0 712 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2167
timestamp 1569139307
transform 1 0 904 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2168
timestamp 1569139307
transform 1 0 776 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2169
timestamp 1569139307
transform 1 0 712 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2170
timestamp 1569139307
transform 1 0 904 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2171
timestamp 1569139307
transform 1 0 904 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2172
timestamp 1569139307
transform 1 0 840 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2173
timestamp 1569139307
transform 1 0 904 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2174
timestamp 1569139307
transform 1 0 840 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2175
timestamp 1569139307
transform 1 0 712 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2176
timestamp 1569139307
transform 1 0 712 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2177
timestamp 1569139307
transform 1 0 776 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2178
timestamp 1569139307
transform 1 0 840 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2179
timestamp 1569139307
transform 1 0 776 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2180
timestamp 1569139307
transform 1 0 840 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2181
timestamp 1569139307
transform 1 0 712 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2182
timestamp 1569139307
transform 1 0 776 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2183
timestamp 1569139307
transform 1 0 776 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2184
timestamp 1569139307
transform 1 0 904 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2185
timestamp 1569139307
transform 1 0 1160 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2186
timestamp 1569139307
transform 1 0 1032 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2187
timestamp 1569139307
transform 1 0 1160 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2188
timestamp 1569139307
transform 1 0 1160 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2189
timestamp 1569139307
transform 1 0 1096 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2190
timestamp 1569139307
transform 1 0 968 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2191
timestamp 1569139307
transform 1 0 1032 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2192
timestamp 1569139307
transform 1 0 1096 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2193
timestamp 1569139307
transform 1 0 1160 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2194
timestamp 1569139307
transform 1 0 968 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2195
timestamp 1569139307
transform 1 0 1224 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2196
timestamp 1569139307
transform 1 0 1224 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2197
timestamp 1569139307
transform 1 0 968 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2198
timestamp 1569139307
transform 1 0 1032 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2199
timestamp 1569139307
transform 1 0 1224 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2200
timestamp 1569139307
transform 1 0 968 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2201
timestamp 1569139307
transform 1 0 1032 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2202
timestamp 1569139307
transform 1 0 1096 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2203
timestamp 1569139307
transform 1 0 1160 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2204
timestamp 1569139307
transform 1 0 1032 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2205
timestamp 1569139307
transform 1 0 968 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2206
timestamp 1569139307
transform 1 0 1096 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2207
timestamp 1569139307
transform 1 0 1224 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2208
timestamp 1569139307
transform 1 0 1096 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2209
timestamp 1569139307
transform 1 0 1224 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2210
timestamp 1569139307
transform 1 0 584 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2211
timestamp 1569139307
transform 1 0 520 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2212
timestamp 1569139307
transform 1 0 392 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2213
timestamp 1569139307
transform 1 0 584 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2214
timestamp 1569139307
transform 1 0 520 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2215
timestamp 1569139307
transform 1 0 392 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2216
timestamp 1569139307
transform 1 0 584 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2217
timestamp 1569139307
transform 1 0 456 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2218
timestamp 1569139307
transform 1 0 392 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2219
timestamp 1569139307
transform 1 0 456 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2220
timestamp 1569139307
transform 1 0 520 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2221
timestamp 1569139307
transform 1 0 520 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2222
timestamp 1569139307
transform 1 0 392 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2223
timestamp 1569139307
transform 1 0 456 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2224
timestamp 1569139307
transform 1 0 456 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2225
timestamp 1569139307
transform 1 0 584 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2226
timestamp 1569139307
transform 1 0 72 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2227
timestamp 1569139307
transform 1 0 328 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2228
timestamp 1569139307
transform 1 0 72 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2229
timestamp 1569139307
transform 1 0 264 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2230
timestamp 1569139307
transform 1 0 264 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2231
timestamp 1569139307
transform 1 0 136 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2232
timestamp 1569139307
transform 1 0 328 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2233
timestamp 1569139307
transform 1 0 200 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2234
timestamp 1569139307
transform 1 0 136 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2235
timestamp 1569139307
transform 1 0 264 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2236
timestamp 1569139307
transform 1 0 328 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2237
timestamp 1569139307
transform 1 0 72 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2238
timestamp 1569139307
transform 1 0 200 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2239
timestamp 1569139307
transform 1 0 72 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2240
timestamp 1569139307
transform 1 0 200 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2241
timestamp 1569139307
transform 1 0 136 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2242
timestamp 1569139307
transform 1 0 264 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2243
timestamp 1569139307
transform 1 0 136 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2244
timestamp 1569139307
transform 1 0 328 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2245
timestamp 1569139307
transform 1 0 200 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2246
timestamp 1569139307
transform 1 0 264 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2247
timestamp 1569139307
transform 1 0 264 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2248
timestamp 1569139307
transform 1 0 136 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2249
timestamp 1569139307
transform 1 0 264 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2250
timestamp 1569139307
transform 1 0 264 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2251
timestamp 1569139307
transform 1 0 200 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2252
timestamp 1569139307
transform 1 0 136 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2253
timestamp 1569139307
transform 1 0 328 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2254
timestamp 1569139307
transform 1 0 136 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2255
timestamp 1569139307
transform 1 0 72 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2256
timestamp 1569139307
transform 1 0 200 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2257
timestamp 1569139307
transform 1 0 136 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2258
timestamp 1569139307
transform 1 0 72 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2259
timestamp 1569139307
transform 1 0 328 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2260
timestamp 1569139307
transform 1 0 328 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2261
timestamp 1569139307
transform 1 0 328 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2262
timestamp 1569139307
transform 1 0 72 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2263
timestamp 1569139307
transform 1 0 328 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2264
timestamp 1569139307
transform 1 0 72 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2265
timestamp 1569139307
transform 1 0 200 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2266
timestamp 1569139307
transform 1 0 200 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2267
timestamp 1569139307
transform 1 0 136 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2268
timestamp 1569139307
transform 1 0 264 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2269
timestamp 1569139307
transform 1 0 200 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2270
timestamp 1569139307
transform 1 0 72 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2271
timestamp 1569139307
transform 1 0 520 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2272
timestamp 1569139307
transform 1 0 392 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2273
timestamp 1569139307
transform 1 0 392 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2274
timestamp 1569139307
transform 1 0 392 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2275
timestamp 1569139307
transform 1 0 520 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2276
timestamp 1569139307
transform 1 0 584 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2277
timestamp 1569139307
transform 1 0 584 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2278
timestamp 1569139307
transform 1 0 456 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2279
timestamp 1569139307
transform 1 0 456 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2280
timestamp 1569139307
transform 1 0 520 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2281
timestamp 1569139307
transform 1 0 520 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2282
timestamp 1569139307
transform 1 0 520 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2283
timestamp 1569139307
transform 1 0 456 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2284
timestamp 1569139307
transform 1 0 392 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2285
timestamp 1569139307
transform 1 0 584 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2286
timestamp 1569139307
transform 1 0 584 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2287
timestamp 1569139307
transform 1 0 584 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2288
timestamp 1569139307
transform 1 0 456 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2289
timestamp 1569139307
transform 1 0 456 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2290
timestamp 1569139307
transform 1 0 392 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2291
timestamp 1569139307
transform 1 0 392 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2292
timestamp 1569139307
transform 1 0 584 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2293
timestamp 1569139307
transform 1 0 520 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2294
timestamp 1569139307
transform 1 0 392 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2295
timestamp 1569139307
transform 1 0 584 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2296
timestamp 1569139307
transform 1 0 392 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2297
timestamp 1569139307
transform 1 0 456 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2298
timestamp 1569139307
transform 1 0 456 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2299
timestamp 1569139307
transform 1 0 456 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2300
timestamp 1569139307
transform 1 0 392 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2301
timestamp 1569139307
transform 1 0 584 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2302
timestamp 1569139307
transform 1 0 520 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2303
timestamp 1569139307
transform 1 0 520 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2304
timestamp 1569139307
transform 1 0 456 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2305
timestamp 1569139307
transform 1 0 584 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2306
timestamp 1569139307
transform 1 0 520 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2307
timestamp 1569139307
transform 1 0 584 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2308
timestamp 1569139307
transform 1 0 520 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2309
timestamp 1569139307
transform 1 0 456 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2310
timestamp 1569139307
transform 1 0 392 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2311
timestamp 1569139307
transform 1 0 264 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2312
timestamp 1569139307
transform 1 0 200 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2313
timestamp 1569139307
transform 1 0 72 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2314
timestamp 1569139307
transform 1 0 72 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2315
timestamp 1569139307
transform 1 0 264 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2316
timestamp 1569139307
transform 1 0 264 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2317
timestamp 1569139307
transform 1 0 200 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2318
timestamp 1569139307
transform 1 0 200 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2319
timestamp 1569139307
transform 1 0 72 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2320
timestamp 1569139307
transform 1 0 328 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2321
timestamp 1569139307
transform 1 0 200 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2322
timestamp 1569139307
transform 1 0 136 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2323
timestamp 1569139307
transform 1 0 136 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2324
timestamp 1569139307
transform 1 0 328 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2325
timestamp 1569139307
transform 1 0 72 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2326
timestamp 1569139307
transform 1 0 136 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2327
timestamp 1569139307
transform 1 0 328 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2328
timestamp 1569139307
transform 1 0 72 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2329
timestamp 1569139307
transform 1 0 136 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2330
timestamp 1569139307
transform 1 0 136 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2331
timestamp 1569139307
transform 1 0 328 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2332
timestamp 1569139307
transform 1 0 200 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2333
timestamp 1569139307
transform 1 0 264 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2334
timestamp 1569139307
transform 1 0 264 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2335
timestamp 1569139307
transform 1 0 328 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2336
timestamp 1569139307
transform 1 0 328 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2337
timestamp 1569139307
transform 1 0 328 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2338
timestamp 1569139307
transform 1 0 72 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2339
timestamp 1569139307
transform 1 0 200 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2340
timestamp 1569139307
transform 1 0 72 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2341
timestamp 1569139307
transform 1 0 136 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2342
timestamp 1569139307
transform 1 0 136 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2343
timestamp 1569139307
transform 1 0 72 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2344
timestamp 1569139307
transform 1 0 136 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2345
timestamp 1569139307
transform 1 0 72 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2346
timestamp 1569139307
transform 1 0 136 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2347
timestamp 1569139307
transform 1 0 328 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2348
timestamp 1569139307
transform 1 0 200 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2349
timestamp 1569139307
transform 1 0 136 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2350
timestamp 1569139307
transform 1 0 72 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2351
timestamp 1569139307
transform 1 0 200 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2352
timestamp 1569139307
transform 1 0 328 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2353
timestamp 1569139307
transform 1 0 264 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2354
timestamp 1569139307
transform 1 0 264 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2355
timestamp 1569139307
transform 1 0 264 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2356
timestamp 1569139307
transform 1 0 264 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2357
timestamp 1569139307
transform 1 0 264 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2358
timestamp 1569139307
transform 1 0 200 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2359
timestamp 1569139307
transform 1 0 200 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2360
timestamp 1569139307
transform 1 0 328 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2361
timestamp 1569139307
transform 1 0 392 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2362
timestamp 1569139307
transform 1 0 456 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2363
timestamp 1569139307
transform 1 0 392 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2364
timestamp 1569139307
transform 1 0 456 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2365
timestamp 1569139307
transform 1 0 584 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2366
timestamp 1569139307
transform 1 0 456 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2367
timestamp 1569139307
transform 1 0 456 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2368
timestamp 1569139307
transform 1 0 456 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2369
timestamp 1569139307
transform 1 0 584 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2370
timestamp 1569139307
transform 1 0 584 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2371
timestamp 1569139307
transform 1 0 520 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2372
timestamp 1569139307
transform 1 0 520 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2373
timestamp 1569139307
transform 1 0 520 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2374
timestamp 1569139307
transform 1 0 520 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2375
timestamp 1569139307
transform 1 0 584 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2376
timestamp 1569139307
transform 1 0 392 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2377
timestamp 1569139307
transform 1 0 584 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2378
timestamp 1569139307
transform 1 0 520 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2379
timestamp 1569139307
transform 1 0 392 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2380
timestamp 1569139307
transform 1 0 392 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2381
timestamp 1569139307
transform 1 0 1224 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2382
timestamp 1569139307
transform 1 0 968 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2383
timestamp 1569139307
transform 1 0 1096 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2384
timestamp 1569139307
transform 1 0 968 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2385
timestamp 1569139307
transform 1 0 968 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2386
timestamp 1569139307
transform 1 0 968 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2387
timestamp 1569139307
transform 1 0 1224 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2388
timestamp 1569139307
transform 1 0 1160 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2389
timestamp 1569139307
transform 1 0 1032 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2390
timestamp 1569139307
transform 1 0 1160 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2391
timestamp 1569139307
transform 1 0 1160 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2392
timestamp 1569139307
transform 1 0 1096 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2393
timestamp 1569139307
transform 1 0 1160 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2394
timestamp 1569139307
transform 1 0 1032 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2395
timestamp 1569139307
transform 1 0 1032 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2396
timestamp 1569139307
transform 1 0 1160 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2397
timestamp 1569139307
transform 1 0 1032 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2398
timestamp 1569139307
transform 1 0 1224 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2399
timestamp 1569139307
transform 1 0 968 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2400
timestamp 1569139307
transform 1 0 1096 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2401
timestamp 1569139307
transform 1 0 1096 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2402
timestamp 1569139307
transform 1 0 1224 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2403
timestamp 1569139307
transform 1 0 1032 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2404
timestamp 1569139307
transform 1 0 1224 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2405
timestamp 1569139307
transform 1 0 1096 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2406
timestamp 1569139307
transform 1 0 840 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2407
timestamp 1569139307
transform 1 0 840 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2408
timestamp 1569139307
transform 1 0 840 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2409
timestamp 1569139307
transform 1 0 712 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2410
timestamp 1569139307
transform 1 0 904 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2411
timestamp 1569139307
transform 1 0 904 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2412
timestamp 1569139307
transform 1 0 904 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2413
timestamp 1569139307
transform 1 0 904 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2414
timestamp 1569139307
transform 1 0 712 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2415
timestamp 1569139307
transform 1 0 776 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2416
timestamp 1569139307
transform 1 0 840 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2417
timestamp 1569139307
transform 1 0 776 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2418
timestamp 1569139307
transform 1 0 776 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2419
timestamp 1569139307
transform 1 0 776 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2420
timestamp 1569139307
transform 1 0 776 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2421
timestamp 1569139307
transform 1 0 712 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2422
timestamp 1569139307
transform 1 0 904 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2423
timestamp 1569139307
transform 1 0 712 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2424
timestamp 1569139307
transform 1 0 840 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2425
timestamp 1569139307
transform 1 0 712 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2426
timestamp 1569139307
transform 1 0 712 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2427
timestamp 1569139307
transform 1 0 712 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2428
timestamp 1569139307
transform 1 0 712 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2429
timestamp 1569139307
transform 1 0 712 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2430
timestamp 1569139307
transform 1 0 776 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2431
timestamp 1569139307
transform 1 0 776 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2432
timestamp 1569139307
transform 1 0 712 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2433
timestamp 1569139307
transform 1 0 840 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2434
timestamp 1569139307
transform 1 0 840 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2435
timestamp 1569139307
transform 1 0 776 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2436
timestamp 1569139307
transform 1 0 776 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2437
timestamp 1569139307
transform 1 0 776 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2438
timestamp 1569139307
transform 1 0 904 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2439
timestamp 1569139307
transform 1 0 840 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2440
timestamp 1569139307
transform 1 0 840 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2441
timestamp 1569139307
transform 1 0 904 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2442
timestamp 1569139307
transform 1 0 840 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2443
timestamp 1569139307
transform 1 0 904 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2444
timestamp 1569139307
transform 1 0 904 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2445
timestamp 1569139307
transform 1 0 904 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2446
timestamp 1569139307
transform 1 0 1096 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2447
timestamp 1569139307
transform 1 0 1096 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2448
timestamp 1569139307
transform 1 0 1096 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2449
timestamp 1569139307
transform 1 0 1224 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2450
timestamp 1569139307
transform 1 0 1096 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2451
timestamp 1569139307
transform 1 0 1096 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2452
timestamp 1569139307
transform 1 0 1224 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2453
timestamp 1569139307
transform 1 0 1160 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2454
timestamp 1569139307
transform 1 0 1160 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2455
timestamp 1569139307
transform 1 0 1160 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2456
timestamp 1569139307
transform 1 0 968 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2457
timestamp 1569139307
transform 1 0 968 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2458
timestamp 1569139307
transform 1 0 968 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2459
timestamp 1569139307
transform 1 0 1032 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2460
timestamp 1569139307
transform 1 0 1032 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2461
timestamp 1569139307
transform 1 0 1032 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2462
timestamp 1569139307
transform 1 0 1224 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2463
timestamp 1569139307
transform 1 0 1224 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2464
timestamp 1569139307
transform 1 0 1224 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2465
timestamp 1569139307
transform 1 0 1160 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2466
timestamp 1569139307
transform 1 0 968 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2467
timestamp 1569139307
transform 1 0 968 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2468
timestamp 1569139307
transform 1 0 1160 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2469
timestamp 1569139307
transform 1 0 1032 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2470
timestamp 1569139307
transform 1 0 1032 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2471
timestamp 1569139307
transform 1 0 648 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2472
timestamp 1569139307
transform 1 0 648 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_2473
timestamp 1569139307
transform 1 0 648 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2474
timestamp 1569139307
transform 1 0 648 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2475
timestamp 1569139307
transform 1 0 648 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2476
timestamp 1569139307
transform 1 0 648 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2477
timestamp 1569139307
transform 1 0 648 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_2478
timestamp 1569139307
transform 1 0 648 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_2479
timestamp 1569139307
transform 1 0 648 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2480
timestamp 1569139307
transform 1 0 648 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_2481
timestamp 1569139307
transform 1 0 648 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2482
timestamp 1569139307
transform 1 0 648 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2483
timestamp 1569139307
transform 1 0 648 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_2484
timestamp 1569139307
transform 1 0 648 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_2485
timestamp 1569139307
transform 1 0 648 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_2486
timestamp 1569139307
transform 1 0 648 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_2487
timestamp 1569139307
transform 1 0 648 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2488
timestamp 1569139307
transform 1 0 648 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_2489
timestamp 1569139307
transform 1 0 648 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_2490
timestamp 1569139307
transform 1 0 1096 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2491
timestamp 1569139307
transform 1 0 1032 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2492
timestamp 1569139307
transform 1 0 1096 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2493
timestamp 1569139307
transform 1 0 1032 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2494
timestamp 1569139307
transform 1 0 968 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2495
timestamp 1569139307
transform 1 0 1160 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2496
timestamp 1569139307
transform 1 0 1160 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2497
timestamp 1569139307
transform 1 0 1096 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2498
timestamp 1569139307
transform 1 0 1096 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2499
timestamp 1569139307
transform 1 0 1224 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2500
timestamp 1569139307
transform 1 0 1224 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2501
timestamp 1569139307
transform 1 0 1224 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2502
timestamp 1569139307
transform 1 0 1160 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2503
timestamp 1569139307
transform 1 0 1224 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2504
timestamp 1569139307
transform 1 0 1224 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2505
timestamp 1569139307
transform 1 0 968 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2506
timestamp 1569139307
transform 1 0 968 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2507
timestamp 1569139307
transform 1 0 968 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2508
timestamp 1569139307
transform 1 0 1032 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2509
timestamp 1569139307
transform 1 0 968 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2510
timestamp 1569139307
transform 1 0 1160 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2511
timestamp 1569139307
transform 1 0 1160 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2512
timestamp 1569139307
transform 1 0 1032 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2513
timestamp 1569139307
transform 1 0 1096 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2514
timestamp 1569139307
transform 1 0 1032 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2515
timestamp 1569139307
transform 1 0 712 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2516
timestamp 1569139307
transform 1 0 840 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2517
timestamp 1569139307
transform 1 0 840 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2518
timestamp 1569139307
transform 1 0 776 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2519
timestamp 1569139307
transform 1 0 776 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2520
timestamp 1569139307
transform 1 0 840 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2521
timestamp 1569139307
transform 1 0 712 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2522
timestamp 1569139307
transform 1 0 904 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2523
timestamp 1569139307
transform 1 0 904 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2524
timestamp 1569139307
transform 1 0 712 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2525
timestamp 1569139307
transform 1 0 904 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2526
timestamp 1569139307
transform 1 0 904 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2527
timestamp 1569139307
transform 1 0 776 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2528
timestamp 1569139307
transform 1 0 712 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2529
timestamp 1569139307
transform 1 0 840 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2530
timestamp 1569139307
transform 1 0 904 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2531
timestamp 1569139307
transform 1 0 776 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2532
timestamp 1569139307
transform 1 0 712 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2533
timestamp 1569139307
transform 1 0 776 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2534
timestamp 1569139307
transform 1 0 840 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2535
timestamp 1569139307
transform 1 0 840 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2536
timestamp 1569139307
transform 1 0 840 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2537
timestamp 1569139307
transform 1 0 712 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2538
timestamp 1569139307
transform 1 0 840 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2539
timestamp 1569139307
transform 1 0 840 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2540
timestamp 1569139307
transform 1 0 712 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2541
timestamp 1569139307
transform 1 0 712 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2542
timestamp 1569139307
transform 1 0 776 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2543
timestamp 1569139307
transform 1 0 776 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2544
timestamp 1569139307
transform 1 0 776 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2545
timestamp 1569139307
transform 1 0 904 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2546
timestamp 1569139307
transform 1 0 776 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2547
timestamp 1569139307
transform 1 0 904 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2548
timestamp 1569139307
transform 1 0 904 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2549
timestamp 1569139307
transform 1 0 712 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2550
timestamp 1569139307
transform 1 0 904 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2551
timestamp 1569139307
transform 1 0 1032 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2552
timestamp 1569139307
transform 1 0 1032 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2553
timestamp 1569139307
transform 1 0 1160 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2554
timestamp 1569139307
transform 1 0 1160 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2555
timestamp 1569139307
transform 1 0 1224 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2556
timestamp 1569139307
transform 1 0 1160 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2557
timestamp 1569139307
transform 1 0 1096 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2558
timestamp 1569139307
transform 1 0 1160 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2559
timestamp 1569139307
transform 1 0 1224 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2560
timestamp 1569139307
transform 1 0 1096 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2561
timestamp 1569139307
transform 1 0 1224 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2562
timestamp 1569139307
transform 1 0 1096 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2563
timestamp 1569139307
transform 1 0 1224 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2564
timestamp 1569139307
transform 1 0 1096 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2565
timestamp 1569139307
transform 1 0 968 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2566
timestamp 1569139307
transform 1 0 968 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2567
timestamp 1569139307
transform 1 0 968 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2568
timestamp 1569139307
transform 1 0 968 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2569
timestamp 1569139307
transform 1 0 1032 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2570
timestamp 1569139307
transform 1 0 1032 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2571
timestamp 1569139307
transform 1 0 392 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2572
timestamp 1569139307
transform 1 0 584 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2573
timestamp 1569139307
transform 1 0 584 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2574
timestamp 1569139307
transform 1 0 392 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2575
timestamp 1569139307
transform 1 0 456 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2576
timestamp 1569139307
transform 1 0 584 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2577
timestamp 1569139307
transform 1 0 392 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2578
timestamp 1569139307
transform 1 0 520 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2579
timestamp 1569139307
transform 1 0 520 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2580
timestamp 1569139307
transform 1 0 392 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2581
timestamp 1569139307
transform 1 0 584 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2582
timestamp 1569139307
transform 1 0 520 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2583
timestamp 1569139307
transform 1 0 456 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2584
timestamp 1569139307
transform 1 0 392 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2585
timestamp 1569139307
transform 1 0 584 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2586
timestamp 1569139307
transform 1 0 520 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2587
timestamp 1569139307
transform 1 0 456 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2588
timestamp 1569139307
transform 1 0 520 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2589
timestamp 1569139307
transform 1 0 456 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2590
timestamp 1569139307
transform 1 0 456 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2591
timestamp 1569139307
transform 1 0 200 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2592
timestamp 1569139307
transform 1 0 72 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2593
timestamp 1569139307
transform 1 0 200 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2594
timestamp 1569139307
transform 1 0 72 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2595
timestamp 1569139307
transform 1 0 72 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2596
timestamp 1569139307
transform 1 0 136 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2597
timestamp 1569139307
transform 1 0 264 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2598
timestamp 1569139307
transform 1 0 136 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2599
timestamp 1569139307
transform 1 0 72 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2600
timestamp 1569139307
transform 1 0 328 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2601
timestamp 1569139307
transform 1 0 264 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2602
timestamp 1569139307
transform 1 0 136 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2603
timestamp 1569139307
transform 1 0 72 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2604
timestamp 1569139307
transform 1 0 136 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2605
timestamp 1569139307
transform 1 0 264 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2606
timestamp 1569139307
transform 1 0 264 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2607
timestamp 1569139307
transform 1 0 136 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2608
timestamp 1569139307
transform 1 0 264 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2609
timestamp 1569139307
transform 1 0 200 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2610
timestamp 1569139307
transform 1 0 328 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2611
timestamp 1569139307
transform 1 0 328 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2612
timestamp 1569139307
transform 1 0 200 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2613
timestamp 1569139307
transform 1 0 200 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2614
timestamp 1569139307
transform 1 0 328 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2615
timestamp 1569139307
transform 1 0 328 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2616
timestamp 1569139307
transform 1 0 136 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2617
timestamp 1569139307
transform 1 0 136 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2618
timestamp 1569139307
transform 1 0 136 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2619
timestamp 1569139307
transform 1 0 136 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2620
timestamp 1569139307
transform 1 0 72 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2621
timestamp 1569139307
transform 1 0 72 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2622
timestamp 1569139307
transform 1 0 200 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2623
timestamp 1569139307
transform 1 0 200 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2624
timestamp 1569139307
transform 1 0 200 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2625
timestamp 1569139307
transform 1 0 200 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2626
timestamp 1569139307
transform 1 0 72 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2627
timestamp 1569139307
transform 1 0 264 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2628
timestamp 1569139307
transform 1 0 264 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2629
timestamp 1569139307
transform 1 0 264 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2630
timestamp 1569139307
transform 1 0 264 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2631
timestamp 1569139307
transform 1 0 328 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2632
timestamp 1569139307
transform 1 0 328 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2633
timestamp 1569139307
transform 1 0 328 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2634
timestamp 1569139307
transform 1 0 328 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2635
timestamp 1569139307
transform 1 0 72 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2636
timestamp 1569139307
transform 1 0 520 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2637
timestamp 1569139307
transform 1 0 520 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2638
timestamp 1569139307
transform 1 0 456 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2639
timestamp 1569139307
transform 1 0 456 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2640
timestamp 1569139307
transform 1 0 392 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2641
timestamp 1569139307
transform 1 0 392 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2642
timestamp 1569139307
transform 1 0 392 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2643
timestamp 1569139307
transform 1 0 392 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2644
timestamp 1569139307
transform 1 0 456 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2645
timestamp 1569139307
transform 1 0 456 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2646
timestamp 1569139307
transform 1 0 584 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2647
timestamp 1569139307
transform 1 0 584 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2648
timestamp 1569139307
transform 1 0 584 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2649
timestamp 1569139307
transform 1 0 520 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2650
timestamp 1569139307
transform 1 0 520 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2651
timestamp 1569139307
transform 1 0 584 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2652
timestamp 1569139307
transform 1 0 584 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2653
timestamp 1569139307
transform 1 0 392 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2654
timestamp 1569139307
transform 1 0 520 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2655
timestamp 1569139307
transform 1 0 520 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2656
timestamp 1569139307
transform 1 0 584 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2657
timestamp 1569139307
transform 1 0 520 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2658
timestamp 1569139307
transform 1 0 456 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2659
timestamp 1569139307
transform 1 0 456 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2660
timestamp 1569139307
transform 1 0 584 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2661
timestamp 1569139307
transform 1 0 520 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2662
timestamp 1569139307
transform 1 0 392 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2663
timestamp 1569139307
transform 1 0 584 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2664
timestamp 1569139307
transform 1 0 392 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2665
timestamp 1569139307
transform 1 0 456 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2666
timestamp 1569139307
transform 1 0 456 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2667
timestamp 1569139307
transform 1 0 392 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2668
timestamp 1569139307
transform 1 0 136 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2669
timestamp 1569139307
transform 1 0 328 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2670
timestamp 1569139307
transform 1 0 264 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2671
timestamp 1569139307
transform 1 0 264 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2672
timestamp 1569139307
transform 1 0 72 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2673
timestamp 1569139307
transform 1 0 200 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2674
timestamp 1569139307
transform 1 0 328 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2675
timestamp 1569139307
transform 1 0 136 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2676
timestamp 1569139307
transform 1 0 328 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2677
timestamp 1569139307
transform 1 0 72 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2678
timestamp 1569139307
transform 1 0 264 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2679
timestamp 1569139307
transform 1 0 328 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2680
timestamp 1569139307
transform 1 0 136 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2681
timestamp 1569139307
transform 1 0 264 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2682
timestamp 1569139307
transform 1 0 136 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2683
timestamp 1569139307
transform 1 0 72 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2684
timestamp 1569139307
transform 1 0 200 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2685
timestamp 1569139307
transform 1 0 200 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2686
timestamp 1569139307
transform 1 0 200 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2687
timestamp 1569139307
transform 1 0 72 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2688
timestamp 1569139307
transform 1 0 264 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2689
timestamp 1569139307
transform 1 0 264 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2690
timestamp 1569139307
transform 1 0 200 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2691
timestamp 1569139307
transform 1 0 136 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2692
timestamp 1569139307
transform 1 0 136 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2693
timestamp 1569139307
transform 1 0 136 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2694
timestamp 1569139307
transform 1 0 136 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2695
timestamp 1569139307
transform 1 0 72 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2696
timestamp 1569139307
transform 1 0 328 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2697
timestamp 1569139307
transform 1 0 328 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2698
timestamp 1569139307
transform 1 0 328 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2699
timestamp 1569139307
transform 1 0 328 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2700
timestamp 1569139307
transform 1 0 72 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2701
timestamp 1569139307
transform 1 0 72 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2702
timestamp 1569139307
transform 1 0 264 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2703
timestamp 1569139307
transform 1 0 200 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2704
timestamp 1569139307
transform 1 0 200 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2705
timestamp 1569139307
transform 1 0 200 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2706
timestamp 1569139307
transform 1 0 264 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2707
timestamp 1569139307
transform 1 0 72 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2708
timestamp 1569139307
transform 1 0 392 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2709
timestamp 1569139307
transform 1 0 392 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2710
timestamp 1569139307
transform 1 0 392 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2711
timestamp 1569139307
transform 1 0 392 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2712
timestamp 1569139307
transform 1 0 456 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2713
timestamp 1569139307
transform 1 0 456 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2714
timestamp 1569139307
transform 1 0 456 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2715
timestamp 1569139307
transform 1 0 456 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2716
timestamp 1569139307
transform 1 0 520 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2717
timestamp 1569139307
transform 1 0 520 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2718
timestamp 1569139307
transform 1 0 520 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2719
timestamp 1569139307
transform 1 0 520 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2720
timestamp 1569139307
transform 1 0 584 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2721
timestamp 1569139307
transform 1 0 584 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2722
timestamp 1569139307
transform 1 0 584 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2723
timestamp 1569139307
transform 1 0 584 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2724
timestamp 1569139307
transform 1 0 1096 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2725
timestamp 1569139307
transform 1 0 1160 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2726
timestamp 1569139307
transform 1 0 968 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2727
timestamp 1569139307
transform 1 0 1096 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2728
timestamp 1569139307
transform 1 0 1224 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2729
timestamp 1569139307
transform 1 0 968 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2730
timestamp 1569139307
transform 1 0 1096 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2731
timestamp 1569139307
transform 1 0 1224 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2732
timestamp 1569139307
transform 1 0 1096 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2733
timestamp 1569139307
transform 1 0 1224 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2734
timestamp 1569139307
transform 1 0 968 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2735
timestamp 1569139307
transform 1 0 968 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2736
timestamp 1569139307
transform 1 0 1160 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2737
timestamp 1569139307
transform 1 0 1160 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2738
timestamp 1569139307
transform 1 0 1032 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2739
timestamp 1569139307
transform 1 0 1032 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2740
timestamp 1569139307
transform 1 0 1032 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2741
timestamp 1569139307
transform 1 0 1032 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2742
timestamp 1569139307
transform 1 0 1224 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2743
timestamp 1569139307
transform 1 0 1160 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2744
timestamp 1569139307
transform 1 0 712 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2745
timestamp 1569139307
transform 1 0 840 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2746
timestamp 1569139307
transform 1 0 776 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2747
timestamp 1569139307
transform 1 0 776 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2748
timestamp 1569139307
transform 1 0 904 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2749
timestamp 1569139307
transform 1 0 776 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2750
timestamp 1569139307
transform 1 0 904 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2751
timestamp 1569139307
transform 1 0 840 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2752
timestamp 1569139307
transform 1 0 840 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2753
timestamp 1569139307
transform 1 0 840 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2754
timestamp 1569139307
transform 1 0 904 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2755
timestamp 1569139307
transform 1 0 776 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2756
timestamp 1569139307
transform 1 0 904 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2757
timestamp 1569139307
transform 1 0 712 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2758
timestamp 1569139307
transform 1 0 712 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2759
timestamp 1569139307
transform 1 0 712 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2760
timestamp 1569139307
transform 1 0 904 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2761
timestamp 1569139307
transform 1 0 904 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2762
timestamp 1569139307
transform 1 0 904 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2763
timestamp 1569139307
transform 1 0 776 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2764
timestamp 1569139307
transform 1 0 840 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2765
timestamp 1569139307
transform 1 0 776 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2766
timestamp 1569139307
transform 1 0 776 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2767
timestamp 1569139307
transform 1 0 776 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2768
timestamp 1569139307
transform 1 0 840 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2769
timestamp 1569139307
transform 1 0 712 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2770
timestamp 1569139307
transform 1 0 712 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2771
timestamp 1569139307
transform 1 0 840 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2772
timestamp 1569139307
transform 1 0 712 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2773
timestamp 1569139307
transform 1 0 712 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2774
timestamp 1569139307
transform 1 0 904 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2775
timestamp 1569139307
transform 1 0 840 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2776
timestamp 1569139307
transform 1 0 968 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2777
timestamp 1569139307
transform 1 0 968 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2778
timestamp 1569139307
transform 1 0 968 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2779
timestamp 1569139307
transform 1 0 968 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2780
timestamp 1569139307
transform 1 0 1032 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2781
timestamp 1569139307
transform 1 0 1032 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2782
timestamp 1569139307
transform 1 0 1032 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2783
timestamp 1569139307
transform 1 0 1032 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2784
timestamp 1569139307
transform 1 0 1096 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2785
timestamp 1569139307
transform 1 0 1096 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2786
timestamp 1569139307
transform 1 0 1096 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2787
timestamp 1569139307
transform 1 0 1096 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2788
timestamp 1569139307
transform 1 0 1160 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2789
timestamp 1569139307
transform 1 0 1160 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2790
timestamp 1569139307
transform 1 0 1160 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2791
timestamp 1569139307
transform 1 0 1160 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2792
timestamp 1569139307
transform 1 0 1224 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2793
timestamp 1569139307
transform 1 0 1224 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2794
timestamp 1569139307
transform 1 0 1224 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2795
timestamp 1569139307
transform 1 0 1224 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2796
timestamp 1569139307
transform 1 0 456 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2797
timestamp 1569139307
transform 1 0 1096 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2798
timestamp 1569139307
transform 1 0 136 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2799
timestamp 1569139307
transform 1 0 776 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2800
timestamp 1569139307
transform 1 0 520 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2801
timestamp 1569139307
transform 1 0 1160 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2802
timestamp 1569139307
transform 1 0 200 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2803
timestamp 1569139307
transform 1 0 840 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2804
timestamp 1569139307
transform 1 0 264 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2805
timestamp 1569139307
transform 1 0 904 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2806
timestamp 1569139307
transform 1 0 328 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2807
timestamp 1569139307
transform 1 0 968 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2808
timestamp 1569139307
transform 1 0 392 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2809
timestamp 1569139307
transform 1 0 1032 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2810
timestamp 1569139307
transform 1 0 648 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2811
timestamp 1569139307
transform 1 0 584 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2812
timestamp 1569139307
transform 1 0 1224 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2813
timestamp 1569139307
transform 1 0 648 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2814
timestamp 1569139307
transform 1 0 648 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2815
timestamp 1569139307
transform 1 0 648 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2816
timestamp 1569139307
transform 1 0 648 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2817
timestamp 1569139307
transform 1 0 648 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2818
timestamp 1569139307
transform 1 0 648 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2819
timestamp 1569139307
transform 1 0 648 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2820
timestamp 1569139307
transform 1 0 648 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2821
timestamp 1569139307
transform 1 0 648 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2822
timestamp 1569139307
transform 1 0 648 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2823
timestamp 1569139307
transform 1 0 648 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2824
timestamp 1569139307
transform 1 0 648 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2825
timestamp 1569139307
transform 1 0 72 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2826
timestamp 1569139307
transform 1 0 712 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2827
timestamp 1569139307
transform 1 0 648 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2828
timestamp 1569139307
transform 1 0 648 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2829
timestamp 1569139307
transform 1 0 648 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2830
timestamp 1569139307
transform 1 0 648 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2831
timestamp 1569139307
transform 1 0 648 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2832
timestamp 1569139307
transform 1 0 2376 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2833
timestamp 1569139307
transform 1 0 2440 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2834
timestamp 1569139307
transform 1 0 2376 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2835
timestamp 1569139307
transform 1 0 2376 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2836
timestamp 1569139307
transform 1 0 2376 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2837
timestamp 1569139307
transform 1 0 2376 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2838
timestamp 1569139307
transform 1 0 2376 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2839
timestamp 1569139307
transform 1 0 2376 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2840
timestamp 1569139307
transform 1 0 2440 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2841
timestamp 1569139307
transform 1 0 2440 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2842
timestamp 1569139307
transform 1 0 2312 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2843
timestamp 1569139307
transform 1 0 2312 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2844
timestamp 1569139307
transform 1 0 2312 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2845
timestamp 1569139307
transform 1 0 2312 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2846
timestamp 1569139307
transform 1 0 2312 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2847
timestamp 1569139307
transform 1 0 2440 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2848
timestamp 1569139307
transform 1 0 2440 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2849
timestamp 1569139307
transform 1 0 2440 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2850
timestamp 1569139307
transform 1 0 2440 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2851
timestamp 1569139307
transform 1 0 2440 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2852
timestamp 1569139307
transform 1 0 2312 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2853
timestamp 1569139307
transform 1 0 2312 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2854
timestamp 1569139307
transform 1 0 2312 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2855
timestamp 1569139307
transform 1 0 2312 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2856
timestamp 1569139307
transform 1 0 2440 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2857
timestamp 1569139307
transform 1 0 2376 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2858
timestamp 1569139307
transform 1 0 2376 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2859
timestamp 1569139307
transform 1 0 1352 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2860
timestamp 1569139307
transform 1 0 1352 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2861
timestamp 1569139307
transform 1 0 1352 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2862
timestamp 1569139307
transform 1 0 1352 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2863
timestamp 1569139307
transform 1 0 1288 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2864
timestamp 1569139307
transform 1 0 1352 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2865
timestamp 1569139307
transform 1 0 1352 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2866
timestamp 1569139307
transform 1 0 1416 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2867
timestamp 1569139307
transform 1 0 1352 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2868
timestamp 1569139307
transform 1 0 1416 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2869
timestamp 1569139307
transform 1 0 1416 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2870
timestamp 1569139307
transform 1 0 1416 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2871
timestamp 1569139307
transform 1 0 1416 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2872
timestamp 1569139307
transform 1 0 1480 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2873
timestamp 1569139307
transform 1 0 1480 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2874
timestamp 1569139307
transform 1 0 1288 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2875
timestamp 1569139307
transform 1 0 1480 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2876
timestamp 1569139307
transform 1 0 1480 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2877
timestamp 1569139307
transform 1 0 1352 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2878
timestamp 1569139307
transform 1 0 1288 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2879
timestamp 1569139307
transform 1 0 1416 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2880
timestamp 1569139307
transform 1 0 1416 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2881
timestamp 1569139307
transform 1 0 1416 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2882
timestamp 1569139307
transform 1 0 1416 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2883
timestamp 1569139307
transform 1 0 1288 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2884
timestamp 1569139307
transform 1 0 1480 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_2885
timestamp 1569139307
transform 1 0 1480 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_2886
timestamp 1569139307
transform 1 0 1480 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_2887
timestamp 1569139307
transform 1 0 1480 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_2888
timestamp 1569139307
transform 1 0 1352 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2889
timestamp 1569139307
transform 1 0 1288 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2890
timestamp 1569139307
transform 1 0 1480 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_2891
timestamp 1569139307
transform 1 0 1288 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_2892
timestamp 1569139307
transform 1 0 1288 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_2893
timestamp 1569139307
transform 1 0 1288 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_2894
timestamp 1569139307
transform 1 0 1288 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_2895
timestamp 1569139307
transform 1 0 1352 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2896
timestamp 1569139307
transform 1 0 1480 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2897
timestamp 1569139307
transform 1 0 1480 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2898
timestamp 1569139307
transform 1 0 1416 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2899
timestamp 1569139307
transform 1 0 1416 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2900
timestamp 1569139307
transform 1 0 1480 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2901
timestamp 1569139307
transform 1 0 1480 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2902
timestamp 1569139307
transform 1 0 1352 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2903
timestamp 1569139307
transform 1 0 1352 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2904
timestamp 1569139307
transform 1 0 1352 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2905
timestamp 1569139307
transform 1 0 1352 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2906
timestamp 1569139307
transform 1 0 1352 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2907
timestamp 1569139307
transform 1 0 1480 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2908
timestamp 1569139307
transform 1 0 1352 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2909
timestamp 1569139307
transform 1 0 1480 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2910
timestamp 1569139307
transform 1 0 1352 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2911
timestamp 1569139307
transform 1 0 1416 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2912
timestamp 1569139307
transform 1 0 1416 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2913
timestamp 1569139307
transform 1 0 1480 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2914
timestamp 1569139307
transform 1 0 1416 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2915
timestamp 1569139307
transform 1 0 1416 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2916
timestamp 1569139307
transform 1 0 1416 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2917
timestamp 1569139307
transform 1 0 1288 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2918
timestamp 1569139307
transform 1 0 1288 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2919
timestamp 1569139307
transform 1 0 1416 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2920
timestamp 1569139307
transform 1 0 1288 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2921
timestamp 1569139307
transform 1 0 1288 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2922
timestamp 1569139307
transform 1 0 1288 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2923
timestamp 1569139307
transform 1 0 1288 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2924
timestamp 1569139307
transform 1 0 1288 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2925
timestamp 1569139307
transform 1 0 1288 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2926
timestamp 1569139307
transform 1 0 1480 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2927
timestamp 1569139307
transform 1 0 2376 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2928
timestamp 1569139307
transform 1 0 2312 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2929
timestamp 1569139307
transform 1 0 2312 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2930
timestamp 1569139307
transform 1 0 2312 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2931
timestamp 1569139307
transform 1 0 2312 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2932
timestamp 1569139307
transform 1 0 2312 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2933
timestamp 1569139307
transform 1 0 2312 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2934
timestamp 1569139307
transform 1 0 2376 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2935
timestamp 1569139307
transform 1 0 2376 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2936
timestamp 1569139307
transform 1 0 2376 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2937
timestamp 1569139307
transform 1 0 2376 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2938
timestamp 1569139307
transform 1 0 2376 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2939
timestamp 1569139307
transform 1 0 2440 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_2940
timestamp 1569139307
transform 1 0 2440 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_2941
timestamp 1569139307
transform 1 0 2440 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_2942
timestamp 1569139307
transform 1 0 2440 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_2943
timestamp 1569139307
transform 1 0 2440 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_2944
timestamp 1569139307
transform 1 0 2312 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2945
timestamp 1569139307
transform 1 0 2440 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_2946
timestamp 1569139307
transform 1 0 2376 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2947
timestamp 1569139307
transform 1 0 2312 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2948
timestamp 1569139307
transform 1 0 2440 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_2949
timestamp 1569139307
transform 1 0 2376 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2950
timestamp 1569139307
transform 1 0 2440 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_2951
timestamp 1569139307
transform 1 0 1416 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2952
timestamp 1569139307
transform 1 0 1480 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2953
timestamp 1569139307
transform 1 0 2312 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2954
timestamp 1569139307
transform 1 0 2376 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2955
timestamp 1569139307
transform 1 0 2440 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2956
timestamp 1569139307
transform 1 0 1288 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2957
timestamp 1569139307
transform 1 0 1352 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_2958
timestamp 1569139307
transform 1 0 4680 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2959
timestamp 1569139307
transform 1 0 4744 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2960
timestamp 1569139307
transform 1 0 4872 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2961
timestamp 1569139307
transform 1 0 4872 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2962
timestamp 1569139307
transform 1 0 4744 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2963
timestamp 1569139307
transform 1 0 4680 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2964
timestamp 1569139307
transform 1 0 4680 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2965
timestamp 1569139307
transform 1 0 4744 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2966
timestamp 1569139307
transform 1 0 4680 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2967
timestamp 1569139307
transform 1 0 4808 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2968
timestamp 1569139307
transform 1 0 4744 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2969
timestamp 1569139307
transform 1 0 4872 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2970
timestamp 1569139307
transform 1 0 4808 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2971
timestamp 1569139307
transform 1 0 4808 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2972
timestamp 1569139307
transform 1 0 4808 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2973
timestamp 1569139307
transform 1 0 4872 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2974
timestamp 1569139307
transform 1 0 4616 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2975
timestamp 1569139307
transform 1 0 4488 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2976
timestamp 1569139307
transform 1 0 4424 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2977
timestamp 1569139307
transform 1 0 4424 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2978
timestamp 1569139307
transform 1 0 4488 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2979
timestamp 1569139307
transform 1 0 4616 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2980
timestamp 1569139307
transform 1 0 4488 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2981
timestamp 1569139307
transform 1 0 4616 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2982
timestamp 1569139307
transform 1 0 4616 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2983
timestamp 1569139307
transform 1 0 4552 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2984
timestamp 1569139307
transform 1 0 4552 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_2985
timestamp 1569139307
transform 1 0 4552 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2986
timestamp 1569139307
transform 1 0 4424 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2987
timestamp 1569139307
transform 1 0 4552 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_2988
timestamp 1569139307
transform 1 0 4424 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_2989
timestamp 1569139307
transform 1 0 4488 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_2990
timestamp 1569139307
transform 1 0 4616 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_2991
timestamp 1569139307
transform 1 0 4552 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2992
timestamp 1569139307
transform 1 0 4424 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2993
timestamp 1569139307
transform 1 0 4616 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_2994
timestamp 1569139307
transform 1 0 4488 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_2995
timestamp 1569139307
transform 1 0 4616 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2996
timestamp 1569139307
transform 1 0 4616 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2997
timestamp 1569139307
transform 1 0 4488 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_2998
timestamp 1569139307
transform 1 0 4488 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_2999
timestamp 1569139307
transform 1 0 4488 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3000
timestamp 1569139307
transform 1 0 4552 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3001
timestamp 1569139307
transform 1 0 4424 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3002
timestamp 1569139307
transform 1 0 4424 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3003
timestamp 1569139307
transform 1 0 4488 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3004
timestamp 1569139307
transform 1 0 4424 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3005
timestamp 1569139307
transform 1 0 4552 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3006
timestamp 1569139307
transform 1 0 4424 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3007
timestamp 1569139307
transform 1 0 4552 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3008
timestamp 1569139307
transform 1 0 4552 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3009
timestamp 1569139307
transform 1 0 4616 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3010
timestamp 1569139307
transform 1 0 4872 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3011
timestamp 1569139307
transform 1 0 4744 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3012
timestamp 1569139307
transform 1 0 4872 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3013
timestamp 1569139307
transform 1 0 4744 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3014
timestamp 1569139307
transform 1 0 4872 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3015
timestamp 1569139307
transform 1 0 4808 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3016
timestamp 1569139307
transform 1 0 4744 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3017
timestamp 1569139307
transform 1 0 4680 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3018
timestamp 1569139307
transform 1 0 4808 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3019
timestamp 1569139307
transform 1 0 4680 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3020
timestamp 1569139307
transform 1 0 4808 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3021
timestamp 1569139307
transform 1 0 4808 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3022
timestamp 1569139307
transform 1 0 4680 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3023
timestamp 1569139307
transform 1 0 4872 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3024
timestamp 1569139307
transform 1 0 4872 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3025
timestamp 1569139307
transform 1 0 4680 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3026
timestamp 1569139307
transform 1 0 4680 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3027
timestamp 1569139307
transform 1 0 4744 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3028
timestamp 1569139307
transform 1 0 4808 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3029
timestamp 1569139307
transform 1 0 4744 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3030
timestamp 1569139307
transform 1 0 4104 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3031
timestamp 1569139307
transform 1 0 4232 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3032
timestamp 1569139307
transform 1 0 4104 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3033
timestamp 1569139307
transform 1 0 4232 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3034
timestamp 1569139307
transform 1 0 4168 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3035
timestamp 1569139307
transform 1 0 4296 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3036
timestamp 1569139307
transform 1 0 4296 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3037
timestamp 1569139307
transform 1 0 4168 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3038
timestamp 1569139307
transform 1 0 4296 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3039
timestamp 1569139307
transform 1 0 4104 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3040
timestamp 1569139307
transform 1 0 4232 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3041
timestamp 1569139307
transform 1 0 4168 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3042
timestamp 1569139307
transform 1 0 4168 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3043
timestamp 1569139307
transform 1 0 4232 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3044
timestamp 1569139307
transform 1 0 4104 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3045
timestamp 1569139307
transform 1 0 4296 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3046
timestamp 1569139307
transform 1 0 3848 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3047
timestamp 1569139307
transform 1 0 3976 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3048
timestamp 1569139307
transform 1 0 3912 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3049
timestamp 1569139307
transform 1 0 3976 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3050
timestamp 1569139307
transform 1 0 3784 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3051
timestamp 1569139307
transform 1 0 3848 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3052
timestamp 1569139307
transform 1 0 3976 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3053
timestamp 1569139307
transform 1 0 3784 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3054
timestamp 1569139307
transform 1 0 4040 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3055
timestamp 1569139307
transform 1 0 3976 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3056
timestamp 1569139307
transform 1 0 3912 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3057
timestamp 1569139307
transform 1 0 3912 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3058
timestamp 1569139307
transform 1 0 3848 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3059
timestamp 1569139307
transform 1 0 3848 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3060
timestamp 1569139307
transform 1 0 3784 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3061
timestamp 1569139307
transform 1 0 4040 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3062
timestamp 1569139307
transform 1 0 4040 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3063
timestamp 1569139307
transform 1 0 3912 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3064
timestamp 1569139307
transform 1 0 4040 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3065
timestamp 1569139307
transform 1 0 3784 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3066
timestamp 1569139307
transform 1 0 3912 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3067
timestamp 1569139307
transform 1 0 3784 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3068
timestamp 1569139307
transform 1 0 3848 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3069
timestamp 1569139307
transform 1 0 4040 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3070
timestamp 1569139307
transform 1 0 3848 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3071
timestamp 1569139307
transform 1 0 3976 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3072
timestamp 1569139307
transform 1 0 3976 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3073
timestamp 1569139307
transform 1 0 3848 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3074
timestamp 1569139307
transform 1 0 3976 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3075
timestamp 1569139307
transform 1 0 3912 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3076
timestamp 1569139307
transform 1 0 3784 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3077
timestamp 1569139307
transform 1 0 3976 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3078
timestamp 1569139307
transform 1 0 4040 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3079
timestamp 1569139307
transform 1 0 3784 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3080
timestamp 1569139307
transform 1 0 3912 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3081
timestamp 1569139307
transform 1 0 4040 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3082
timestamp 1569139307
transform 1 0 3784 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3083
timestamp 1569139307
transform 1 0 3848 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3084
timestamp 1569139307
transform 1 0 4040 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3085
timestamp 1569139307
transform 1 0 4040 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3086
timestamp 1569139307
transform 1 0 3912 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3087
timestamp 1569139307
transform 1 0 3848 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3088
timestamp 1569139307
transform 1 0 3784 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3089
timestamp 1569139307
transform 1 0 3976 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3090
timestamp 1569139307
transform 1 0 3912 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3091
timestamp 1569139307
transform 1 0 4104 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3092
timestamp 1569139307
transform 1 0 4104 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3093
timestamp 1569139307
transform 1 0 4232 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3094
timestamp 1569139307
transform 1 0 4104 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3095
timestamp 1569139307
transform 1 0 4232 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3096
timestamp 1569139307
transform 1 0 4168 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3097
timestamp 1569139307
transform 1 0 4296 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3098
timestamp 1569139307
transform 1 0 4168 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3099
timestamp 1569139307
transform 1 0 4232 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3100
timestamp 1569139307
transform 1 0 4296 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3101
timestamp 1569139307
transform 1 0 4168 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3102
timestamp 1569139307
transform 1 0 4104 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3103
timestamp 1569139307
transform 1 0 4104 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3104
timestamp 1569139307
transform 1 0 4168 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3105
timestamp 1569139307
transform 1 0 4168 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3106
timestamp 1569139307
transform 1 0 4232 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3107
timestamp 1569139307
transform 1 0 4232 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3108
timestamp 1569139307
transform 1 0 4296 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3109
timestamp 1569139307
transform 1 0 4296 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3110
timestamp 1569139307
transform 1 0 4296 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3111
timestamp 1569139307
transform 1 0 4168 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3112
timestamp 1569139307
transform 1 0 4232 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3113
timestamp 1569139307
transform 1 0 4104 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3114
timestamp 1569139307
transform 1 0 4104 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3115
timestamp 1569139307
transform 1 0 4232 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3116
timestamp 1569139307
transform 1 0 4168 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3117
timestamp 1569139307
transform 1 0 4232 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3118
timestamp 1569139307
transform 1 0 4104 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3119
timestamp 1569139307
transform 1 0 4104 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3120
timestamp 1569139307
transform 1 0 4168 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3121
timestamp 1569139307
transform 1 0 4104 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3122
timestamp 1569139307
transform 1 0 4296 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3123
timestamp 1569139307
transform 1 0 4232 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3124
timestamp 1569139307
transform 1 0 4168 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3125
timestamp 1569139307
transform 1 0 4232 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3126
timestamp 1569139307
transform 1 0 4296 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3127
timestamp 1569139307
transform 1 0 4296 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3128
timestamp 1569139307
transform 1 0 4296 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3129
timestamp 1569139307
transform 1 0 4296 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3130
timestamp 1569139307
transform 1 0 4168 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3131
timestamp 1569139307
transform 1 0 3848 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3132
timestamp 1569139307
transform 1 0 4040 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3133
timestamp 1569139307
transform 1 0 3912 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3134
timestamp 1569139307
transform 1 0 3848 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3135
timestamp 1569139307
transform 1 0 3784 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3136
timestamp 1569139307
transform 1 0 3784 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3137
timestamp 1569139307
transform 1 0 3848 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3138
timestamp 1569139307
transform 1 0 3784 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3139
timestamp 1569139307
transform 1 0 3912 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3140
timestamp 1569139307
transform 1 0 3976 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3141
timestamp 1569139307
transform 1 0 3912 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3142
timestamp 1569139307
transform 1 0 3848 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3143
timestamp 1569139307
transform 1 0 3976 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3144
timestamp 1569139307
transform 1 0 3976 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3145
timestamp 1569139307
transform 1 0 3784 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3146
timestamp 1569139307
transform 1 0 3976 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3147
timestamp 1569139307
transform 1 0 3976 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3148
timestamp 1569139307
transform 1 0 3784 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3149
timestamp 1569139307
transform 1 0 4040 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3150
timestamp 1569139307
transform 1 0 3912 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3151
timestamp 1569139307
transform 1 0 4040 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3152
timestamp 1569139307
transform 1 0 3848 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3153
timestamp 1569139307
transform 1 0 4040 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3154
timestamp 1569139307
transform 1 0 3912 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3155
timestamp 1569139307
transform 1 0 4040 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3156
timestamp 1569139307
transform 1 0 4040 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3157
timestamp 1569139307
transform 1 0 3784 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3158
timestamp 1569139307
transform 1 0 3784 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3159
timestamp 1569139307
transform 1 0 3784 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3160
timestamp 1569139307
transform 1 0 3784 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3161
timestamp 1569139307
transform 1 0 4040 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3162
timestamp 1569139307
transform 1 0 3912 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3163
timestamp 1569139307
transform 1 0 3912 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3164
timestamp 1569139307
transform 1 0 3976 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3165
timestamp 1569139307
transform 1 0 3976 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3166
timestamp 1569139307
transform 1 0 3976 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3167
timestamp 1569139307
transform 1 0 3848 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3168
timestamp 1569139307
transform 1 0 3976 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3169
timestamp 1569139307
transform 1 0 3976 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3170
timestamp 1569139307
transform 1 0 3848 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3171
timestamp 1569139307
transform 1 0 3848 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3172
timestamp 1569139307
transform 1 0 3848 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3173
timestamp 1569139307
transform 1 0 4040 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3174
timestamp 1569139307
transform 1 0 3912 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3175
timestamp 1569139307
transform 1 0 4040 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3176
timestamp 1569139307
transform 1 0 3912 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3177
timestamp 1569139307
transform 1 0 3912 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3178
timestamp 1569139307
transform 1 0 3848 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3179
timestamp 1569139307
transform 1 0 4040 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3180
timestamp 1569139307
transform 1 0 3784 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3181
timestamp 1569139307
transform 1 0 4232 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3182
timestamp 1569139307
transform 1 0 4232 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3183
timestamp 1569139307
transform 1 0 4232 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3184
timestamp 1569139307
transform 1 0 4104 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3185
timestamp 1569139307
transform 1 0 4296 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3186
timestamp 1569139307
transform 1 0 4296 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3187
timestamp 1569139307
transform 1 0 4296 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3188
timestamp 1569139307
transform 1 0 4104 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3189
timestamp 1569139307
transform 1 0 4168 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3190
timestamp 1569139307
transform 1 0 4104 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3191
timestamp 1569139307
transform 1 0 4104 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3192
timestamp 1569139307
transform 1 0 4296 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3193
timestamp 1569139307
transform 1 0 4296 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3194
timestamp 1569139307
transform 1 0 4168 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3195
timestamp 1569139307
transform 1 0 4168 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3196
timestamp 1569139307
transform 1 0 4232 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3197
timestamp 1569139307
transform 1 0 4232 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3198
timestamp 1569139307
transform 1 0 4168 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3199
timestamp 1569139307
transform 1 0 4168 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3200
timestamp 1569139307
transform 1 0 4104 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3201
timestamp 1569139307
transform 1 0 4744 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3202
timestamp 1569139307
transform 1 0 4744 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3203
timestamp 1569139307
transform 1 0 4744 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3204
timestamp 1569139307
transform 1 0 4744 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3205
timestamp 1569139307
transform 1 0 4744 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3206
timestamp 1569139307
transform 1 0 4808 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3207
timestamp 1569139307
transform 1 0 4808 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3208
timestamp 1569139307
transform 1 0 4808 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3209
timestamp 1569139307
transform 1 0 4872 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3210
timestamp 1569139307
transform 1 0 4680 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3211
timestamp 1569139307
transform 1 0 4808 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3212
timestamp 1569139307
transform 1 0 4808 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3213
timestamp 1569139307
transform 1 0 4872 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3214
timestamp 1569139307
transform 1 0 4680 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3215
timestamp 1569139307
transform 1 0 4680 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3216
timestamp 1569139307
transform 1 0 4872 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3217
timestamp 1569139307
transform 1 0 4680 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3218
timestamp 1569139307
transform 1 0 4680 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3219
timestamp 1569139307
transform 1 0 4872 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3220
timestamp 1569139307
transform 1 0 4872 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3221
timestamp 1569139307
transform 1 0 4552 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3222
timestamp 1569139307
transform 1 0 4488 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3223
timestamp 1569139307
transform 1 0 4488 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3224
timestamp 1569139307
transform 1 0 4488 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3225
timestamp 1569139307
transform 1 0 4616 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3226
timestamp 1569139307
transform 1 0 4552 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3227
timestamp 1569139307
transform 1 0 4424 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3228
timestamp 1569139307
transform 1 0 4616 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3229
timestamp 1569139307
transform 1 0 4616 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3230
timestamp 1569139307
transform 1 0 4616 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3231
timestamp 1569139307
transform 1 0 4616 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3232
timestamp 1569139307
transform 1 0 4552 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3233
timestamp 1569139307
transform 1 0 4552 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3234
timestamp 1569139307
transform 1 0 4552 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3235
timestamp 1569139307
transform 1 0 4424 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3236
timestamp 1569139307
transform 1 0 4424 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3237
timestamp 1569139307
transform 1 0 4424 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3238
timestamp 1569139307
transform 1 0 4424 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3239
timestamp 1569139307
transform 1 0 4488 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3240
timestamp 1569139307
transform 1 0 4488 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3241
timestamp 1569139307
transform 1 0 4552 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3242
timestamp 1569139307
transform 1 0 4616 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3243
timestamp 1569139307
transform 1 0 4616 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3244
timestamp 1569139307
transform 1 0 4424 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3245
timestamp 1569139307
transform 1 0 4424 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3246
timestamp 1569139307
transform 1 0 4424 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3247
timestamp 1569139307
transform 1 0 4424 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3248
timestamp 1569139307
transform 1 0 4424 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3249
timestamp 1569139307
transform 1 0 4488 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3250
timestamp 1569139307
transform 1 0 4616 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3251
timestamp 1569139307
transform 1 0 4616 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3252
timestamp 1569139307
transform 1 0 4616 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3253
timestamp 1569139307
transform 1 0 4488 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3254
timestamp 1569139307
transform 1 0 4488 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3255
timestamp 1569139307
transform 1 0 4488 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3256
timestamp 1569139307
transform 1 0 4488 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3257
timestamp 1569139307
transform 1 0 4552 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3258
timestamp 1569139307
transform 1 0 4552 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3259
timestamp 1569139307
transform 1 0 4552 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3260
timestamp 1569139307
transform 1 0 4552 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3261
timestamp 1569139307
transform 1 0 4680 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3262
timestamp 1569139307
transform 1 0 4680 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3263
timestamp 1569139307
transform 1 0 4744 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3264
timestamp 1569139307
transform 1 0 4744 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3265
timestamp 1569139307
transform 1 0 4808 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3266
timestamp 1569139307
transform 1 0 4808 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3267
timestamp 1569139307
transform 1 0 4872 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3268
timestamp 1569139307
transform 1 0 4872 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3269
timestamp 1569139307
transform 1 0 4680 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3270
timestamp 1569139307
transform 1 0 4680 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3271
timestamp 1569139307
transform 1 0 4680 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3272
timestamp 1569139307
transform 1 0 4744 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3273
timestamp 1569139307
transform 1 0 4744 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3274
timestamp 1569139307
transform 1 0 4744 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3275
timestamp 1569139307
transform 1 0 4808 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3276
timestamp 1569139307
transform 1 0 4808 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3277
timestamp 1569139307
transform 1 0 4808 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3278
timestamp 1569139307
transform 1 0 4872 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3279
timestamp 1569139307
transform 1 0 4872 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3280
timestamp 1569139307
transform 1 0 4872 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3281
timestamp 1569139307
transform 1 0 4360 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3282
timestamp 1569139307
transform 1 0 4360 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3283
timestamp 1569139307
transform 1 0 4360 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3284
timestamp 1569139307
transform 1 0 4360 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3285
timestamp 1569139307
transform 1 0 4360 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3286
timestamp 1569139307
transform 1 0 4360 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3287
timestamp 1569139307
transform 1 0 4360 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3288
timestamp 1569139307
transform 1 0 4360 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3289
timestamp 1569139307
transform 1 0 4360 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3290
timestamp 1569139307
transform 1 0 4360 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3291
timestamp 1569139307
transform 1 0 4360 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3292
timestamp 1569139307
transform 1 0 4360 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3293
timestamp 1569139307
transform 1 0 4360 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3294
timestamp 1569139307
transform 1 0 4360 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3295
timestamp 1569139307
transform 1 0 4360 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3296
timestamp 1569139307
transform 1 0 4360 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3297
timestamp 1569139307
transform 1 0 4360 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3298
timestamp 1569139307
transform 1 0 4360 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3299
timestamp 1569139307
transform 1 0 4360 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3300
timestamp 1569139307
transform 1 0 3464 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3301
timestamp 1569139307
transform 1 0 3720 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3302
timestamp 1569139307
transform 1 0 3592 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3303
timestamp 1569139307
transform 1 0 3720 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3304
timestamp 1569139307
transform 1 0 3464 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3305
timestamp 1569139307
transform 1 0 3592 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3306
timestamp 1569139307
transform 1 0 3464 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3307
timestamp 1569139307
transform 1 0 3656 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3308
timestamp 1569139307
transform 1 0 3528 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3309
timestamp 1569139307
transform 1 0 3656 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3310
timestamp 1569139307
transform 1 0 3720 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3311
timestamp 1569139307
transform 1 0 3528 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3312
timestamp 1569139307
transform 1 0 3592 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3313
timestamp 1569139307
transform 1 0 3528 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3314
timestamp 1569139307
transform 1 0 3528 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3315
timestamp 1569139307
transform 1 0 3656 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3316
timestamp 1569139307
transform 1 0 3656 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3317
timestamp 1569139307
transform 1 0 3592 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3318
timestamp 1569139307
transform 1 0 3464 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3319
timestamp 1569139307
transform 1 0 3720 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3320
timestamp 1569139307
transform 1 0 3336 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3321
timestamp 1569139307
transform 1 0 3336 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3322
timestamp 1569139307
transform 1 0 3208 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3323
timestamp 1569139307
transform 1 0 3336 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3324
timestamp 1569139307
transform 1 0 3400 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3325
timestamp 1569139307
transform 1 0 3144 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3326
timestamp 1569139307
transform 1 0 3400 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3327
timestamp 1569139307
transform 1 0 3208 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3328
timestamp 1569139307
transform 1 0 3272 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3329
timestamp 1569139307
transform 1 0 3400 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3330
timestamp 1569139307
transform 1 0 3144 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3331
timestamp 1569139307
transform 1 0 3144 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3332
timestamp 1569139307
transform 1 0 3208 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3333
timestamp 1569139307
transform 1 0 3144 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3334
timestamp 1569139307
transform 1 0 3400 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3335
timestamp 1569139307
transform 1 0 3272 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3336
timestamp 1569139307
transform 1 0 3208 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3337
timestamp 1569139307
transform 1 0 3272 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3338
timestamp 1569139307
transform 1 0 3336 0 1 2568
box -8 -8 8 8
use VIA1  VIA1_3339
timestamp 1569139307
transform 1 0 3272 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3340
timestamp 1569139307
transform 1 0 3336 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3341
timestamp 1569139307
transform 1 0 3208 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3342
timestamp 1569139307
transform 1 0 3272 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3343
timestamp 1569139307
transform 1 0 3208 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3344
timestamp 1569139307
transform 1 0 3144 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3345
timestamp 1569139307
transform 1 0 3400 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3346
timestamp 1569139307
transform 1 0 3400 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3347
timestamp 1569139307
transform 1 0 3272 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3348
timestamp 1569139307
transform 1 0 3336 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3349
timestamp 1569139307
transform 1 0 3272 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3350
timestamp 1569139307
transform 1 0 3208 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3351
timestamp 1569139307
transform 1 0 3336 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3352
timestamp 1569139307
transform 1 0 3272 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3353
timestamp 1569139307
transform 1 0 3336 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3354
timestamp 1569139307
transform 1 0 3208 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3355
timestamp 1569139307
transform 1 0 3400 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3356
timestamp 1569139307
transform 1 0 3400 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3357
timestamp 1569139307
transform 1 0 3144 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3358
timestamp 1569139307
transform 1 0 3144 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3359
timestamp 1569139307
transform 1 0 3400 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3360
timestamp 1569139307
transform 1 0 3144 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3361
timestamp 1569139307
transform 1 0 3336 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3362
timestamp 1569139307
transform 1 0 3144 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3363
timestamp 1569139307
transform 1 0 3272 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3364
timestamp 1569139307
transform 1 0 3208 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3365
timestamp 1569139307
transform 1 0 3592 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3366
timestamp 1569139307
transform 1 0 3720 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3367
timestamp 1569139307
transform 1 0 3464 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3368
timestamp 1569139307
transform 1 0 3720 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3369
timestamp 1569139307
transform 1 0 3464 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3370
timestamp 1569139307
transform 1 0 3656 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3371
timestamp 1569139307
transform 1 0 3528 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3372
timestamp 1569139307
transform 1 0 3528 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3373
timestamp 1569139307
transform 1 0 3592 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3374
timestamp 1569139307
transform 1 0 3592 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3375
timestamp 1569139307
transform 1 0 3528 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3376
timestamp 1569139307
transform 1 0 3656 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3377
timestamp 1569139307
transform 1 0 3656 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3378
timestamp 1569139307
transform 1 0 3656 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3379
timestamp 1569139307
transform 1 0 3528 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3380
timestamp 1569139307
transform 1 0 3528 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3381
timestamp 1569139307
transform 1 0 3464 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3382
timestamp 1569139307
transform 1 0 3720 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3383
timestamp 1569139307
transform 1 0 3592 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3384
timestamp 1569139307
transform 1 0 3464 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3385
timestamp 1569139307
transform 1 0 3720 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3386
timestamp 1569139307
transform 1 0 3464 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3387
timestamp 1569139307
transform 1 0 3720 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3388
timestamp 1569139307
transform 1 0 3656 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3389
timestamp 1569139307
transform 1 0 3592 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3390
timestamp 1569139307
transform 1 0 3080 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3391
timestamp 1569139307
transform 1 0 3080 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3392
timestamp 1569139307
transform 1 0 2952 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3393
timestamp 1569139307
transform 1 0 2696 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3394
timestamp 1569139307
transform 1 0 2952 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3395
timestamp 1569139307
transform 1 0 3016 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3396
timestamp 1569139307
transform 1 0 2888 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3397
timestamp 1569139307
transform 1 0 3016 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3398
timestamp 1569139307
transform 1 0 2760 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3399
timestamp 1569139307
transform 1 0 3016 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3400
timestamp 1569139307
transform 1 0 2952 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3401
timestamp 1569139307
transform 1 0 3080 0 1 2696
box -8 -8 8 8
use VIA1  VIA1_3402
timestamp 1569139307
transform 1 0 2824 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3403
timestamp 1569139307
transform 1 0 3080 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3404
timestamp 1569139307
transform 1 0 2824 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3405
timestamp 1569139307
transform 1 0 3080 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3406
timestamp 1569139307
transform 1 0 2952 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3407
timestamp 1569139307
transform 1 0 2952 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3408
timestamp 1569139307
transform 1 0 2888 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3409
timestamp 1569139307
transform 1 0 2888 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3410
timestamp 1569139307
transform 1 0 2632 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3411
timestamp 1569139307
transform 1 0 2952 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3412
timestamp 1569139307
transform 1 0 2696 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3413
timestamp 1569139307
transform 1 0 2888 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3414
timestamp 1569139307
transform 1 0 3016 0 1 2760
box -8 -8 8 8
use VIA1  VIA1_3415
timestamp 1569139307
transform 1 0 3016 0 1 2824
box -8 -8 8 8
use VIA1  VIA1_3416
timestamp 1569139307
transform 1 0 3016 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3417
timestamp 1569139307
transform 1 0 2760 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3418
timestamp 1569139307
transform 1 0 3016 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3419
timestamp 1569139307
transform 1 0 2760 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3420
timestamp 1569139307
transform 1 0 2888 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3421
timestamp 1569139307
transform 1 0 3080 0 1 2888
box -8 -8 8 8
use VIA1  VIA1_3422
timestamp 1569139307
transform 1 0 2824 0 1 2952
box -8 -8 8 8
use VIA1  VIA1_3423
timestamp 1569139307
transform 1 0 3080 0 1 3016
box -8 -8 8 8
use VIA1  VIA1_3424
timestamp 1569139307
transform 1 0 2824 0 1 3080
box -8 -8 8 8
use VIA1  VIA1_3425
timestamp 1569139307
transform 1 0 3080 0 1 2632
box -8 -8 8 8
use VIA1  VIA1_3426
timestamp 1569139307
transform 1 0 2888 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3427
timestamp 1569139307
transform 1 0 3016 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3428
timestamp 1569139307
transform 1 0 3080 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3429
timestamp 1569139307
transform 1 0 2888 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3430
timestamp 1569139307
transform 1 0 2824 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3431
timestamp 1569139307
transform 1 0 2888 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3432
timestamp 1569139307
transform 1 0 2888 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3433
timestamp 1569139307
transform 1 0 2888 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3434
timestamp 1569139307
transform 1 0 3016 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3435
timestamp 1569139307
transform 1 0 3080 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3436
timestamp 1569139307
transform 1 0 3080 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3437
timestamp 1569139307
transform 1 0 2952 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3438
timestamp 1569139307
transform 1 0 2952 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3439
timestamp 1569139307
transform 1 0 2952 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3440
timestamp 1569139307
transform 1 0 2952 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3441
timestamp 1569139307
transform 1 0 3016 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3442
timestamp 1569139307
transform 1 0 3016 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3443
timestamp 1569139307
transform 1 0 3080 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3444
timestamp 1569139307
transform 1 0 2824 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3445
timestamp 1569139307
transform 1 0 2824 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3446
timestamp 1569139307
transform 1 0 3016 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3447
timestamp 1569139307
transform 1 0 2824 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3448
timestamp 1569139307
transform 1 0 2824 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3449
timestamp 1569139307
transform 1 0 2952 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3450
timestamp 1569139307
transform 1 0 3080 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3451
timestamp 1569139307
transform 1 0 2696 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3452
timestamp 1569139307
transform 1 0 2568 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3453
timestamp 1569139307
transform 1 0 2760 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3454
timestamp 1569139307
transform 1 0 2632 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3455
timestamp 1569139307
transform 1 0 2696 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3456
timestamp 1569139307
transform 1 0 2696 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3457
timestamp 1569139307
transform 1 0 2696 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3458
timestamp 1569139307
transform 1 0 2696 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3459
timestamp 1569139307
transform 1 0 2632 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3460
timestamp 1569139307
transform 1 0 2632 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3461
timestamp 1569139307
transform 1 0 2568 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3462
timestamp 1569139307
transform 1 0 2760 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3463
timestamp 1569139307
transform 1 0 2760 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3464
timestamp 1569139307
transform 1 0 2760 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3465
timestamp 1569139307
transform 1 0 2632 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3466
timestamp 1569139307
transform 1 0 2760 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3467
timestamp 1569139307
transform 1 0 2568 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3468
timestamp 1569139307
transform 1 0 2568 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3469
timestamp 1569139307
transform 1 0 2568 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3470
timestamp 1569139307
transform 1 0 2632 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3471
timestamp 1569139307
transform 1 0 2568 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3472
timestamp 1569139307
transform 1 0 2632 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3473
timestamp 1569139307
transform 1 0 2632 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3474
timestamp 1569139307
transform 1 0 2632 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3475
timestamp 1569139307
transform 1 0 2760 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3476
timestamp 1569139307
transform 1 0 2760 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3477
timestamp 1569139307
transform 1 0 2696 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3478
timestamp 1569139307
transform 1 0 2696 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3479
timestamp 1569139307
transform 1 0 2760 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3480
timestamp 1569139307
transform 1 0 2760 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3481
timestamp 1569139307
transform 1 0 2760 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3482
timestamp 1569139307
transform 1 0 2632 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3483
timestamp 1569139307
transform 1 0 2568 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3484
timestamp 1569139307
transform 1 0 2632 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3485
timestamp 1569139307
transform 1 0 2568 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3486
timestamp 1569139307
transform 1 0 2568 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3487
timestamp 1569139307
transform 1 0 2568 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3488
timestamp 1569139307
transform 1 0 2696 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3489
timestamp 1569139307
transform 1 0 2696 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3490
timestamp 1569139307
transform 1 0 2696 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3491
timestamp 1569139307
transform 1 0 3080 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3492
timestamp 1569139307
transform 1 0 3016 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3493
timestamp 1569139307
transform 1 0 3080 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3494
timestamp 1569139307
transform 1 0 3016 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3495
timestamp 1569139307
transform 1 0 2824 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3496
timestamp 1569139307
transform 1 0 2824 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3497
timestamp 1569139307
transform 1 0 2888 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3498
timestamp 1569139307
transform 1 0 2888 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3499
timestamp 1569139307
transform 1 0 3080 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3500
timestamp 1569139307
transform 1 0 2952 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3501
timestamp 1569139307
transform 1 0 2952 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3502
timestamp 1569139307
transform 1 0 3080 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3503
timestamp 1569139307
transform 1 0 3016 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3504
timestamp 1569139307
transform 1 0 3080 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3505
timestamp 1569139307
transform 1 0 2824 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3506
timestamp 1569139307
transform 1 0 2824 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3507
timestamp 1569139307
transform 1 0 2824 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3508
timestamp 1569139307
transform 1 0 2888 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3509
timestamp 1569139307
transform 1 0 2888 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3510
timestamp 1569139307
transform 1 0 2888 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3511
timestamp 1569139307
transform 1 0 3016 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3512
timestamp 1569139307
transform 1 0 2952 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3513
timestamp 1569139307
transform 1 0 2952 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3514
timestamp 1569139307
transform 1 0 2952 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3515
timestamp 1569139307
transform 1 0 3016 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3516
timestamp 1569139307
transform 1 0 3656 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3517
timestamp 1569139307
transform 1 0 3720 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3518
timestamp 1569139307
transform 1 0 3720 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3519
timestamp 1569139307
transform 1 0 3720 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3520
timestamp 1569139307
transform 1 0 3720 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3521
timestamp 1569139307
transform 1 0 3720 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3522
timestamp 1569139307
transform 1 0 3464 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3523
timestamp 1569139307
transform 1 0 3464 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3524
timestamp 1569139307
transform 1 0 3464 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3525
timestamp 1569139307
transform 1 0 3464 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3526
timestamp 1569139307
transform 1 0 3464 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3527
timestamp 1569139307
transform 1 0 3528 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3528
timestamp 1569139307
transform 1 0 3528 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3529
timestamp 1569139307
transform 1 0 3528 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3530
timestamp 1569139307
transform 1 0 3528 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3531
timestamp 1569139307
transform 1 0 3528 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3532
timestamp 1569139307
transform 1 0 3592 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3533
timestamp 1569139307
transform 1 0 3592 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3534
timestamp 1569139307
transform 1 0 3592 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3535
timestamp 1569139307
transform 1 0 3592 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3536
timestamp 1569139307
transform 1 0 3592 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3537
timestamp 1569139307
transform 1 0 3656 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3538
timestamp 1569139307
transform 1 0 3656 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3539
timestamp 1569139307
transform 1 0 3656 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3540
timestamp 1569139307
transform 1 0 3656 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3541
timestamp 1569139307
transform 1 0 3208 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3542
timestamp 1569139307
transform 1 0 3272 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3543
timestamp 1569139307
transform 1 0 3336 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3544
timestamp 1569139307
transform 1 0 3400 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3545
timestamp 1569139307
transform 1 0 3336 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3546
timestamp 1569139307
transform 1 0 3336 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3547
timestamp 1569139307
transform 1 0 3336 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3548
timestamp 1569139307
transform 1 0 3336 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3549
timestamp 1569139307
transform 1 0 3144 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3550
timestamp 1569139307
transform 1 0 3400 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3551
timestamp 1569139307
transform 1 0 3400 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3552
timestamp 1569139307
transform 1 0 3400 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3553
timestamp 1569139307
transform 1 0 3400 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3554
timestamp 1569139307
transform 1 0 3208 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3555
timestamp 1569139307
transform 1 0 3208 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3556
timestamp 1569139307
transform 1 0 3208 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3557
timestamp 1569139307
transform 1 0 3208 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3558
timestamp 1569139307
transform 1 0 3144 0 1 3144
box -8 -8 8 8
use VIA1  VIA1_3559
timestamp 1569139307
transform 1 0 3272 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3560
timestamp 1569139307
transform 1 0 3272 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3561
timestamp 1569139307
transform 1 0 3272 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3562
timestamp 1569139307
transform 1 0 3272 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_3563
timestamp 1569139307
transform 1 0 3144 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_3564
timestamp 1569139307
transform 1 0 3144 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_3565
timestamp 1569139307
transform 1 0 3144 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_3566
timestamp 1569139307
transform 1 0 3336 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3567
timestamp 1569139307
transform 1 0 3336 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3568
timestamp 1569139307
transform 1 0 3400 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3569
timestamp 1569139307
transform 1 0 3400 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3570
timestamp 1569139307
transform 1 0 3272 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3571
timestamp 1569139307
transform 1 0 3272 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3572
timestamp 1569139307
transform 1 0 3336 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3573
timestamp 1569139307
transform 1 0 3336 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3574
timestamp 1569139307
transform 1 0 3336 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3575
timestamp 1569139307
transform 1 0 3272 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3576
timestamp 1569139307
transform 1 0 3272 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3577
timestamp 1569139307
transform 1 0 3400 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3578
timestamp 1569139307
transform 1 0 3400 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3579
timestamp 1569139307
transform 1 0 3400 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3580
timestamp 1569139307
transform 1 0 3272 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3581
timestamp 1569139307
transform 1 0 3144 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3582
timestamp 1569139307
transform 1 0 3144 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3583
timestamp 1569139307
transform 1 0 3144 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3584
timestamp 1569139307
transform 1 0 3208 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3585
timestamp 1569139307
transform 1 0 3208 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3586
timestamp 1569139307
transform 1 0 3208 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3587
timestamp 1569139307
transform 1 0 3144 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3588
timestamp 1569139307
transform 1 0 3144 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3589
timestamp 1569139307
transform 1 0 3208 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3590
timestamp 1569139307
transform 1 0 3208 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3591
timestamp 1569139307
transform 1 0 3464 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3592
timestamp 1569139307
transform 1 0 3464 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3593
timestamp 1569139307
transform 1 0 3528 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3594
timestamp 1569139307
transform 1 0 3528 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3595
timestamp 1569139307
transform 1 0 3592 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3596
timestamp 1569139307
transform 1 0 3592 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3597
timestamp 1569139307
transform 1 0 3720 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3598
timestamp 1569139307
transform 1 0 3464 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3599
timestamp 1569139307
transform 1 0 3464 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3600
timestamp 1569139307
transform 1 0 3464 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3601
timestamp 1569139307
transform 1 0 3528 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3602
timestamp 1569139307
transform 1 0 3528 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3603
timestamp 1569139307
transform 1 0 3528 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3604
timestamp 1569139307
transform 1 0 3592 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3605
timestamp 1569139307
transform 1 0 3592 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3606
timestamp 1569139307
transform 1 0 3592 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3607
timestamp 1569139307
transform 1 0 3720 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3608
timestamp 1569139307
transform 1 0 3720 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3609
timestamp 1569139307
transform 1 0 3656 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3610
timestamp 1569139307
transform 1 0 3656 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3611
timestamp 1569139307
transform 1 0 3720 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_3612
timestamp 1569139307
transform 1 0 3720 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_3613
timestamp 1569139307
transform 1 0 3656 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_3614
timestamp 1569139307
transform 1 0 3656 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_3615
timestamp 1569139307
transform 1 0 3656 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_3616
timestamp 1569139307
transform 1 0 3592 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3617
timestamp 1569139307
transform 1 0 3720 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3618
timestamp 1569139307
transform 1 0 3720 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3619
timestamp 1569139307
transform 1 0 3720 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3620
timestamp 1569139307
transform 1 0 3592 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3621
timestamp 1569139307
transform 1 0 3592 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3622
timestamp 1569139307
transform 1 0 3656 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3623
timestamp 1569139307
transform 1 0 3720 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3624
timestamp 1569139307
transform 1 0 3656 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3625
timestamp 1569139307
transform 1 0 3592 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3626
timestamp 1569139307
transform 1 0 3528 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3627
timestamp 1569139307
transform 1 0 3464 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3628
timestamp 1569139307
transform 1 0 3464 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3629
timestamp 1569139307
transform 1 0 3464 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3630
timestamp 1569139307
transform 1 0 3656 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3631
timestamp 1569139307
transform 1 0 3464 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3632
timestamp 1569139307
transform 1 0 3656 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3633
timestamp 1569139307
transform 1 0 3464 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3634
timestamp 1569139307
transform 1 0 3528 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3635
timestamp 1569139307
transform 1 0 3720 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3636
timestamp 1569139307
transform 1 0 3528 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3637
timestamp 1569139307
transform 1 0 3528 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3638
timestamp 1569139307
transform 1 0 3528 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3639
timestamp 1569139307
transform 1 0 3656 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3640
timestamp 1569139307
transform 1 0 3592 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3641
timestamp 1569139307
transform 1 0 3336 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3642
timestamp 1569139307
transform 1 0 3336 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3643
timestamp 1569139307
transform 1 0 3336 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3644
timestamp 1569139307
transform 1 0 3272 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3645
timestamp 1569139307
transform 1 0 3336 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3646
timestamp 1569139307
transform 1 0 3272 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3647
timestamp 1569139307
transform 1 0 3400 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3648
timestamp 1569139307
transform 1 0 3144 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3649
timestamp 1569139307
transform 1 0 3400 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3650
timestamp 1569139307
transform 1 0 3400 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3651
timestamp 1569139307
transform 1 0 3272 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3652
timestamp 1569139307
transform 1 0 3144 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3653
timestamp 1569139307
transform 1 0 3400 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3654
timestamp 1569139307
transform 1 0 3400 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3655
timestamp 1569139307
transform 1 0 3144 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3656
timestamp 1569139307
transform 1 0 3144 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3657
timestamp 1569139307
transform 1 0 3272 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3658
timestamp 1569139307
transform 1 0 3208 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3659
timestamp 1569139307
transform 1 0 3208 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3660
timestamp 1569139307
transform 1 0 3336 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3661
timestamp 1569139307
transform 1 0 3208 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3662
timestamp 1569139307
transform 1 0 3208 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3663
timestamp 1569139307
transform 1 0 3208 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3664
timestamp 1569139307
transform 1 0 3272 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3665
timestamp 1569139307
transform 1 0 3144 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3666
timestamp 1569139307
transform 1 0 3272 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3667
timestamp 1569139307
transform 1 0 3272 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3668
timestamp 1569139307
transform 1 0 3272 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3669
timestamp 1569139307
transform 1 0 3272 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3670
timestamp 1569139307
transform 1 0 3144 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3671
timestamp 1569139307
transform 1 0 3336 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3672
timestamp 1569139307
transform 1 0 3336 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3673
timestamp 1569139307
transform 1 0 3336 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3674
timestamp 1569139307
transform 1 0 3336 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3675
timestamp 1569139307
transform 1 0 3208 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3676
timestamp 1569139307
transform 1 0 3144 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3677
timestamp 1569139307
transform 1 0 3400 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3678
timestamp 1569139307
transform 1 0 3400 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3679
timestamp 1569139307
transform 1 0 3400 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3680
timestamp 1569139307
transform 1 0 3400 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3681
timestamp 1569139307
transform 1 0 3208 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3682
timestamp 1569139307
transform 1 0 3208 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3683
timestamp 1569139307
transform 1 0 3144 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3684
timestamp 1569139307
transform 1 0 3144 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3685
timestamp 1569139307
transform 1 0 3208 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3686
timestamp 1569139307
transform 1 0 3592 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3687
timestamp 1569139307
transform 1 0 3656 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3688
timestamp 1569139307
transform 1 0 3656 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3689
timestamp 1569139307
transform 1 0 3656 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3690
timestamp 1569139307
transform 1 0 3464 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3691
timestamp 1569139307
transform 1 0 3656 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3692
timestamp 1569139307
transform 1 0 3464 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3693
timestamp 1569139307
transform 1 0 3464 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3694
timestamp 1569139307
transform 1 0 3464 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3695
timestamp 1569139307
transform 1 0 3720 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3696
timestamp 1569139307
transform 1 0 3528 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3697
timestamp 1569139307
transform 1 0 3720 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3698
timestamp 1569139307
transform 1 0 3528 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3699
timestamp 1569139307
transform 1 0 3528 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3700
timestamp 1569139307
transform 1 0 3720 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3701
timestamp 1569139307
transform 1 0 3528 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3702
timestamp 1569139307
transform 1 0 3720 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3703
timestamp 1569139307
transform 1 0 3592 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3704
timestamp 1569139307
transform 1 0 3592 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3705
timestamp 1569139307
transform 1 0 3592 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3706
timestamp 1569139307
transform 1 0 2824 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3707
timestamp 1569139307
transform 1 0 3080 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3708
timestamp 1569139307
transform 1 0 2824 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3709
timestamp 1569139307
transform 1 0 2824 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3710
timestamp 1569139307
transform 1 0 2824 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3711
timestamp 1569139307
transform 1 0 2824 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3712
timestamp 1569139307
transform 1 0 2888 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3713
timestamp 1569139307
transform 1 0 2888 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3714
timestamp 1569139307
transform 1 0 2888 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3715
timestamp 1569139307
transform 1 0 2888 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3716
timestamp 1569139307
transform 1 0 2952 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3717
timestamp 1569139307
transform 1 0 2952 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3718
timestamp 1569139307
transform 1 0 2952 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3719
timestamp 1569139307
transform 1 0 2952 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3720
timestamp 1569139307
transform 1 0 2888 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3721
timestamp 1569139307
transform 1 0 3016 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3722
timestamp 1569139307
transform 1 0 3016 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3723
timestamp 1569139307
transform 1 0 3016 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3724
timestamp 1569139307
transform 1 0 3016 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3725
timestamp 1569139307
transform 1 0 3016 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3726
timestamp 1569139307
transform 1 0 3080 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3727
timestamp 1569139307
transform 1 0 3080 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3728
timestamp 1569139307
transform 1 0 2952 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3729
timestamp 1569139307
transform 1 0 3080 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3730
timestamp 1569139307
transform 1 0 3080 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3731
timestamp 1569139307
transform 1 0 2696 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3732
timestamp 1569139307
transform 1 0 2696 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3733
timestamp 1569139307
transform 1 0 2696 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3734
timestamp 1569139307
transform 1 0 2696 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3735
timestamp 1569139307
transform 1 0 2760 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3736
timestamp 1569139307
transform 1 0 2760 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3737
timestamp 1569139307
transform 1 0 2760 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3738
timestamp 1569139307
transform 1 0 2760 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3739
timestamp 1569139307
transform 1 0 2696 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3740
timestamp 1569139307
transform 1 0 2568 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3741
timestamp 1569139307
transform 1 0 2568 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3742
timestamp 1569139307
transform 1 0 2760 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3743
timestamp 1569139307
transform 1 0 2568 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3744
timestamp 1569139307
transform 1 0 2568 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3745
timestamp 1569139307
transform 1 0 2632 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3746
timestamp 1569139307
transform 1 0 2568 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3747
timestamp 1569139307
transform 1 0 2632 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3748
timestamp 1569139307
transform 1 0 2632 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3749
timestamp 1569139307
transform 1 0 2632 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3750
timestamp 1569139307
transform 1 0 2632 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3751
timestamp 1569139307
transform 1 0 2696 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3752
timestamp 1569139307
transform 1 0 2696 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3753
timestamp 1569139307
transform 1 0 2696 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3754
timestamp 1569139307
transform 1 0 2696 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3755
timestamp 1569139307
transform 1 0 2760 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3756
timestamp 1569139307
transform 1 0 2760 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3757
timestamp 1569139307
transform 1 0 2760 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3758
timestamp 1569139307
transform 1 0 2760 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3759
timestamp 1569139307
transform 1 0 2632 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3760
timestamp 1569139307
transform 1 0 2632 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3761
timestamp 1569139307
transform 1 0 2632 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3762
timestamp 1569139307
transform 1 0 2632 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3763
timestamp 1569139307
transform 1 0 2568 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3764
timestamp 1569139307
transform 1 0 2568 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3765
timestamp 1569139307
transform 1 0 2568 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3766
timestamp 1569139307
transform 1 0 2568 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3767
timestamp 1569139307
transform 1 0 2824 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3768
timestamp 1569139307
transform 1 0 2824 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3769
timestamp 1569139307
transform 1 0 2824 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3770
timestamp 1569139307
transform 1 0 2824 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3771
timestamp 1569139307
transform 1 0 2888 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3772
timestamp 1569139307
transform 1 0 2888 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3773
timestamp 1569139307
transform 1 0 2888 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3774
timestamp 1569139307
transform 1 0 2888 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3775
timestamp 1569139307
transform 1 0 2952 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3776
timestamp 1569139307
transform 1 0 2952 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3777
timestamp 1569139307
transform 1 0 2952 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3778
timestamp 1569139307
transform 1 0 2952 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3779
timestamp 1569139307
transform 1 0 3016 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3780
timestamp 1569139307
transform 1 0 3016 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3781
timestamp 1569139307
transform 1 0 3016 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3782
timestamp 1569139307
transform 1 0 3016 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3783
timestamp 1569139307
transform 1 0 3080 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3784
timestamp 1569139307
transform 1 0 3080 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3785
timestamp 1569139307
transform 1 0 3080 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_3786
timestamp 1569139307
transform 1 0 3080 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3787
timestamp 1569139307
transform 1 0 3016 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3788
timestamp 1569139307
transform 1 0 2888 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3789
timestamp 1569139307
transform 1 0 3080 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3790
timestamp 1569139307
transform 1 0 2952 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3791
timestamp 1569139307
transform 1 0 2824 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3792
timestamp 1569139307
transform 1 0 2824 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3793
timestamp 1569139307
transform 1 0 3080 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3794
timestamp 1569139307
transform 1 0 3080 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3795
timestamp 1569139307
transform 1 0 3016 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3796
timestamp 1569139307
transform 1 0 2888 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3797
timestamp 1569139307
transform 1 0 2824 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3798
timestamp 1569139307
transform 1 0 2888 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3799
timestamp 1569139307
transform 1 0 3016 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3800
timestamp 1569139307
transform 1 0 2952 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3801
timestamp 1569139307
transform 1 0 2952 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3802
timestamp 1569139307
transform 1 0 2888 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3803
timestamp 1569139307
transform 1 0 2824 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3804
timestamp 1569139307
transform 1 0 2952 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3805
timestamp 1569139307
transform 1 0 3016 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3806
timestamp 1569139307
transform 1 0 3080 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3807
timestamp 1569139307
transform 1 0 2760 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3808
timestamp 1569139307
transform 1 0 2696 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3809
timestamp 1569139307
transform 1 0 2632 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3810
timestamp 1569139307
transform 1 0 2568 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3811
timestamp 1569139307
transform 1 0 2632 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3812
timestamp 1569139307
transform 1 0 2760 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3813
timestamp 1569139307
transform 1 0 2632 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3814
timestamp 1569139307
transform 1 0 2696 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3815
timestamp 1569139307
transform 1 0 2760 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3816
timestamp 1569139307
transform 1 0 2568 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3817
timestamp 1569139307
transform 1 0 2568 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3818
timestamp 1569139307
transform 1 0 2696 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3819
timestamp 1569139307
transform 1 0 2696 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3820
timestamp 1569139307
transform 1 0 2760 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3821
timestamp 1569139307
transform 1 0 2568 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3822
timestamp 1569139307
transform 1 0 2632 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3823
timestamp 1569139307
transform 1 0 2696 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3824
timestamp 1569139307
transform 1 0 2632 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3825
timestamp 1569139307
transform 1 0 2760 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3826
timestamp 1569139307
transform 1 0 2760 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3827
timestamp 1569139307
transform 1 0 2760 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3828
timestamp 1569139307
transform 1 0 2696 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3829
timestamp 1569139307
transform 1 0 2696 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3830
timestamp 1569139307
transform 1 0 2760 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3831
timestamp 1569139307
transform 1 0 2696 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3832
timestamp 1569139307
transform 1 0 2568 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3833
timestamp 1569139307
transform 1 0 2568 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3834
timestamp 1569139307
transform 1 0 2568 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3835
timestamp 1569139307
transform 1 0 2632 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3836
timestamp 1569139307
transform 1 0 2568 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3837
timestamp 1569139307
transform 1 0 2632 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3838
timestamp 1569139307
transform 1 0 2632 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3839
timestamp 1569139307
transform 1 0 2824 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3840
timestamp 1569139307
transform 1 0 2952 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3841
timestamp 1569139307
transform 1 0 2952 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3842
timestamp 1569139307
transform 1 0 2824 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3843
timestamp 1569139307
transform 1 0 2952 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3844
timestamp 1569139307
transform 1 0 2952 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3845
timestamp 1569139307
transform 1 0 2824 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3846
timestamp 1569139307
transform 1 0 3016 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3847
timestamp 1569139307
transform 1 0 3016 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3848
timestamp 1569139307
transform 1 0 2824 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3849
timestamp 1569139307
transform 1 0 3016 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3850
timestamp 1569139307
transform 1 0 3016 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3851
timestamp 1569139307
transform 1 0 3080 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3852
timestamp 1569139307
transform 1 0 3080 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3853
timestamp 1569139307
transform 1 0 3080 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3854
timestamp 1569139307
transform 1 0 3080 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3855
timestamp 1569139307
transform 1 0 2888 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3856
timestamp 1569139307
transform 1 0 2888 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3857
timestamp 1569139307
transform 1 0 2888 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3858
timestamp 1569139307
transform 1 0 2888 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3859
timestamp 1569139307
transform 1 0 3464 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3860
timestamp 1569139307
transform 1 0 3656 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3861
timestamp 1569139307
transform 1 0 3464 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3862
timestamp 1569139307
transform 1 0 3464 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3863
timestamp 1569139307
transform 1 0 3528 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3864
timestamp 1569139307
transform 1 0 3592 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3865
timestamp 1569139307
transform 1 0 3720 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3866
timestamp 1569139307
transform 1 0 3592 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3867
timestamp 1569139307
transform 1 0 3592 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3868
timestamp 1569139307
transform 1 0 3720 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3869
timestamp 1569139307
transform 1 0 3528 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3870
timestamp 1569139307
transform 1 0 3464 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3871
timestamp 1569139307
transform 1 0 3592 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3872
timestamp 1569139307
transform 1 0 3528 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3873
timestamp 1569139307
transform 1 0 3656 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3874
timestamp 1569139307
transform 1 0 3656 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3875
timestamp 1569139307
transform 1 0 3720 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3876
timestamp 1569139307
transform 1 0 3656 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3877
timestamp 1569139307
transform 1 0 3528 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3878
timestamp 1569139307
transform 1 0 3720 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3879
timestamp 1569139307
transform 1 0 3336 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3880
timestamp 1569139307
transform 1 0 3208 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3881
timestamp 1569139307
transform 1 0 3400 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3882
timestamp 1569139307
transform 1 0 3336 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3883
timestamp 1569139307
transform 1 0 3208 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3884
timestamp 1569139307
transform 1 0 3336 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3885
timestamp 1569139307
transform 1 0 3208 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3886
timestamp 1569139307
transform 1 0 3272 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3887
timestamp 1569139307
transform 1 0 3400 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3888
timestamp 1569139307
transform 1 0 3144 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3889
timestamp 1569139307
transform 1 0 3272 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3890
timestamp 1569139307
transform 1 0 3272 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3891
timestamp 1569139307
transform 1 0 3272 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3892
timestamp 1569139307
transform 1 0 3144 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3893
timestamp 1569139307
transform 1 0 3400 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3894
timestamp 1569139307
transform 1 0 3400 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3895
timestamp 1569139307
transform 1 0 3144 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_3896
timestamp 1569139307
transform 1 0 3336 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3897
timestamp 1569139307
transform 1 0 3208 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_3898
timestamp 1569139307
transform 1 0 3144 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3899
timestamp 1569139307
transform 1 0 3272 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3900
timestamp 1569139307
transform 1 0 3272 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3901
timestamp 1569139307
transform 1 0 3272 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3902
timestamp 1569139307
transform 1 0 3336 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3903
timestamp 1569139307
transform 1 0 3336 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3904
timestamp 1569139307
transform 1 0 3336 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3905
timestamp 1569139307
transform 1 0 3336 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3906
timestamp 1569139307
transform 1 0 3400 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3907
timestamp 1569139307
transform 1 0 3400 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3908
timestamp 1569139307
transform 1 0 3400 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3909
timestamp 1569139307
transform 1 0 3144 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3910
timestamp 1569139307
transform 1 0 3144 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3911
timestamp 1569139307
transform 1 0 3400 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3912
timestamp 1569139307
transform 1 0 3144 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3913
timestamp 1569139307
transform 1 0 3144 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3914
timestamp 1569139307
transform 1 0 3208 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3915
timestamp 1569139307
transform 1 0 3208 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3916
timestamp 1569139307
transform 1 0 3208 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3917
timestamp 1569139307
transform 1 0 3208 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3918
timestamp 1569139307
transform 1 0 3272 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3919
timestamp 1569139307
transform 1 0 3464 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3920
timestamp 1569139307
transform 1 0 3592 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3921
timestamp 1569139307
transform 1 0 3592 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3922
timestamp 1569139307
transform 1 0 3592 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3923
timestamp 1569139307
transform 1 0 3592 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3924
timestamp 1569139307
transform 1 0 3656 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3925
timestamp 1569139307
transform 1 0 3656 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3926
timestamp 1569139307
transform 1 0 3656 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3927
timestamp 1569139307
transform 1 0 3656 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3928
timestamp 1569139307
transform 1 0 3720 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3929
timestamp 1569139307
transform 1 0 3720 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3930
timestamp 1569139307
transform 1 0 3720 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3931
timestamp 1569139307
transform 1 0 3464 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3932
timestamp 1569139307
transform 1 0 3720 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3933
timestamp 1569139307
transform 1 0 3464 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3934
timestamp 1569139307
transform 1 0 3528 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3935
timestamp 1569139307
transform 1 0 3528 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3936
timestamp 1569139307
transform 1 0 3528 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3937
timestamp 1569139307
transform 1 0 3528 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3938
timestamp 1569139307
transform 1 0 3464 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3939
timestamp 1569139307
transform 1 0 2696 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3940
timestamp 1569139307
transform 1 0 3336 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3941
timestamp 1569139307
transform 1 0 2760 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3942
timestamp 1569139307
transform 1 0 3400 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3943
timestamp 1569139307
transform 1 0 2824 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3944
timestamp 1569139307
transform 1 0 3464 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3945
timestamp 1569139307
transform 1 0 2888 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3946
timestamp 1569139307
transform 1 0 3528 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3947
timestamp 1569139307
transform 1 0 2952 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3948
timestamp 1569139307
transform 1 0 3592 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3949
timestamp 1569139307
transform 1 0 3016 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3950
timestamp 1569139307
transform 1 0 3656 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3951
timestamp 1569139307
transform 1 0 3080 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3952
timestamp 1569139307
transform 1 0 3720 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3953
timestamp 1569139307
transform 1 0 3144 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3954
timestamp 1569139307
transform 1 0 2568 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3955
timestamp 1569139307
transform 1 0 3208 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3956
timestamp 1569139307
transform 1 0 2632 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3957
timestamp 1569139307
transform 1 0 3272 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_3958
timestamp 1569139307
transform 1 0 4616 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3959
timestamp 1569139307
transform 1 0 4680 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3960
timestamp 1569139307
transform 1 0 4744 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3961
timestamp 1569139307
transform 1 0 4808 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3962
timestamp 1569139307
transform 1 0 4872 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3963
timestamp 1569139307
transform 1 0 4488 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3964
timestamp 1569139307
transform 1 0 4552 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_3965
timestamp 1569139307
transform 1 0 3976 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3966
timestamp 1569139307
transform 1 0 3976 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3967
timestamp 1569139307
transform 1 0 3976 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3968
timestamp 1569139307
transform 1 0 3976 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3969
timestamp 1569139307
transform 1 0 4040 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3970
timestamp 1569139307
transform 1 0 4040 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3971
timestamp 1569139307
transform 1 0 4040 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3972
timestamp 1569139307
transform 1 0 4104 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3973
timestamp 1569139307
transform 1 0 4104 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3974
timestamp 1569139307
transform 1 0 4168 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3975
timestamp 1569139307
transform 1 0 3848 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3976
timestamp 1569139307
transform 1 0 3848 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3977
timestamp 1569139307
transform 1 0 3912 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3978
timestamp 1569139307
transform 1 0 3912 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3979
timestamp 1569139307
transform 1 0 3912 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3980
timestamp 1569139307
transform 1 0 3912 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3981
timestamp 1569139307
transform 1 0 3784 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3982
timestamp 1569139307
transform 1 0 3784 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3983
timestamp 1569139307
transform 1 0 3784 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_3984
timestamp 1569139307
transform 1 0 3848 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3985
timestamp 1569139307
transform 1 0 3848 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_3986
timestamp 1569139307
transform 1 0 3912 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_3987
timestamp 1569139307
transform 1 0 3784 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3988
timestamp 1569139307
transform 1 0 3784 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3989
timestamp 1569139307
transform 1 0 3784 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_3990
timestamp 1569139307
transform 1 0 3784 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_3991
timestamp 1569139307
transform 1 0 3848 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_3992
timestamp 1569139307
transform 1 0 3848 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_3993
timestamp 1569139307
transform 1 0 4296 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_3994
timestamp 1569139307
transform 1 0 4296 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_3995
timestamp 1569139307
transform 1 0 4296 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_3996
timestamp 1569139307
transform 1 0 4296 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_3997
timestamp 1569139307
transform 1 0 4296 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_3998
timestamp 1569139307
transform 1 0 4296 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_3999
timestamp 1569139307
transform 1 0 4296 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_4000
timestamp 1569139307
transform 1 0 4616 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4001
timestamp 1569139307
transform 1 0 4680 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4002
timestamp 1569139307
transform 1 0 4744 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4003
timestamp 1569139307
transform 1 0 4808 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4004
timestamp 1569139307
transform 1 0 4872 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4005
timestamp 1569139307
transform 1 0 4936 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_4006
timestamp 1569139307
transform 1 0 4936 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_4007
timestamp 1569139307
transform 1 0 4936 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_4008
timestamp 1569139307
transform 1 0 4936 0 1 4936
box -8 -8 8 8
use VIA1  VIA1_4009
timestamp 1569139307
transform 1 0 4424 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_4010
timestamp 1569139307
transform 1 0 4488 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_4011
timestamp 1569139307
transform 1 0 4424 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_4012
timestamp 1569139307
transform 1 0 4424 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_4013
timestamp 1569139307
transform 1 0 4424 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_4014
timestamp 1569139307
transform 1 0 4424 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_4015
timestamp 1569139307
transform 1 0 4424 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_4016
timestamp 1569139307
transform 1 0 4488 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_4017
timestamp 1569139307
transform 1 0 4616 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_4018
timestamp 1569139307
transform 1 0 4552 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_4019
timestamp 1569139307
transform 1 0 4488 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_4020
timestamp 1569139307
transform 1 0 4424 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4021
timestamp 1569139307
transform 1 0 4488 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4022
timestamp 1569139307
transform 1 0 4552 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4023
timestamp 1569139307
transform 1 0 4744 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_4024
timestamp 1569139307
transform 1 0 4744 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_4025
timestamp 1569139307
transform 1 0 4744 0 1 4936
box -8 -8 8 8
use VIA1  VIA1_4026
timestamp 1569139307
transform 1 0 4808 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_4027
timestamp 1569139307
transform 1 0 4808 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_4028
timestamp 1569139307
transform 1 0 4808 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_4029
timestamp 1569139307
transform 1 0 4808 0 1 4936
box -8 -8 8 8
use VIA1  VIA1_4030
timestamp 1569139307
transform 1 0 4424 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_4031
timestamp 1569139307
transform 1 0 4552 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_4032
timestamp 1569139307
transform 1 0 4872 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_4033
timestamp 1569139307
transform 1 0 4872 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_4034
timestamp 1569139307
transform 1 0 4872 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_4035
timestamp 1569139307
transform 1 0 4872 0 1 4936
box -8 -8 8 8
use VIA1  VIA1_4036
timestamp 1569139307
transform 1 0 4616 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4037
timestamp 1569139307
transform 1 0 4680 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4038
timestamp 1569139307
transform 1 0 4744 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4039
timestamp 1569139307
transform 1 0 4808 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4040
timestamp 1569139307
transform 1 0 4872 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4041
timestamp 1569139307
transform 1 0 4360 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_4042
timestamp 1569139307
transform 1 0 4360 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_4043
timestamp 1569139307
transform 1 0 4360 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_4044
timestamp 1569139307
transform 1 0 4360 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_4045
timestamp 1569139307
transform 1 0 4360 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_4046
timestamp 1569139307
transform 1 0 4360 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_4047
timestamp 1569139307
transform 1 0 4360 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_4048
timestamp 1569139307
transform 1 0 4360 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4049
timestamp 1569139307
transform 1 0 4424 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4050
timestamp 1569139307
transform 1 0 4488 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4051
timestamp 1569139307
transform 1 0 4552 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4052
timestamp 1569139307
transform 1 0 2504 0 1 4616
box -8 -8 8 8
use VIA1  VIA1_4053
timestamp 1569139307
transform 1 0 2504 0 1 4680
box -8 -8 8 8
use VIA1  VIA1_4054
timestamp 1569139307
transform 1 0 2504 0 1 4744
box -8 -8 8 8
use VIA1  VIA1_4055
timestamp 1569139307
transform 1 0 2504 0 1 4808
box -8 -8 8 8
use VIA1  VIA1_4056
timestamp 1569139307
transform 1 0 2504 0 1 4872
box -8 -8 8 8
use VIA1  VIA1_4057
timestamp 1569139307
transform 1 0 2504 0 1 136
box -8 -8 8 8
use VIA1  VIA1_4058
timestamp 1569139307
transform 1 0 2504 0 1 200
box -8 -8 8 8
use VIA1  VIA1_4059
timestamp 1569139307
transform 1 0 2504 0 1 264
box -8 -8 8 8
use VIA1  VIA1_4060
timestamp 1569139307
transform 1 0 2504 0 1 328
box -8 -8 8 8
use VIA1  VIA1_4061
timestamp 1569139307
transform 1 0 2504 0 1 392
box -8 -8 8 8
use VIA1  VIA1_4062
timestamp 1569139307
transform 1 0 2504 0 1 456
box -8 -8 8 8
use VIA1  VIA1_4063
timestamp 1569139307
transform 1 0 2504 0 1 520
box -8 -8 8 8
use VIA1  VIA1_4064
timestamp 1569139307
transform 1 0 2504 0 1 584
box -8 -8 8 8
use VIA1  VIA1_4065
timestamp 1569139307
transform 1 0 2504 0 1 648
box -8 -8 8 8
use VIA1  VIA1_4066
timestamp 1569139307
transform 1 0 2504 0 1 712
box -8 -8 8 8
use VIA1  VIA1_4067
timestamp 1569139307
transform 1 0 2504 0 1 776
box -8 -8 8 8
use VIA1  VIA1_4068
timestamp 1569139307
transform 1 0 2504 0 1 840
box -8 -8 8 8
use VIA1  VIA1_4069
timestamp 1569139307
transform 1 0 2504 0 1 904
box -8 -8 8 8
use VIA1  VIA1_4070
timestamp 1569139307
transform 1 0 2504 0 1 968
box -8 -8 8 8
use VIA1  VIA1_4071
timestamp 1569139307
transform 1 0 2504 0 1 1032
box -8 -8 8 8
use VIA1  VIA1_4072
timestamp 1569139307
transform 1 0 2504 0 1 1096
box -8 -8 8 8
use VIA1  VIA1_4073
timestamp 1569139307
transform 1 0 2504 0 1 1160
box -8 -8 8 8
use VIA1  VIA1_4074
timestamp 1569139307
transform 1 0 2504 0 1 1224
box -8 -8 8 8
use VIA1  VIA1_4075
timestamp 1569139307
transform 1 0 2504 0 1 1288
box -8 -8 8 8
use VIA1  VIA1_4076
timestamp 1569139307
transform 1 0 2504 0 1 1352
box -8 -8 8 8
use VIA1  VIA1_4077
timestamp 1569139307
transform 1 0 2504 0 1 1416
box -8 -8 8 8
use VIA1  VIA1_4078
timestamp 1569139307
transform 1 0 2504 0 1 1480
box -8 -8 8 8
use VIA1  VIA1_4079
timestamp 1569139307
transform 1 0 2504 0 1 1544
box -8 -8 8 8
use VIA1  VIA1_4080
timestamp 1569139307
transform 1 0 2504 0 1 1608
box -8 -8 8 8
use VIA1  VIA1_4081
timestamp 1569139307
transform 1 0 2504 0 1 1672
box -8 -8 8 8
use VIA1  VIA1_4082
timestamp 1569139307
transform 1 0 2504 0 1 1736
box -8 -8 8 8
use VIA1  VIA1_4083
timestamp 1569139307
transform 1 0 2504 0 1 1800
box -8 -8 8 8
use VIA1  VIA1_4084
timestamp 1569139307
transform 1 0 2504 0 1 1864
box -8 -8 8 8
use VIA1  VIA1_4085
timestamp 1569139307
transform 1 0 2504 0 1 1928
box -8 -8 8 8
use VIA1  VIA1_4086
timestamp 1569139307
transform 1 0 392 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4087
timestamp 1569139307
transform 1 0 1160 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4088
timestamp 1569139307
transform 1 0 1928 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4089
timestamp 1569139307
transform 1 0 3464 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4090
timestamp 1569139307
transform 1 0 4232 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4091
timestamp 1569139307
transform 1 0 456 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4092
timestamp 1569139307
transform 1 0 1224 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4093
timestamp 1569139307
transform 1 0 3528 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4094
timestamp 1569139307
transform 1 0 4296 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4095
timestamp 1569139307
transform 1 0 520 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4096
timestamp 1569139307
transform 1 0 1288 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4097
timestamp 1569139307
transform 1 0 3592 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4098
timestamp 1569139307
transform 1 0 4360 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4099
timestamp 1569139307
transform 1 0 584 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4100
timestamp 1569139307
transform 1 0 1352 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4101
timestamp 1569139307
transform 1 0 3656 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4102
timestamp 1569139307
transform 1 0 4424 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4103
timestamp 1569139307
transform 1 0 648 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4104
timestamp 1569139307
transform 1 0 1416 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4105
timestamp 1569139307
transform 1 0 3720 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4106
timestamp 1569139307
transform 1 0 4488 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4107
timestamp 1569139307
transform 1 0 712 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4108
timestamp 1569139307
transform 1 0 1480 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4109
timestamp 1569139307
transform 1 0 3784 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4110
timestamp 1569139307
transform 1 0 4552 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4111
timestamp 1569139307
transform 1 0 2504 0 1 3208
box -8 -8 8 8
use VIA1  VIA1_4112
timestamp 1569139307
transform 1 0 2504 0 1 3272
box -8 -8 8 8
use VIA1  VIA1_4113
timestamp 1569139307
transform 1 0 2504 0 1 3336
box -8 -8 8 8
use VIA1  VIA1_4114
timestamp 1569139307
transform 1 0 2504 0 1 3400
box -8 -8 8 8
use VIA1  VIA1_4115
timestamp 1569139307
transform 1 0 2504 0 1 3464
box -8 -8 8 8
use VIA1  VIA1_4116
timestamp 1569139307
transform 1 0 2504 0 1 3528
box -8 -8 8 8
use VIA1  VIA1_4117
timestamp 1569139307
transform 1 0 2504 0 1 3592
box -8 -8 8 8
use VIA1  VIA1_4118
timestamp 1569139307
transform 1 0 2504 0 1 3656
box -8 -8 8 8
use VIA1  VIA1_4119
timestamp 1569139307
transform 1 0 2504 0 1 3720
box -8 -8 8 8
use VIA1  VIA1_4120
timestamp 1569139307
transform 1 0 2504 0 1 3784
box -8 -8 8 8
use VIA1  VIA1_4121
timestamp 1569139307
transform 1 0 2504 0 1 3848
box -8 -8 8 8
use VIA1  VIA1_4122
timestamp 1569139307
transform 1 0 2504 0 1 3912
box -8 -8 8 8
use VIA1  VIA1_4123
timestamp 1569139307
transform 1 0 2504 0 1 3976
box -8 -8 8 8
use VIA1  VIA1_4124
timestamp 1569139307
transform 1 0 2504 0 1 4040
box -8 -8 8 8
use VIA1  VIA1_4125
timestamp 1569139307
transform 1 0 2504 0 1 4104
box -8 -8 8 8
use VIA1  VIA1_4126
timestamp 1569139307
transform 1 0 2504 0 1 4168
box -8 -8 8 8
use VIA1  VIA1_4127
timestamp 1569139307
transform 1 0 2504 0 1 4232
box -8 -8 8 8
use VIA1  VIA1_4128
timestamp 1569139307
transform 1 0 2504 0 1 4296
box -8 -8 8 8
use VIA1  VIA1_4129
timestamp 1569139307
transform 1 0 2504 0 1 4360
box -8 -8 8 8
use VIA1  VIA1_4130
timestamp 1569139307
transform 1 0 2504 0 1 4424
box -8 -8 8 8
use VIA1  VIA1_4131
timestamp 1569139307
transform 1 0 2504 0 1 4488
box -8 -8 8 8
use VIA1  VIA1_4132
timestamp 1569139307
transform 1 0 2504 0 1 4552
box -8 -8 8 8
use VIA1  VIA1_4133
timestamp 1569139307
transform 1 0 2504 0 1 72
box -8 -8 8 8
use VIA1  VIA1_4134
timestamp 1569139307
transform 1 0 776 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4135
timestamp 1569139307
transform 1 0 1544 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4136
timestamp 1569139307
transform 1 0 3848 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4137
timestamp 1569139307
transform 1 0 4616 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4138
timestamp 1569139307
transform 1 0 72 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4139
timestamp 1569139307
transform 1 0 840 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4140
timestamp 1569139307
transform 1 0 1608 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4141
timestamp 1569139307
transform 1 0 3912 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4142
timestamp 1569139307
transform 1 0 4680 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4143
timestamp 1569139307
transform 1 0 136 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4144
timestamp 1569139307
transform 1 0 904 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4145
timestamp 1569139307
transform 1 0 1672 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4146
timestamp 1569139307
transform 1 0 3208 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4147
timestamp 1569139307
transform 1 0 3976 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4148
timestamp 1569139307
transform 1 0 4744 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4149
timestamp 1569139307
transform 1 0 200 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4150
timestamp 1569139307
transform 1 0 968 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4151
timestamp 1569139307
transform 1 0 1736 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4152
timestamp 1569139307
transform 1 0 3272 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4153
timestamp 1569139307
transform 1 0 4040 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4154
timestamp 1569139307
transform 1 0 4808 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4155
timestamp 1569139307
transform 1 0 264 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4156
timestamp 1569139307
transform 1 0 1032 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4157
timestamp 1569139307
transform 1 0 1800 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4158
timestamp 1569139307
transform 1 0 3336 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4159
timestamp 1569139307
transform 1 0 4104 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4160
timestamp 1569139307
transform 1 0 4872 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4161
timestamp 1569139307
transform 1 0 328 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4162
timestamp 1569139307
transform 1 0 1096 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4163
timestamp 1569139307
transform 1 0 1864 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4164
timestamp 1569139307
transform 1 0 3400 0 1 2504
box -8 -8 8 8
use VIA1  VIA1_4165
timestamp 1569139307
transform 1 0 4168 0 1 2504
box -8 -8 8 8
use VIA2  VIA2_0
timestamp 1569139307
transform 1 0 4840 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1
timestamp 1569139307
transform 1 0 4776 0 1 104
box -8 -8 8 8
use VIA2  VIA2_2
timestamp 1569139307
transform 1 0 4712 0 1 232
box -8 -8 8 8
use VIA2  VIA2_3
timestamp 1569139307
transform 1 0 4712 0 1 168
box -8 -8 8 8
use VIA2  VIA2_4
timestamp 1569139307
transform 1 0 4712 0 1 296
box -8 -8 8 8
use VIA2  VIA2_5
timestamp 1569139307
transform 1 0 4776 0 1 296
box -8 -8 8 8
use VIA2  VIA2_6
timestamp 1569139307
transform 1 0 4904 0 1 40
box -8 -8 8 8
use VIA2  VIA2_7
timestamp 1569139307
transform 1 0 4776 0 1 168
box -8 -8 8 8
use VIA2  VIA2_8
timestamp 1569139307
transform 1 0 4904 0 1 232
box -8 -8 8 8
use VIA2  VIA2_9
timestamp 1569139307
transform 1 0 4712 0 1 104
box -8 -8 8 8
use VIA2  VIA2_10
timestamp 1569139307
transform 1 0 4904 0 1 104
box -8 -8 8 8
use VIA2  VIA2_11
timestamp 1569139307
transform 1 0 4840 0 1 104
box -8 -8 8 8
use VIA2  VIA2_12
timestamp 1569139307
transform 1 0 4712 0 1 40
box -8 -8 8 8
use VIA2  VIA2_13
timestamp 1569139307
transform 1 0 4776 0 1 40
box -8 -8 8 8
use VIA2  VIA2_14
timestamp 1569139307
transform 1 0 4904 0 1 168
box -8 -8 8 8
use VIA2  VIA2_15
timestamp 1569139307
transform 1 0 4840 0 1 296
box -8 -8 8 8
use VIA2  VIA2_16
timestamp 1569139307
transform 1 0 4904 0 1 296
box -8 -8 8 8
use VIA2  VIA2_17
timestamp 1569139307
transform 1 0 4776 0 1 232
box -8 -8 8 8
use VIA2  VIA2_18
timestamp 1569139307
transform 1 0 4840 0 1 232
box -8 -8 8 8
use VIA2  VIA2_19
timestamp 1569139307
transform 1 0 4840 0 1 168
box -8 -8 8 8
use VIA2  VIA2_20
timestamp 1569139307
transform 1 0 4584 0 1 40
box -8 -8 8 8
use VIA2  VIA2_21
timestamp 1569139307
transform 1 0 4520 0 1 232
box -8 -8 8 8
use VIA2  VIA2_22
timestamp 1569139307
transform 1 0 4584 0 1 232
box -8 -8 8 8
use VIA2  VIA2_23
timestamp 1569139307
transform 1 0 4456 0 1 232
box -8 -8 8 8
use VIA2  VIA2_24
timestamp 1569139307
transform 1 0 4648 0 1 232
box -8 -8 8 8
use VIA2  VIA2_25
timestamp 1569139307
transform 1 0 4648 0 1 104
box -8 -8 8 8
use VIA2  VIA2_26
timestamp 1569139307
transform 1 0 4456 0 1 104
box -8 -8 8 8
use VIA2  VIA2_27
timestamp 1569139307
transform 1 0 4456 0 1 168
box -8 -8 8 8
use VIA2  VIA2_28
timestamp 1569139307
transform 1 0 4584 0 1 104
box -8 -8 8 8
use VIA2  VIA2_29
timestamp 1569139307
transform 1 0 4392 0 1 168
box -8 -8 8 8
use VIA2  VIA2_30
timestamp 1569139307
transform 1 0 4520 0 1 296
box -8 -8 8 8
use VIA2  VIA2_31
timestamp 1569139307
transform 1 0 4648 0 1 296
box -8 -8 8 8
use VIA2  VIA2_32
timestamp 1569139307
transform 1 0 4584 0 1 296
box -8 -8 8 8
use VIA2  VIA2_33
timestamp 1569139307
transform 1 0 4520 0 1 168
box -8 -8 8 8
use VIA2  VIA2_34
timestamp 1569139307
transform 1 0 4520 0 1 104
box -8 -8 8 8
use VIA2  VIA2_35
timestamp 1569139307
transform 1 0 4584 0 1 168
box -8 -8 8 8
use VIA2  VIA2_36
timestamp 1569139307
transform 1 0 4392 0 1 104
box -8 -8 8 8
use VIA2  VIA2_37
timestamp 1569139307
transform 1 0 4456 0 1 296
box -8 -8 8 8
use VIA2  VIA2_38
timestamp 1569139307
transform 1 0 4392 0 1 232
box -8 -8 8 8
use VIA2  VIA2_39
timestamp 1569139307
transform 1 0 4392 0 1 40
box -8 -8 8 8
use VIA2  VIA2_40
timestamp 1569139307
transform 1 0 4648 0 1 168
box -8 -8 8 8
use VIA2  VIA2_41
timestamp 1569139307
transform 1 0 4520 0 1 40
box -8 -8 8 8
use VIA2  VIA2_42
timestamp 1569139307
transform 1 0 4648 0 1 40
box -8 -8 8 8
use VIA2  VIA2_43
timestamp 1569139307
transform 1 0 4456 0 1 40
box -8 -8 8 8
use VIA2  VIA2_44
timestamp 1569139307
transform 1 0 4392 0 1 296
box -8 -8 8 8
use VIA2  VIA2_45
timestamp 1569139307
transform 1 0 4584 0 1 616
box -8 -8 8 8
use VIA2  VIA2_46
timestamp 1569139307
transform 1 0 4456 0 1 424
box -8 -8 8 8
use VIA2  VIA2_47
timestamp 1569139307
transform 1 0 4520 0 1 488
box -8 -8 8 8
use VIA2  VIA2_48
timestamp 1569139307
transform 1 0 4456 0 1 488
box -8 -8 8 8
use VIA2  VIA2_49
timestamp 1569139307
transform 1 0 4584 0 1 360
box -8 -8 8 8
use VIA2  VIA2_50
timestamp 1569139307
transform 1 0 4392 0 1 616
box -8 -8 8 8
use VIA2  VIA2_51
timestamp 1569139307
transform 1 0 4584 0 1 552
box -8 -8 8 8
use VIA2  VIA2_52
timestamp 1569139307
transform 1 0 4648 0 1 616
box -8 -8 8 8
use VIA2  VIA2_53
timestamp 1569139307
transform 1 0 4520 0 1 616
box -8 -8 8 8
use VIA2  VIA2_54
timestamp 1569139307
transform 1 0 4456 0 1 552
box -8 -8 8 8
use VIA2  VIA2_55
timestamp 1569139307
transform 1 0 4520 0 1 552
box -8 -8 8 8
use VIA2  VIA2_56
timestamp 1569139307
transform 1 0 4456 0 1 616
box -8 -8 8 8
use VIA2  VIA2_57
timestamp 1569139307
transform 1 0 4648 0 1 552
box -8 -8 8 8
use VIA2  VIA2_58
timestamp 1569139307
transform 1 0 4648 0 1 360
box -8 -8 8 8
use VIA2  VIA2_59
timestamp 1569139307
transform 1 0 4520 0 1 360
box -8 -8 8 8
use VIA2  VIA2_60
timestamp 1569139307
transform 1 0 4584 0 1 424
box -8 -8 8 8
use VIA2  VIA2_61
timestamp 1569139307
transform 1 0 4648 0 1 424
box -8 -8 8 8
use VIA2  VIA2_62
timestamp 1569139307
transform 1 0 4392 0 1 360
box -8 -8 8 8
use VIA2  VIA2_63
timestamp 1569139307
transform 1 0 4520 0 1 424
box -8 -8 8 8
use VIA2  VIA2_64
timestamp 1569139307
transform 1 0 4392 0 1 424
box -8 -8 8 8
use VIA2  VIA2_65
timestamp 1569139307
transform 1 0 4648 0 1 488
box -8 -8 8 8
use VIA2  VIA2_66
timestamp 1569139307
transform 1 0 4392 0 1 488
box -8 -8 8 8
use VIA2  VIA2_67
timestamp 1569139307
transform 1 0 4456 0 1 360
box -8 -8 8 8
use VIA2  VIA2_68
timestamp 1569139307
transform 1 0 4392 0 1 552
box -8 -8 8 8
use VIA2  VIA2_69
timestamp 1569139307
transform 1 0 4584 0 1 488
box -8 -8 8 8
use VIA2  VIA2_70
timestamp 1569139307
transform 1 0 4776 0 1 552
box -8 -8 8 8
use VIA2  VIA2_71
timestamp 1569139307
transform 1 0 4712 0 1 616
box -8 -8 8 8
use VIA2  VIA2_72
timestamp 1569139307
transform 1 0 4840 0 1 552
box -8 -8 8 8
use VIA2  VIA2_73
timestamp 1569139307
transform 1 0 4904 0 1 488
box -8 -8 8 8
use VIA2  VIA2_74
timestamp 1569139307
transform 1 0 4904 0 1 616
box -8 -8 8 8
use VIA2  VIA2_75
timestamp 1569139307
transform 1 0 4904 0 1 360
box -8 -8 8 8
use VIA2  VIA2_76
timestamp 1569139307
transform 1 0 4840 0 1 616
box -8 -8 8 8
use VIA2  VIA2_77
timestamp 1569139307
transform 1 0 4776 0 1 360
box -8 -8 8 8
use VIA2  VIA2_78
timestamp 1569139307
transform 1 0 4904 0 1 552
box -8 -8 8 8
use VIA2  VIA2_79
timestamp 1569139307
transform 1 0 4776 0 1 424
box -8 -8 8 8
use VIA2  VIA2_80
timestamp 1569139307
transform 1 0 4840 0 1 360
box -8 -8 8 8
use VIA2  VIA2_81
timestamp 1569139307
transform 1 0 4712 0 1 552
box -8 -8 8 8
use VIA2  VIA2_82
timestamp 1569139307
transform 1 0 4712 0 1 424
box -8 -8 8 8
use VIA2  VIA2_83
timestamp 1569139307
transform 1 0 4840 0 1 424
box -8 -8 8 8
use VIA2  VIA2_84
timestamp 1569139307
transform 1 0 4904 0 1 424
box -8 -8 8 8
use VIA2  VIA2_85
timestamp 1569139307
transform 1 0 4776 0 1 488
box -8 -8 8 8
use VIA2  VIA2_86
timestamp 1569139307
transform 1 0 4712 0 1 488
box -8 -8 8 8
use VIA2  VIA2_87
timestamp 1569139307
transform 1 0 4840 0 1 488
box -8 -8 8 8
use VIA2  VIA2_88
timestamp 1569139307
transform 1 0 4712 0 1 360
box -8 -8 8 8
use VIA2  VIA2_89
timestamp 1569139307
transform 1 0 4776 0 1 616
box -8 -8 8 8
use VIA2  VIA2_90
timestamp 1569139307
transform 1 0 4136 0 1 232
box -8 -8 8 8
use VIA2  VIA2_91
timestamp 1569139307
transform 1 0 4264 0 1 296
box -8 -8 8 8
use VIA2  VIA2_92
timestamp 1569139307
transform 1 0 4200 0 1 40
box -8 -8 8 8
use VIA2  VIA2_93
timestamp 1569139307
transform 1 0 4200 0 1 104
box -8 -8 8 8
use VIA2  VIA2_94
timestamp 1569139307
transform 1 0 4200 0 1 232
box -8 -8 8 8
use VIA2  VIA2_95
timestamp 1569139307
transform 1 0 4072 0 1 168
box -8 -8 8 8
use VIA2  VIA2_96
timestamp 1569139307
transform 1 0 4072 0 1 40
box -8 -8 8 8
use VIA2  VIA2_97
timestamp 1569139307
transform 1 0 4136 0 1 296
box -8 -8 8 8
use VIA2  VIA2_98
timestamp 1569139307
transform 1 0 4200 0 1 168
box -8 -8 8 8
use VIA2  VIA2_99
timestamp 1569139307
transform 1 0 4072 0 1 232
box -8 -8 8 8
use VIA2  VIA2_100
timestamp 1569139307
transform 1 0 4072 0 1 104
box -8 -8 8 8
use VIA2  VIA2_101
timestamp 1569139307
transform 1 0 4328 0 1 40
box -8 -8 8 8
use VIA2  VIA2_102
timestamp 1569139307
transform 1 0 4136 0 1 40
box -8 -8 8 8
use VIA2  VIA2_103
timestamp 1569139307
transform 1 0 4328 0 1 232
box -8 -8 8 8
use VIA2  VIA2_104
timestamp 1569139307
transform 1 0 4264 0 1 104
box -8 -8 8 8
use VIA2  VIA2_105
timestamp 1569139307
transform 1 0 4200 0 1 296
box -8 -8 8 8
use VIA2  VIA2_106
timestamp 1569139307
transform 1 0 4136 0 1 168
box -8 -8 8 8
use VIA2  VIA2_107
timestamp 1569139307
transform 1 0 4328 0 1 104
box -8 -8 8 8
use VIA2  VIA2_108
timestamp 1569139307
transform 1 0 4328 0 1 168
box -8 -8 8 8
use VIA2  VIA2_109
timestamp 1569139307
transform 1 0 4264 0 1 232
box -8 -8 8 8
use VIA2  VIA2_110
timestamp 1569139307
transform 1 0 4264 0 1 40
box -8 -8 8 8
use VIA2  VIA2_111
timestamp 1569139307
transform 1 0 4264 0 1 168
box -8 -8 8 8
use VIA2  VIA2_112
timestamp 1569139307
transform 1 0 4072 0 1 296
box -8 -8 8 8
use VIA2  VIA2_113
timestamp 1569139307
transform 1 0 4136 0 1 104
box -8 -8 8 8
use VIA2  VIA2_114
timestamp 1569139307
transform 1 0 4328 0 1 296
box -8 -8 8 8
use VIA2  VIA2_115
timestamp 1569139307
transform 1 0 3816 0 1 232
box -8 -8 8 8
use VIA2  VIA2_116
timestamp 1569139307
transform 1 0 3880 0 1 296
box -8 -8 8 8
use VIA2  VIA2_117
timestamp 1569139307
transform 1 0 4008 0 1 168
box -8 -8 8 8
use VIA2  VIA2_118
timestamp 1569139307
transform 1 0 3816 0 1 104
box -8 -8 8 8
use VIA2  VIA2_119
timestamp 1569139307
transform 1 0 3944 0 1 104
box -8 -8 8 8
use VIA2  VIA2_120
timestamp 1569139307
transform 1 0 3752 0 1 104
box -8 -8 8 8
use VIA2  VIA2_121
timestamp 1569139307
transform 1 0 3944 0 1 232
box -8 -8 8 8
use VIA2  VIA2_122
timestamp 1569139307
transform 1 0 3880 0 1 232
box -8 -8 8 8
use VIA2  VIA2_123
timestamp 1569139307
transform 1 0 4008 0 1 232
box -8 -8 8 8
use VIA2  VIA2_124
timestamp 1569139307
transform 1 0 3944 0 1 168
box -8 -8 8 8
use VIA2  VIA2_125
timestamp 1569139307
transform 1 0 3944 0 1 40
box -8 -8 8 8
use VIA2  VIA2_126
timestamp 1569139307
transform 1 0 3880 0 1 40
box -8 -8 8 8
use VIA2  VIA2_127
timestamp 1569139307
transform 1 0 3752 0 1 40
box -8 -8 8 8
use VIA2  VIA2_128
timestamp 1569139307
transform 1 0 4008 0 1 296
box -8 -8 8 8
use VIA2  VIA2_129
timestamp 1569139307
transform 1 0 3752 0 1 232
box -8 -8 8 8
use VIA2  VIA2_130
timestamp 1569139307
transform 1 0 4008 0 1 40
box -8 -8 8 8
use VIA2  VIA2_131
timestamp 1569139307
transform 1 0 3944 0 1 296
box -8 -8 8 8
use VIA2  VIA2_132
timestamp 1569139307
transform 1 0 3880 0 1 168
box -8 -8 8 8
use VIA2  VIA2_133
timestamp 1569139307
transform 1 0 3816 0 1 168
box -8 -8 8 8
use VIA2  VIA2_134
timestamp 1569139307
transform 1 0 4008 0 1 104
box -8 -8 8 8
use VIA2  VIA2_135
timestamp 1569139307
transform 1 0 3752 0 1 296
box -8 -8 8 8
use VIA2  VIA2_136
timestamp 1569139307
transform 1 0 3752 0 1 168
box -8 -8 8 8
use VIA2  VIA2_137
timestamp 1569139307
transform 1 0 3816 0 1 296
box -8 -8 8 8
use VIA2  VIA2_138
timestamp 1569139307
transform 1 0 3880 0 1 104
box -8 -8 8 8
use VIA2  VIA2_139
timestamp 1569139307
transform 1 0 3816 0 1 40
box -8 -8 8 8
use VIA2  VIA2_140
timestamp 1569139307
transform 1 0 3752 0 1 488
box -8 -8 8 8
use VIA2  VIA2_141
timestamp 1569139307
transform 1 0 3880 0 1 616
box -8 -8 8 8
use VIA2  VIA2_142
timestamp 1569139307
transform 1 0 3944 0 1 552
box -8 -8 8 8
use VIA2  VIA2_143
timestamp 1569139307
transform 1 0 3752 0 1 552
box -8 -8 8 8
use VIA2  VIA2_144
timestamp 1569139307
transform 1 0 3816 0 1 616
box -8 -8 8 8
use VIA2  VIA2_145
timestamp 1569139307
transform 1 0 3752 0 1 616
box -8 -8 8 8
use VIA2  VIA2_146
timestamp 1569139307
transform 1 0 3944 0 1 616
box -8 -8 8 8
use VIA2  VIA2_147
timestamp 1569139307
transform 1 0 4008 0 1 360
box -8 -8 8 8
use VIA2  VIA2_148
timestamp 1569139307
transform 1 0 4008 0 1 552
box -8 -8 8 8
use VIA2  VIA2_149
timestamp 1569139307
transform 1 0 3880 0 1 360
box -8 -8 8 8
use VIA2  VIA2_150
timestamp 1569139307
transform 1 0 4008 0 1 424
box -8 -8 8 8
use VIA2  VIA2_151
timestamp 1569139307
transform 1 0 3944 0 1 360
box -8 -8 8 8
use VIA2  VIA2_152
timestamp 1569139307
transform 1 0 3880 0 1 424
box -8 -8 8 8
use VIA2  VIA2_153
timestamp 1569139307
transform 1 0 4008 0 1 616
box -8 -8 8 8
use VIA2  VIA2_154
timestamp 1569139307
transform 1 0 3880 0 1 552
box -8 -8 8 8
use VIA2  VIA2_155
timestamp 1569139307
transform 1 0 3752 0 1 424
box -8 -8 8 8
use VIA2  VIA2_156
timestamp 1569139307
transform 1 0 3816 0 1 360
box -8 -8 8 8
use VIA2  VIA2_157
timestamp 1569139307
transform 1 0 4008 0 1 488
box -8 -8 8 8
use VIA2  VIA2_158
timestamp 1569139307
transform 1 0 3944 0 1 424
box -8 -8 8 8
use VIA2  VIA2_159
timestamp 1569139307
transform 1 0 3816 0 1 424
box -8 -8 8 8
use VIA2  VIA2_160
timestamp 1569139307
transform 1 0 3816 0 1 488
box -8 -8 8 8
use VIA2  VIA2_161
timestamp 1569139307
transform 1 0 3944 0 1 488
box -8 -8 8 8
use VIA2  VIA2_162
timestamp 1569139307
transform 1 0 3752 0 1 360
box -8 -8 8 8
use VIA2  VIA2_163
timestamp 1569139307
transform 1 0 3816 0 1 552
box -8 -8 8 8
use VIA2  VIA2_164
timestamp 1569139307
transform 1 0 3880 0 1 488
box -8 -8 8 8
use VIA2  VIA2_165
timestamp 1569139307
transform 1 0 4200 0 1 360
box -8 -8 8 8
use VIA2  VIA2_166
timestamp 1569139307
transform 1 0 4072 0 1 616
box -8 -8 8 8
use VIA2  VIA2_167
timestamp 1569139307
transform 1 0 4200 0 1 424
box -8 -8 8 8
use VIA2  VIA2_168
timestamp 1569139307
transform 1 0 4264 0 1 552
box -8 -8 8 8
use VIA2  VIA2_169
timestamp 1569139307
transform 1 0 4072 0 1 424
box -8 -8 8 8
use VIA2  VIA2_170
timestamp 1569139307
transform 1 0 4136 0 1 360
box -8 -8 8 8
use VIA2  VIA2_171
timestamp 1569139307
transform 1 0 4200 0 1 488
box -8 -8 8 8
use VIA2  VIA2_172
timestamp 1569139307
transform 1 0 4264 0 1 360
box -8 -8 8 8
use VIA2  VIA2_173
timestamp 1569139307
transform 1 0 4328 0 1 360
box -8 -8 8 8
use VIA2  VIA2_174
timestamp 1569139307
transform 1 0 4136 0 1 424
box -8 -8 8 8
use VIA2  VIA2_175
timestamp 1569139307
transform 1 0 4136 0 1 488
box -8 -8 8 8
use VIA2  VIA2_176
timestamp 1569139307
transform 1 0 4328 0 1 424
box -8 -8 8 8
use VIA2  VIA2_177
timestamp 1569139307
transform 1 0 4072 0 1 552
box -8 -8 8 8
use VIA2  VIA2_178
timestamp 1569139307
transform 1 0 4328 0 1 488
box -8 -8 8 8
use VIA2  VIA2_179
timestamp 1569139307
transform 1 0 4200 0 1 552
box -8 -8 8 8
use VIA2  VIA2_180
timestamp 1569139307
transform 1 0 4328 0 1 552
box -8 -8 8 8
use VIA2  VIA2_181
timestamp 1569139307
transform 1 0 4264 0 1 616
box -8 -8 8 8
use VIA2  VIA2_182
timestamp 1569139307
transform 1 0 4328 0 1 616
box -8 -8 8 8
use VIA2  VIA2_183
timestamp 1569139307
transform 1 0 4200 0 1 616
box -8 -8 8 8
use VIA2  VIA2_184
timestamp 1569139307
transform 1 0 4264 0 1 424
box -8 -8 8 8
use VIA2  VIA2_185
timestamp 1569139307
transform 1 0 4072 0 1 360
box -8 -8 8 8
use VIA2  VIA2_186
timestamp 1569139307
transform 1 0 4136 0 1 552
box -8 -8 8 8
use VIA2  VIA2_187
timestamp 1569139307
transform 1 0 4264 0 1 488
box -8 -8 8 8
use VIA2  VIA2_188
timestamp 1569139307
transform 1 0 4072 0 1 488
box -8 -8 8 8
use VIA2  VIA2_189
timestamp 1569139307
transform 1 0 4136 0 1 616
box -8 -8 8 8
use VIA2  VIA2_190
timestamp 1569139307
transform 1 0 4136 0 1 744
box -8 -8 8 8
use VIA2  VIA2_191
timestamp 1569139307
transform 1 0 4264 0 1 808
box -8 -8 8 8
use VIA2  VIA2_192
timestamp 1569139307
transform 1 0 4200 0 1 680
box -8 -8 8 8
use VIA2  VIA2_193
timestamp 1569139307
transform 1 0 4072 0 1 808
box -8 -8 8 8
use VIA2  VIA2_194
timestamp 1569139307
transform 1 0 4264 0 1 936
box -8 -8 8 8
use VIA2  VIA2_195
timestamp 1569139307
transform 1 0 4328 0 1 872
box -8 -8 8 8
use VIA2  VIA2_196
timestamp 1569139307
transform 1 0 4072 0 1 744
box -8 -8 8 8
use VIA2  VIA2_197
timestamp 1569139307
transform 1 0 4328 0 1 680
box -8 -8 8 8
use VIA2  VIA2_198
timestamp 1569139307
transform 1 0 4136 0 1 680
box -8 -8 8 8
use VIA2  VIA2_199
timestamp 1569139307
transform 1 0 4200 0 1 936
box -8 -8 8 8
use VIA2  VIA2_200
timestamp 1569139307
transform 1 0 4136 0 1 872
box -8 -8 8 8
use VIA2  VIA2_201
timestamp 1569139307
transform 1 0 4264 0 1 872
box -8 -8 8 8
use VIA2  VIA2_202
timestamp 1569139307
transform 1 0 4328 0 1 744
box -8 -8 8 8
use VIA2  VIA2_203
timestamp 1569139307
transform 1 0 4200 0 1 744
box -8 -8 8 8
use VIA2  VIA2_204
timestamp 1569139307
transform 1 0 4072 0 1 936
box -8 -8 8 8
use VIA2  VIA2_205
timestamp 1569139307
transform 1 0 4136 0 1 936
box -8 -8 8 8
use VIA2  VIA2_206
timestamp 1569139307
transform 1 0 4200 0 1 872
box -8 -8 8 8
use VIA2  VIA2_207
timestamp 1569139307
transform 1 0 4264 0 1 680
box -8 -8 8 8
use VIA2  VIA2_208
timestamp 1569139307
transform 1 0 4072 0 1 872
box -8 -8 8 8
use VIA2  VIA2_209
timestamp 1569139307
transform 1 0 4136 0 1 808
box -8 -8 8 8
use VIA2  VIA2_210
timestamp 1569139307
transform 1 0 4328 0 1 808
box -8 -8 8 8
use VIA2  VIA2_211
timestamp 1569139307
transform 1 0 4264 0 1 744
box -8 -8 8 8
use VIA2  VIA2_212
timestamp 1569139307
transform 1 0 4328 0 1 936
box -8 -8 8 8
use VIA2  VIA2_213
timestamp 1569139307
transform 1 0 4072 0 1 680
box -8 -8 8 8
use VIA2  VIA2_214
timestamp 1569139307
transform 1 0 4200 0 1 808
box -8 -8 8 8
use VIA2  VIA2_215
timestamp 1569139307
transform 1 0 3816 0 1 872
box -8 -8 8 8
use VIA2  VIA2_216
timestamp 1569139307
transform 1 0 4008 0 1 744
box -8 -8 8 8
use VIA2  VIA2_217
timestamp 1569139307
transform 1 0 4008 0 1 808
box -8 -8 8 8
use VIA2  VIA2_218
timestamp 1569139307
transform 1 0 3752 0 1 744
box -8 -8 8 8
use VIA2  VIA2_219
timestamp 1569139307
transform 1 0 3880 0 1 936
box -8 -8 8 8
use VIA2  VIA2_220
timestamp 1569139307
transform 1 0 3816 0 1 936
box -8 -8 8 8
use VIA2  VIA2_221
timestamp 1569139307
transform 1 0 3944 0 1 936
box -8 -8 8 8
use VIA2  VIA2_222
timestamp 1569139307
transform 1 0 3752 0 1 808
box -8 -8 8 8
use VIA2  VIA2_223
timestamp 1569139307
transform 1 0 3944 0 1 808
box -8 -8 8 8
use VIA2  VIA2_224
timestamp 1569139307
transform 1 0 3816 0 1 680
box -8 -8 8 8
use VIA2  VIA2_225
timestamp 1569139307
transform 1 0 3816 0 1 808
box -8 -8 8 8
use VIA2  VIA2_226
timestamp 1569139307
transform 1 0 3752 0 1 872
box -8 -8 8 8
use VIA2  VIA2_227
timestamp 1569139307
transform 1 0 3752 0 1 936
box -8 -8 8 8
use VIA2  VIA2_228
timestamp 1569139307
transform 1 0 3944 0 1 872
box -8 -8 8 8
use VIA2  VIA2_229
timestamp 1569139307
transform 1 0 4008 0 1 936
box -8 -8 8 8
use VIA2  VIA2_230
timestamp 1569139307
transform 1 0 3880 0 1 680
box -8 -8 8 8
use VIA2  VIA2_231
timestamp 1569139307
transform 1 0 4008 0 1 872
box -8 -8 8 8
use VIA2  VIA2_232
timestamp 1569139307
transform 1 0 4008 0 1 680
box -8 -8 8 8
use VIA2  VIA2_233
timestamp 1569139307
transform 1 0 3816 0 1 744
box -8 -8 8 8
use VIA2  VIA2_234
timestamp 1569139307
transform 1 0 3880 0 1 744
box -8 -8 8 8
use VIA2  VIA2_235
timestamp 1569139307
transform 1 0 3944 0 1 680
box -8 -8 8 8
use VIA2  VIA2_236
timestamp 1569139307
transform 1 0 3944 0 1 744
box -8 -8 8 8
use VIA2  VIA2_237
timestamp 1569139307
transform 1 0 3880 0 1 808
box -8 -8 8 8
use VIA2  VIA2_238
timestamp 1569139307
transform 1 0 3752 0 1 680
box -8 -8 8 8
use VIA2  VIA2_239
timestamp 1569139307
transform 1 0 3880 0 1 872
box -8 -8 8 8
use VIA2  VIA2_240
timestamp 1569139307
transform 1 0 3816 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_241
timestamp 1569139307
transform 1 0 4008 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_242
timestamp 1569139307
transform 1 0 3880 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_243
timestamp 1569139307
transform 1 0 3944 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_244
timestamp 1569139307
transform 1 0 3944 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_245
timestamp 1569139307
transform 1 0 3816 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_246
timestamp 1569139307
transform 1 0 3880 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_247
timestamp 1569139307
transform 1 0 4008 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_248
timestamp 1569139307
transform 1 0 3880 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_249
timestamp 1569139307
transform 1 0 3816 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_250
timestamp 1569139307
transform 1 0 3816 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_251
timestamp 1569139307
transform 1 0 4008 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_252
timestamp 1569139307
transform 1 0 3944 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_253
timestamp 1569139307
transform 1 0 3944 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_254
timestamp 1569139307
transform 1 0 3944 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_255
timestamp 1569139307
transform 1 0 3752 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_256
timestamp 1569139307
transform 1 0 3816 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_257
timestamp 1569139307
transform 1 0 3752 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_258
timestamp 1569139307
transform 1 0 4008 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_259
timestamp 1569139307
transform 1 0 3752 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_260
timestamp 1569139307
transform 1 0 3752 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_261
timestamp 1569139307
transform 1 0 3752 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_262
timestamp 1569139307
transform 1 0 4008 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_263
timestamp 1569139307
transform 1 0 3880 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_264
timestamp 1569139307
transform 1 0 3880 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_265
timestamp 1569139307
transform 1 0 4328 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_266
timestamp 1569139307
transform 1 0 4200 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_267
timestamp 1569139307
transform 1 0 4264 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_268
timestamp 1569139307
transform 1 0 4200 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_269
timestamp 1569139307
transform 1 0 4328 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_270
timestamp 1569139307
transform 1 0 4072 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_271
timestamp 1569139307
transform 1 0 4136 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_272
timestamp 1569139307
transform 1 0 4328 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_273
timestamp 1569139307
transform 1 0 4072 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_274
timestamp 1569139307
transform 1 0 4264 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_275
timestamp 1569139307
transform 1 0 4136 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_276
timestamp 1569139307
transform 1 0 4072 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_277
timestamp 1569139307
transform 1 0 4264 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_278
timestamp 1569139307
transform 1 0 4200 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_279
timestamp 1569139307
transform 1 0 4136 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_280
timestamp 1569139307
transform 1 0 4136 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_281
timestamp 1569139307
transform 1 0 4328 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_282
timestamp 1569139307
transform 1 0 4136 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_283
timestamp 1569139307
transform 1 0 4200 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_284
timestamp 1569139307
transform 1 0 4072 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_285
timestamp 1569139307
transform 1 0 4328 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_286
timestamp 1569139307
transform 1 0 4264 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_287
timestamp 1569139307
transform 1 0 4200 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_288
timestamp 1569139307
transform 1 0 4264 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_289
timestamp 1569139307
transform 1 0 4072 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_290
timestamp 1569139307
transform 1 0 4712 0 1 808
box -8 -8 8 8
use VIA2  VIA2_291
timestamp 1569139307
transform 1 0 4712 0 1 936
box -8 -8 8 8
use VIA2  VIA2_292
timestamp 1569139307
transform 1 0 4904 0 1 936
box -8 -8 8 8
use VIA2  VIA2_293
timestamp 1569139307
transform 1 0 4776 0 1 680
box -8 -8 8 8
use VIA2  VIA2_294
timestamp 1569139307
transform 1 0 4776 0 1 872
box -8 -8 8 8
use VIA2  VIA2_295
timestamp 1569139307
transform 1 0 4904 0 1 872
box -8 -8 8 8
use VIA2  VIA2_296
timestamp 1569139307
transform 1 0 4840 0 1 872
box -8 -8 8 8
use VIA2  VIA2_297
timestamp 1569139307
transform 1 0 4904 0 1 680
box -8 -8 8 8
use VIA2  VIA2_298
timestamp 1569139307
transform 1 0 4840 0 1 680
box -8 -8 8 8
use VIA2  VIA2_299
timestamp 1569139307
transform 1 0 4904 0 1 808
box -8 -8 8 8
use VIA2  VIA2_300
timestamp 1569139307
transform 1 0 4840 0 1 936
box -8 -8 8 8
use VIA2  VIA2_301
timestamp 1569139307
transform 1 0 4776 0 1 744
box -8 -8 8 8
use VIA2  VIA2_302
timestamp 1569139307
transform 1 0 4840 0 1 744
box -8 -8 8 8
use VIA2  VIA2_303
timestamp 1569139307
transform 1 0 4776 0 1 936
box -8 -8 8 8
use VIA2  VIA2_304
timestamp 1569139307
transform 1 0 4904 0 1 744
box -8 -8 8 8
use VIA2  VIA2_305
timestamp 1569139307
transform 1 0 4712 0 1 872
box -8 -8 8 8
use VIA2  VIA2_306
timestamp 1569139307
transform 1 0 4712 0 1 744
box -8 -8 8 8
use VIA2  VIA2_307
timestamp 1569139307
transform 1 0 4776 0 1 808
box -8 -8 8 8
use VIA2  VIA2_308
timestamp 1569139307
transform 1 0 4712 0 1 680
box -8 -8 8 8
use VIA2  VIA2_309
timestamp 1569139307
transform 1 0 4840 0 1 808
box -8 -8 8 8
use VIA2  VIA2_310
timestamp 1569139307
transform 1 0 4520 0 1 744
box -8 -8 8 8
use VIA2  VIA2_311
timestamp 1569139307
transform 1 0 4520 0 1 808
box -8 -8 8 8
use VIA2  VIA2_312
timestamp 1569139307
transform 1 0 4520 0 1 872
box -8 -8 8 8
use VIA2  VIA2_313
timestamp 1569139307
transform 1 0 4520 0 1 936
box -8 -8 8 8
use VIA2  VIA2_314
timestamp 1569139307
transform 1 0 4392 0 1 680
box -8 -8 8 8
use VIA2  VIA2_315
timestamp 1569139307
transform 1 0 4392 0 1 744
box -8 -8 8 8
use VIA2  VIA2_316
timestamp 1569139307
transform 1 0 4392 0 1 808
box -8 -8 8 8
use VIA2  VIA2_317
timestamp 1569139307
transform 1 0 4392 0 1 872
box -8 -8 8 8
use VIA2  VIA2_318
timestamp 1569139307
transform 1 0 4392 0 1 936
box -8 -8 8 8
use VIA2  VIA2_319
timestamp 1569139307
transform 1 0 4584 0 1 680
box -8 -8 8 8
use VIA2  VIA2_320
timestamp 1569139307
transform 1 0 4584 0 1 744
box -8 -8 8 8
use VIA2  VIA2_321
timestamp 1569139307
transform 1 0 4648 0 1 680
box -8 -8 8 8
use VIA2  VIA2_322
timestamp 1569139307
transform 1 0 4648 0 1 808
box -8 -8 8 8
use VIA2  VIA2_323
timestamp 1569139307
transform 1 0 4648 0 1 872
box -8 -8 8 8
use VIA2  VIA2_324
timestamp 1569139307
transform 1 0 4584 0 1 808
box -8 -8 8 8
use VIA2  VIA2_325
timestamp 1569139307
transform 1 0 4456 0 1 680
box -8 -8 8 8
use VIA2  VIA2_326
timestamp 1569139307
transform 1 0 4456 0 1 744
box -8 -8 8 8
use VIA2  VIA2_327
timestamp 1569139307
transform 1 0 4456 0 1 808
box -8 -8 8 8
use VIA2  VIA2_328
timestamp 1569139307
transform 1 0 4648 0 1 936
box -8 -8 8 8
use VIA2  VIA2_329
timestamp 1569139307
transform 1 0 4584 0 1 872
box -8 -8 8 8
use VIA2  VIA2_330
timestamp 1569139307
transform 1 0 4456 0 1 872
box -8 -8 8 8
use VIA2  VIA2_331
timestamp 1569139307
transform 1 0 4456 0 1 936
box -8 -8 8 8
use VIA2  VIA2_332
timestamp 1569139307
transform 1 0 4648 0 1 744
box -8 -8 8 8
use VIA2  VIA2_333
timestamp 1569139307
transform 1 0 4584 0 1 936
box -8 -8 8 8
use VIA2  VIA2_334
timestamp 1569139307
transform 1 0 4520 0 1 680
box -8 -8 8 8
use VIA2  VIA2_335
timestamp 1569139307
transform 1 0 4648 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_336
timestamp 1569139307
transform 1 0 4456 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_337
timestamp 1569139307
transform 1 0 4520 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_338
timestamp 1569139307
transform 1 0 4584 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_339
timestamp 1569139307
transform 1 0 4456 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_340
timestamp 1569139307
transform 1 0 4520 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_341
timestamp 1569139307
transform 1 0 4392 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_342
timestamp 1569139307
transform 1 0 4520 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_343
timestamp 1569139307
transform 1 0 4648 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_344
timestamp 1569139307
transform 1 0 4456 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_345
timestamp 1569139307
transform 1 0 4520 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_346
timestamp 1569139307
transform 1 0 4584 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_347
timestamp 1569139307
transform 1 0 4392 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_348
timestamp 1569139307
transform 1 0 4648 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_349
timestamp 1569139307
transform 1 0 4520 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_350
timestamp 1569139307
transform 1 0 4392 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_351
timestamp 1569139307
transform 1 0 4392 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_352
timestamp 1569139307
transform 1 0 4584 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_353
timestamp 1569139307
transform 1 0 4456 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_354
timestamp 1569139307
transform 1 0 4648 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_355
timestamp 1569139307
transform 1 0 4584 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_356
timestamp 1569139307
transform 1 0 4392 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_357
timestamp 1569139307
transform 1 0 4456 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_358
timestamp 1569139307
transform 1 0 4584 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_359
timestamp 1569139307
transform 1 0 4648 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_360
timestamp 1569139307
transform 1 0 4712 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_361
timestamp 1569139307
transform 1 0 4840 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_362
timestamp 1569139307
transform 1 0 4904 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_363
timestamp 1569139307
transform 1 0 4776 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_364
timestamp 1569139307
transform 1 0 4776 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_365
timestamp 1569139307
transform 1 0 4712 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_366
timestamp 1569139307
transform 1 0 4904 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_367
timestamp 1569139307
transform 1 0 4840 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_368
timestamp 1569139307
transform 1 0 4776 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_369
timestamp 1569139307
transform 1 0 4712 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_370
timestamp 1569139307
transform 1 0 4904 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_371
timestamp 1569139307
transform 1 0 4840 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_372
timestamp 1569139307
transform 1 0 4840 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_373
timestamp 1569139307
transform 1 0 4712 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_374
timestamp 1569139307
transform 1 0 4840 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_375
timestamp 1569139307
transform 1 0 4712 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_376
timestamp 1569139307
transform 1 0 4904 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_377
timestamp 1569139307
transform 1 0 4776 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_378
timestamp 1569139307
transform 1 0 4776 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_379
timestamp 1569139307
transform 1 0 4904 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_380
timestamp 1569139307
transform 1 0 3688 0 1 232
box -8 -8 8 8
use VIA2  VIA2_381
timestamp 1569139307
transform 1 0 3560 0 1 104
box -8 -8 8 8
use VIA2  VIA2_382
timestamp 1569139307
transform 1 0 3624 0 1 40
box -8 -8 8 8
use VIA2  VIA2_383
timestamp 1569139307
transform 1 0 3496 0 1 296
box -8 -8 8 8
use VIA2  VIA2_384
timestamp 1569139307
transform 1 0 3560 0 1 232
box -8 -8 8 8
use VIA2  VIA2_385
timestamp 1569139307
transform 1 0 3560 0 1 40
box -8 -8 8 8
use VIA2  VIA2_386
timestamp 1569139307
transform 1 0 3496 0 1 232
box -8 -8 8 8
use VIA2  VIA2_387
timestamp 1569139307
transform 1 0 3624 0 1 104
box -8 -8 8 8
use VIA2  VIA2_388
timestamp 1569139307
transform 1 0 3688 0 1 104
box -8 -8 8 8
use VIA2  VIA2_389
timestamp 1569139307
transform 1 0 3688 0 1 40
box -8 -8 8 8
use VIA2  VIA2_390
timestamp 1569139307
transform 1 0 3688 0 1 296
box -8 -8 8 8
use VIA2  VIA2_391
timestamp 1569139307
transform 1 0 3496 0 1 104
box -8 -8 8 8
use VIA2  VIA2_392
timestamp 1569139307
transform 1 0 3496 0 1 40
box -8 -8 8 8
use VIA2  VIA2_393
timestamp 1569139307
transform 1 0 3688 0 1 168
box -8 -8 8 8
use VIA2  VIA2_394
timestamp 1569139307
transform 1 0 3560 0 1 168
box -8 -8 8 8
use VIA2  VIA2_395
timestamp 1569139307
transform 1 0 3624 0 1 232
box -8 -8 8 8
use VIA2  VIA2_396
timestamp 1569139307
transform 1 0 3624 0 1 296
box -8 -8 8 8
use VIA2  VIA2_397
timestamp 1569139307
transform 1 0 3496 0 1 168
box -8 -8 8 8
use VIA2  VIA2_398
timestamp 1569139307
transform 1 0 3624 0 1 168
box -8 -8 8 8
use VIA2  VIA2_399
timestamp 1569139307
transform 1 0 3560 0 1 296
box -8 -8 8 8
use VIA2  VIA2_400
timestamp 1569139307
transform 1 0 3368 0 1 104
box -8 -8 8 8
use VIA2  VIA2_401
timestamp 1569139307
transform 1 0 3240 0 1 168
box -8 -8 8 8
use VIA2  VIA2_402
timestamp 1569139307
transform 1 0 3176 0 1 296
box -8 -8 8 8
use VIA2  VIA2_403
timestamp 1569139307
transform 1 0 3368 0 1 232
box -8 -8 8 8
use VIA2  VIA2_404
timestamp 1569139307
transform 1 0 3304 0 1 104
box -8 -8 8 8
use VIA2  VIA2_405
timestamp 1569139307
transform 1 0 3240 0 1 296
box -8 -8 8 8
use VIA2  VIA2_406
timestamp 1569139307
transform 1 0 3304 0 1 168
box -8 -8 8 8
use VIA2  VIA2_407
timestamp 1569139307
transform 1 0 3368 0 1 168
box -8 -8 8 8
use VIA2  VIA2_408
timestamp 1569139307
transform 1 0 3176 0 1 232
box -8 -8 8 8
use VIA2  VIA2_409
timestamp 1569139307
transform 1 0 3240 0 1 40
box -8 -8 8 8
use VIA2  VIA2_410
timestamp 1569139307
transform 1 0 3176 0 1 40
box -8 -8 8 8
use VIA2  VIA2_411
timestamp 1569139307
transform 1 0 3304 0 1 232
box -8 -8 8 8
use VIA2  VIA2_412
timestamp 1569139307
transform 1 0 3176 0 1 168
box -8 -8 8 8
use VIA2  VIA2_413
timestamp 1569139307
transform 1 0 3368 0 1 40
box -8 -8 8 8
use VIA2  VIA2_414
timestamp 1569139307
transform 1 0 3304 0 1 296
box -8 -8 8 8
use VIA2  VIA2_415
timestamp 1569139307
transform 1 0 3304 0 1 40
box -8 -8 8 8
use VIA2  VIA2_416
timestamp 1569139307
transform 1 0 3176 0 1 104
box -8 -8 8 8
use VIA2  VIA2_417
timestamp 1569139307
transform 1 0 3240 0 1 104
box -8 -8 8 8
use VIA2  VIA2_418
timestamp 1569139307
transform 1 0 3368 0 1 296
box -8 -8 8 8
use VIA2  VIA2_419
timestamp 1569139307
transform 1 0 3240 0 1 232
box -8 -8 8 8
use VIA2  VIA2_420
timestamp 1569139307
transform 1 0 3240 0 1 424
box -8 -8 8 8
use VIA2  VIA2_421
timestamp 1569139307
transform 1 0 3240 0 1 488
box -8 -8 8 8
use VIA2  VIA2_422
timestamp 1569139307
transform 1 0 3176 0 1 360
box -8 -8 8 8
use VIA2  VIA2_423
timestamp 1569139307
transform 1 0 3176 0 1 424
box -8 -8 8 8
use VIA2  VIA2_424
timestamp 1569139307
transform 1 0 3368 0 1 360
box -8 -8 8 8
use VIA2  VIA2_425
timestamp 1569139307
transform 1 0 3176 0 1 488
box -8 -8 8 8
use VIA2  VIA2_426
timestamp 1569139307
transform 1 0 3240 0 1 552
box -8 -8 8 8
use VIA2  VIA2_427
timestamp 1569139307
transform 1 0 3176 0 1 552
box -8 -8 8 8
use VIA2  VIA2_428
timestamp 1569139307
transform 1 0 3176 0 1 616
box -8 -8 8 8
use VIA2  VIA2_429
timestamp 1569139307
transform 1 0 3368 0 1 616
box -8 -8 8 8
use VIA2  VIA2_430
timestamp 1569139307
transform 1 0 3240 0 1 616
box -8 -8 8 8
use VIA2  VIA2_431
timestamp 1569139307
transform 1 0 3368 0 1 424
box -8 -8 8 8
use VIA2  VIA2_432
timestamp 1569139307
transform 1 0 3368 0 1 488
box -8 -8 8 8
use VIA2  VIA2_433
timestamp 1569139307
transform 1 0 3368 0 1 552
box -8 -8 8 8
use VIA2  VIA2_434
timestamp 1569139307
transform 1 0 3304 0 1 424
box -8 -8 8 8
use VIA2  VIA2_435
timestamp 1569139307
transform 1 0 3304 0 1 616
box -8 -8 8 8
use VIA2  VIA2_436
timestamp 1569139307
transform 1 0 3304 0 1 488
box -8 -8 8 8
use VIA2  VIA2_437
timestamp 1569139307
transform 1 0 3240 0 1 360
box -8 -8 8 8
use VIA2  VIA2_438
timestamp 1569139307
transform 1 0 3304 0 1 360
box -8 -8 8 8
use VIA2  VIA2_439
timestamp 1569139307
transform 1 0 3304 0 1 552
box -8 -8 8 8
use VIA2  VIA2_440
timestamp 1569139307
transform 1 0 3560 0 1 552
box -8 -8 8 8
use VIA2  VIA2_441
timestamp 1569139307
transform 1 0 3624 0 1 360
box -8 -8 8 8
use VIA2  VIA2_442
timestamp 1569139307
transform 1 0 3496 0 1 552
box -8 -8 8 8
use VIA2  VIA2_443
timestamp 1569139307
transform 1 0 3560 0 1 616
box -8 -8 8 8
use VIA2  VIA2_444
timestamp 1569139307
transform 1 0 3688 0 1 360
box -8 -8 8 8
use VIA2  VIA2_445
timestamp 1569139307
transform 1 0 3688 0 1 424
box -8 -8 8 8
use VIA2  VIA2_446
timestamp 1569139307
transform 1 0 3624 0 1 424
box -8 -8 8 8
use VIA2  VIA2_447
timestamp 1569139307
transform 1 0 3560 0 1 360
box -8 -8 8 8
use VIA2  VIA2_448
timestamp 1569139307
transform 1 0 3688 0 1 488
box -8 -8 8 8
use VIA2  VIA2_449
timestamp 1569139307
transform 1 0 3560 0 1 424
box -8 -8 8 8
use VIA2  VIA2_450
timestamp 1569139307
transform 1 0 3624 0 1 488
box -8 -8 8 8
use VIA2  VIA2_451
timestamp 1569139307
transform 1 0 3688 0 1 552
box -8 -8 8 8
use VIA2  VIA2_452
timestamp 1569139307
transform 1 0 3688 0 1 616
box -8 -8 8 8
use VIA2  VIA2_453
timestamp 1569139307
transform 1 0 3496 0 1 424
box -8 -8 8 8
use VIA2  VIA2_454
timestamp 1569139307
transform 1 0 3560 0 1 488
box -8 -8 8 8
use VIA2  VIA2_455
timestamp 1569139307
transform 1 0 3624 0 1 552
box -8 -8 8 8
use VIA2  VIA2_456
timestamp 1569139307
transform 1 0 3496 0 1 488
box -8 -8 8 8
use VIA2  VIA2_457
timestamp 1569139307
transform 1 0 3496 0 1 616
box -8 -8 8 8
use VIA2  VIA2_458
timestamp 1569139307
transform 1 0 3624 0 1 616
box -8 -8 8 8
use VIA2  VIA2_459
timestamp 1569139307
transform 1 0 3496 0 1 360
box -8 -8 8 8
use VIA2  VIA2_460
timestamp 1569139307
transform 1 0 3432 0 1 360
box -8 -8 8 8
use VIA2  VIA2_461
timestamp 1569139307
transform 1 0 3432 0 1 424
box -8 -8 8 8
use VIA2  VIA2_462
timestamp 1569139307
transform 1 0 3432 0 1 488
box -8 -8 8 8
use VIA2  VIA2_463
timestamp 1569139307
transform 1 0 3432 0 1 40
box -8 -8 8 8
use VIA2  VIA2_464
timestamp 1569139307
transform 1 0 3432 0 1 552
box -8 -8 8 8
use VIA2  VIA2_465
timestamp 1569139307
transform 1 0 3432 0 1 104
box -8 -8 8 8
use VIA2  VIA2_466
timestamp 1569139307
transform 1 0 3432 0 1 296
box -8 -8 8 8
use VIA2  VIA2_467
timestamp 1569139307
transform 1 0 3432 0 1 616
box -8 -8 8 8
use VIA2  VIA2_468
timestamp 1569139307
transform 1 0 3432 0 1 168
box -8 -8 8 8
use VIA2  VIA2_469
timestamp 1569139307
transform 1 0 3432 0 1 232
box -8 -8 8 8
use VIA2  VIA2_470
timestamp 1569139307
transform 1 0 3048 0 1 104
box -8 -8 8 8
use VIA2  VIA2_471
timestamp 1569139307
transform 1 0 2920 0 1 40
box -8 -8 8 8
use VIA2  VIA2_472
timestamp 1569139307
transform 1 0 3048 0 1 168
box -8 -8 8 8
use VIA2  VIA2_473
timestamp 1569139307
transform 1 0 3048 0 1 40
box -8 -8 8 8
use VIA2  VIA2_474
timestamp 1569139307
transform 1 0 2920 0 1 104
box -8 -8 8 8
use VIA2  VIA2_475
timestamp 1569139307
transform 1 0 2984 0 1 40
box -8 -8 8 8
use VIA2  VIA2_476
timestamp 1569139307
transform 1 0 2984 0 1 104
box -8 -8 8 8
use VIA2  VIA2_477
timestamp 1569139307
transform 1 0 2920 0 1 296
box -8 -8 8 8
use VIA2  VIA2_478
timestamp 1569139307
transform 1 0 2984 0 1 296
box -8 -8 8 8
use VIA2  VIA2_479
timestamp 1569139307
transform 1 0 2920 0 1 168
box -8 -8 8 8
use VIA2  VIA2_480
timestamp 1569139307
transform 1 0 2856 0 1 104
box -8 -8 8 8
use VIA2  VIA2_481
timestamp 1569139307
transform 1 0 3048 0 1 296
box -8 -8 8 8
use VIA2  VIA2_482
timestamp 1569139307
transform 1 0 3112 0 1 296
box -8 -8 8 8
use VIA2  VIA2_483
timestamp 1569139307
transform 1 0 2856 0 1 168
box -8 -8 8 8
use VIA2  VIA2_484
timestamp 1569139307
transform 1 0 3048 0 1 232
box -8 -8 8 8
use VIA2  VIA2_485
timestamp 1569139307
transform 1 0 3112 0 1 232
box -8 -8 8 8
use VIA2  VIA2_486
timestamp 1569139307
transform 1 0 2920 0 1 232
box -8 -8 8 8
use VIA2  VIA2_487
timestamp 1569139307
transform 1 0 3112 0 1 168
box -8 -8 8 8
use VIA2  VIA2_488
timestamp 1569139307
transform 1 0 3112 0 1 40
box -8 -8 8 8
use VIA2  VIA2_489
timestamp 1569139307
transform 1 0 2856 0 1 40
box -8 -8 8 8
use VIA2  VIA2_490
timestamp 1569139307
transform 1 0 2984 0 1 168
box -8 -8 8 8
use VIA2  VIA2_491
timestamp 1569139307
transform 1 0 2856 0 1 232
box -8 -8 8 8
use VIA2  VIA2_492
timestamp 1569139307
transform 1 0 3112 0 1 104
box -8 -8 8 8
use VIA2  VIA2_493
timestamp 1569139307
transform 1 0 2984 0 1 232
box -8 -8 8 8
use VIA2  VIA2_494
timestamp 1569139307
transform 1 0 2856 0 1 296
box -8 -8 8 8
use VIA2  VIA2_495
timestamp 1569139307
transform 1 0 2792 0 1 40
box -8 -8 8 8
use VIA2  VIA2_496
timestamp 1569139307
transform 1 0 2664 0 1 104
box -8 -8 8 8
use VIA2  VIA2_497
timestamp 1569139307
transform 1 0 2728 0 1 296
box -8 -8 8 8
use VIA2  VIA2_498
timestamp 1569139307
transform 1 0 2792 0 1 104
box -8 -8 8 8
use VIA2  VIA2_499
timestamp 1569139307
transform 1 0 2728 0 1 40
box -8 -8 8 8
use VIA2  VIA2_500
timestamp 1569139307
transform 1 0 2664 0 1 168
box -8 -8 8 8
use VIA2  VIA2_501
timestamp 1569139307
transform 1 0 2536 0 1 40
box -8 -8 8 8
use VIA2  VIA2_502
timestamp 1569139307
transform 1 0 2536 0 1 168
box -8 -8 8 8
use VIA2  VIA2_503
timestamp 1569139307
transform 1 0 2664 0 1 40
box -8 -8 8 8
use VIA2  VIA2_504
timestamp 1569139307
transform 1 0 2664 0 1 232
box -8 -8 8 8
use VIA2  VIA2_505
timestamp 1569139307
transform 1 0 2536 0 1 232
box -8 -8 8 8
use VIA2  VIA2_506
timestamp 1569139307
transform 1 0 2792 0 1 168
box -8 -8 8 8
use VIA2  VIA2_507
timestamp 1569139307
transform 1 0 2728 0 1 104
box -8 -8 8 8
use VIA2  VIA2_508
timestamp 1569139307
transform 1 0 2600 0 1 104
box -8 -8 8 8
use VIA2  VIA2_509
timestamp 1569139307
transform 1 0 2664 0 1 296
box -8 -8 8 8
use VIA2  VIA2_510
timestamp 1569139307
transform 1 0 2792 0 1 232
box -8 -8 8 8
use VIA2  VIA2_511
timestamp 1569139307
transform 1 0 2728 0 1 168
box -8 -8 8 8
use VIA2  VIA2_512
timestamp 1569139307
transform 1 0 2600 0 1 40
box -8 -8 8 8
use VIA2  VIA2_513
timestamp 1569139307
transform 1 0 2600 0 1 296
box -8 -8 8 8
use VIA2  VIA2_514
timestamp 1569139307
transform 1 0 2536 0 1 104
box -8 -8 8 8
use VIA2  VIA2_515
timestamp 1569139307
transform 1 0 2600 0 1 232
box -8 -8 8 8
use VIA2  VIA2_516
timestamp 1569139307
transform 1 0 2600 0 1 168
box -8 -8 8 8
use VIA2  VIA2_517
timestamp 1569139307
transform 1 0 2728 0 1 232
box -8 -8 8 8
use VIA2  VIA2_518
timestamp 1569139307
transform 1 0 2536 0 1 296
box -8 -8 8 8
use VIA2  VIA2_519
timestamp 1569139307
transform 1 0 2792 0 1 296
box -8 -8 8 8
use VIA2  VIA2_520
timestamp 1569139307
transform 1 0 2728 0 1 424
box -8 -8 8 8
use VIA2  VIA2_521
timestamp 1569139307
transform 1 0 2792 0 1 360
box -8 -8 8 8
use VIA2  VIA2_522
timestamp 1569139307
transform 1 0 2728 0 1 488
box -8 -8 8 8
use VIA2  VIA2_523
timestamp 1569139307
transform 1 0 2792 0 1 424
box -8 -8 8 8
use VIA2  VIA2_524
timestamp 1569139307
transform 1 0 2728 0 1 552
box -8 -8 8 8
use VIA2  VIA2_525
timestamp 1569139307
transform 1 0 2792 0 1 488
box -8 -8 8 8
use VIA2  VIA2_526
timestamp 1569139307
transform 1 0 2664 0 1 360
box -8 -8 8 8
use VIA2  VIA2_527
timestamp 1569139307
transform 1 0 2664 0 1 424
box -8 -8 8 8
use VIA2  VIA2_528
timestamp 1569139307
transform 1 0 2792 0 1 552
box -8 -8 8 8
use VIA2  VIA2_529
timestamp 1569139307
transform 1 0 2792 0 1 616
box -8 -8 8 8
use VIA2  VIA2_530
timestamp 1569139307
transform 1 0 2664 0 1 488
box -8 -8 8 8
use VIA2  VIA2_531
timestamp 1569139307
transform 1 0 2536 0 1 424
box -8 -8 8 8
use VIA2  VIA2_532
timestamp 1569139307
transform 1 0 2664 0 1 552
box -8 -8 8 8
use VIA2  VIA2_533
timestamp 1569139307
transform 1 0 2664 0 1 616
box -8 -8 8 8
use VIA2  VIA2_534
timestamp 1569139307
transform 1 0 2536 0 1 488
box -8 -8 8 8
use VIA2  VIA2_535
timestamp 1569139307
transform 1 0 2536 0 1 552
box -8 -8 8 8
use VIA2  VIA2_536
timestamp 1569139307
transform 1 0 2536 0 1 616
box -8 -8 8 8
use VIA2  VIA2_537
timestamp 1569139307
transform 1 0 2600 0 1 424
box -8 -8 8 8
use VIA2  VIA2_538
timestamp 1569139307
transform 1 0 2728 0 1 616
box -8 -8 8 8
use VIA2  VIA2_539
timestamp 1569139307
transform 1 0 2600 0 1 488
box -8 -8 8 8
use VIA2  VIA2_540
timestamp 1569139307
transform 1 0 2728 0 1 360
box -8 -8 8 8
use VIA2  VIA2_541
timestamp 1569139307
transform 1 0 2600 0 1 552
box -8 -8 8 8
use VIA2  VIA2_542
timestamp 1569139307
transform 1 0 2600 0 1 616
box -8 -8 8 8
use VIA2  VIA2_543
timestamp 1569139307
transform 1 0 2600 0 1 360
box -8 -8 8 8
use VIA2  VIA2_544
timestamp 1569139307
transform 1 0 2536 0 1 360
box -8 -8 8 8
use VIA2  VIA2_545
timestamp 1569139307
transform 1 0 2856 0 1 360
box -8 -8 8 8
use VIA2  VIA2_546
timestamp 1569139307
transform 1 0 3048 0 1 360
box -8 -8 8 8
use VIA2  VIA2_547
timestamp 1569139307
transform 1 0 3048 0 1 424
box -8 -8 8 8
use VIA2  VIA2_548
timestamp 1569139307
transform 1 0 3048 0 1 488
box -8 -8 8 8
use VIA2  VIA2_549
timestamp 1569139307
transform 1 0 3048 0 1 552
box -8 -8 8 8
use VIA2  VIA2_550
timestamp 1569139307
transform 1 0 3048 0 1 616
box -8 -8 8 8
use VIA2  VIA2_551
timestamp 1569139307
transform 1 0 2856 0 1 424
box -8 -8 8 8
use VIA2  VIA2_552
timestamp 1569139307
transform 1 0 2984 0 1 360
box -8 -8 8 8
use VIA2  VIA2_553
timestamp 1569139307
transform 1 0 2856 0 1 552
box -8 -8 8 8
use VIA2  VIA2_554
timestamp 1569139307
transform 1 0 2856 0 1 616
box -8 -8 8 8
use VIA2  VIA2_555
timestamp 1569139307
transform 1 0 3112 0 1 360
box -8 -8 8 8
use VIA2  VIA2_556
timestamp 1569139307
transform 1 0 3112 0 1 424
box -8 -8 8 8
use VIA2  VIA2_557
timestamp 1569139307
transform 1 0 2920 0 1 360
box -8 -8 8 8
use VIA2  VIA2_558
timestamp 1569139307
transform 1 0 3112 0 1 488
box -8 -8 8 8
use VIA2  VIA2_559
timestamp 1569139307
transform 1 0 3112 0 1 552
box -8 -8 8 8
use VIA2  VIA2_560
timestamp 1569139307
transform 1 0 2984 0 1 424
box -8 -8 8 8
use VIA2  VIA2_561
timestamp 1569139307
transform 1 0 3112 0 1 616
box -8 -8 8 8
use VIA2  VIA2_562
timestamp 1569139307
transform 1 0 2920 0 1 424
box -8 -8 8 8
use VIA2  VIA2_563
timestamp 1569139307
transform 1 0 2984 0 1 488
box -8 -8 8 8
use VIA2  VIA2_564
timestamp 1569139307
transform 1 0 2856 0 1 488
box -8 -8 8 8
use VIA2  VIA2_565
timestamp 1569139307
transform 1 0 2920 0 1 488
box -8 -8 8 8
use VIA2  VIA2_566
timestamp 1569139307
transform 1 0 2984 0 1 552
box -8 -8 8 8
use VIA2  VIA2_567
timestamp 1569139307
transform 1 0 2920 0 1 552
box -8 -8 8 8
use VIA2  VIA2_568
timestamp 1569139307
transform 1 0 2920 0 1 616
box -8 -8 8 8
use VIA2  VIA2_569
timestamp 1569139307
transform 1 0 2984 0 1 616
box -8 -8 8 8
use VIA2  VIA2_570
timestamp 1569139307
transform 1 0 3048 0 1 744
box -8 -8 8 8
use VIA2  VIA2_571
timestamp 1569139307
transform 1 0 2920 0 1 936
box -8 -8 8 8
use VIA2  VIA2_572
timestamp 1569139307
transform 1 0 3112 0 1 680
box -8 -8 8 8
use VIA2  VIA2_573
timestamp 1569139307
transform 1 0 2984 0 1 872
box -8 -8 8 8
use VIA2  VIA2_574
timestamp 1569139307
transform 1 0 3048 0 1 808
box -8 -8 8 8
use VIA2  VIA2_575
timestamp 1569139307
transform 1 0 3112 0 1 744
box -8 -8 8 8
use VIA2  VIA2_576
timestamp 1569139307
transform 1 0 2856 0 1 744
box -8 -8 8 8
use VIA2  VIA2_577
timestamp 1569139307
transform 1 0 2920 0 1 744
box -8 -8 8 8
use VIA2  VIA2_578
timestamp 1569139307
transform 1 0 2856 0 1 936
box -8 -8 8 8
use VIA2  VIA2_579
timestamp 1569139307
transform 1 0 3112 0 1 808
box -8 -8 8 8
use VIA2  VIA2_580
timestamp 1569139307
transform 1 0 2984 0 1 808
box -8 -8 8 8
use VIA2  VIA2_581
timestamp 1569139307
transform 1 0 3048 0 1 872
box -8 -8 8 8
use VIA2  VIA2_582
timestamp 1569139307
transform 1 0 2984 0 1 744
box -8 -8 8 8
use VIA2  VIA2_583
timestamp 1569139307
transform 1 0 2920 0 1 808
box -8 -8 8 8
use VIA2  VIA2_584
timestamp 1569139307
transform 1 0 2856 0 1 808
box -8 -8 8 8
use VIA2  VIA2_585
timestamp 1569139307
transform 1 0 3112 0 1 872
box -8 -8 8 8
use VIA2  VIA2_586
timestamp 1569139307
transform 1 0 2856 0 1 680
box -8 -8 8 8
use VIA2  VIA2_587
timestamp 1569139307
transform 1 0 2920 0 1 872
box -8 -8 8 8
use VIA2  VIA2_588
timestamp 1569139307
transform 1 0 3048 0 1 936
box -8 -8 8 8
use VIA2  VIA2_589
timestamp 1569139307
transform 1 0 2920 0 1 680
box -8 -8 8 8
use VIA2  VIA2_590
timestamp 1569139307
transform 1 0 3112 0 1 936
box -8 -8 8 8
use VIA2  VIA2_591
timestamp 1569139307
transform 1 0 2984 0 1 936
box -8 -8 8 8
use VIA2  VIA2_592
timestamp 1569139307
transform 1 0 3048 0 1 680
box -8 -8 8 8
use VIA2  VIA2_593
timestamp 1569139307
transform 1 0 2856 0 1 872
box -8 -8 8 8
use VIA2  VIA2_594
timestamp 1569139307
transform 1 0 2984 0 1 680
box -8 -8 8 8
use VIA2  VIA2_595
timestamp 1569139307
transform 1 0 2728 0 1 936
box -8 -8 8 8
use VIA2  VIA2_596
timestamp 1569139307
transform 1 0 2664 0 1 808
box -8 -8 8 8
use VIA2  VIA2_597
timestamp 1569139307
transform 1 0 2536 0 1 936
box -8 -8 8 8
use VIA2  VIA2_598
timestamp 1569139307
transform 1 0 2728 0 1 808
box -8 -8 8 8
use VIA2  VIA2_599
timestamp 1569139307
transform 1 0 2728 0 1 744
box -8 -8 8 8
use VIA2  VIA2_600
timestamp 1569139307
transform 1 0 2600 0 1 680
box -8 -8 8 8
use VIA2  VIA2_601
timestamp 1569139307
transform 1 0 2792 0 1 680
box -8 -8 8 8
use VIA2  VIA2_602
timestamp 1569139307
transform 1 0 2600 0 1 744
box -8 -8 8 8
use VIA2  VIA2_603
timestamp 1569139307
transform 1 0 2792 0 1 872
box -8 -8 8 8
use VIA2  VIA2_604
timestamp 1569139307
transform 1 0 2600 0 1 808
box -8 -8 8 8
use VIA2  VIA2_605
timestamp 1569139307
transform 1 0 2664 0 1 680
box -8 -8 8 8
use VIA2  VIA2_606
timestamp 1569139307
transform 1 0 2600 0 1 872
box -8 -8 8 8
use VIA2  VIA2_607
timestamp 1569139307
transform 1 0 2728 0 1 680
box -8 -8 8 8
use VIA2  VIA2_608
timestamp 1569139307
transform 1 0 2792 0 1 808
box -8 -8 8 8
use VIA2  VIA2_609
timestamp 1569139307
transform 1 0 2728 0 1 872
box -8 -8 8 8
use VIA2  VIA2_610
timestamp 1569139307
transform 1 0 2600 0 1 936
box -8 -8 8 8
use VIA2  VIA2_611
timestamp 1569139307
transform 1 0 2664 0 1 936
box -8 -8 8 8
use VIA2  VIA2_612
timestamp 1569139307
transform 1 0 2792 0 1 744
box -8 -8 8 8
use VIA2  VIA2_613
timestamp 1569139307
transform 1 0 2536 0 1 680
box -8 -8 8 8
use VIA2  VIA2_614
timestamp 1569139307
transform 1 0 2664 0 1 744
box -8 -8 8 8
use VIA2  VIA2_615
timestamp 1569139307
transform 1 0 2536 0 1 744
box -8 -8 8 8
use VIA2  VIA2_616
timestamp 1569139307
transform 1 0 2664 0 1 872
box -8 -8 8 8
use VIA2  VIA2_617
timestamp 1569139307
transform 1 0 2536 0 1 808
box -8 -8 8 8
use VIA2  VIA2_618
timestamp 1569139307
transform 1 0 2792 0 1 936
box -8 -8 8 8
use VIA2  VIA2_619
timestamp 1569139307
transform 1 0 2536 0 1 872
box -8 -8 8 8
use VIA2  VIA2_620
timestamp 1569139307
transform 1 0 2792 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_621
timestamp 1569139307
transform 1 0 2664 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_622
timestamp 1569139307
transform 1 0 2536 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_623
timestamp 1569139307
transform 1 0 2664 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_624
timestamp 1569139307
transform 1 0 2792 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_625
timestamp 1569139307
transform 1 0 2536 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_626
timestamp 1569139307
transform 1 0 2600 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_627
timestamp 1569139307
transform 1 0 2792 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_628
timestamp 1569139307
transform 1 0 2792 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_629
timestamp 1569139307
transform 1 0 2536 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_630
timestamp 1569139307
transform 1 0 2728 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_631
timestamp 1569139307
transform 1 0 2600 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_632
timestamp 1569139307
transform 1 0 2600 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_633
timestamp 1569139307
transform 1 0 2664 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_634
timestamp 1569139307
transform 1 0 2536 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_635
timestamp 1569139307
transform 1 0 2728 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_636
timestamp 1569139307
transform 1 0 2664 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_637
timestamp 1569139307
transform 1 0 2728 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_638
timestamp 1569139307
transform 1 0 2792 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_639
timestamp 1569139307
transform 1 0 2664 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_640
timestamp 1569139307
transform 1 0 2728 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_641
timestamp 1569139307
transform 1 0 2600 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_642
timestamp 1569139307
transform 1 0 2600 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_643
timestamp 1569139307
transform 1 0 2536 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_644
timestamp 1569139307
transform 1 0 2728 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_645
timestamp 1569139307
transform 1 0 2920 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_646
timestamp 1569139307
transform 1 0 2856 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_647
timestamp 1569139307
transform 1 0 2920 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_648
timestamp 1569139307
transform 1 0 2920 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_649
timestamp 1569139307
transform 1 0 2856 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_650
timestamp 1569139307
transform 1 0 3112 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_651
timestamp 1569139307
transform 1 0 3112 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_652
timestamp 1569139307
transform 1 0 3048 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_653
timestamp 1569139307
transform 1 0 2856 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_654
timestamp 1569139307
transform 1 0 3112 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_655
timestamp 1569139307
transform 1 0 2856 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_656
timestamp 1569139307
transform 1 0 3112 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_657
timestamp 1569139307
transform 1 0 2984 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_658
timestamp 1569139307
transform 1 0 3048 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_659
timestamp 1569139307
transform 1 0 2856 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_660
timestamp 1569139307
transform 1 0 2984 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_661
timestamp 1569139307
transform 1 0 2984 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_662
timestamp 1569139307
transform 1 0 2984 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_663
timestamp 1569139307
transform 1 0 2920 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_664
timestamp 1569139307
transform 1 0 2984 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_665
timestamp 1569139307
transform 1 0 2920 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_666
timestamp 1569139307
transform 1 0 3048 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_667
timestamp 1569139307
transform 1 0 3112 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_668
timestamp 1569139307
transform 1 0 3048 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_669
timestamp 1569139307
transform 1 0 3048 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_670
timestamp 1569139307
transform 1 0 3496 0 1 680
box -8 -8 8 8
use VIA2  VIA2_671
timestamp 1569139307
transform 1 0 3624 0 1 680
box -8 -8 8 8
use VIA2  VIA2_672
timestamp 1569139307
transform 1 0 3560 0 1 872
box -8 -8 8 8
use VIA2  VIA2_673
timestamp 1569139307
transform 1 0 3496 0 1 744
box -8 -8 8 8
use VIA2  VIA2_674
timestamp 1569139307
transform 1 0 3624 0 1 808
box -8 -8 8 8
use VIA2  VIA2_675
timestamp 1569139307
transform 1 0 3560 0 1 936
box -8 -8 8 8
use VIA2  VIA2_676
timestamp 1569139307
transform 1 0 3496 0 1 808
box -8 -8 8 8
use VIA2  VIA2_677
timestamp 1569139307
transform 1 0 3560 0 1 680
box -8 -8 8 8
use VIA2  VIA2_678
timestamp 1569139307
transform 1 0 3688 0 1 680
box -8 -8 8 8
use VIA2  VIA2_679
timestamp 1569139307
transform 1 0 3496 0 1 872
box -8 -8 8 8
use VIA2  VIA2_680
timestamp 1569139307
transform 1 0 3688 0 1 744
box -8 -8 8 8
use VIA2  VIA2_681
timestamp 1569139307
transform 1 0 3624 0 1 744
box -8 -8 8 8
use VIA2  VIA2_682
timestamp 1569139307
transform 1 0 3688 0 1 808
box -8 -8 8 8
use VIA2  VIA2_683
timestamp 1569139307
transform 1 0 3496 0 1 936
box -8 -8 8 8
use VIA2  VIA2_684
timestamp 1569139307
transform 1 0 3560 0 1 744
box -8 -8 8 8
use VIA2  VIA2_685
timestamp 1569139307
transform 1 0 3688 0 1 872
box -8 -8 8 8
use VIA2  VIA2_686
timestamp 1569139307
transform 1 0 3560 0 1 808
box -8 -8 8 8
use VIA2  VIA2_687
timestamp 1569139307
transform 1 0 3688 0 1 936
box -8 -8 8 8
use VIA2  VIA2_688
timestamp 1569139307
transform 1 0 3624 0 1 936
box -8 -8 8 8
use VIA2  VIA2_689
timestamp 1569139307
transform 1 0 3624 0 1 872
box -8 -8 8 8
use VIA2  VIA2_690
timestamp 1569139307
transform 1 0 3240 0 1 872
box -8 -8 8 8
use VIA2  VIA2_691
timestamp 1569139307
transform 1 0 3240 0 1 936
box -8 -8 8 8
use VIA2  VIA2_692
timestamp 1569139307
transform 1 0 3368 0 1 808
box -8 -8 8 8
use VIA2  VIA2_693
timestamp 1569139307
transform 1 0 3304 0 1 680
box -8 -8 8 8
use VIA2  VIA2_694
timestamp 1569139307
transform 1 0 3304 0 1 744
box -8 -8 8 8
use VIA2  VIA2_695
timestamp 1569139307
transform 1 0 3304 0 1 808
box -8 -8 8 8
use VIA2  VIA2_696
timestamp 1569139307
transform 1 0 3304 0 1 872
box -8 -8 8 8
use VIA2  VIA2_697
timestamp 1569139307
transform 1 0 3304 0 1 936
box -8 -8 8 8
use VIA2  VIA2_698
timestamp 1569139307
transform 1 0 3368 0 1 872
box -8 -8 8 8
use VIA2  VIA2_699
timestamp 1569139307
transform 1 0 3368 0 1 744
box -8 -8 8 8
use VIA2  VIA2_700
timestamp 1569139307
transform 1 0 3368 0 1 936
box -8 -8 8 8
use VIA2  VIA2_701
timestamp 1569139307
transform 1 0 3176 0 1 680
box -8 -8 8 8
use VIA2  VIA2_702
timestamp 1569139307
transform 1 0 3176 0 1 744
box -8 -8 8 8
use VIA2  VIA2_703
timestamp 1569139307
transform 1 0 3176 0 1 808
box -8 -8 8 8
use VIA2  VIA2_704
timestamp 1569139307
transform 1 0 3176 0 1 872
box -8 -8 8 8
use VIA2  VIA2_705
timestamp 1569139307
transform 1 0 3176 0 1 936
box -8 -8 8 8
use VIA2  VIA2_706
timestamp 1569139307
transform 1 0 3368 0 1 680
box -8 -8 8 8
use VIA2  VIA2_707
timestamp 1569139307
transform 1 0 3240 0 1 680
box -8 -8 8 8
use VIA2  VIA2_708
timestamp 1569139307
transform 1 0 3240 0 1 744
box -8 -8 8 8
use VIA2  VIA2_709
timestamp 1569139307
transform 1 0 3240 0 1 808
box -8 -8 8 8
use VIA2  VIA2_710
timestamp 1569139307
transform 1 0 3368 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_711
timestamp 1569139307
transform 1 0 3176 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_712
timestamp 1569139307
transform 1 0 3368 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_713
timestamp 1569139307
transform 1 0 3176 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_714
timestamp 1569139307
transform 1 0 3368 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_715
timestamp 1569139307
transform 1 0 3368 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_716
timestamp 1569139307
transform 1 0 3240 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_717
timestamp 1569139307
transform 1 0 3304 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_718
timestamp 1569139307
transform 1 0 3176 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_719
timestamp 1569139307
transform 1 0 3240 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_720
timestamp 1569139307
transform 1 0 3368 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_721
timestamp 1569139307
transform 1 0 3240 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_722
timestamp 1569139307
transform 1 0 3304 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_723
timestamp 1569139307
transform 1 0 3176 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_724
timestamp 1569139307
transform 1 0 3304 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_725
timestamp 1569139307
transform 1 0 3240 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_726
timestamp 1569139307
transform 1 0 3304 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_727
timestamp 1569139307
transform 1 0 3240 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_728
timestamp 1569139307
transform 1 0 3304 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_729
timestamp 1569139307
transform 1 0 3176 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_730
timestamp 1569139307
transform 1 0 3624 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_731
timestamp 1569139307
transform 1 0 3624 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_732
timestamp 1569139307
transform 1 0 3496 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_733
timestamp 1569139307
transform 1 0 3624 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_734
timestamp 1569139307
transform 1 0 3560 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_735
timestamp 1569139307
transform 1 0 3688 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_736
timestamp 1569139307
transform 1 0 3560 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_737
timestamp 1569139307
transform 1 0 3560 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_738
timestamp 1569139307
transform 1 0 3688 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_739
timestamp 1569139307
transform 1 0 3624 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_740
timestamp 1569139307
transform 1 0 3688 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_741
timestamp 1569139307
transform 1 0 3624 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_742
timestamp 1569139307
transform 1 0 3496 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_743
timestamp 1569139307
transform 1 0 3560 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_744
timestamp 1569139307
transform 1 0 3496 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_745
timestamp 1569139307
transform 1 0 3496 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_746
timestamp 1569139307
transform 1 0 3688 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_747
timestamp 1569139307
transform 1 0 3496 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_748
timestamp 1569139307
transform 1 0 3560 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_749
timestamp 1569139307
transform 1 0 3688 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_750
timestamp 1569139307
transform 1 0 3432 0 1 680
box -8 -8 8 8
use VIA2  VIA2_751
timestamp 1569139307
transform 1 0 3432 0 1 744
box -8 -8 8 8
use VIA2  VIA2_752
timestamp 1569139307
transform 1 0 3432 0 1 808
box -8 -8 8 8
use VIA2  VIA2_753
timestamp 1569139307
transform 1 0 3432 0 1 872
box -8 -8 8 8
use VIA2  VIA2_754
timestamp 1569139307
transform 1 0 3432 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_755
timestamp 1569139307
transform 1 0 3432 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_756
timestamp 1569139307
transform 1 0 3432 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_757
timestamp 1569139307
transform 1 0 3432 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_758
timestamp 1569139307
transform 1 0 3432 0 1 936
box -8 -8 8 8
use VIA2  VIA2_759
timestamp 1569139307
transform 1 0 3432 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_760
timestamp 1569139307
transform 1 0 3688 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_761
timestamp 1569139307
transform 1 0 3368 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_762
timestamp 1569139307
transform 1 0 3624 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_763
timestamp 1569139307
transform 1 0 3496 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_764
timestamp 1569139307
transform 1 0 3432 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_765
timestamp 1569139307
transform 1 0 3304 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_766
timestamp 1569139307
transform 1 0 3176 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_767
timestamp 1569139307
transform 1 0 3688 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_768
timestamp 1569139307
transform 1 0 3432 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_769
timestamp 1569139307
transform 1 0 3432 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_770
timestamp 1569139307
transform 1 0 3624 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_771
timestamp 1569139307
transform 1 0 3176 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_772
timestamp 1569139307
transform 1 0 3240 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_773
timestamp 1569139307
transform 1 0 3240 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_774
timestamp 1569139307
transform 1 0 3176 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_775
timestamp 1569139307
transform 1 0 3560 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_776
timestamp 1569139307
transform 1 0 3496 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_777
timestamp 1569139307
transform 1 0 3432 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_778
timestamp 1569139307
transform 1 0 3560 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_779
timestamp 1569139307
transform 1 0 3624 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_780
timestamp 1569139307
transform 1 0 3624 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_781
timestamp 1569139307
transform 1 0 3240 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_782
timestamp 1569139307
transform 1 0 3176 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_783
timestamp 1569139307
transform 1 0 3688 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_784
timestamp 1569139307
transform 1 0 3304 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_785
timestamp 1569139307
transform 1 0 3240 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_786
timestamp 1569139307
transform 1 0 3304 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_787
timestamp 1569139307
transform 1 0 3688 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_788
timestamp 1569139307
transform 1 0 3496 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_789
timestamp 1569139307
transform 1 0 3304 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_790
timestamp 1569139307
transform 1 0 3368 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_791
timestamp 1569139307
transform 1 0 3496 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_792
timestamp 1569139307
transform 1 0 3368 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_793
timestamp 1569139307
transform 1 0 3560 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_794
timestamp 1569139307
transform 1 0 3560 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_795
timestamp 1569139307
transform 1 0 3368 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_796
timestamp 1569139307
transform 1 0 3112 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_797
timestamp 1569139307
transform 1 0 3048 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_798
timestamp 1569139307
transform 1 0 2920 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_799
timestamp 1569139307
transform 1 0 3112 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_800
timestamp 1569139307
transform 1 0 2984 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_801
timestamp 1569139307
transform 1 0 2984 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_802
timestamp 1569139307
transform 1 0 2920 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_803
timestamp 1569139307
transform 1 0 2856 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_804
timestamp 1569139307
transform 1 0 3048 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_805
timestamp 1569139307
transform 1 0 2920 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_806
timestamp 1569139307
transform 1 0 2984 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_807
timestamp 1569139307
transform 1 0 2920 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_808
timestamp 1569139307
transform 1 0 3112 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_809
timestamp 1569139307
transform 1 0 2856 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_810
timestamp 1569139307
transform 1 0 3112 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_811
timestamp 1569139307
transform 1 0 3048 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_812
timestamp 1569139307
transform 1 0 2984 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_813
timestamp 1569139307
transform 1 0 2856 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_814
timestamp 1569139307
transform 1 0 3048 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_815
timestamp 1569139307
transform 1 0 2856 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_816
timestamp 1569139307
transform 1 0 2664 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_817
timestamp 1569139307
transform 1 0 2600 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_818
timestamp 1569139307
transform 1 0 2792 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_819
timestamp 1569139307
transform 1 0 2664 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_820
timestamp 1569139307
transform 1 0 2728 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_821
timestamp 1569139307
transform 1 0 2536 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_822
timestamp 1569139307
transform 1 0 2728 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_823
timestamp 1569139307
transform 1 0 2728 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_824
timestamp 1569139307
transform 1 0 2664 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_825
timestamp 1569139307
transform 1 0 2600 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_826
timestamp 1569139307
transform 1 0 2792 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_827
timestamp 1569139307
transform 1 0 2536 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_828
timestamp 1569139307
transform 1 0 2728 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_829
timestamp 1569139307
transform 1 0 2792 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_830
timestamp 1569139307
transform 1 0 2792 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_831
timestamp 1569139307
transform 1 0 2600 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_832
timestamp 1569139307
transform 1 0 2536 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_833
timestamp 1569139307
transform 1 0 2664 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_834
timestamp 1569139307
transform 1 0 2600 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_835
timestamp 1569139307
transform 1 0 2536 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_836
timestamp 1569139307
transform 1 0 2664 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_837
timestamp 1569139307
transform 1 0 2600 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_838
timestamp 1569139307
transform 1 0 2536 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_839
timestamp 1569139307
transform 1 0 2728 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_840
timestamp 1569139307
transform 1 0 2536 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_841
timestamp 1569139307
transform 1 0 2600 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_842
timestamp 1569139307
transform 1 0 2600 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_843
timestamp 1569139307
transform 1 0 2600 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_844
timestamp 1569139307
transform 1 0 2792 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_845
timestamp 1569139307
transform 1 0 2664 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_846
timestamp 1569139307
transform 1 0 2664 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_847
timestamp 1569139307
transform 1 0 2536 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_848
timestamp 1569139307
transform 1 0 2536 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_849
timestamp 1569139307
transform 1 0 2728 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_850
timestamp 1569139307
transform 1 0 2664 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_851
timestamp 1569139307
transform 1 0 2536 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_852
timestamp 1569139307
transform 1 0 2600 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_853
timestamp 1569139307
transform 1 0 2728 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_854
timestamp 1569139307
transform 1 0 2792 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_855
timestamp 1569139307
transform 1 0 2856 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_856
timestamp 1569139307
transform 1 0 2536 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_857
timestamp 1569139307
transform 1 0 3688 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_858
timestamp 1569139307
transform 1 0 3624 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_859
timestamp 1569139307
transform 1 0 3688 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_860
timestamp 1569139307
transform 1 0 3688 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_861
timestamp 1569139307
transform 1 0 3240 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_862
timestamp 1569139307
transform 1 0 3432 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_863
timestamp 1569139307
transform 1 0 3432 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_864
timestamp 1569139307
transform 1 0 3432 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_865
timestamp 1569139307
transform 1 0 3496 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_866
timestamp 1569139307
transform 1 0 3496 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_867
timestamp 1569139307
transform 1 0 3496 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_868
timestamp 1569139307
transform 1 0 3304 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_869
timestamp 1569139307
transform 1 0 3304 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_870
timestamp 1569139307
transform 1 0 3560 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_871
timestamp 1569139307
transform 1 0 3560 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_872
timestamp 1569139307
transform 1 0 3560 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_873
timestamp 1569139307
transform 1 0 3368 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_874
timestamp 1569139307
transform 1 0 3368 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_875
timestamp 1569139307
transform 1 0 3624 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_876
timestamp 1569139307
transform 1 0 3368 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_877
timestamp 1569139307
transform 1 0 3624 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_878
timestamp 1569139307
transform 1 0 4648 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_879
timestamp 1569139307
transform 1 0 4712 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_880
timestamp 1569139307
transform 1 0 4392 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_881
timestamp 1569139307
transform 1 0 4904 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_882
timestamp 1569139307
transform 1 0 4712 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_883
timestamp 1569139307
transform 1 0 4584 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_884
timestamp 1569139307
transform 1 0 4456 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_885
timestamp 1569139307
transform 1 0 4584 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_886
timestamp 1569139307
transform 1 0 4712 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_887
timestamp 1569139307
transform 1 0 4456 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_888
timestamp 1569139307
transform 1 0 4840 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_889
timestamp 1569139307
transform 1 0 4776 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_890
timestamp 1569139307
transform 1 0 4648 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_891
timestamp 1569139307
transform 1 0 4840 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_892
timestamp 1569139307
transform 1 0 4776 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_893
timestamp 1569139307
transform 1 0 4456 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_894
timestamp 1569139307
transform 1 0 4584 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_895
timestamp 1569139307
transform 1 0 4520 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_896
timestamp 1569139307
transform 1 0 4840 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_897
timestamp 1569139307
transform 1 0 4776 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_898
timestamp 1569139307
transform 1 0 4776 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_899
timestamp 1569139307
transform 1 0 4520 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_900
timestamp 1569139307
transform 1 0 4392 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_901
timestamp 1569139307
transform 1 0 4904 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_902
timestamp 1569139307
transform 1 0 4520 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_903
timestamp 1569139307
transform 1 0 4520 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_904
timestamp 1569139307
transform 1 0 4648 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_905
timestamp 1569139307
transform 1 0 4648 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_906
timestamp 1569139307
transform 1 0 4712 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_907
timestamp 1569139307
transform 1 0 4584 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_908
timestamp 1569139307
transform 1 0 4456 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_909
timestamp 1569139307
transform 1 0 4392 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_910
timestamp 1569139307
transform 1 0 4904 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_911
timestamp 1569139307
transform 1 0 4392 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_912
timestamp 1569139307
transform 1 0 4904 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_913
timestamp 1569139307
transform 1 0 4840 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_914
timestamp 1569139307
transform 1 0 4072 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_915
timestamp 1569139307
transform 1 0 3944 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_916
timestamp 1569139307
transform 1 0 3880 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_917
timestamp 1569139307
transform 1 0 4136 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_918
timestamp 1569139307
transform 1 0 3880 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_919
timestamp 1569139307
transform 1 0 3944 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_920
timestamp 1569139307
transform 1 0 4200 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_921
timestamp 1569139307
transform 1 0 4200 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_922
timestamp 1569139307
transform 1 0 3880 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_923
timestamp 1569139307
transform 1 0 3944 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_924
timestamp 1569139307
transform 1 0 4200 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_925
timestamp 1569139307
transform 1 0 3944 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_926
timestamp 1569139307
transform 1 0 3752 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_927
timestamp 1569139307
transform 1 0 4136 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_928
timestamp 1569139307
transform 1 0 4200 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_929
timestamp 1569139307
transform 1 0 4264 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_930
timestamp 1569139307
transform 1 0 4008 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_931
timestamp 1569139307
transform 1 0 4008 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_932
timestamp 1569139307
transform 1 0 3752 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_933
timestamp 1569139307
transform 1 0 4264 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_934
timestamp 1569139307
transform 1 0 3880 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_935
timestamp 1569139307
transform 1 0 4008 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_936
timestamp 1569139307
transform 1 0 3816 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_937
timestamp 1569139307
transform 1 0 3752 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_938
timestamp 1569139307
transform 1 0 4264 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_939
timestamp 1569139307
transform 1 0 4328 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_940
timestamp 1569139307
transform 1 0 4264 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_941
timestamp 1569139307
transform 1 0 3752 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_942
timestamp 1569139307
transform 1 0 4072 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_943
timestamp 1569139307
transform 1 0 4136 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_944
timestamp 1569139307
transform 1 0 3816 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_945
timestamp 1569139307
transform 1 0 4328 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_946
timestamp 1569139307
transform 1 0 4072 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_947
timestamp 1569139307
transform 1 0 3816 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_948
timestamp 1569139307
transform 1 0 4328 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_949
timestamp 1569139307
transform 1 0 4072 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_950
timestamp 1569139307
transform 1 0 3816 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_951
timestamp 1569139307
transform 1 0 4328 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_952
timestamp 1569139307
transform 1 0 4008 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_953
timestamp 1569139307
transform 1 0 4136 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_954
timestamp 1569139307
transform 1 0 4072 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_955
timestamp 1569139307
transform 1 0 4072 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_956
timestamp 1569139307
transform 1 0 3752 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_957
timestamp 1569139307
transform 1 0 4072 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_958
timestamp 1569139307
transform 1 0 3880 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_959
timestamp 1569139307
transform 1 0 3816 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_960
timestamp 1569139307
transform 1 0 3880 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_961
timestamp 1569139307
transform 1 0 4136 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_962
timestamp 1569139307
transform 1 0 3880 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_963
timestamp 1569139307
transform 1 0 3752 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_964
timestamp 1569139307
transform 1 0 4136 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_965
timestamp 1569139307
transform 1 0 4136 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_966
timestamp 1569139307
transform 1 0 3944 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_967
timestamp 1569139307
transform 1 0 4328 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_968
timestamp 1569139307
transform 1 0 4200 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_969
timestamp 1569139307
transform 1 0 3944 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_970
timestamp 1569139307
transform 1 0 4200 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_971
timestamp 1569139307
transform 1 0 3944 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_972
timestamp 1569139307
transform 1 0 4328 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_973
timestamp 1569139307
transform 1 0 4200 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_974
timestamp 1569139307
transform 1 0 4328 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_975
timestamp 1569139307
transform 1 0 4264 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_976
timestamp 1569139307
transform 1 0 3816 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_977
timestamp 1569139307
transform 1 0 4264 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_978
timestamp 1569139307
transform 1 0 4264 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_979
timestamp 1569139307
transform 1 0 4008 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_980
timestamp 1569139307
transform 1 0 4008 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_981
timestamp 1569139307
transform 1 0 3816 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_982
timestamp 1569139307
transform 1 0 4008 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_983
timestamp 1569139307
transform 1 0 3752 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_984
timestamp 1569139307
transform 1 0 4520 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_985
timestamp 1569139307
transform 1 0 4520 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_986
timestamp 1569139307
transform 1 0 4520 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_987
timestamp 1569139307
transform 1 0 4584 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_988
timestamp 1569139307
transform 1 0 4584 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_989
timestamp 1569139307
transform 1 0 4584 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_990
timestamp 1569139307
transform 1 0 4456 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_991
timestamp 1569139307
transform 1 0 4648 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_992
timestamp 1569139307
transform 1 0 4648 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_993
timestamp 1569139307
transform 1 0 4648 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_994
timestamp 1569139307
transform 1 0 4712 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_995
timestamp 1569139307
transform 1 0 4712 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_996
timestamp 1569139307
transform 1 0 4712 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_997
timestamp 1569139307
transform 1 0 4776 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_998
timestamp 1569139307
transform 1 0 4776 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_999
timestamp 1569139307
transform 1 0 4776 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1000
timestamp 1569139307
transform 1 0 4840 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1001
timestamp 1569139307
transform 1 0 4840 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1002
timestamp 1569139307
transform 1 0 4840 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1003
timestamp 1569139307
transform 1 0 4904 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1004
timestamp 1569139307
transform 1 0 4904 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1005
timestamp 1569139307
transform 1 0 4904 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1006
timestamp 1569139307
transform 1 0 4392 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1007
timestamp 1569139307
transform 1 0 4392 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1008
timestamp 1569139307
transform 1 0 4392 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1009
timestamp 1569139307
transform 1 0 4456 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1010
timestamp 1569139307
transform 1 0 4456 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1011
timestamp 1569139307
transform 1 0 2472 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1012
timestamp 1569139307
transform 1 0 2472 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1013
timestamp 1569139307
transform 1 0 2344 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1014
timestamp 1569139307
transform 1 0 2216 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1015
timestamp 1569139307
transform 1 0 2408 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1016
timestamp 1569139307
transform 1 0 2344 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1017
timestamp 1569139307
transform 1 0 2216 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1018
timestamp 1569139307
transform 1 0 2344 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1019
timestamp 1569139307
transform 1 0 2472 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1020
timestamp 1569139307
transform 1 0 2280 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1021
timestamp 1569139307
transform 1 0 2408 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1022
timestamp 1569139307
transform 1 0 2216 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1023
timestamp 1569139307
transform 1 0 2344 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1024
timestamp 1569139307
transform 1 0 2344 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1025
timestamp 1569139307
transform 1 0 2408 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1026
timestamp 1569139307
transform 1 0 2280 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1027
timestamp 1569139307
transform 1 0 2280 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1028
timestamp 1569139307
transform 1 0 2408 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1029
timestamp 1569139307
transform 1 0 2408 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1030
timestamp 1569139307
transform 1 0 2280 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1031
timestamp 1569139307
transform 1 0 2472 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1032
timestamp 1569139307
transform 1 0 2216 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1033
timestamp 1569139307
transform 1 0 2216 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1034
timestamp 1569139307
transform 1 0 2472 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1035
timestamp 1569139307
transform 1 0 2280 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1036
timestamp 1569139307
transform 1 0 2088 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1037
timestamp 1569139307
transform 1 0 2088 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1038
timestamp 1569139307
transform 1 0 1960 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1039
timestamp 1569139307
transform 1 0 2088 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1040
timestamp 1569139307
transform 1 0 2088 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1041
timestamp 1569139307
transform 1 0 2152 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1042
timestamp 1569139307
transform 1 0 2152 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1043
timestamp 1569139307
transform 1 0 1960 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1044
timestamp 1569139307
transform 1 0 2152 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1045
timestamp 1569139307
transform 1 0 1960 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1046
timestamp 1569139307
transform 1 0 1960 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1047
timestamp 1569139307
transform 1 0 1960 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1048
timestamp 1569139307
transform 1 0 2024 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1049
timestamp 1569139307
transform 1 0 2024 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1050
timestamp 1569139307
transform 1 0 2024 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1051
timestamp 1569139307
transform 1 0 1896 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1052
timestamp 1569139307
transform 1 0 2152 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1053
timestamp 1569139307
transform 1 0 1896 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1054
timestamp 1569139307
transform 1 0 2024 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1055
timestamp 1569139307
transform 1 0 2024 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1056
timestamp 1569139307
transform 1 0 1896 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1057
timestamp 1569139307
transform 1 0 2152 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1058
timestamp 1569139307
transform 1 0 1896 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1059
timestamp 1569139307
transform 1 0 2088 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1060
timestamp 1569139307
transform 1 0 1896 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1061
timestamp 1569139307
transform 1 0 1896 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1062
timestamp 1569139307
transform 1 0 2152 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1063
timestamp 1569139307
transform 1 0 1960 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1064
timestamp 1569139307
transform 1 0 1960 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1065
timestamp 1569139307
transform 1 0 1960 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1066
timestamp 1569139307
transform 1 0 1960 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1067
timestamp 1569139307
transform 1 0 2152 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1068
timestamp 1569139307
transform 1 0 1960 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1069
timestamp 1569139307
transform 1 0 2152 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1070
timestamp 1569139307
transform 1 0 2024 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1071
timestamp 1569139307
transform 1 0 2024 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1072
timestamp 1569139307
transform 1 0 2024 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1073
timestamp 1569139307
transform 1 0 2024 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1074
timestamp 1569139307
transform 1 0 2024 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1075
timestamp 1569139307
transform 1 0 2152 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1076
timestamp 1569139307
transform 1 0 2152 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1077
timestamp 1569139307
transform 1 0 1896 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1078
timestamp 1569139307
transform 1 0 2088 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1079
timestamp 1569139307
transform 1 0 1896 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1080
timestamp 1569139307
transform 1 0 1896 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1081
timestamp 1569139307
transform 1 0 2088 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1082
timestamp 1569139307
transform 1 0 2088 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1083
timestamp 1569139307
transform 1 0 2088 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1084
timestamp 1569139307
transform 1 0 1896 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1085
timestamp 1569139307
transform 1 0 2088 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1086
timestamp 1569139307
transform 1 0 2344 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1087
timestamp 1569139307
transform 1 0 2344 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1088
timestamp 1569139307
transform 1 0 2344 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1089
timestamp 1569139307
transform 1 0 2472 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1090
timestamp 1569139307
transform 1 0 2472 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1091
timestamp 1569139307
transform 1 0 2472 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1092
timestamp 1569139307
transform 1 0 2472 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1093
timestamp 1569139307
transform 1 0 2472 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1094
timestamp 1569139307
transform 1 0 2344 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1095
timestamp 1569139307
transform 1 0 2216 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1096
timestamp 1569139307
transform 1 0 2216 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1097
timestamp 1569139307
transform 1 0 2216 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1098
timestamp 1569139307
transform 1 0 2216 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1099
timestamp 1569139307
transform 1 0 2344 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1100
timestamp 1569139307
transform 1 0 2216 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1101
timestamp 1569139307
transform 1 0 2408 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1102
timestamp 1569139307
transform 1 0 2408 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1103
timestamp 1569139307
transform 1 0 2408 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1104
timestamp 1569139307
transform 1 0 2408 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1105
timestamp 1569139307
transform 1 0 2408 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1106
timestamp 1569139307
transform 1 0 2280 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1107
timestamp 1569139307
transform 1 0 2280 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1108
timestamp 1569139307
transform 1 0 2280 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1109
timestamp 1569139307
transform 1 0 2280 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1110
timestamp 1569139307
transform 1 0 2280 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1111
timestamp 1569139307
transform 1 0 1832 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1112
timestamp 1569139307
transform 1 0 1768 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1113
timestamp 1569139307
transform 1 0 1768 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1114
timestamp 1569139307
transform 1 0 1768 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1115
timestamp 1569139307
transform 1 0 1768 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1116
timestamp 1569139307
transform 1 0 1640 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1117
timestamp 1569139307
transform 1 0 1832 0 1 40
box -8 -8 8 8
use VIA2  VIA2_1118
timestamp 1569139307
transform 1 0 1832 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1119
timestamp 1569139307
transform 1 0 1832 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1120
timestamp 1569139307
transform 1 0 1768 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1121
timestamp 1569139307
transform 1 0 1832 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1122
timestamp 1569139307
transform 1 0 1704 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1123
timestamp 1569139307
transform 1 0 1704 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1124
timestamp 1569139307
transform 1 0 1640 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1125
timestamp 1569139307
transform 1 0 1640 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1126
timestamp 1569139307
transform 1 0 1704 0 1 104
box -8 -8 8 8
use VIA2  VIA2_1127
timestamp 1569139307
transform 1 0 1704 0 1 168
box -8 -8 8 8
use VIA2  VIA2_1128
timestamp 1569139307
transform 1 0 1512 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1129
timestamp 1569139307
transform 1 0 1320 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1130
timestamp 1569139307
transform 1 0 1320 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1131
timestamp 1569139307
transform 1 0 1320 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1132
timestamp 1569139307
transform 1 0 1512 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1133
timestamp 1569139307
transform 1 0 1512 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1134
timestamp 1569139307
transform 1 0 1448 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1135
timestamp 1569139307
transform 1 0 1448 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1136
timestamp 1569139307
transform 1 0 1384 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1137
timestamp 1569139307
transform 1 0 1384 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1138
timestamp 1569139307
transform 1 0 1384 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1139
timestamp 1569139307
transform 1 0 1384 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1140
timestamp 1569139307
transform 1 0 1512 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1141
timestamp 1569139307
transform 1 0 1512 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1142
timestamp 1569139307
transform 1 0 1448 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1143
timestamp 1569139307
transform 1 0 1512 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1144
timestamp 1569139307
transform 1 0 1448 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1145
timestamp 1569139307
transform 1 0 1448 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1146
timestamp 1569139307
transform 1 0 1640 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1147
timestamp 1569139307
transform 1 0 1640 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1148
timestamp 1569139307
transform 1 0 1704 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1149
timestamp 1569139307
transform 1 0 1704 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1150
timestamp 1569139307
transform 1 0 1832 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1151
timestamp 1569139307
transform 1 0 1832 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1152
timestamp 1569139307
transform 1 0 1832 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1153
timestamp 1569139307
transform 1 0 1832 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1154
timestamp 1569139307
transform 1 0 1832 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1155
timestamp 1569139307
transform 1 0 1768 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1156
timestamp 1569139307
transform 1 0 1768 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1157
timestamp 1569139307
transform 1 0 1768 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1158
timestamp 1569139307
transform 1 0 1704 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1159
timestamp 1569139307
transform 1 0 1640 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1160
timestamp 1569139307
transform 1 0 1640 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1161
timestamp 1569139307
transform 1 0 1640 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1162
timestamp 1569139307
transform 1 0 1704 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1163
timestamp 1569139307
transform 1 0 1704 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1164
timestamp 1569139307
transform 1 0 1768 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1165
timestamp 1569139307
transform 1 0 1768 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1166
timestamp 1569139307
transform 1 0 1576 0 1 296
box -8 -8 8 8
use VIA2  VIA2_1167
timestamp 1569139307
transform 1 0 1576 0 1 360
box -8 -8 8 8
use VIA2  VIA2_1168
timestamp 1569139307
transform 1 0 1576 0 1 424
box -8 -8 8 8
use VIA2  VIA2_1169
timestamp 1569139307
transform 1 0 1576 0 1 488
box -8 -8 8 8
use VIA2  VIA2_1170
timestamp 1569139307
transform 1 0 1576 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1171
timestamp 1569139307
transform 1 0 1576 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1172
timestamp 1569139307
transform 1 0 1576 0 1 232
box -8 -8 8 8
use VIA2  VIA2_1173
timestamp 1569139307
transform 1 0 1640 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1174
timestamp 1569139307
transform 1 0 1704 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1175
timestamp 1569139307
transform 1 0 1640 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1176
timestamp 1569139307
transform 1 0 1704 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1177
timestamp 1569139307
transform 1 0 1768 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1178
timestamp 1569139307
transform 1 0 1832 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1179
timestamp 1569139307
transform 1 0 1704 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1180
timestamp 1569139307
transform 1 0 1832 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1181
timestamp 1569139307
transform 1 0 1640 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1182
timestamp 1569139307
transform 1 0 1768 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1183
timestamp 1569139307
transform 1 0 1832 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1184
timestamp 1569139307
transform 1 0 1768 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1185
timestamp 1569139307
transform 1 0 1640 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1186
timestamp 1569139307
transform 1 0 1832 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1187
timestamp 1569139307
transform 1 0 1768 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1188
timestamp 1569139307
transform 1 0 1704 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1189
timestamp 1569139307
transform 1 0 1704 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1190
timestamp 1569139307
transform 1 0 1832 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1191
timestamp 1569139307
transform 1 0 1768 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1192
timestamp 1569139307
transform 1 0 1640 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1193
timestamp 1569139307
transform 1 0 1512 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1194
timestamp 1569139307
transform 1 0 1512 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1195
timestamp 1569139307
transform 1 0 1320 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1196
timestamp 1569139307
transform 1 0 1320 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1197
timestamp 1569139307
transform 1 0 1320 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1198
timestamp 1569139307
transform 1 0 1320 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1199
timestamp 1569139307
transform 1 0 1320 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1200
timestamp 1569139307
transform 1 0 1384 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1201
timestamp 1569139307
transform 1 0 1384 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1202
timestamp 1569139307
transform 1 0 1448 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1203
timestamp 1569139307
transform 1 0 1384 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1204
timestamp 1569139307
transform 1 0 1384 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1205
timestamp 1569139307
transform 1 0 1448 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1206
timestamp 1569139307
transform 1 0 1384 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1207
timestamp 1569139307
transform 1 0 1512 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1208
timestamp 1569139307
transform 1 0 1448 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1209
timestamp 1569139307
transform 1 0 1448 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1210
timestamp 1569139307
transform 1 0 1512 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1211
timestamp 1569139307
transform 1 0 1448 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1212
timestamp 1569139307
transform 1 0 1512 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1213
timestamp 1569139307
transform 1 0 1320 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1214
timestamp 1569139307
transform 1 0 1320 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1215
timestamp 1569139307
transform 1 0 1384 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1216
timestamp 1569139307
transform 1 0 1448 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1217
timestamp 1569139307
transform 1 0 1512 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1218
timestamp 1569139307
transform 1 0 1384 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1219
timestamp 1569139307
transform 1 0 1512 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1220
timestamp 1569139307
transform 1 0 1512 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1221
timestamp 1569139307
transform 1 0 1384 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1222
timestamp 1569139307
transform 1 0 1448 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1223
timestamp 1569139307
transform 1 0 1384 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1224
timestamp 1569139307
transform 1 0 1512 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1225
timestamp 1569139307
transform 1 0 1320 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1226
timestamp 1569139307
transform 1 0 1448 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1227
timestamp 1569139307
transform 1 0 1320 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1228
timestamp 1569139307
transform 1 0 1448 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1229
timestamp 1569139307
transform 1 0 1512 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1230
timestamp 1569139307
transform 1 0 1448 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1231
timestamp 1569139307
transform 1 0 1384 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1232
timestamp 1569139307
transform 1 0 1320 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1233
timestamp 1569139307
transform 1 0 1832 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1234
timestamp 1569139307
transform 1 0 1768 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1235
timestamp 1569139307
transform 1 0 1768 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1236
timestamp 1569139307
transform 1 0 1768 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1237
timestamp 1569139307
transform 1 0 1640 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1238
timestamp 1569139307
transform 1 0 1640 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1239
timestamp 1569139307
transform 1 0 1832 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1240
timestamp 1569139307
transform 1 0 1704 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1241
timestamp 1569139307
transform 1 0 1832 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1242
timestamp 1569139307
transform 1 0 1832 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1243
timestamp 1569139307
transform 1 0 1832 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1244
timestamp 1569139307
transform 1 0 1704 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1245
timestamp 1569139307
transform 1 0 1768 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1246
timestamp 1569139307
transform 1 0 1768 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1247
timestamp 1569139307
transform 1 0 1640 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1248
timestamp 1569139307
transform 1 0 1640 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1249
timestamp 1569139307
transform 1 0 1704 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1250
timestamp 1569139307
transform 1 0 1704 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1251
timestamp 1569139307
transform 1 0 1704 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1252
timestamp 1569139307
transform 1 0 1640 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1253
timestamp 1569139307
transform 1 0 1576 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1254
timestamp 1569139307
transform 1 0 1576 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1255
timestamp 1569139307
transform 1 0 1576 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1256
timestamp 1569139307
transform 1 0 1576 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1257
timestamp 1569139307
transform 1 0 1576 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1258
timestamp 1569139307
transform 1 0 1576 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1259
timestamp 1569139307
transform 1 0 1576 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1260
timestamp 1569139307
transform 1 0 1576 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1261
timestamp 1569139307
transform 1 0 1576 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1262
timestamp 1569139307
transform 1 0 1576 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1263
timestamp 1569139307
transform 1 0 2280 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1264
timestamp 1569139307
transform 1 0 2344 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1265
timestamp 1569139307
transform 1 0 2472 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1266
timestamp 1569139307
transform 1 0 2472 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1267
timestamp 1569139307
transform 1 0 2472 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1268
timestamp 1569139307
transform 1 0 2344 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1269
timestamp 1569139307
transform 1 0 2216 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1270
timestamp 1569139307
transform 1 0 2216 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1271
timestamp 1569139307
transform 1 0 2216 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1272
timestamp 1569139307
transform 1 0 2408 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1273
timestamp 1569139307
transform 1 0 2216 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1274
timestamp 1569139307
transform 1 0 2216 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1275
timestamp 1569139307
transform 1 0 2408 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1276
timestamp 1569139307
transform 1 0 2472 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1277
timestamp 1569139307
transform 1 0 2344 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1278
timestamp 1569139307
transform 1 0 2408 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1279
timestamp 1569139307
transform 1 0 2344 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1280
timestamp 1569139307
transform 1 0 2344 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1281
timestamp 1569139307
transform 1 0 2408 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1282
timestamp 1569139307
transform 1 0 2408 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1283
timestamp 1569139307
transform 1 0 2472 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1284
timestamp 1569139307
transform 1 0 2280 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1285
timestamp 1569139307
transform 1 0 2280 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1286
timestamp 1569139307
transform 1 0 2280 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1287
timestamp 1569139307
transform 1 0 2280 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1288
timestamp 1569139307
transform 1 0 1896 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1289
timestamp 1569139307
transform 1 0 1896 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1290
timestamp 1569139307
transform 1 0 1896 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1291
timestamp 1569139307
transform 1 0 1896 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1292
timestamp 1569139307
transform 1 0 2152 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1293
timestamp 1569139307
transform 1 0 1896 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1294
timestamp 1569139307
transform 1 0 1960 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1295
timestamp 1569139307
transform 1 0 1960 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1296
timestamp 1569139307
transform 1 0 1960 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1297
timestamp 1569139307
transform 1 0 1960 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1298
timestamp 1569139307
transform 1 0 1960 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1299
timestamp 1569139307
transform 1 0 2024 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1300
timestamp 1569139307
transform 1 0 2024 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1301
timestamp 1569139307
transform 1 0 2024 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1302
timestamp 1569139307
transform 1 0 2024 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1303
timestamp 1569139307
transform 1 0 2024 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1304
timestamp 1569139307
transform 1 0 2088 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1305
timestamp 1569139307
transform 1 0 2088 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1306
timestamp 1569139307
transform 1 0 2088 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1307
timestamp 1569139307
transform 1 0 2088 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1308
timestamp 1569139307
transform 1 0 2088 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1309
timestamp 1569139307
transform 1 0 2152 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1310
timestamp 1569139307
transform 1 0 2152 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1311
timestamp 1569139307
transform 1 0 2152 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1312
timestamp 1569139307
transform 1 0 2152 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1313
timestamp 1569139307
transform 1 0 2152 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1314
timestamp 1569139307
transform 1 0 1960 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1315
timestamp 1569139307
transform 1 0 2024 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1316
timestamp 1569139307
transform 1 0 2024 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1317
timestamp 1569139307
transform 1 0 1896 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1318
timestamp 1569139307
transform 1 0 2088 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1319
timestamp 1569139307
transform 1 0 2088 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1320
timestamp 1569139307
transform 1 0 2152 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1321
timestamp 1569139307
transform 1 0 1896 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1322
timestamp 1569139307
transform 1 0 2088 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1323
timestamp 1569139307
transform 1 0 2024 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1324
timestamp 1569139307
transform 1 0 2152 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1325
timestamp 1569139307
transform 1 0 2088 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1326
timestamp 1569139307
transform 1 0 2088 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1327
timestamp 1569139307
transform 1 0 2024 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1328
timestamp 1569139307
transform 1 0 2024 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1329
timestamp 1569139307
transform 1 0 1896 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1330
timestamp 1569139307
transform 1 0 2152 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1331
timestamp 1569139307
transform 1 0 1896 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1332
timestamp 1569139307
transform 1 0 2152 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1333
timestamp 1569139307
transform 1 0 1896 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1334
timestamp 1569139307
transform 1 0 1960 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1335
timestamp 1569139307
transform 1 0 1960 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1336
timestamp 1569139307
transform 1 0 1960 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1337
timestamp 1569139307
transform 1 0 1960 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1338
timestamp 1569139307
transform 1 0 2280 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1339
timestamp 1569139307
transform 1 0 2280 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1340
timestamp 1569139307
transform 1 0 2280 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1341
timestamp 1569139307
transform 1 0 2408 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1342
timestamp 1569139307
transform 1 0 2408 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1343
timestamp 1569139307
transform 1 0 2344 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1344
timestamp 1569139307
transform 1 0 2344 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1345
timestamp 1569139307
transform 1 0 2344 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1346
timestamp 1569139307
transform 1 0 2408 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1347
timestamp 1569139307
transform 1 0 2408 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1348
timestamp 1569139307
transform 1 0 2408 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1349
timestamp 1569139307
transform 1 0 2472 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1350
timestamp 1569139307
transform 1 0 2216 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1351
timestamp 1569139307
transform 1 0 2472 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1352
timestamp 1569139307
transform 1 0 2216 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1353
timestamp 1569139307
transform 1 0 2472 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1354
timestamp 1569139307
transform 1 0 2216 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1355
timestamp 1569139307
transform 1 0 2472 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1356
timestamp 1569139307
transform 1 0 2216 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1357
timestamp 1569139307
transform 1 0 2472 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1358
timestamp 1569139307
transform 1 0 2216 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1359
timestamp 1569139307
transform 1 0 2344 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1360
timestamp 1569139307
transform 1 0 2344 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1361
timestamp 1569139307
transform 1 0 2280 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1362
timestamp 1569139307
transform 1 0 2280 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1363
timestamp 1569139307
transform 1 0 1192 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1364
timestamp 1569139307
transform 1 0 1256 0 1 552
box -8 -8 8 8
use VIA2  VIA2_1365
timestamp 1569139307
transform 1 0 1256 0 1 616
box -8 -8 8 8
use VIA2  VIA2_1366
timestamp 1569139307
transform 1 0 616 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1367
timestamp 1569139307
transform 1 0 552 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1368
timestamp 1569139307
transform 1 0 616 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1369
timestamp 1569139307
transform 1 0 1256 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1370
timestamp 1569139307
transform 1 0 1256 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1371
timestamp 1569139307
transform 1 0 1256 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1372
timestamp 1569139307
transform 1 0 1256 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1373
timestamp 1569139307
transform 1 0 1256 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1374
timestamp 1569139307
transform 1 0 1064 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1375
timestamp 1569139307
transform 1 0 1064 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1376
timestamp 1569139307
transform 1 0 1192 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1377
timestamp 1569139307
transform 1 0 1192 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1378
timestamp 1569139307
transform 1 0 1192 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1379
timestamp 1569139307
transform 1 0 1192 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1380
timestamp 1569139307
transform 1 0 1064 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1381
timestamp 1569139307
transform 1 0 1128 0 1 744
box -8 -8 8 8
use VIA2  VIA2_1382
timestamp 1569139307
transform 1 0 1128 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1383
timestamp 1569139307
transform 1 0 1128 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1384
timestamp 1569139307
transform 1 0 1128 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1385
timestamp 1569139307
transform 1 0 1128 0 1 680
box -8 -8 8 8
use VIA2  VIA2_1386
timestamp 1569139307
transform 1 0 1064 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1387
timestamp 1569139307
transform 1 0 1000 0 1 808
box -8 -8 8 8
use VIA2  VIA2_1388
timestamp 1569139307
transform 1 0 1192 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1389
timestamp 1569139307
transform 1 0 1000 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1390
timestamp 1569139307
transform 1 0 1000 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1391
timestamp 1569139307
transform 1 0 936 0 1 872
box -8 -8 8 8
use VIA2  VIA2_1392
timestamp 1569139307
transform 1 0 936 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1393
timestamp 1569139307
transform 1 0 872 0 1 936
box -8 -8 8 8
use VIA2  VIA2_1394
timestamp 1569139307
transform 1 0 872 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1395
timestamp 1569139307
transform 1 0 744 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1396
timestamp 1569139307
transform 1 0 744 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1397
timestamp 1569139307
transform 1 0 872 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1398
timestamp 1569139307
transform 1 0 808 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1399
timestamp 1569139307
transform 1 0 872 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1400
timestamp 1569139307
transform 1 0 808 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1401
timestamp 1569139307
transform 1 0 936 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1402
timestamp 1569139307
transform 1 0 808 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1403
timestamp 1569139307
transform 1 0 680 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1404
timestamp 1569139307
transform 1 0 744 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1405
timestamp 1569139307
transform 1 0 936 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1406
timestamp 1569139307
transform 1 0 936 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1407
timestamp 1569139307
transform 1 0 808 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1408
timestamp 1569139307
transform 1 0 680 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1409
timestamp 1569139307
transform 1 0 744 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1410
timestamp 1569139307
transform 1 0 808 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1411
timestamp 1569139307
transform 1 0 936 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1412
timestamp 1569139307
transform 1 0 680 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1413
timestamp 1569139307
transform 1 0 872 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1414
timestamp 1569139307
transform 1 0 936 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1415
timestamp 1569139307
transform 1 0 872 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1416
timestamp 1569139307
transform 1 0 1128 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1417
timestamp 1569139307
transform 1 0 1000 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1418
timestamp 1569139307
transform 1 0 1256 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1419
timestamp 1569139307
transform 1 0 1000 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1420
timestamp 1569139307
transform 1 0 1256 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1421
timestamp 1569139307
transform 1 0 1128 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1422
timestamp 1569139307
transform 1 0 1000 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1423
timestamp 1569139307
transform 1 0 1064 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1424
timestamp 1569139307
transform 1 0 1064 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1425
timestamp 1569139307
transform 1 0 1256 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1426
timestamp 1569139307
transform 1 0 1064 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1427
timestamp 1569139307
transform 1 0 1064 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1428
timestamp 1569139307
transform 1 0 1128 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1429
timestamp 1569139307
transform 1 0 1128 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1430
timestamp 1569139307
transform 1 0 1064 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1431
timestamp 1569139307
transform 1 0 1192 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1432
timestamp 1569139307
transform 1 0 1192 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1433
timestamp 1569139307
transform 1 0 1192 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1434
timestamp 1569139307
transform 1 0 1192 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1435
timestamp 1569139307
transform 1 0 1192 0 1 1000
box -8 -8 8 8
use VIA2  VIA2_1436
timestamp 1569139307
transform 1 0 1128 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1437
timestamp 1569139307
transform 1 0 1256 0 1 1064
box -8 -8 8 8
use VIA2  VIA2_1438
timestamp 1569139307
transform 1 0 1000 0 1 1128
box -8 -8 8 8
use VIA2  VIA2_1439
timestamp 1569139307
transform 1 0 1256 0 1 1192
box -8 -8 8 8
use VIA2  VIA2_1440
timestamp 1569139307
transform 1 0 1000 0 1 1256
box -8 -8 8 8
use VIA2  VIA2_1441
timestamp 1569139307
transform 1 0 1000 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1442
timestamp 1569139307
transform 1 0 1256 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1443
timestamp 1569139307
transform 1 0 1128 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1444
timestamp 1569139307
transform 1 0 1064 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1445
timestamp 1569139307
transform 1 0 1000 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1446
timestamp 1569139307
transform 1 0 1256 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1447
timestamp 1569139307
transform 1 0 1000 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1448
timestamp 1569139307
transform 1 0 1192 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1449
timestamp 1569139307
transform 1 0 1064 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1450
timestamp 1569139307
transform 1 0 1064 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1451
timestamp 1569139307
transform 1 0 1192 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1452
timestamp 1569139307
transform 1 0 1192 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1453
timestamp 1569139307
transform 1 0 1128 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1454
timestamp 1569139307
transform 1 0 1064 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1455
timestamp 1569139307
transform 1 0 1256 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1456
timestamp 1569139307
transform 1 0 1256 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1457
timestamp 1569139307
transform 1 0 1192 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1458
timestamp 1569139307
transform 1 0 1000 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1459
timestamp 1569139307
transform 1 0 1128 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1460
timestamp 1569139307
transform 1 0 1128 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1461
timestamp 1569139307
transform 1 0 744 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1462
timestamp 1569139307
transform 1 0 680 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1463
timestamp 1569139307
transform 1 0 936 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1464
timestamp 1569139307
transform 1 0 744 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1465
timestamp 1569139307
transform 1 0 680 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1466
timestamp 1569139307
transform 1 0 936 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1467
timestamp 1569139307
transform 1 0 808 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1468
timestamp 1569139307
transform 1 0 936 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1469
timestamp 1569139307
transform 1 0 872 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1470
timestamp 1569139307
transform 1 0 808 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1471
timestamp 1569139307
transform 1 0 744 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1472
timestamp 1569139307
transform 1 0 872 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1473
timestamp 1569139307
transform 1 0 872 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1474
timestamp 1569139307
transform 1 0 808 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1475
timestamp 1569139307
transform 1 0 936 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1476
timestamp 1569139307
transform 1 0 680 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1477
timestamp 1569139307
transform 1 0 872 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1478
timestamp 1569139307
transform 1 0 808 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1479
timestamp 1569139307
transform 1 0 680 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1480
timestamp 1569139307
transform 1 0 744 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1481
timestamp 1569139307
transform 1 0 808 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1482
timestamp 1569139307
transform 1 0 936 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1483
timestamp 1569139307
transform 1 0 872 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1484
timestamp 1569139307
transform 1 0 808 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1485
timestamp 1569139307
transform 1 0 808 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1486
timestamp 1569139307
transform 1 0 936 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1487
timestamp 1569139307
transform 1 0 936 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1488
timestamp 1569139307
transform 1 0 872 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1489
timestamp 1569139307
transform 1 0 680 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1490
timestamp 1569139307
transform 1 0 744 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1491
timestamp 1569139307
transform 1 0 680 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1492
timestamp 1569139307
transform 1 0 680 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1493
timestamp 1569139307
transform 1 0 872 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1494
timestamp 1569139307
transform 1 0 744 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1495
timestamp 1569139307
transform 1 0 744 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1496
timestamp 1569139307
transform 1 0 808 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1497
timestamp 1569139307
transform 1 0 936 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1498
timestamp 1569139307
transform 1 0 744 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1499
timestamp 1569139307
transform 1 0 680 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1500
timestamp 1569139307
transform 1 0 872 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1501
timestamp 1569139307
transform 1 0 1000 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1502
timestamp 1569139307
transform 1 0 1256 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1503
timestamp 1569139307
transform 1 0 1128 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1504
timestamp 1569139307
transform 1 0 1064 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1505
timestamp 1569139307
transform 1 0 1256 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1506
timestamp 1569139307
transform 1 0 1256 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1507
timestamp 1569139307
transform 1 0 1000 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1508
timestamp 1569139307
transform 1 0 1128 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1509
timestamp 1569139307
transform 1 0 1192 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1510
timestamp 1569139307
transform 1 0 1192 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1511
timestamp 1569139307
transform 1 0 1000 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1512
timestamp 1569139307
transform 1 0 1000 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1513
timestamp 1569139307
transform 1 0 1256 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1514
timestamp 1569139307
transform 1 0 1064 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1515
timestamp 1569139307
transform 1 0 1064 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1516
timestamp 1569139307
transform 1 0 1064 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1517
timestamp 1569139307
transform 1 0 1128 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1518
timestamp 1569139307
transform 1 0 1128 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1519
timestamp 1569139307
transform 1 0 1192 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1520
timestamp 1569139307
transform 1 0 1192 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1521
timestamp 1569139307
transform 1 0 872 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1522
timestamp 1569139307
transform 1 0 1128 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1523
timestamp 1569139307
transform 1 0 936 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1524
timestamp 1569139307
transform 1 0 808 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1525
timestamp 1569139307
transform 1 0 1064 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1526
timestamp 1569139307
transform 1 0 680 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1527
timestamp 1569139307
transform 1 0 1000 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1528
timestamp 1569139307
transform 1 0 1192 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1529
timestamp 1569139307
transform 1 0 1256 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1530
timestamp 1569139307
transform 1 0 744 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1531
timestamp 1569139307
transform 1 0 488 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1532
timestamp 1569139307
transform 1 0 488 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1533
timestamp 1569139307
transform 1 0 424 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1534
timestamp 1569139307
transform 1 0 616 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1535
timestamp 1569139307
transform 1 0 552 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1536
timestamp 1569139307
transform 1 0 616 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1537
timestamp 1569139307
transform 1 0 552 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1538
timestamp 1569139307
transform 1 0 424 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1539
timestamp 1569139307
transform 1 0 616 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1540
timestamp 1569139307
transform 1 0 552 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1541
timestamp 1569139307
transform 1 0 616 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1542
timestamp 1569139307
transform 1 0 360 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1543
timestamp 1569139307
transform 1 0 488 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1544
timestamp 1569139307
transform 1 0 360 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1545
timestamp 1569139307
transform 1 0 488 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1546
timestamp 1569139307
transform 1 0 424 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1547
timestamp 1569139307
transform 1 0 552 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1548
timestamp 1569139307
transform 1 0 296 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1549
timestamp 1569139307
transform 1 0 40 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1550
timestamp 1569139307
transform 1 0 296 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1551
timestamp 1569139307
transform 1 0 40 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1552
timestamp 1569139307
transform 1 0 232 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1553
timestamp 1569139307
transform 1 0 168 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1554
timestamp 1569139307
transform 1 0 232 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1555
timestamp 1569139307
transform 1 0 232 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1556
timestamp 1569139307
transform 1 0 104 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1557
timestamp 1569139307
transform 1 0 296 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1558
timestamp 1569139307
transform 1 0 296 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1559
timestamp 1569139307
transform 1 0 168 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1560
timestamp 1569139307
transform 1 0 296 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1561
timestamp 1569139307
transform 1 0 168 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1562
timestamp 1569139307
transform 1 0 104 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1563
timestamp 1569139307
transform 1 0 168 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1564
timestamp 1569139307
transform 1 0 232 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1565
timestamp 1569139307
transform 1 0 104 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1566
timestamp 1569139307
transform 1 0 360 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1567
timestamp 1569139307
transform 1 0 360 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1568
timestamp 1569139307
transform 1 0 616 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1569
timestamp 1569139307
transform 1 0 552 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1570
timestamp 1569139307
transform 1 0 424 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1571
timestamp 1569139307
transform 1 0 360 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1572
timestamp 1569139307
transform 1 0 616 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1573
timestamp 1569139307
transform 1 0 424 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1574
timestamp 1569139307
transform 1 0 488 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1575
timestamp 1569139307
transform 1 0 552 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1576
timestamp 1569139307
transform 1 0 424 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1577
timestamp 1569139307
transform 1 0 424 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1578
timestamp 1569139307
transform 1 0 488 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1579
timestamp 1569139307
transform 1 0 488 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1580
timestamp 1569139307
transform 1 0 360 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1581
timestamp 1569139307
transform 1 0 552 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1582
timestamp 1569139307
transform 1 0 552 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1583
timestamp 1569139307
transform 1 0 488 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1584
timestamp 1569139307
transform 1 0 616 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1585
timestamp 1569139307
transform 1 0 616 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1586
timestamp 1569139307
transform 1 0 488 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1587
timestamp 1569139307
transform 1 0 552 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1588
timestamp 1569139307
transform 1 0 616 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1589
timestamp 1569139307
transform 1 0 232 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1590
timestamp 1569139307
transform 1 0 296 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1591
timestamp 1569139307
transform 1 0 424 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1592
timestamp 1569139307
transform 1 0 360 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1593
timestamp 1569139307
transform 1 0 552 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1594
timestamp 1569139307
transform 1 0 488 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1595
timestamp 1569139307
transform 1 0 424 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1596
timestamp 1569139307
transform 1 0 552 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1597
timestamp 1569139307
transform 1 0 360 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1598
timestamp 1569139307
transform 1 0 616 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1599
timestamp 1569139307
transform 1 0 488 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1600
timestamp 1569139307
transform 1 0 424 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1601
timestamp 1569139307
transform 1 0 360 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1602
timestamp 1569139307
transform 1 0 488 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1603
timestamp 1569139307
transform 1 0 616 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1604
timestamp 1569139307
transform 1 0 360 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1605
timestamp 1569139307
transform 1 0 616 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1606
timestamp 1569139307
transform 1 0 552 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1607
timestamp 1569139307
transform 1 0 424 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1608
timestamp 1569139307
transform 1 0 488 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1609
timestamp 1569139307
transform 1 0 424 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1610
timestamp 1569139307
transform 1 0 488 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1611
timestamp 1569139307
transform 1 0 552 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1612
timestamp 1569139307
transform 1 0 552 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1613
timestamp 1569139307
transform 1 0 360 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1614
timestamp 1569139307
transform 1 0 360 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1615
timestamp 1569139307
transform 1 0 616 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1616
timestamp 1569139307
transform 1 0 424 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1617
timestamp 1569139307
transform 1 0 616 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1618
timestamp 1569139307
transform 1 0 40 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1619
timestamp 1569139307
transform 1 0 168 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1620
timestamp 1569139307
transform 1 0 296 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1621
timestamp 1569139307
transform 1 0 40 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1622
timestamp 1569139307
transform 1 0 232 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1623
timestamp 1569139307
transform 1 0 296 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1624
timestamp 1569139307
transform 1 0 168 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1625
timestamp 1569139307
transform 1 0 296 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1626
timestamp 1569139307
transform 1 0 104 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1627
timestamp 1569139307
transform 1 0 168 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1628
timestamp 1569139307
transform 1 0 168 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1629
timestamp 1569139307
transform 1 0 40 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1630
timestamp 1569139307
transform 1 0 296 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1631
timestamp 1569139307
transform 1 0 168 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1632
timestamp 1569139307
transform 1 0 104 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1633
timestamp 1569139307
transform 1 0 232 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1634
timestamp 1569139307
transform 1 0 104 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1635
timestamp 1569139307
transform 1 0 232 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1636
timestamp 1569139307
transform 1 0 40 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1637
timestamp 1569139307
transform 1 0 296 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1638
timestamp 1569139307
transform 1 0 232 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1639
timestamp 1569139307
transform 1 0 104 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1640
timestamp 1569139307
transform 1 0 232 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1641
timestamp 1569139307
transform 1 0 40 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1642
timestamp 1569139307
transform 1 0 104 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1643
timestamp 1569139307
transform 1 0 296 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1644
timestamp 1569139307
transform 1 0 40 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1645
timestamp 1569139307
transform 1 0 296 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1646
timestamp 1569139307
transform 1 0 296 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1647
timestamp 1569139307
transform 1 0 40 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1648
timestamp 1569139307
transform 1 0 168 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1649
timestamp 1569139307
transform 1 0 232 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1650
timestamp 1569139307
transform 1 0 40 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1651
timestamp 1569139307
transform 1 0 168 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1652
timestamp 1569139307
transform 1 0 104 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1653
timestamp 1569139307
transform 1 0 40 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1654
timestamp 1569139307
transform 1 0 232 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1655
timestamp 1569139307
transform 1 0 104 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1656
timestamp 1569139307
transform 1 0 168 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1657
timestamp 1569139307
transform 1 0 232 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1658
timestamp 1569139307
transform 1 0 40 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1659
timestamp 1569139307
transform 1 0 104 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1660
timestamp 1569139307
transform 1 0 104 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1661
timestamp 1569139307
transform 1 0 296 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1662
timestamp 1569139307
transform 1 0 104 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1663
timestamp 1569139307
transform 1 0 168 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1664
timestamp 1569139307
transform 1 0 232 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1665
timestamp 1569139307
transform 1 0 168 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1666
timestamp 1569139307
transform 1 0 296 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1667
timestamp 1569139307
transform 1 0 232 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1668
timestamp 1569139307
transform 1 0 424 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1669
timestamp 1569139307
transform 1 0 488 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1670
timestamp 1569139307
transform 1 0 424 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1671
timestamp 1569139307
transform 1 0 424 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1672
timestamp 1569139307
transform 1 0 488 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1673
timestamp 1569139307
transform 1 0 616 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1674
timestamp 1569139307
transform 1 0 424 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1675
timestamp 1569139307
transform 1 0 360 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1676
timestamp 1569139307
transform 1 0 616 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1677
timestamp 1569139307
transform 1 0 552 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1678
timestamp 1569139307
transform 1 0 552 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1679
timestamp 1569139307
transform 1 0 616 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1680
timestamp 1569139307
transform 1 0 552 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1681
timestamp 1569139307
transform 1 0 552 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1682
timestamp 1569139307
transform 1 0 488 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1683
timestamp 1569139307
transform 1 0 360 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1684
timestamp 1569139307
transform 1 0 552 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1685
timestamp 1569139307
transform 1 0 616 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1686
timestamp 1569139307
transform 1 0 488 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1687
timestamp 1569139307
transform 1 0 360 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1688
timestamp 1569139307
transform 1 0 616 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1689
timestamp 1569139307
transform 1 0 360 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1690
timestamp 1569139307
transform 1 0 424 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1691
timestamp 1569139307
transform 1 0 360 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1692
timestamp 1569139307
transform 1 0 488 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1693
timestamp 1569139307
transform 1 0 1192 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1694
timestamp 1569139307
transform 1 0 1192 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1695
timestamp 1569139307
transform 1 0 1256 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1696
timestamp 1569139307
transform 1 0 1128 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1697
timestamp 1569139307
transform 1 0 1064 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1698
timestamp 1569139307
transform 1 0 1128 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1699
timestamp 1569139307
transform 1 0 1192 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1700
timestamp 1569139307
transform 1 0 1128 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1701
timestamp 1569139307
transform 1 0 1192 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1702
timestamp 1569139307
transform 1 0 1128 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1703
timestamp 1569139307
transform 1 0 1256 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1704
timestamp 1569139307
transform 1 0 1064 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1705
timestamp 1569139307
transform 1 0 1000 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1706
timestamp 1569139307
transform 1 0 1256 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1707
timestamp 1569139307
transform 1 0 1000 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1708
timestamp 1569139307
transform 1 0 1256 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1709
timestamp 1569139307
transform 1 0 1000 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1710
timestamp 1569139307
transform 1 0 1256 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1711
timestamp 1569139307
transform 1 0 1128 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1712
timestamp 1569139307
transform 1 0 1000 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1713
timestamp 1569139307
transform 1 0 1064 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1714
timestamp 1569139307
transform 1 0 1064 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1715
timestamp 1569139307
transform 1 0 1192 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1716
timestamp 1569139307
transform 1 0 1064 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1717
timestamp 1569139307
transform 1 0 1000 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1718
timestamp 1569139307
transform 1 0 808 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1719
timestamp 1569139307
transform 1 0 680 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1720
timestamp 1569139307
transform 1 0 872 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1721
timestamp 1569139307
transform 1 0 936 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1722
timestamp 1569139307
transform 1 0 872 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1723
timestamp 1569139307
transform 1 0 936 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1724
timestamp 1569139307
transform 1 0 744 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1725
timestamp 1569139307
transform 1 0 744 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1726
timestamp 1569139307
transform 1 0 744 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1727
timestamp 1569139307
transform 1 0 872 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1728
timestamp 1569139307
transform 1 0 744 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1729
timestamp 1569139307
transform 1 0 744 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1730
timestamp 1569139307
transform 1 0 680 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1731
timestamp 1569139307
transform 1 0 808 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1732
timestamp 1569139307
transform 1 0 808 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1733
timestamp 1569139307
transform 1 0 808 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1734
timestamp 1569139307
transform 1 0 808 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1735
timestamp 1569139307
transform 1 0 872 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1736
timestamp 1569139307
transform 1 0 680 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1737
timestamp 1569139307
transform 1 0 680 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1738
timestamp 1569139307
transform 1 0 936 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1739
timestamp 1569139307
transform 1 0 872 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1740
timestamp 1569139307
transform 1 0 936 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1741
timestamp 1569139307
transform 1 0 680 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1742
timestamp 1569139307
transform 1 0 936 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1743
timestamp 1569139307
transform 1 0 936 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1744
timestamp 1569139307
transform 1 0 936 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1745
timestamp 1569139307
transform 1 0 808 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1746
timestamp 1569139307
transform 1 0 680 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1747
timestamp 1569139307
transform 1 0 680 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1748
timestamp 1569139307
transform 1 0 680 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1749
timestamp 1569139307
transform 1 0 872 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1750
timestamp 1569139307
transform 1 0 680 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1751
timestamp 1569139307
transform 1 0 808 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1752
timestamp 1569139307
transform 1 0 744 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1753
timestamp 1569139307
transform 1 0 872 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1754
timestamp 1569139307
transform 1 0 808 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1755
timestamp 1569139307
transform 1 0 872 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1756
timestamp 1569139307
transform 1 0 872 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1757
timestamp 1569139307
transform 1 0 872 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1758
timestamp 1569139307
transform 1 0 936 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1759
timestamp 1569139307
transform 1 0 744 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1760
timestamp 1569139307
transform 1 0 744 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1761
timestamp 1569139307
transform 1 0 936 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1762
timestamp 1569139307
transform 1 0 744 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1763
timestamp 1569139307
transform 1 0 936 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1764
timestamp 1569139307
transform 1 0 808 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1765
timestamp 1569139307
transform 1 0 680 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1766
timestamp 1569139307
transform 1 0 744 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1767
timestamp 1569139307
transform 1 0 808 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1768
timestamp 1569139307
transform 1 0 1064 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1769
timestamp 1569139307
transform 1 0 1064 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1770
timestamp 1569139307
transform 1 0 1128 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1771
timestamp 1569139307
transform 1 0 1000 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1772
timestamp 1569139307
transform 1 0 1192 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1773
timestamp 1569139307
transform 1 0 1192 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1774
timestamp 1569139307
transform 1 0 1192 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1775
timestamp 1569139307
transform 1 0 1192 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1776
timestamp 1569139307
transform 1 0 1192 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1777
timestamp 1569139307
transform 1 0 1064 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1778
timestamp 1569139307
transform 1 0 1000 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1779
timestamp 1569139307
transform 1 0 1064 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1780
timestamp 1569139307
transform 1 0 1000 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1781
timestamp 1569139307
transform 1 0 1064 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1782
timestamp 1569139307
transform 1 0 1128 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1783
timestamp 1569139307
transform 1 0 1000 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1784
timestamp 1569139307
transform 1 0 1128 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1785
timestamp 1569139307
transform 1 0 1000 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1786
timestamp 1569139307
transform 1 0 1256 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1787
timestamp 1569139307
transform 1 0 1256 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1788
timestamp 1569139307
transform 1 0 1256 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_1789
timestamp 1569139307
transform 1 0 1128 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_1790
timestamp 1569139307
transform 1 0 1256 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_1791
timestamp 1569139307
transform 1 0 1256 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_1792
timestamp 1569139307
transform 1 0 1128 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_1793
timestamp 1569139307
transform 1 0 2280 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1794
timestamp 1569139307
transform 1 0 2280 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1795
timestamp 1569139307
transform 1 0 2472 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1796
timestamp 1569139307
transform 1 0 2344 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1797
timestamp 1569139307
transform 1 0 2216 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1798
timestamp 1569139307
transform 1 0 2472 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1799
timestamp 1569139307
transform 1 0 2344 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1800
timestamp 1569139307
transform 1 0 2216 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1801
timestamp 1569139307
transform 1 0 2408 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1802
timestamp 1569139307
transform 1 0 2408 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1803
timestamp 1569139307
transform 1 0 2408 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1804
timestamp 1569139307
transform 1 0 2344 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1805
timestamp 1569139307
transform 1 0 2344 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1806
timestamp 1569139307
transform 1 0 2408 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1807
timestamp 1569139307
transform 1 0 2216 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1808
timestamp 1569139307
transform 1 0 2280 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1809
timestamp 1569139307
transform 1 0 2472 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1810
timestamp 1569139307
transform 1 0 2216 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1811
timestamp 1569139307
transform 1 0 2472 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1812
timestamp 1569139307
transform 1 0 2280 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1813
timestamp 1569139307
transform 1 0 2024 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1814
timestamp 1569139307
transform 1 0 1896 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1815
timestamp 1569139307
transform 1 0 2024 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1816
timestamp 1569139307
transform 1 0 2088 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1817
timestamp 1569139307
transform 1 0 2088 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1818
timestamp 1569139307
transform 1 0 2024 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1819
timestamp 1569139307
transform 1 0 2088 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1820
timestamp 1569139307
transform 1 0 2152 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1821
timestamp 1569139307
transform 1 0 1896 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1822
timestamp 1569139307
transform 1 0 1896 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1823
timestamp 1569139307
transform 1 0 2152 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1824
timestamp 1569139307
transform 1 0 1896 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1825
timestamp 1569139307
transform 1 0 1960 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1826
timestamp 1569139307
transform 1 0 1960 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1827
timestamp 1569139307
transform 1 0 1960 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1828
timestamp 1569139307
transform 1 0 2152 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1829
timestamp 1569139307
transform 1 0 1960 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1830
timestamp 1569139307
transform 1 0 2088 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1831
timestamp 1569139307
transform 1 0 2024 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1832
timestamp 1569139307
transform 1 0 2152 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1833
timestamp 1569139307
transform 1 0 1896 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1834
timestamp 1569139307
transform 1 0 2024 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1835
timestamp 1569139307
transform 1 0 2088 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1836
timestamp 1569139307
transform 1 0 2024 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1837
timestamp 1569139307
transform 1 0 2152 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1838
timestamp 1569139307
transform 1 0 2152 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1839
timestamp 1569139307
transform 1 0 1896 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1840
timestamp 1569139307
transform 1 0 1960 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1841
timestamp 1569139307
transform 1 0 1960 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1842
timestamp 1569139307
transform 1 0 1960 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1843
timestamp 1569139307
transform 1 0 2024 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1844
timestamp 1569139307
transform 1 0 2024 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1845
timestamp 1569139307
transform 1 0 1896 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1846
timestamp 1569139307
transform 1 0 2088 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1847
timestamp 1569139307
transform 1 0 2088 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1848
timestamp 1569139307
transform 1 0 1960 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1849
timestamp 1569139307
transform 1 0 2152 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1850
timestamp 1569139307
transform 1 0 2152 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1851
timestamp 1569139307
transform 1 0 2088 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1852
timestamp 1569139307
transform 1 0 1896 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1853
timestamp 1569139307
transform 1 0 2344 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1854
timestamp 1569139307
transform 1 0 2280 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1855
timestamp 1569139307
transform 1 0 2344 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1856
timestamp 1569139307
transform 1 0 2408 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1857
timestamp 1569139307
transform 1 0 2408 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1858
timestamp 1569139307
transform 1 0 2472 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1859
timestamp 1569139307
transform 1 0 2472 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1860
timestamp 1569139307
transform 1 0 2344 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1861
timestamp 1569139307
transform 1 0 2344 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1862
timestamp 1569139307
transform 1 0 2408 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1863
timestamp 1569139307
transform 1 0 2408 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1864
timestamp 1569139307
transform 1 0 2280 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1865
timestamp 1569139307
transform 1 0 2472 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1866
timestamp 1569139307
transform 1 0 2472 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1867
timestamp 1569139307
transform 1 0 2216 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1868
timestamp 1569139307
transform 1 0 2280 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1869
timestamp 1569139307
transform 1 0 2280 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1870
timestamp 1569139307
transform 1 0 2216 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1871
timestamp 1569139307
transform 1 0 2216 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1872
timestamp 1569139307
transform 1 0 2216 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1873
timestamp 1569139307
transform 1 0 1896 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1874
timestamp 1569139307
transform 1 0 2344 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1875
timestamp 1569139307
transform 1 0 2408 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1876
timestamp 1569139307
transform 1 0 1960 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1877
timestamp 1569139307
transform 1 0 2472 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1878
timestamp 1569139307
transform 1 0 2024 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1879
timestamp 1569139307
transform 1 0 2088 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1880
timestamp 1569139307
transform 1 0 2152 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1881
timestamp 1569139307
transform 1 0 2216 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1882
timestamp 1569139307
transform 1 0 2280 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1883
timestamp 1569139307
transform 1 0 1768 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1884
timestamp 1569139307
transform 1 0 1768 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1885
timestamp 1569139307
transform 1 0 1832 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1886
timestamp 1569139307
transform 1 0 1704 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1887
timestamp 1569139307
transform 1 0 1768 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1888
timestamp 1569139307
transform 1 0 1832 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1889
timestamp 1569139307
transform 1 0 1640 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1890
timestamp 1569139307
transform 1 0 1640 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1891
timestamp 1569139307
transform 1 0 1640 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1892
timestamp 1569139307
transform 1 0 1704 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1893
timestamp 1569139307
transform 1 0 1704 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1894
timestamp 1569139307
transform 1 0 1704 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1895
timestamp 1569139307
transform 1 0 1832 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1896
timestamp 1569139307
transform 1 0 1640 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1897
timestamp 1569139307
transform 1 0 1832 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1898
timestamp 1569139307
transform 1 0 1768 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1899
timestamp 1569139307
transform 1 0 1512 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1900
timestamp 1569139307
transform 1 0 1512 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1901
timestamp 1569139307
transform 1 0 1320 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1902
timestamp 1569139307
transform 1 0 1320 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1903
timestamp 1569139307
transform 1 0 1384 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1904
timestamp 1569139307
transform 1 0 1384 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1905
timestamp 1569139307
transform 1 0 1448 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1906
timestamp 1569139307
transform 1 0 1448 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1907
timestamp 1569139307
transform 1 0 1512 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1908
timestamp 1569139307
transform 1 0 1320 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1909
timestamp 1569139307
transform 1 0 1320 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1910
timestamp 1569139307
transform 1 0 1512 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1911
timestamp 1569139307
transform 1 0 1448 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1912
timestamp 1569139307
transform 1 0 1384 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1913
timestamp 1569139307
transform 1 0 1448 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1914
timestamp 1569139307
transform 1 0 1384 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1915
timestamp 1569139307
transform 1 0 1384 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1916
timestamp 1569139307
transform 1 0 1448 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1917
timestamp 1569139307
transform 1 0 1448 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1918
timestamp 1569139307
transform 1 0 1512 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1919
timestamp 1569139307
transform 1 0 1320 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1920
timestamp 1569139307
transform 1 0 1448 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1921
timestamp 1569139307
transform 1 0 1448 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1922
timestamp 1569139307
transform 1 0 1384 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1923
timestamp 1569139307
transform 1 0 1512 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1924
timestamp 1569139307
transform 1 0 1512 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1925
timestamp 1569139307
transform 1 0 1384 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1926
timestamp 1569139307
transform 1 0 1320 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1927
timestamp 1569139307
transform 1 0 1320 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1928
timestamp 1569139307
transform 1 0 1384 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1929
timestamp 1569139307
transform 1 0 1320 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1930
timestamp 1569139307
transform 1 0 1512 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1931
timestamp 1569139307
transform 1 0 1704 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1932
timestamp 1569139307
transform 1 0 1768 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1933
timestamp 1569139307
transform 1 0 1832 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1934
timestamp 1569139307
transform 1 0 1704 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1935
timestamp 1569139307
transform 1 0 1704 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1936
timestamp 1569139307
transform 1 0 1768 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1937
timestamp 1569139307
transform 1 0 1768 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1938
timestamp 1569139307
transform 1 0 1832 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1939
timestamp 1569139307
transform 1 0 1832 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1940
timestamp 1569139307
transform 1 0 1640 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1941
timestamp 1569139307
transform 1 0 1640 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1942
timestamp 1569139307
transform 1 0 1832 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1943
timestamp 1569139307
transform 1 0 1640 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1944
timestamp 1569139307
transform 1 0 1640 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1945
timestamp 1569139307
transform 1 0 1704 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1946
timestamp 1569139307
transform 1 0 1768 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1947
timestamp 1569139307
transform 1 0 1576 0 1 1320
box -8 -8 8 8
use VIA2  VIA2_1948
timestamp 1569139307
transform 1 0 1576 0 1 1448
box -8 -8 8 8
use VIA2  VIA2_1949
timestamp 1569139307
transform 1 0 1320 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1950
timestamp 1569139307
transform 1 0 1640 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1951
timestamp 1569139307
transform 1 0 1448 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1952
timestamp 1569139307
transform 1 0 1704 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1953
timestamp 1569139307
transform 1 0 1576 0 1 1640
box -8 -8 8 8
use VIA2  VIA2_1954
timestamp 1569139307
transform 1 0 1576 0 1 1768
box -8 -8 8 8
use VIA2  VIA2_1955
timestamp 1569139307
transform 1 0 1768 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1956
timestamp 1569139307
transform 1 0 1512 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1957
timestamp 1569139307
transform 1 0 1832 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1958
timestamp 1569139307
transform 1 0 1384 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1959
timestamp 1569139307
transform 1 0 1576 0 1 1576
box -8 -8 8 8
use VIA2  VIA2_1960
timestamp 1569139307
transform 1 0 1576 0 1 1832
box -8 -8 8 8
use VIA2  VIA2_1961
timestamp 1569139307
transform 1 0 1576 0 1 1384
box -8 -8 8 8
use VIA2  VIA2_1962
timestamp 1569139307
transform 1 0 1576 0 1 1512
box -8 -8 8 8
use VIA2  VIA2_1963
timestamp 1569139307
transform 1 0 1576 0 1 1704
box -8 -8 8 8
use VIA2  VIA2_1964
timestamp 1569139307
transform 1 0 1704 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1965
timestamp 1569139307
transform 1 0 1768 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1966
timestamp 1569139307
transform 1 0 1704 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1967
timestamp 1569139307
transform 1 0 1832 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1968
timestamp 1569139307
transform 1 0 1768 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1969
timestamp 1569139307
transform 1 0 1768 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1970
timestamp 1569139307
transform 1 0 1768 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1971
timestamp 1569139307
transform 1 0 1640 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1972
timestamp 1569139307
transform 1 0 1640 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1973
timestamp 1569139307
transform 1 0 1704 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1974
timestamp 1569139307
transform 1 0 1768 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1975
timestamp 1569139307
transform 1 0 1832 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1976
timestamp 1569139307
transform 1 0 1640 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1977
timestamp 1569139307
transform 1 0 1832 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1978
timestamp 1569139307
transform 1 0 1832 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1979
timestamp 1569139307
transform 1 0 1832 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1980
timestamp 1569139307
transform 1 0 1640 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1981
timestamp 1569139307
transform 1 0 1640 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1982
timestamp 1569139307
transform 1 0 1704 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1983
timestamp 1569139307
transform 1 0 1704 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1984
timestamp 1569139307
transform 1 0 1384 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1985
timestamp 1569139307
transform 1 0 1512 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1986
timestamp 1569139307
transform 1 0 1448 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1987
timestamp 1569139307
transform 1 0 1512 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1988
timestamp 1569139307
transform 1 0 1512 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1989
timestamp 1569139307
transform 1 0 1512 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1990
timestamp 1569139307
transform 1 0 1320 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_1991
timestamp 1569139307
transform 1 0 1320 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1992
timestamp 1569139307
transform 1 0 1384 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1993
timestamp 1569139307
transform 1 0 1320 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1994
timestamp 1569139307
transform 1 0 1384 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_1995
timestamp 1569139307
transform 1 0 1320 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_1996
timestamp 1569139307
transform 1 0 1512 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1997
timestamp 1569139307
transform 1 0 1448 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_1998
timestamp 1569139307
transform 1 0 1448 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_1999
timestamp 1569139307
transform 1 0 1448 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2000
timestamp 1569139307
transform 1 0 1448 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2001
timestamp 1569139307
transform 1 0 1320 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2002
timestamp 1569139307
transform 1 0 1384 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2003
timestamp 1569139307
transform 1 0 1384 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2004
timestamp 1569139307
transform 1 0 1384 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2005
timestamp 1569139307
transform 1 0 1320 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2006
timestamp 1569139307
transform 1 0 1512 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2007
timestamp 1569139307
transform 1 0 1384 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2008
timestamp 1569139307
transform 1 0 1320 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2009
timestamp 1569139307
transform 1 0 1512 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2010
timestamp 1569139307
transform 1 0 1320 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2011
timestamp 1569139307
transform 1 0 1384 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2012
timestamp 1569139307
transform 1 0 1320 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2013
timestamp 1569139307
transform 1 0 1448 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2014
timestamp 1569139307
transform 1 0 1384 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2015
timestamp 1569139307
transform 1 0 1448 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2016
timestamp 1569139307
transform 1 0 1384 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2017
timestamp 1569139307
transform 1 0 1448 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2018
timestamp 1569139307
transform 1 0 1320 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2019
timestamp 1569139307
transform 1 0 1512 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2020
timestamp 1569139307
transform 1 0 1448 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2021
timestamp 1569139307
transform 1 0 1512 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2022
timestamp 1569139307
transform 1 0 1448 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2023
timestamp 1569139307
transform 1 0 1512 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2024
timestamp 1569139307
transform 1 0 1704 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2025
timestamp 1569139307
transform 1 0 1704 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2026
timestamp 1569139307
transform 1 0 1768 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2027
timestamp 1569139307
transform 1 0 1768 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2028
timestamp 1569139307
transform 1 0 1704 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2029
timestamp 1569139307
transform 1 0 1768 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2030
timestamp 1569139307
transform 1 0 1832 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2031
timestamp 1569139307
transform 1 0 1832 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2032
timestamp 1569139307
transform 1 0 1832 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2033
timestamp 1569139307
transform 1 0 1832 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2034
timestamp 1569139307
transform 1 0 1832 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2035
timestamp 1569139307
transform 1 0 1704 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2036
timestamp 1569139307
transform 1 0 1704 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2037
timestamp 1569139307
transform 1 0 1768 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2038
timestamp 1569139307
transform 1 0 1768 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2039
timestamp 1569139307
transform 1 0 1640 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2040
timestamp 1569139307
transform 1 0 1640 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2041
timestamp 1569139307
transform 1 0 1640 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2042
timestamp 1569139307
transform 1 0 1640 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2043
timestamp 1569139307
transform 1 0 1640 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2044
timestamp 1569139307
transform 1 0 1576 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2045
timestamp 1569139307
transform 1 0 1576 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2046
timestamp 1569139307
transform 1 0 1576 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2047
timestamp 1569139307
transform 1 0 1576 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2048
timestamp 1569139307
transform 1 0 1576 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2049
timestamp 1569139307
transform 1 0 1576 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2050
timestamp 1569139307
transform 1 0 1576 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2051
timestamp 1569139307
transform 1 0 1576 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2052
timestamp 1569139307
transform 1 0 1576 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2053
timestamp 1569139307
transform 1 0 1576 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2054
timestamp 1569139307
transform 1 0 2344 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2055
timestamp 1569139307
transform 1 0 2408 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2056
timestamp 1569139307
transform 1 0 2472 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2057
timestamp 1569139307
transform 1 0 2408 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2058
timestamp 1569139307
transform 1 0 2280 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2059
timestamp 1569139307
transform 1 0 2280 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2060
timestamp 1569139307
transform 1 0 2280 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2061
timestamp 1569139307
transform 1 0 2344 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2062
timestamp 1569139307
transform 1 0 2344 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2063
timestamp 1569139307
transform 1 0 2216 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2064
timestamp 1569139307
transform 1 0 2344 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2065
timestamp 1569139307
transform 1 0 2280 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2066
timestamp 1569139307
transform 1 0 2280 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2067
timestamp 1569139307
transform 1 0 2216 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2068
timestamp 1569139307
transform 1 0 2216 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2069
timestamp 1569139307
transform 1 0 2216 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2070
timestamp 1569139307
transform 1 0 2408 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2071
timestamp 1569139307
transform 1 0 2472 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2072
timestamp 1569139307
transform 1 0 2216 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2073
timestamp 1569139307
transform 1 0 1896 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2074
timestamp 1569139307
transform 1 0 2024 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2075
timestamp 1569139307
transform 1 0 2024 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2076
timestamp 1569139307
transform 1 0 2024 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2077
timestamp 1569139307
transform 1 0 1960 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2078
timestamp 1569139307
transform 1 0 2088 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2079
timestamp 1569139307
transform 1 0 2088 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2080
timestamp 1569139307
transform 1 0 2088 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2081
timestamp 1569139307
transform 1 0 1896 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2082
timestamp 1569139307
transform 1 0 1960 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2083
timestamp 1569139307
transform 1 0 2152 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2084
timestamp 1569139307
transform 1 0 2024 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2085
timestamp 1569139307
transform 1 0 2088 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2086
timestamp 1569139307
transform 1 0 2024 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2087
timestamp 1569139307
transform 1 0 1960 0 1 2152
box -8 -8 8 8
use VIA2  VIA2_2088
timestamp 1569139307
transform 1 0 2088 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2089
timestamp 1569139307
transform 1 0 2152 0 1 1896
box -8 -8 8 8
use VIA2  VIA2_2090
timestamp 1569139307
transform 1 0 1896 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2091
timestamp 1569139307
transform 1 0 2152 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2092
timestamp 1569139307
transform 1 0 1896 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2093
timestamp 1569139307
transform 1 0 2152 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2094
timestamp 1569139307
transform 1 0 1896 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2095
timestamp 1569139307
transform 1 0 2152 0 1 2088
box -8 -8 8 8
use VIA2  VIA2_2096
timestamp 1569139307
transform 1 0 1960 0 1 1960
box -8 -8 8 8
use VIA2  VIA2_2097
timestamp 1569139307
transform 1 0 1960 0 1 2024
box -8 -8 8 8
use VIA2  VIA2_2098
timestamp 1569139307
transform 1 0 1896 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2099
timestamp 1569139307
transform 1 0 1896 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2100
timestamp 1569139307
transform 1 0 1896 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2101
timestamp 1569139307
transform 1 0 1896 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2102
timestamp 1569139307
transform 1 0 1896 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2103
timestamp 1569139307
transform 1 0 1960 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2104
timestamp 1569139307
transform 1 0 1960 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2105
timestamp 1569139307
transform 1 0 1960 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2106
timestamp 1569139307
transform 1 0 1960 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2107
timestamp 1569139307
transform 1 0 1960 0 1 2472
box -8 -8 8 8
use VIA2  VIA2_2108
timestamp 1569139307
transform 1 0 2152 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2109
timestamp 1569139307
transform 1 0 2152 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2110
timestamp 1569139307
transform 1 0 2024 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2111
timestamp 1569139307
transform 1 0 2024 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2112
timestamp 1569139307
transform 1 0 2024 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2113
timestamp 1569139307
transform 1 0 2024 0 1 2408
box -8 -8 8 8
use VIA2  VIA2_2114
timestamp 1569139307
transform 1 0 2088 0 1 2344
box -8 -8 8 8
use VIA2  VIA2_2115
timestamp 1569139307
transform 1 0 2088 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2116
timestamp 1569139307
transform 1 0 2088 0 1 2280
box -8 -8 8 8
use VIA2  VIA2_2117
timestamp 1569139307
transform 1 0 2216 0 1 2216
box -8 -8 8 8
use VIA2  VIA2_2118
timestamp 1569139307
transform 1 0 1896 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2119
timestamp 1569139307
transform 1 0 1640 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2120
timestamp 1569139307
transform 1 0 1768 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2121
timestamp 1569139307
transform 1 0 1704 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2122
timestamp 1569139307
transform 1 0 1768 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2123
timestamp 1569139307
transform 1 0 1832 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2124
timestamp 1569139307
transform 1 0 1704 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2125
timestamp 1569139307
transform 1 0 1640 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2126
timestamp 1569139307
transform 1 0 1704 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2127
timestamp 1569139307
transform 1 0 1768 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2128
timestamp 1569139307
transform 1 0 1640 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2129
timestamp 1569139307
transform 1 0 1640 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2130
timestamp 1569139307
transform 1 0 1704 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2131
timestamp 1569139307
transform 1 0 1832 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2132
timestamp 1569139307
transform 1 0 1640 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2133
timestamp 1569139307
transform 1 0 1384 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2134
timestamp 1569139307
transform 1 0 1448 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2135
timestamp 1569139307
transform 1 0 1512 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2136
timestamp 1569139307
transform 1 0 1512 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2137
timestamp 1569139307
transform 1 0 1448 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2138
timestamp 1569139307
transform 1 0 1384 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2139
timestamp 1569139307
transform 1 0 1320 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2140
timestamp 1569139307
transform 1 0 1448 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2141
timestamp 1569139307
transform 1 0 1320 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2142
timestamp 1569139307
transform 1 0 1448 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2143
timestamp 1569139307
transform 1 0 1320 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2144
timestamp 1569139307
transform 1 0 1384 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2145
timestamp 1569139307
transform 1 0 1512 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2146
timestamp 1569139307
transform 1 0 1512 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2147
timestamp 1569139307
transform 1 0 1448 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2148
timestamp 1569139307
transform 1 0 1384 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2149
timestamp 1569139307
transform 1 0 1384 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2150
timestamp 1569139307
transform 1 0 1320 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2151
timestamp 1569139307
transform 1 0 1320 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2152
timestamp 1569139307
transform 1 0 1512 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2153
timestamp 1569139307
transform 1 0 1512 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2154
timestamp 1569139307
transform 1 0 1448 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2155
timestamp 1569139307
transform 1 0 1384 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2156
timestamp 1569139307
transform 1 0 1512 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2157
timestamp 1569139307
transform 1 0 1512 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2158
timestamp 1569139307
transform 1 0 1384 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2159
timestamp 1569139307
transform 1 0 1384 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2160
timestamp 1569139307
transform 1 0 1448 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2161
timestamp 1569139307
transform 1 0 1512 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2162
timestamp 1569139307
transform 1 0 1512 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2163
timestamp 1569139307
transform 1 0 1384 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2164
timestamp 1569139307
transform 1 0 1320 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2165
timestamp 1569139307
transform 1 0 1320 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2166
timestamp 1569139307
transform 1 0 1384 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2167
timestamp 1569139307
transform 1 0 1448 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2168
timestamp 1569139307
transform 1 0 1448 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2169
timestamp 1569139307
transform 1 0 1448 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2170
timestamp 1569139307
transform 1 0 1320 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2171
timestamp 1569139307
transform 1 0 1320 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2172
timestamp 1569139307
transform 1 0 1320 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2173
timestamp 1569139307
transform 1 0 1576 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2174
timestamp 1569139307
transform 1 0 1576 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2175
timestamp 1569139307
transform 1 0 1576 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2176
timestamp 1569139307
transform 1 0 1576 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2177
timestamp 1569139307
transform 1 0 1576 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2178
timestamp 1569139307
transform 1 0 1576 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2179
timestamp 1569139307
transform 1 0 1320 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2180
timestamp 1569139307
transform 1 0 1384 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2181
timestamp 1569139307
transform 1 0 1320 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2182
timestamp 1569139307
transform 1 0 1512 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2183
timestamp 1569139307
transform 1 0 1384 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2184
timestamp 1569139307
transform 1 0 1320 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2185
timestamp 1569139307
transform 1 0 1512 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2186
timestamp 1569139307
transform 1 0 1384 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2187
timestamp 1569139307
transform 1 0 1320 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2188
timestamp 1569139307
transform 1 0 1512 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2189
timestamp 1569139307
transform 1 0 1448 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2190
timestamp 1569139307
transform 1 0 1512 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2191
timestamp 1569139307
transform 1 0 1384 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2192
timestamp 1569139307
transform 1 0 1320 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2193
timestamp 1569139307
transform 1 0 1448 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2194
timestamp 1569139307
transform 1 0 1384 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2195
timestamp 1569139307
transform 1 0 1320 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2196
timestamp 1569139307
transform 1 0 1384 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2197
timestamp 1569139307
transform 1 0 1384 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2198
timestamp 1569139307
transform 1 0 1384 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2199
timestamp 1569139307
transform 1 0 1320 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2200
timestamp 1569139307
transform 1 0 1512 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2201
timestamp 1569139307
transform 1 0 1448 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2202
timestamp 1569139307
transform 1 0 1512 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2203
timestamp 1569139307
transform 1 0 1320 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2204
timestamp 1569139307
transform 1 0 1384 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2205
timestamp 1569139307
transform 1 0 1448 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2206
timestamp 1569139307
transform 1 0 1448 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2207
timestamp 1569139307
transform 1 0 1512 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2208
timestamp 1569139307
transform 1 0 1512 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2209
timestamp 1569139307
transform 1 0 1448 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2210
timestamp 1569139307
transform 1 0 1320 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2211
timestamp 1569139307
transform 1 0 1512 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2212
timestamp 1569139307
transform 1 0 1448 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2213
timestamp 1569139307
transform 1 0 1448 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2214
timestamp 1569139307
transform 1 0 1448 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2215
timestamp 1569139307
transform 1 0 2472 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2216
timestamp 1569139307
transform 1 0 2344 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2217
timestamp 1569139307
transform 1 0 2344 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2218
timestamp 1569139307
transform 1 0 2472 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2219
timestamp 1569139307
transform 1 0 2472 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2220
timestamp 1569139307
transform 1 0 2472 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2221
timestamp 1569139307
transform 1 0 2472 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2222
timestamp 1569139307
transform 1 0 2344 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2223
timestamp 1569139307
transform 1 0 2408 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2224
timestamp 1569139307
transform 1 0 2472 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2225
timestamp 1569139307
transform 1 0 2408 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2226
timestamp 1569139307
transform 1 0 2472 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2227
timestamp 1569139307
transform 1 0 2408 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2228
timestamp 1569139307
transform 1 0 2344 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2229
timestamp 1569139307
transform 1 0 2408 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2230
timestamp 1569139307
transform 1 0 2408 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2231
timestamp 1569139307
transform 1 0 2408 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2232
timestamp 1569139307
transform 1 0 2344 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2233
timestamp 1569139307
transform 1 0 2408 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2234
timestamp 1569139307
transform 1 0 2344 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2235
timestamp 1569139307
transform 1 0 2472 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2236
timestamp 1569139307
transform 1 0 1256 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2237
timestamp 1569139307
transform 1 0 1064 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2238
timestamp 1569139307
transform 1 0 1000 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2239
timestamp 1569139307
transform 1 0 1256 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2240
timestamp 1569139307
transform 1 0 1000 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2241
timestamp 1569139307
transform 1 0 1128 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2242
timestamp 1569139307
transform 1 0 1064 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2243
timestamp 1569139307
transform 1 0 1192 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2244
timestamp 1569139307
transform 1 0 1064 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2245
timestamp 1569139307
transform 1 0 1192 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2246
timestamp 1569139307
transform 1 0 1256 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2247
timestamp 1569139307
transform 1 0 1064 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2248
timestamp 1569139307
transform 1 0 1000 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2249
timestamp 1569139307
transform 1 0 1128 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2250
timestamp 1569139307
transform 1 0 1000 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2251
timestamp 1569139307
transform 1 0 1192 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2252
timestamp 1569139307
transform 1 0 1128 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2253
timestamp 1569139307
transform 1 0 1256 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2254
timestamp 1569139307
transform 1 0 1192 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2255
timestamp 1569139307
transform 1 0 1256 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2256
timestamp 1569139307
transform 1 0 1064 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2257
timestamp 1569139307
transform 1 0 1128 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2258
timestamp 1569139307
transform 1 0 1128 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2259
timestamp 1569139307
transform 1 0 1192 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2260
timestamp 1569139307
transform 1 0 1000 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2261
timestamp 1569139307
transform 1 0 680 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2262
timestamp 1569139307
transform 1 0 936 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2263
timestamp 1569139307
transform 1 0 808 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2264
timestamp 1569139307
transform 1 0 680 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2265
timestamp 1569139307
transform 1 0 744 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2266
timestamp 1569139307
transform 1 0 744 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2267
timestamp 1569139307
transform 1 0 744 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2268
timestamp 1569139307
transform 1 0 936 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2269
timestamp 1569139307
transform 1 0 680 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2270
timestamp 1569139307
transform 1 0 808 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2271
timestamp 1569139307
transform 1 0 808 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2272
timestamp 1569139307
transform 1 0 808 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2273
timestamp 1569139307
transform 1 0 872 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2274
timestamp 1569139307
transform 1 0 872 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2275
timestamp 1569139307
transform 1 0 936 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2276
timestamp 1569139307
transform 1 0 872 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2277
timestamp 1569139307
transform 1 0 936 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2278
timestamp 1569139307
transform 1 0 680 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2279
timestamp 1569139307
transform 1 0 808 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2280
timestamp 1569139307
transform 1 0 744 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2281
timestamp 1569139307
transform 1 0 680 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2282
timestamp 1569139307
transform 1 0 872 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2283
timestamp 1569139307
transform 1 0 936 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2284
timestamp 1569139307
transform 1 0 744 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2285
timestamp 1569139307
transform 1 0 872 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2286
timestamp 1569139307
transform 1 0 936 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2287
timestamp 1569139307
transform 1 0 808 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2288
timestamp 1569139307
transform 1 0 872 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2289
timestamp 1569139307
transform 1 0 680 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2290
timestamp 1569139307
transform 1 0 872 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2291
timestamp 1569139307
transform 1 0 680 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2292
timestamp 1569139307
transform 1 0 744 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2293
timestamp 1569139307
transform 1 0 744 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2294
timestamp 1569139307
transform 1 0 808 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2295
timestamp 1569139307
transform 1 0 808 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2296
timestamp 1569139307
transform 1 0 936 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2297
timestamp 1569139307
transform 1 0 872 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2298
timestamp 1569139307
transform 1 0 936 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2299
timestamp 1569139307
transform 1 0 808 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2300
timestamp 1569139307
transform 1 0 744 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2301
timestamp 1569139307
transform 1 0 744 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2302
timestamp 1569139307
transform 1 0 808 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2303
timestamp 1569139307
transform 1 0 936 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2304
timestamp 1569139307
transform 1 0 680 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2305
timestamp 1569139307
transform 1 0 680 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2306
timestamp 1569139307
transform 1 0 936 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2307
timestamp 1569139307
transform 1 0 872 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2308
timestamp 1569139307
transform 1 0 744 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2309
timestamp 1569139307
transform 1 0 872 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2310
timestamp 1569139307
transform 1 0 680 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2311
timestamp 1569139307
transform 1 0 1000 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2312
timestamp 1569139307
transform 1 0 1128 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2313
timestamp 1569139307
transform 1 0 1192 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2314
timestamp 1569139307
transform 1 0 1000 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2315
timestamp 1569139307
transform 1 0 1000 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2316
timestamp 1569139307
transform 1 0 1064 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2317
timestamp 1569139307
transform 1 0 1256 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2318
timestamp 1569139307
transform 1 0 1256 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2319
timestamp 1569139307
transform 1 0 1128 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2320
timestamp 1569139307
transform 1 0 1256 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2321
timestamp 1569139307
transform 1 0 1000 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2322
timestamp 1569139307
transform 1 0 1256 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2323
timestamp 1569139307
transform 1 0 1000 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2324
timestamp 1569139307
transform 1 0 1064 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2325
timestamp 1569139307
transform 1 0 1192 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2326
timestamp 1569139307
transform 1 0 1192 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2327
timestamp 1569139307
transform 1 0 1128 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2328
timestamp 1569139307
transform 1 0 1064 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2329
timestamp 1569139307
transform 1 0 1128 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2330
timestamp 1569139307
transform 1 0 1192 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2331
timestamp 1569139307
transform 1 0 1192 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2332
timestamp 1569139307
transform 1 0 1064 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2333
timestamp 1569139307
transform 1 0 1064 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2334
timestamp 1569139307
transform 1 0 1256 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2335
timestamp 1569139307
transform 1 0 1128 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2336
timestamp 1569139307
transform 1 0 488 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2337
timestamp 1569139307
transform 1 0 616 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2338
timestamp 1569139307
transform 1 0 552 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2339
timestamp 1569139307
transform 1 0 616 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2340
timestamp 1569139307
transform 1 0 616 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2341
timestamp 1569139307
transform 1 0 552 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2342
timestamp 1569139307
transform 1 0 488 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2343
timestamp 1569139307
transform 1 0 616 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2344
timestamp 1569139307
transform 1 0 552 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2345
timestamp 1569139307
transform 1 0 552 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2346
timestamp 1569139307
transform 1 0 488 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2347
timestamp 1569139307
transform 1 0 360 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2348
timestamp 1569139307
transform 1 0 424 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2349
timestamp 1569139307
transform 1 0 360 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2350
timestamp 1569139307
transform 1 0 488 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2351
timestamp 1569139307
transform 1 0 552 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2352
timestamp 1569139307
transform 1 0 424 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2353
timestamp 1569139307
transform 1 0 424 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2354
timestamp 1569139307
transform 1 0 360 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2355
timestamp 1569139307
transform 1 0 488 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2356
timestamp 1569139307
transform 1 0 424 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2357
timestamp 1569139307
transform 1 0 360 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2358
timestamp 1569139307
transform 1 0 616 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2359
timestamp 1569139307
transform 1 0 424 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2360
timestamp 1569139307
transform 1 0 360 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2361
timestamp 1569139307
transform 1 0 232 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2362
timestamp 1569139307
transform 1 0 232 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2363
timestamp 1569139307
transform 1 0 296 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2364
timestamp 1569139307
transform 1 0 296 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2365
timestamp 1569139307
transform 1 0 104 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2366
timestamp 1569139307
transform 1 0 232 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2367
timestamp 1569139307
transform 1 0 168 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2368
timestamp 1569139307
transform 1 0 104 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2369
timestamp 1569139307
transform 1 0 296 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2370
timestamp 1569139307
transform 1 0 104 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2371
timestamp 1569139307
transform 1 0 40 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2372
timestamp 1569139307
transform 1 0 232 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2373
timestamp 1569139307
transform 1 0 40 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2374
timestamp 1569139307
transform 1 0 104 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2375
timestamp 1569139307
transform 1 0 168 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2376
timestamp 1569139307
transform 1 0 168 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2377
timestamp 1569139307
transform 1 0 40 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2378
timestamp 1569139307
transform 1 0 296 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2379
timestamp 1569139307
transform 1 0 168 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2380
timestamp 1569139307
transform 1 0 40 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_2381
timestamp 1569139307
transform 1 0 296 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2382
timestamp 1569139307
transform 1 0 104 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_2383
timestamp 1569139307
transform 1 0 40 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_2384
timestamp 1569139307
transform 1 0 232 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_2385
timestamp 1569139307
transform 1 0 168 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_2386
timestamp 1569139307
transform 1 0 232 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2387
timestamp 1569139307
transform 1 0 168 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2388
timestamp 1569139307
transform 1 0 232 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2389
timestamp 1569139307
transform 1 0 232 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2390
timestamp 1569139307
transform 1 0 232 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2391
timestamp 1569139307
transform 1 0 168 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2392
timestamp 1569139307
transform 1 0 40 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2393
timestamp 1569139307
transform 1 0 40 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2394
timestamp 1569139307
transform 1 0 296 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2395
timestamp 1569139307
transform 1 0 232 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2396
timestamp 1569139307
transform 1 0 296 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2397
timestamp 1569139307
transform 1 0 40 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2398
timestamp 1569139307
transform 1 0 168 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2399
timestamp 1569139307
transform 1 0 104 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2400
timestamp 1569139307
transform 1 0 168 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2401
timestamp 1569139307
transform 1 0 104 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2402
timestamp 1569139307
transform 1 0 104 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2403
timestamp 1569139307
transform 1 0 40 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2404
timestamp 1569139307
transform 1 0 296 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2405
timestamp 1569139307
transform 1 0 296 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2406
timestamp 1569139307
transform 1 0 296 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2407
timestamp 1569139307
transform 1 0 104 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2408
timestamp 1569139307
transform 1 0 40 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2409
timestamp 1569139307
transform 1 0 104 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2410
timestamp 1569139307
transform 1 0 168 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2411
timestamp 1569139307
transform 1 0 616 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2412
timestamp 1569139307
transform 1 0 360 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2413
timestamp 1569139307
transform 1 0 616 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2414
timestamp 1569139307
transform 1 0 616 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2415
timestamp 1569139307
transform 1 0 488 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2416
timestamp 1569139307
transform 1 0 616 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2417
timestamp 1569139307
transform 1 0 360 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2418
timestamp 1569139307
transform 1 0 616 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2419
timestamp 1569139307
transform 1 0 488 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2420
timestamp 1569139307
transform 1 0 360 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2421
timestamp 1569139307
transform 1 0 424 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2422
timestamp 1569139307
transform 1 0 552 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2423
timestamp 1569139307
transform 1 0 488 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2424
timestamp 1569139307
transform 1 0 360 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2425
timestamp 1569139307
transform 1 0 424 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2426
timestamp 1569139307
transform 1 0 488 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2427
timestamp 1569139307
transform 1 0 552 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2428
timestamp 1569139307
transform 1 0 488 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2429
timestamp 1569139307
transform 1 0 424 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2430
timestamp 1569139307
transform 1 0 424 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2431
timestamp 1569139307
transform 1 0 552 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_2432
timestamp 1569139307
transform 1 0 552 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_2433
timestamp 1569139307
transform 1 0 552 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_2434
timestamp 1569139307
transform 1 0 360 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_2435
timestamp 1569139307
transform 1 0 424 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_2436
timestamp 1569139307
transform 1 0 616 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2437
timestamp 1569139307
transform 1 0 552 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2438
timestamp 1569139307
transform 1 0 616 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2439
timestamp 1569139307
transform 1 0 424 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2440
timestamp 1569139307
transform 1 0 360 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2441
timestamp 1569139307
transform 1 0 488 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2442
timestamp 1569139307
transform 1 0 552 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2443
timestamp 1569139307
transform 1 0 360 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2444
timestamp 1569139307
transform 1 0 424 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2445
timestamp 1569139307
transform 1 0 424 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2446
timestamp 1569139307
transform 1 0 488 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2447
timestamp 1569139307
transform 1 0 360 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2448
timestamp 1569139307
transform 1 0 488 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2449
timestamp 1569139307
transform 1 0 552 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2450
timestamp 1569139307
transform 1 0 616 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2451
timestamp 1569139307
transform 1 0 424 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2452
timestamp 1569139307
transform 1 0 616 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2453
timestamp 1569139307
transform 1 0 552 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2454
timestamp 1569139307
transform 1 0 488 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2455
timestamp 1569139307
transform 1 0 360 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2456
timestamp 1569139307
transform 1 0 232 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2457
timestamp 1569139307
transform 1 0 104 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2458
timestamp 1569139307
transform 1 0 168 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2459
timestamp 1569139307
transform 1 0 40 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2460
timestamp 1569139307
transform 1 0 168 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2461
timestamp 1569139307
transform 1 0 296 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2462
timestamp 1569139307
transform 1 0 40 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2463
timestamp 1569139307
transform 1 0 232 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2464
timestamp 1569139307
transform 1 0 40 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2465
timestamp 1569139307
transform 1 0 40 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2466
timestamp 1569139307
transform 1 0 104 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2467
timestamp 1569139307
transform 1 0 296 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2468
timestamp 1569139307
transform 1 0 232 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2469
timestamp 1569139307
transform 1 0 168 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2470
timestamp 1569139307
transform 1 0 296 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2471
timestamp 1569139307
transform 1 0 104 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2472
timestamp 1569139307
transform 1 0 296 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2473
timestamp 1569139307
transform 1 0 168 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2474
timestamp 1569139307
transform 1 0 232 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2475
timestamp 1569139307
transform 1 0 104 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2476
timestamp 1569139307
transform 1 0 296 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2477
timestamp 1569139307
transform 1 0 232 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2478
timestamp 1569139307
transform 1 0 40 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2479
timestamp 1569139307
transform 1 0 104 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2480
timestamp 1569139307
transform 1 0 232 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2481
timestamp 1569139307
transform 1 0 168 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2482
timestamp 1569139307
transform 1 0 104 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2483
timestamp 1569139307
transform 1 0 168 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2484
timestamp 1569139307
transform 1 0 232 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2485
timestamp 1569139307
transform 1 0 296 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2486
timestamp 1569139307
transform 1 0 168 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2487
timestamp 1569139307
transform 1 0 104 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2488
timestamp 1569139307
transform 1 0 296 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2489
timestamp 1569139307
transform 1 0 296 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2490
timestamp 1569139307
transform 1 0 40 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2491
timestamp 1569139307
transform 1 0 40 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2492
timestamp 1569139307
transform 1 0 40 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2493
timestamp 1569139307
transform 1 0 168 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2494
timestamp 1569139307
transform 1 0 232 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2495
timestamp 1569139307
transform 1 0 104 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2496
timestamp 1569139307
transform 1 0 552 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2497
timestamp 1569139307
transform 1 0 360 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2498
timestamp 1569139307
transform 1 0 552 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2499
timestamp 1569139307
transform 1 0 616 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2500
timestamp 1569139307
transform 1 0 424 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2501
timestamp 1569139307
transform 1 0 488 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2502
timestamp 1569139307
transform 1 0 424 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2503
timestamp 1569139307
transform 1 0 616 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2504
timestamp 1569139307
transform 1 0 488 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2505
timestamp 1569139307
transform 1 0 424 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2506
timestamp 1569139307
transform 1 0 616 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2507
timestamp 1569139307
transform 1 0 488 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2508
timestamp 1569139307
transform 1 0 616 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2509
timestamp 1569139307
transform 1 0 552 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2510
timestamp 1569139307
transform 1 0 360 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2511
timestamp 1569139307
transform 1 0 552 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2512
timestamp 1569139307
transform 1 0 360 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2513
timestamp 1569139307
transform 1 0 424 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2514
timestamp 1569139307
transform 1 0 488 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2515
timestamp 1569139307
transform 1 0 360 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2516
timestamp 1569139307
transform 1 0 424 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2517
timestamp 1569139307
transform 1 0 40 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2518
timestamp 1569139307
transform 1 0 296 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2519
timestamp 1569139307
transform 1 0 168 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2520
timestamp 1569139307
transform 1 0 616 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2521
timestamp 1569139307
transform 1 0 488 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2522
timestamp 1569139307
transform 1 0 360 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2523
timestamp 1569139307
transform 1 0 232 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2524
timestamp 1569139307
transform 1 0 104 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2525
timestamp 1569139307
transform 1 0 552 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2526
timestamp 1569139307
transform 1 0 1064 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2527
timestamp 1569139307
transform 1 0 1128 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2528
timestamp 1569139307
transform 1 0 1192 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2529
timestamp 1569139307
transform 1 0 1064 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2530
timestamp 1569139307
transform 1 0 1192 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2531
timestamp 1569139307
transform 1 0 1256 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2532
timestamp 1569139307
transform 1 0 1000 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2533
timestamp 1569139307
transform 1 0 1256 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2534
timestamp 1569139307
transform 1 0 1256 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2535
timestamp 1569139307
transform 1 0 1192 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2536
timestamp 1569139307
transform 1 0 1000 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2537
timestamp 1569139307
transform 1 0 1128 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2538
timestamp 1569139307
transform 1 0 1000 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2539
timestamp 1569139307
transform 1 0 1192 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2540
timestamp 1569139307
transform 1 0 1256 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2541
timestamp 1569139307
transform 1 0 1064 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2542
timestamp 1569139307
transform 1 0 1128 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2543
timestamp 1569139307
transform 1 0 1000 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2544
timestamp 1569139307
transform 1 0 1064 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2545
timestamp 1569139307
transform 1 0 1128 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2546
timestamp 1569139307
transform 1 0 872 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2547
timestamp 1569139307
transform 1 0 680 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2548
timestamp 1569139307
transform 1 0 808 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2549
timestamp 1569139307
transform 1 0 808 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2550
timestamp 1569139307
transform 1 0 936 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2551
timestamp 1569139307
transform 1 0 680 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2552
timestamp 1569139307
transform 1 0 872 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2553
timestamp 1569139307
transform 1 0 744 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2554
timestamp 1569139307
transform 1 0 744 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2555
timestamp 1569139307
transform 1 0 872 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2556
timestamp 1569139307
transform 1 0 872 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2557
timestamp 1569139307
transform 1 0 680 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2558
timestamp 1569139307
transform 1 0 808 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2559
timestamp 1569139307
transform 1 0 744 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_2560
timestamp 1569139307
transform 1 0 936 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_2561
timestamp 1569139307
transform 1 0 936 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2562
timestamp 1569139307
transform 1 0 808 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2563
timestamp 1569139307
transform 1 0 744 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_2564
timestamp 1569139307
transform 1 0 936 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2565
timestamp 1569139307
transform 1 0 680 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_2566
timestamp 1569139307
transform 1 0 680 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2567
timestamp 1569139307
transform 1 0 680 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2568
timestamp 1569139307
transform 1 0 744 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2569
timestamp 1569139307
transform 1 0 808 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2570
timestamp 1569139307
transform 1 0 744 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2571
timestamp 1569139307
transform 1 0 808 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2572
timestamp 1569139307
transform 1 0 936 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2573
timestamp 1569139307
transform 1 0 808 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2574
timestamp 1569139307
transform 1 0 872 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2575
timestamp 1569139307
transform 1 0 936 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2576
timestamp 1569139307
transform 1 0 808 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2577
timestamp 1569139307
transform 1 0 872 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2578
timestamp 1569139307
transform 1 0 936 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2579
timestamp 1569139307
transform 1 0 936 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2580
timestamp 1569139307
transform 1 0 680 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2581
timestamp 1569139307
transform 1 0 680 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2582
timestamp 1569139307
transform 1 0 872 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2583
timestamp 1569139307
transform 1 0 744 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2584
timestamp 1569139307
transform 1 0 872 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2585
timestamp 1569139307
transform 1 0 744 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2586
timestamp 1569139307
transform 1 0 1064 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2587
timestamp 1569139307
transform 1 0 1192 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2588
timestamp 1569139307
transform 1 0 1064 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2589
timestamp 1569139307
transform 1 0 1128 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2590
timestamp 1569139307
transform 1 0 1000 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2591
timestamp 1569139307
transform 1 0 1256 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2592
timestamp 1569139307
transform 1 0 1256 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2593
timestamp 1569139307
transform 1 0 1000 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2594
timestamp 1569139307
transform 1 0 1064 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2595
timestamp 1569139307
transform 1 0 1000 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2596
timestamp 1569139307
transform 1 0 1256 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2597
timestamp 1569139307
transform 1 0 1192 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2598
timestamp 1569139307
transform 1 0 1064 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2599
timestamp 1569139307
transform 1 0 1256 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2600
timestamp 1569139307
transform 1 0 1128 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2601
timestamp 1569139307
transform 1 0 1192 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2602
timestamp 1569139307
transform 1 0 1192 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_2603
timestamp 1569139307
transform 1 0 1128 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_2604
timestamp 1569139307
transform 1 0 1000 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_2605
timestamp 1569139307
transform 1 0 1128 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_2606
timestamp 1569139307
transform 1 0 872 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2607
timestamp 1569139307
transform 1 0 1256 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2608
timestamp 1569139307
transform 1 0 1000 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2609
timestamp 1569139307
transform 1 0 680 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2610
timestamp 1569139307
transform 1 0 1192 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2611
timestamp 1569139307
transform 1 0 744 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2612
timestamp 1569139307
transform 1 0 808 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2613
timestamp 1569139307
transform 1 0 1064 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2614
timestamp 1569139307
transform 1 0 1128 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2615
timestamp 1569139307
transform 1 0 936 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_2616
timestamp 1569139307
transform 1 0 1192 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2617
timestamp 1569139307
transform 1 0 1000 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2618
timestamp 1569139307
transform 1 0 1256 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2619
timestamp 1569139307
transform 1 0 1128 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2620
timestamp 1569139307
transform 1 0 1064 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2621
timestamp 1569139307
transform 1 0 1192 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2622
timestamp 1569139307
transform 1 0 1000 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2623
timestamp 1569139307
transform 1 0 1000 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2624
timestamp 1569139307
transform 1 0 1128 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2625
timestamp 1569139307
transform 1 0 1192 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2626
timestamp 1569139307
transform 1 0 1256 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2627
timestamp 1569139307
transform 1 0 1064 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2628
timestamp 1569139307
transform 1 0 1256 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2629
timestamp 1569139307
transform 1 0 1064 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2630
timestamp 1569139307
transform 1 0 1192 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2631
timestamp 1569139307
transform 1 0 1064 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2632
timestamp 1569139307
transform 1 0 1256 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2633
timestamp 1569139307
transform 1 0 1000 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2634
timestamp 1569139307
transform 1 0 1128 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2635
timestamp 1569139307
transform 1 0 1000 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2636
timestamp 1569139307
transform 1 0 1256 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2637
timestamp 1569139307
transform 1 0 1064 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2638
timestamp 1569139307
transform 1 0 1128 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2639
timestamp 1569139307
transform 1 0 1192 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2640
timestamp 1569139307
transform 1 0 1128 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2641
timestamp 1569139307
transform 1 0 744 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2642
timestamp 1569139307
transform 1 0 936 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2643
timestamp 1569139307
transform 1 0 936 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2644
timestamp 1569139307
transform 1 0 936 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2645
timestamp 1569139307
transform 1 0 872 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2646
timestamp 1569139307
transform 1 0 680 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2647
timestamp 1569139307
transform 1 0 936 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2648
timestamp 1569139307
transform 1 0 872 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2649
timestamp 1569139307
transform 1 0 744 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2650
timestamp 1569139307
transform 1 0 808 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2651
timestamp 1569139307
transform 1 0 744 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2652
timestamp 1569139307
transform 1 0 872 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2653
timestamp 1569139307
transform 1 0 808 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2654
timestamp 1569139307
transform 1 0 744 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2655
timestamp 1569139307
transform 1 0 680 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2656
timestamp 1569139307
transform 1 0 680 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2657
timestamp 1569139307
transform 1 0 808 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2658
timestamp 1569139307
transform 1 0 680 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2659
timestamp 1569139307
transform 1 0 936 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2660
timestamp 1569139307
transform 1 0 872 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2661
timestamp 1569139307
transform 1 0 808 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2662
timestamp 1569139307
transform 1 0 744 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2663
timestamp 1569139307
transform 1 0 808 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2664
timestamp 1569139307
transform 1 0 872 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2665
timestamp 1569139307
transform 1 0 680 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2666
timestamp 1569139307
transform 1 0 744 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2667
timestamp 1569139307
transform 1 0 936 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2668
timestamp 1569139307
transform 1 0 872 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2669
timestamp 1569139307
transform 1 0 936 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2670
timestamp 1569139307
transform 1 0 808 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2671
timestamp 1569139307
transform 1 0 808 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2672
timestamp 1569139307
transform 1 0 872 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2673
timestamp 1569139307
transform 1 0 872 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2674
timestamp 1569139307
transform 1 0 808 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2675
timestamp 1569139307
transform 1 0 936 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2676
timestamp 1569139307
transform 1 0 680 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2677
timestamp 1569139307
transform 1 0 872 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2678
timestamp 1569139307
transform 1 0 680 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2679
timestamp 1569139307
transform 1 0 744 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2680
timestamp 1569139307
transform 1 0 680 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2681
timestamp 1569139307
transform 1 0 872 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2682
timestamp 1569139307
transform 1 0 680 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2683
timestamp 1569139307
transform 1 0 744 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2684
timestamp 1569139307
transform 1 0 808 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2685
timestamp 1569139307
transform 1 0 936 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2686
timestamp 1569139307
transform 1 0 936 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2687
timestamp 1569139307
transform 1 0 744 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2688
timestamp 1569139307
transform 1 0 744 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2689
timestamp 1569139307
transform 1 0 808 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2690
timestamp 1569139307
transform 1 0 680 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2691
timestamp 1569139307
transform 1 0 1128 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2692
timestamp 1569139307
transform 1 0 1000 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2693
timestamp 1569139307
transform 1 0 1256 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2694
timestamp 1569139307
transform 1 0 1256 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2695
timestamp 1569139307
transform 1 0 1256 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2696
timestamp 1569139307
transform 1 0 1256 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2697
timestamp 1569139307
transform 1 0 1192 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2698
timestamp 1569139307
transform 1 0 1128 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2699
timestamp 1569139307
transform 1 0 1000 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2700
timestamp 1569139307
transform 1 0 1192 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2701
timestamp 1569139307
transform 1 0 1000 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2702
timestamp 1569139307
transform 1 0 1064 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2703
timestamp 1569139307
transform 1 0 1192 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2704
timestamp 1569139307
transform 1 0 1000 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2705
timestamp 1569139307
transform 1 0 1000 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2706
timestamp 1569139307
transform 1 0 1192 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2707
timestamp 1569139307
transform 1 0 1064 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2708
timestamp 1569139307
transform 1 0 1064 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2709
timestamp 1569139307
transform 1 0 1064 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2710
timestamp 1569139307
transform 1 0 1128 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2711
timestamp 1569139307
transform 1 0 1256 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2712
timestamp 1569139307
transform 1 0 1128 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2713
timestamp 1569139307
transform 1 0 1128 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2714
timestamp 1569139307
transform 1 0 1192 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2715
timestamp 1569139307
transform 1 0 1064 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2716
timestamp 1569139307
transform 1 0 424 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2717
timestamp 1569139307
transform 1 0 424 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2718
timestamp 1569139307
transform 1 0 488 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2719
timestamp 1569139307
transform 1 0 616 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2720
timestamp 1569139307
transform 1 0 552 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2721
timestamp 1569139307
transform 1 0 360 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2722
timestamp 1569139307
transform 1 0 488 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2723
timestamp 1569139307
transform 1 0 360 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2724
timestamp 1569139307
transform 1 0 424 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2725
timestamp 1569139307
transform 1 0 488 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2726
timestamp 1569139307
transform 1 0 424 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2727
timestamp 1569139307
transform 1 0 616 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2728
timestamp 1569139307
transform 1 0 488 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2729
timestamp 1569139307
transform 1 0 616 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2730
timestamp 1569139307
transform 1 0 552 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2731
timestamp 1569139307
transform 1 0 360 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2732
timestamp 1569139307
transform 1 0 360 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2733
timestamp 1569139307
transform 1 0 616 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2734
timestamp 1569139307
transform 1 0 552 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2735
timestamp 1569139307
transform 1 0 424 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2736
timestamp 1569139307
transform 1 0 552 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2737
timestamp 1569139307
transform 1 0 616 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2738
timestamp 1569139307
transform 1 0 552 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2739
timestamp 1569139307
transform 1 0 360 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2740
timestamp 1569139307
transform 1 0 488 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2741
timestamp 1569139307
transform 1 0 104 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2742
timestamp 1569139307
transform 1 0 104 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2743
timestamp 1569139307
transform 1 0 40 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2744
timestamp 1569139307
transform 1 0 232 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2745
timestamp 1569139307
transform 1 0 232 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2746
timestamp 1569139307
transform 1 0 40 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2747
timestamp 1569139307
transform 1 0 40 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2748
timestamp 1569139307
transform 1 0 40 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2749
timestamp 1569139307
transform 1 0 104 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2750
timestamp 1569139307
transform 1 0 168 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2751
timestamp 1569139307
transform 1 0 232 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2752
timestamp 1569139307
transform 1 0 296 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_2753
timestamp 1569139307
transform 1 0 232 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2754
timestamp 1569139307
transform 1 0 104 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2755
timestamp 1569139307
transform 1 0 40 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2756
timestamp 1569139307
transform 1 0 168 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2757
timestamp 1569139307
transform 1 0 296 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2758
timestamp 1569139307
transform 1 0 168 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2759
timestamp 1569139307
transform 1 0 232 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2760
timestamp 1569139307
transform 1 0 296 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2761
timestamp 1569139307
transform 1 0 168 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_2762
timestamp 1569139307
transform 1 0 168 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2763
timestamp 1569139307
transform 1 0 296 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2764
timestamp 1569139307
transform 1 0 104 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_2765
timestamp 1569139307
transform 1 0 296 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_2766
timestamp 1569139307
transform 1 0 232 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2767
timestamp 1569139307
transform 1 0 168 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2768
timestamp 1569139307
transform 1 0 168 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2769
timestamp 1569139307
transform 1 0 232 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2770
timestamp 1569139307
transform 1 0 104 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2771
timestamp 1569139307
transform 1 0 232 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2772
timestamp 1569139307
transform 1 0 168 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2773
timestamp 1569139307
transform 1 0 296 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2774
timestamp 1569139307
transform 1 0 104 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2775
timestamp 1569139307
transform 1 0 40 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2776
timestamp 1569139307
transform 1 0 296 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2777
timestamp 1569139307
transform 1 0 296 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2778
timestamp 1569139307
transform 1 0 296 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2779
timestamp 1569139307
transform 1 0 104 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2780
timestamp 1569139307
transform 1 0 232 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2781
timestamp 1569139307
transform 1 0 40 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2782
timestamp 1569139307
transform 1 0 40 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2783
timestamp 1569139307
transform 1 0 40 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2784
timestamp 1569139307
transform 1 0 168 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2785
timestamp 1569139307
transform 1 0 232 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2786
timestamp 1569139307
transform 1 0 104 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2787
timestamp 1569139307
transform 1 0 104 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2788
timestamp 1569139307
transform 1 0 296 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2789
timestamp 1569139307
transform 1 0 40 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2790
timestamp 1569139307
transform 1 0 168 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2791
timestamp 1569139307
transform 1 0 616 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2792
timestamp 1569139307
transform 1 0 616 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2793
timestamp 1569139307
transform 1 0 424 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2794
timestamp 1569139307
transform 1 0 488 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2795
timestamp 1569139307
transform 1 0 488 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2796
timestamp 1569139307
transform 1 0 424 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2797
timestamp 1569139307
transform 1 0 424 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2798
timestamp 1569139307
transform 1 0 552 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2799
timestamp 1569139307
transform 1 0 360 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2800
timestamp 1569139307
transform 1 0 424 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2801
timestamp 1569139307
transform 1 0 552 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2802
timestamp 1569139307
transform 1 0 360 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2803
timestamp 1569139307
transform 1 0 552 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2804
timestamp 1569139307
transform 1 0 360 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2805
timestamp 1569139307
transform 1 0 360 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2806
timestamp 1569139307
transform 1 0 552 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2807
timestamp 1569139307
transform 1 0 616 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2808
timestamp 1569139307
transform 1 0 616 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2809
timestamp 1569139307
transform 1 0 616 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_2810
timestamp 1569139307
transform 1 0 360 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2811
timestamp 1569139307
transform 1 0 424 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_2812
timestamp 1569139307
transform 1 0 488 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2813
timestamp 1569139307
transform 1 0 488 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2814
timestamp 1569139307
transform 1 0 552 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_2815
timestamp 1569139307
transform 1 0 488 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2816
timestamp 1569139307
transform 1 0 424 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2817
timestamp 1569139307
transform 1 0 424 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2818
timestamp 1569139307
transform 1 0 360 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2819
timestamp 1569139307
transform 1 0 616 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2820
timestamp 1569139307
transform 1 0 488 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2821
timestamp 1569139307
transform 1 0 488 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2822
timestamp 1569139307
transform 1 0 424 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2823
timestamp 1569139307
transform 1 0 360 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2824
timestamp 1569139307
transform 1 0 488 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2825
timestamp 1569139307
transform 1 0 552 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2826
timestamp 1569139307
transform 1 0 552 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2827
timestamp 1569139307
transform 1 0 360 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2828
timestamp 1569139307
transform 1 0 616 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2829
timestamp 1569139307
transform 1 0 616 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2830
timestamp 1569139307
transform 1 0 488 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2831
timestamp 1569139307
transform 1 0 360 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2832
timestamp 1569139307
transform 1 0 360 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2833
timestamp 1569139307
transform 1 0 424 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2834
timestamp 1569139307
transform 1 0 616 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2835
timestamp 1569139307
transform 1 0 552 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2836
timestamp 1569139307
transform 1 0 488 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2837
timestamp 1569139307
transform 1 0 552 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2838
timestamp 1569139307
transform 1 0 424 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2839
timestamp 1569139307
transform 1 0 616 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2840
timestamp 1569139307
transform 1 0 552 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2841
timestamp 1569139307
transform 1 0 40 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2842
timestamp 1569139307
transform 1 0 232 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2843
timestamp 1569139307
transform 1 0 104 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2844
timestamp 1569139307
transform 1 0 232 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2845
timestamp 1569139307
transform 1 0 232 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2846
timestamp 1569139307
transform 1 0 168 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2847
timestamp 1569139307
transform 1 0 296 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2848
timestamp 1569139307
transform 1 0 296 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2849
timestamp 1569139307
transform 1 0 232 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2850
timestamp 1569139307
transform 1 0 40 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2851
timestamp 1569139307
transform 1 0 296 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2852
timestamp 1569139307
transform 1 0 104 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2853
timestamp 1569139307
transform 1 0 296 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2854
timestamp 1569139307
transform 1 0 296 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2855
timestamp 1569139307
transform 1 0 104 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2856
timestamp 1569139307
transform 1 0 232 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2857
timestamp 1569139307
transform 1 0 104 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2858
timestamp 1569139307
transform 1 0 168 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2859
timestamp 1569139307
transform 1 0 104 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2860
timestamp 1569139307
transform 1 0 168 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2861
timestamp 1569139307
transform 1 0 40 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2862
timestamp 1569139307
transform 1 0 168 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2863
timestamp 1569139307
transform 1 0 40 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2864
timestamp 1569139307
transform 1 0 40 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2865
timestamp 1569139307
transform 1 0 168 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2866
timestamp 1569139307
transform 1 0 40 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2867
timestamp 1569139307
transform 1 0 232 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2868
timestamp 1569139307
transform 1 0 296 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2869
timestamp 1569139307
transform 1 0 232 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2870
timestamp 1569139307
transform 1 0 168 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2871
timestamp 1569139307
transform 1 0 168 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2872
timestamp 1569139307
transform 1 0 104 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2873
timestamp 1569139307
transform 1 0 232 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2874
timestamp 1569139307
transform 1 0 296 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2875
timestamp 1569139307
transform 1 0 296 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2876
timestamp 1569139307
transform 1 0 104 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2877
timestamp 1569139307
transform 1 0 296 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2878
timestamp 1569139307
transform 1 0 104 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2879
timestamp 1569139307
transform 1 0 232 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2880
timestamp 1569139307
transform 1 0 168 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2881
timestamp 1569139307
transform 1 0 168 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2882
timestamp 1569139307
transform 1 0 40 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2883
timestamp 1569139307
transform 1 0 40 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2884
timestamp 1569139307
transform 1 0 40 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2885
timestamp 1569139307
transform 1 0 104 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2886
timestamp 1569139307
transform 1 0 552 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2887
timestamp 1569139307
transform 1 0 424 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2888
timestamp 1569139307
transform 1 0 488 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2889
timestamp 1569139307
transform 1 0 424 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2890
timestamp 1569139307
transform 1 0 552 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2891
timestamp 1569139307
transform 1 0 360 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2892
timestamp 1569139307
transform 1 0 616 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2893
timestamp 1569139307
transform 1 0 616 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2894
timestamp 1569139307
transform 1 0 552 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2895
timestamp 1569139307
transform 1 0 616 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2896
timestamp 1569139307
transform 1 0 616 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2897
timestamp 1569139307
transform 1 0 488 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2898
timestamp 1569139307
transform 1 0 424 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2899
timestamp 1569139307
transform 1 0 488 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2900
timestamp 1569139307
transform 1 0 360 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2901
timestamp 1569139307
transform 1 0 360 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2902
timestamp 1569139307
transform 1 0 552 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2903
timestamp 1569139307
transform 1 0 424 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2904
timestamp 1569139307
transform 1 0 488 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2905
timestamp 1569139307
transform 1 0 360 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2906
timestamp 1569139307
transform 1 0 1128 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2907
timestamp 1569139307
transform 1 0 1000 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2908
timestamp 1569139307
transform 1 0 1256 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2909
timestamp 1569139307
transform 1 0 1064 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2910
timestamp 1569139307
transform 1 0 1192 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2911
timestamp 1569139307
transform 1 0 1192 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2912
timestamp 1569139307
transform 1 0 1192 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2913
timestamp 1569139307
transform 1 0 1256 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2914
timestamp 1569139307
transform 1 0 1256 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2915
timestamp 1569139307
transform 1 0 1256 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2916
timestamp 1569139307
transform 1 0 1256 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2917
timestamp 1569139307
transform 1 0 1064 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2918
timestamp 1569139307
transform 1 0 1064 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2919
timestamp 1569139307
transform 1 0 1192 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2920
timestamp 1569139307
transform 1 0 1000 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2921
timestamp 1569139307
transform 1 0 1064 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2922
timestamp 1569139307
transform 1 0 1128 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2923
timestamp 1569139307
transform 1 0 1000 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2924
timestamp 1569139307
transform 1 0 1000 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2925
timestamp 1569139307
transform 1 0 1128 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2926
timestamp 1569139307
transform 1 0 1128 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2927
timestamp 1569139307
transform 1 0 1128 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2928
timestamp 1569139307
transform 1 0 1064 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2929
timestamp 1569139307
transform 1 0 1000 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2930
timestamp 1569139307
transform 1 0 1192 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2931
timestamp 1569139307
transform 1 0 936 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2932
timestamp 1569139307
transform 1 0 808 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2933
timestamp 1569139307
transform 1 0 936 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2934
timestamp 1569139307
transform 1 0 808 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2935
timestamp 1569139307
transform 1 0 872 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2936
timestamp 1569139307
transform 1 0 936 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2937
timestamp 1569139307
transform 1 0 872 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2938
timestamp 1569139307
transform 1 0 872 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2939
timestamp 1569139307
transform 1 0 680 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2940
timestamp 1569139307
transform 1 0 680 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2941
timestamp 1569139307
transform 1 0 680 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2942
timestamp 1569139307
transform 1 0 872 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2943
timestamp 1569139307
transform 1 0 680 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2944
timestamp 1569139307
transform 1 0 680 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2945
timestamp 1569139307
transform 1 0 936 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2946
timestamp 1569139307
transform 1 0 744 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_2947
timestamp 1569139307
transform 1 0 808 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2948
timestamp 1569139307
transform 1 0 744 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2949
timestamp 1569139307
transform 1 0 808 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2950
timestamp 1569139307
transform 1 0 744 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_2951
timestamp 1569139307
transform 1 0 808 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2952
timestamp 1569139307
transform 1 0 744 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_2953
timestamp 1569139307
transform 1 0 744 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2954
timestamp 1569139307
transform 1 0 872 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_2955
timestamp 1569139307
transform 1 0 936 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_2956
timestamp 1569139307
transform 1 0 808 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2957
timestamp 1569139307
transform 1 0 872 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2958
timestamp 1569139307
transform 1 0 936 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2959
timestamp 1569139307
transform 1 0 808 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2960
timestamp 1569139307
transform 1 0 872 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2961
timestamp 1569139307
transform 1 0 872 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2962
timestamp 1569139307
transform 1 0 680 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2963
timestamp 1569139307
transform 1 0 680 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2964
timestamp 1569139307
transform 1 0 680 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2965
timestamp 1569139307
transform 1 0 680 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2966
timestamp 1569139307
transform 1 0 872 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2967
timestamp 1569139307
transform 1 0 808 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2968
timestamp 1569139307
transform 1 0 936 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2969
timestamp 1569139307
transform 1 0 744 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2970
timestamp 1569139307
transform 1 0 744 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2971
timestamp 1569139307
transform 1 0 744 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2972
timestamp 1569139307
transform 1 0 744 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2973
timestamp 1569139307
transform 1 0 936 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2974
timestamp 1569139307
transform 1 0 808 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2975
timestamp 1569139307
transform 1 0 936 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2976
timestamp 1569139307
transform 1 0 1192 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2977
timestamp 1569139307
transform 1 0 1064 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2978
timestamp 1569139307
transform 1 0 1256 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2979
timestamp 1569139307
transform 1 0 1256 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2980
timestamp 1569139307
transform 1 0 1256 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2981
timestamp 1569139307
transform 1 0 1256 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2982
timestamp 1569139307
transform 1 0 1192 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2983
timestamp 1569139307
transform 1 0 1128 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2984
timestamp 1569139307
transform 1 0 1064 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2985
timestamp 1569139307
transform 1 0 1000 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2986
timestamp 1569139307
transform 1 0 1000 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2987
timestamp 1569139307
transform 1 0 1128 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2988
timestamp 1569139307
transform 1 0 1192 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2989
timestamp 1569139307
transform 1 0 1064 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2990
timestamp 1569139307
transform 1 0 1192 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2991
timestamp 1569139307
transform 1 0 1000 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2992
timestamp 1569139307
transform 1 0 1128 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_2993
timestamp 1569139307
transform 1 0 1064 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_2994
timestamp 1569139307
transform 1 0 1000 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_2995
timestamp 1569139307
transform 1 0 1128 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_2996
timestamp 1569139307
transform 1 0 2344 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_2997
timestamp 1569139307
transform 1 0 2344 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_2998
timestamp 1569139307
transform 1 0 2344 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_2999
timestamp 1569139307
transform 1 0 2408 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3000
timestamp 1569139307
transform 1 0 2408 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3001
timestamp 1569139307
transform 1 0 2408 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3002
timestamp 1569139307
transform 1 0 2344 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3003
timestamp 1569139307
transform 1 0 2408 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3004
timestamp 1569139307
transform 1 0 2408 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3005
timestamp 1569139307
transform 1 0 2408 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3006
timestamp 1569139307
transform 1 0 2408 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3007
timestamp 1569139307
transform 1 0 2344 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3008
timestamp 1569139307
transform 1 0 2408 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3009
timestamp 1569139307
transform 1 0 2472 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3010
timestamp 1569139307
transform 1 0 2472 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3011
timestamp 1569139307
transform 1 0 2472 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3012
timestamp 1569139307
transform 1 0 2344 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3013
timestamp 1569139307
transform 1 0 2472 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3014
timestamp 1569139307
transform 1 0 2472 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3015
timestamp 1569139307
transform 1 0 2472 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3016
timestamp 1569139307
transform 1 0 2344 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3017
timestamp 1569139307
transform 1 0 2472 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3018
timestamp 1569139307
transform 1 0 2472 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3019
timestamp 1569139307
transform 1 0 2472 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3020
timestamp 1569139307
transform 1 0 2408 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3021
timestamp 1569139307
transform 1 0 2472 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3022
timestamp 1569139307
transform 1 0 2344 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3023
timestamp 1569139307
transform 1 0 2344 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3024
timestamp 1569139307
transform 1 0 2408 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3025
timestamp 1569139307
transform 1 0 2344 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3026
timestamp 1569139307
transform 1 0 1384 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3027
timestamp 1569139307
transform 1 0 1384 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3028
timestamp 1569139307
transform 1 0 1384 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3029
timestamp 1569139307
transform 1 0 1384 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3030
timestamp 1569139307
transform 1 0 1320 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3031
timestamp 1569139307
transform 1 0 1320 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3032
timestamp 1569139307
transform 1 0 1448 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3033
timestamp 1569139307
transform 1 0 1384 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3034
timestamp 1569139307
transform 1 0 1384 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3035
timestamp 1569139307
transform 1 0 1448 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3036
timestamp 1569139307
transform 1 0 1448 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3037
timestamp 1569139307
transform 1 0 1448 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3038
timestamp 1569139307
transform 1 0 1448 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3039
timestamp 1569139307
transform 1 0 1384 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3040
timestamp 1569139307
transform 1 0 1448 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3041
timestamp 1569139307
transform 1 0 1384 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3042
timestamp 1569139307
transform 1 0 1384 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3043
timestamp 1569139307
transform 1 0 1448 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3044
timestamp 1569139307
transform 1 0 1448 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3045
timestamp 1569139307
transform 1 0 1448 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3046
timestamp 1569139307
transform 1 0 1448 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3047
timestamp 1569139307
transform 1 0 1512 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3048
timestamp 1569139307
transform 1 0 1512 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3049
timestamp 1569139307
transform 1 0 1512 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3050
timestamp 1569139307
transform 1 0 1512 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3051
timestamp 1569139307
transform 1 0 1512 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3052
timestamp 1569139307
transform 1 0 1512 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3053
timestamp 1569139307
transform 1 0 1512 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3054
timestamp 1569139307
transform 1 0 1512 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3055
timestamp 1569139307
transform 1 0 1320 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3056
timestamp 1569139307
transform 1 0 1320 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3057
timestamp 1569139307
transform 1 0 1320 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3058
timestamp 1569139307
transform 1 0 1320 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3059
timestamp 1569139307
transform 1 0 1320 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3060
timestamp 1569139307
transform 1 0 1320 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3061
timestamp 1569139307
transform 1 0 1320 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3062
timestamp 1569139307
transform 1 0 1512 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3063
timestamp 1569139307
transform 1 0 1320 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3064
timestamp 1569139307
transform 1 0 1384 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3065
timestamp 1569139307
transform 1 0 1512 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3066
timestamp 1569139307
transform 1 0 1512 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3067
timestamp 1569139307
transform 1 0 1448 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3068
timestamp 1569139307
transform 1 0 1512 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_3069
timestamp 1569139307
transform 1 0 1448 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3070
timestamp 1569139307
transform 1 0 1448 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3071
timestamp 1569139307
transform 1 0 1512 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_3072
timestamp 1569139307
transform 1 0 1320 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3073
timestamp 1569139307
transform 1 0 1320 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3074
timestamp 1569139307
transform 1 0 1320 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3075
timestamp 1569139307
transform 1 0 1320 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3076
timestamp 1569139307
transform 1 0 1320 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3077
timestamp 1569139307
transform 1 0 1512 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_3078
timestamp 1569139307
transform 1 0 1320 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_3079
timestamp 1569139307
transform 1 0 1320 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_3080
timestamp 1569139307
transform 1 0 1320 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_3081
timestamp 1569139307
transform 1 0 1320 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_3082
timestamp 1569139307
transform 1 0 1384 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3083
timestamp 1569139307
transform 1 0 1384 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3084
timestamp 1569139307
transform 1 0 1512 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_3085
timestamp 1569139307
transform 1 0 1384 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3086
timestamp 1569139307
transform 1 0 1448 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3087
timestamp 1569139307
transform 1 0 1384 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3088
timestamp 1569139307
transform 1 0 1384 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3089
timestamp 1569139307
transform 1 0 1384 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_3090
timestamp 1569139307
transform 1 0 1384 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_3091
timestamp 1569139307
transform 1 0 1384 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_3092
timestamp 1569139307
transform 1 0 1384 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_3093
timestamp 1569139307
transform 1 0 1448 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_3094
timestamp 1569139307
transform 1 0 1448 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_3095
timestamp 1569139307
transform 1 0 1448 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_3096
timestamp 1569139307
transform 1 0 1448 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_3097
timestamp 1569139307
transform 1 0 1512 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3098
timestamp 1569139307
transform 1 0 1512 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3099
timestamp 1569139307
transform 1 0 1512 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3100
timestamp 1569139307
transform 1 0 1512 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3101
timestamp 1569139307
transform 1 0 1448 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3102
timestamp 1569139307
transform 1 0 2344 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3103
timestamp 1569139307
transform 1 0 2344 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_3104
timestamp 1569139307
transform 1 0 2344 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_3105
timestamp 1569139307
transform 1 0 2344 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3106
timestamp 1569139307
transform 1 0 2408 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_3107
timestamp 1569139307
transform 1 0 2472 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_3108
timestamp 1569139307
transform 1 0 2344 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_3109
timestamp 1569139307
transform 1 0 2344 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3110
timestamp 1569139307
transform 1 0 2472 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3111
timestamp 1569139307
transform 1 0 2472 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3112
timestamp 1569139307
transform 1 0 2344 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3113
timestamp 1569139307
transform 1 0 2344 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_3114
timestamp 1569139307
transform 1 0 2344 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3115
timestamp 1569139307
transform 1 0 2472 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3116
timestamp 1569139307
transform 1 0 2472 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_3117
timestamp 1569139307
transform 1 0 2408 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3118
timestamp 1569139307
transform 1 0 2408 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3119
timestamp 1569139307
transform 1 0 2408 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3120
timestamp 1569139307
transform 1 0 2408 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3121
timestamp 1569139307
transform 1 0 2408 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3122
timestamp 1569139307
transform 1 0 2408 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_3123
timestamp 1569139307
transform 1 0 2408 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_3124
timestamp 1569139307
transform 1 0 2472 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_3125
timestamp 1569139307
transform 1 0 2408 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_3126
timestamp 1569139307
transform 1 0 2472 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_3127
timestamp 1569139307
transform 1 0 2472 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3128
timestamp 1569139307
transform 1 0 2472 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3129
timestamp 1569139307
transform 1 0 4840 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3130
timestamp 1569139307
transform 1 0 4840 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3131
timestamp 1569139307
transform 1 0 4904 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3132
timestamp 1569139307
transform 1 0 4712 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3133
timestamp 1569139307
transform 1 0 4776 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3134
timestamp 1569139307
transform 1 0 4904 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3135
timestamp 1569139307
transform 1 0 4840 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3136
timestamp 1569139307
transform 1 0 4904 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3137
timestamp 1569139307
transform 1 0 4776 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3138
timestamp 1569139307
transform 1 0 4776 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3139
timestamp 1569139307
transform 1 0 4840 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3140
timestamp 1569139307
transform 1 0 4712 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3141
timestamp 1569139307
transform 1 0 4712 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3142
timestamp 1569139307
transform 1 0 4776 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3143
timestamp 1569139307
transform 1 0 4712 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3144
timestamp 1569139307
transform 1 0 4712 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3145
timestamp 1569139307
transform 1 0 4840 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3146
timestamp 1569139307
transform 1 0 4904 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3147
timestamp 1569139307
transform 1 0 4776 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3148
timestamp 1569139307
transform 1 0 4904 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3149
timestamp 1569139307
transform 1 0 4520 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3150
timestamp 1569139307
transform 1 0 4648 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3151
timestamp 1569139307
transform 1 0 4456 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3152
timestamp 1569139307
transform 1 0 4456 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3153
timestamp 1569139307
transform 1 0 4648 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3154
timestamp 1569139307
transform 1 0 4392 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3155
timestamp 1569139307
transform 1 0 4584 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3156
timestamp 1569139307
transform 1 0 4392 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3157
timestamp 1569139307
transform 1 0 4520 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3158
timestamp 1569139307
transform 1 0 4648 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3159
timestamp 1569139307
transform 1 0 4584 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3160
timestamp 1569139307
transform 1 0 4456 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3161
timestamp 1569139307
transform 1 0 4584 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3162
timestamp 1569139307
transform 1 0 4648 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3163
timestamp 1569139307
transform 1 0 4392 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3164
timestamp 1569139307
transform 1 0 4520 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3165
timestamp 1569139307
transform 1 0 4520 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3166
timestamp 1569139307
transform 1 0 4520 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3167
timestamp 1569139307
transform 1 0 4456 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3168
timestamp 1569139307
transform 1 0 4584 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3169
timestamp 1569139307
transform 1 0 4392 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3170
timestamp 1569139307
transform 1 0 4392 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3171
timestamp 1569139307
transform 1 0 4456 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3172
timestamp 1569139307
transform 1 0 4584 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3173
timestamp 1569139307
transform 1 0 4648 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3174
timestamp 1569139307
transform 1 0 4392 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3175
timestamp 1569139307
transform 1 0 4456 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3176
timestamp 1569139307
transform 1 0 4520 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3177
timestamp 1569139307
transform 1 0 4392 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3178
timestamp 1569139307
transform 1 0 4584 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3179
timestamp 1569139307
transform 1 0 4392 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3180
timestamp 1569139307
transform 1 0 4520 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3181
timestamp 1569139307
transform 1 0 4584 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3182
timestamp 1569139307
transform 1 0 4392 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3183
timestamp 1569139307
transform 1 0 4392 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3184
timestamp 1569139307
transform 1 0 4456 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3185
timestamp 1569139307
transform 1 0 4456 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3186
timestamp 1569139307
transform 1 0 4648 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3187
timestamp 1569139307
transform 1 0 4584 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3188
timestamp 1569139307
transform 1 0 4456 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3189
timestamp 1569139307
transform 1 0 4520 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3190
timestamp 1569139307
transform 1 0 4584 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3191
timestamp 1569139307
transform 1 0 4520 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3192
timestamp 1569139307
transform 1 0 4648 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3193
timestamp 1569139307
transform 1 0 4648 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3194
timestamp 1569139307
transform 1 0 4648 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3195
timestamp 1569139307
transform 1 0 4584 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3196
timestamp 1569139307
transform 1 0 4520 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3197
timestamp 1569139307
transform 1 0 4456 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3198
timestamp 1569139307
transform 1 0 4648 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3199
timestamp 1569139307
transform 1 0 4776 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3200
timestamp 1569139307
transform 1 0 4904 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3201
timestamp 1569139307
transform 1 0 4904 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3202
timestamp 1569139307
transform 1 0 4840 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3203
timestamp 1569139307
transform 1 0 4712 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3204
timestamp 1569139307
transform 1 0 4904 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3205
timestamp 1569139307
transform 1 0 4712 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3206
timestamp 1569139307
transform 1 0 4776 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3207
timestamp 1569139307
transform 1 0 4840 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3208
timestamp 1569139307
transform 1 0 4712 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3209
timestamp 1569139307
transform 1 0 4904 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3210
timestamp 1569139307
transform 1 0 4776 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3211
timestamp 1569139307
transform 1 0 4776 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3212
timestamp 1569139307
transform 1 0 4840 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3213
timestamp 1569139307
transform 1 0 4712 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3214
timestamp 1569139307
transform 1 0 4776 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3215
timestamp 1569139307
transform 1 0 4840 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3216
timestamp 1569139307
transform 1 0 4904 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3217
timestamp 1569139307
transform 1 0 4840 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3218
timestamp 1569139307
transform 1 0 4712 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3219
timestamp 1569139307
transform 1 0 4328 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3220
timestamp 1569139307
transform 1 0 4136 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3221
timestamp 1569139307
transform 1 0 4200 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3222
timestamp 1569139307
transform 1 0 4264 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3223
timestamp 1569139307
transform 1 0 4264 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3224
timestamp 1569139307
transform 1 0 4264 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3225
timestamp 1569139307
transform 1 0 4072 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3226
timestamp 1569139307
transform 1 0 4328 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3227
timestamp 1569139307
transform 1 0 4264 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3228
timestamp 1569139307
transform 1 0 4200 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3229
timestamp 1569139307
transform 1 0 4136 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3230
timestamp 1569139307
transform 1 0 4136 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3231
timestamp 1569139307
transform 1 0 4072 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3232
timestamp 1569139307
transform 1 0 4328 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3233
timestamp 1569139307
transform 1 0 4200 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3234
timestamp 1569139307
transform 1 0 4072 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3235
timestamp 1569139307
transform 1 0 4072 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3236
timestamp 1569139307
transform 1 0 4264 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3237
timestamp 1569139307
transform 1 0 4200 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3238
timestamp 1569139307
transform 1 0 4136 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3239
timestamp 1569139307
transform 1 0 4328 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3240
timestamp 1569139307
transform 1 0 4136 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3241
timestamp 1569139307
transform 1 0 4200 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3242
timestamp 1569139307
transform 1 0 4328 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3243
timestamp 1569139307
transform 1 0 4072 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3244
timestamp 1569139307
transform 1 0 3816 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3245
timestamp 1569139307
transform 1 0 3880 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3246
timestamp 1569139307
transform 1 0 3752 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3247
timestamp 1569139307
transform 1 0 4008 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3248
timestamp 1569139307
transform 1 0 3752 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3249
timestamp 1569139307
transform 1 0 3880 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3250
timestamp 1569139307
transform 1 0 3944 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3251
timestamp 1569139307
transform 1 0 3944 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3252
timestamp 1569139307
transform 1 0 3944 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3253
timestamp 1569139307
transform 1 0 4008 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3254
timestamp 1569139307
transform 1 0 3752 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3255
timestamp 1569139307
transform 1 0 3944 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3256
timestamp 1569139307
transform 1 0 3944 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3257
timestamp 1569139307
transform 1 0 3752 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3258
timestamp 1569139307
transform 1 0 4008 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3259
timestamp 1569139307
transform 1 0 3880 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3260
timestamp 1569139307
transform 1 0 3816 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3261
timestamp 1569139307
transform 1 0 4008 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3262
timestamp 1569139307
transform 1 0 3816 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3263
timestamp 1569139307
transform 1 0 3880 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3264
timestamp 1569139307
transform 1 0 4008 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3265
timestamp 1569139307
transform 1 0 3816 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3266
timestamp 1569139307
transform 1 0 3816 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3267
timestamp 1569139307
transform 1 0 3752 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3268
timestamp 1569139307
transform 1 0 3880 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3269
timestamp 1569139307
transform 1 0 3944 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3270
timestamp 1569139307
transform 1 0 3752 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3271
timestamp 1569139307
transform 1 0 4008 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3272
timestamp 1569139307
transform 1 0 3880 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3273
timestamp 1569139307
transform 1 0 3752 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3274
timestamp 1569139307
transform 1 0 3944 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3275
timestamp 1569139307
transform 1 0 3880 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3276
timestamp 1569139307
transform 1 0 3752 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3277
timestamp 1569139307
transform 1 0 3752 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3278
timestamp 1569139307
transform 1 0 3944 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3279
timestamp 1569139307
transform 1 0 3816 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3280
timestamp 1569139307
transform 1 0 3944 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3281
timestamp 1569139307
transform 1 0 4008 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3282
timestamp 1569139307
transform 1 0 3880 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3283
timestamp 1569139307
transform 1 0 3816 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3284
timestamp 1569139307
transform 1 0 3816 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3285
timestamp 1569139307
transform 1 0 3816 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3286
timestamp 1569139307
transform 1 0 3816 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3287
timestamp 1569139307
transform 1 0 4008 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3288
timestamp 1569139307
transform 1 0 3752 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3289
timestamp 1569139307
transform 1 0 4008 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3290
timestamp 1569139307
transform 1 0 4008 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3291
timestamp 1569139307
transform 1 0 3944 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3292
timestamp 1569139307
transform 1 0 3880 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3293
timestamp 1569139307
transform 1 0 3880 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3294
timestamp 1569139307
transform 1 0 4136 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3295
timestamp 1569139307
transform 1 0 4200 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3296
timestamp 1569139307
transform 1 0 4136 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3297
timestamp 1569139307
transform 1 0 4264 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3298
timestamp 1569139307
transform 1 0 4264 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3299
timestamp 1569139307
transform 1 0 4072 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3300
timestamp 1569139307
transform 1 0 4200 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3301
timestamp 1569139307
transform 1 0 4072 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3302
timestamp 1569139307
transform 1 0 4136 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3303
timestamp 1569139307
transform 1 0 4264 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3304
timestamp 1569139307
transform 1 0 4072 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3305
timestamp 1569139307
transform 1 0 4136 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3306
timestamp 1569139307
transform 1 0 4264 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3307
timestamp 1569139307
transform 1 0 4136 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3308
timestamp 1569139307
transform 1 0 4200 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3309
timestamp 1569139307
transform 1 0 4264 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3310
timestamp 1569139307
transform 1 0 4328 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3311
timestamp 1569139307
transform 1 0 4328 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3312
timestamp 1569139307
transform 1 0 4328 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3313
timestamp 1569139307
transform 1 0 4200 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3314
timestamp 1569139307
transform 1 0 4328 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3315
timestamp 1569139307
transform 1 0 4328 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3316
timestamp 1569139307
transform 1 0 4072 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3317
timestamp 1569139307
transform 1 0 4200 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3318
timestamp 1569139307
transform 1 0 4072 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3319
timestamp 1569139307
transform 1 0 4328 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3320
timestamp 1569139307
transform 1 0 4264 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3321
timestamp 1569139307
transform 1 0 4072 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3322
timestamp 1569139307
transform 1 0 4200 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3323
timestamp 1569139307
transform 1 0 4200 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3324
timestamp 1569139307
transform 1 0 4136 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3325
timestamp 1569139307
transform 1 0 4264 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3326
timestamp 1569139307
transform 1 0 4136 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3327
timestamp 1569139307
transform 1 0 4136 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3328
timestamp 1569139307
transform 1 0 4072 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3329
timestamp 1569139307
transform 1 0 4200 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3330
timestamp 1569139307
transform 1 0 4328 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3331
timestamp 1569139307
transform 1 0 4072 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3332
timestamp 1569139307
transform 1 0 4072 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3333
timestamp 1569139307
transform 1 0 4264 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3334
timestamp 1569139307
transform 1 0 4328 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3335
timestamp 1569139307
transform 1 0 4264 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3336
timestamp 1569139307
transform 1 0 4200 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3337
timestamp 1569139307
transform 1 0 4136 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3338
timestamp 1569139307
transform 1 0 4328 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3339
timestamp 1569139307
transform 1 0 3816 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3340
timestamp 1569139307
transform 1 0 3880 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3341
timestamp 1569139307
transform 1 0 3944 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3342
timestamp 1569139307
transform 1 0 3944 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3343
timestamp 1569139307
transform 1 0 3880 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3344
timestamp 1569139307
transform 1 0 3752 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3345
timestamp 1569139307
transform 1 0 3944 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3346
timestamp 1569139307
transform 1 0 3944 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3347
timestamp 1569139307
transform 1 0 4008 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3348
timestamp 1569139307
transform 1 0 3816 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3349
timestamp 1569139307
transform 1 0 3752 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3350
timestamp 1569139307
transform 1 0 4008 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3351
timestamp 1569139307
transform 1 0 4008 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3352
timestamp 1569139307
transform 1 0 3816 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3353
timestamp 1569139307
transform 1 0 3880 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3354
timestamp 1569139307
transform 1 0 3752 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3355
timestamp 1569139307
transform 1 0 3752 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3356
timestamp 1569139307
transform 1 0 4008 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3357
timestamp 1569139307
transform 1 0 3816 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3358
timestamp 1569139307
transform 1 0 3880 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3359
timestamp 1569139307
transform 1 0 3752 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3360
timestamp 1569139307
transform 1 0 4008 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3361
timestamp 1569139307
transform 1 0 3880 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3362
timestamp 1569139307
transform 1 0 4008 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3363
timestamp 1569139307
transform 1 0 3752 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3364
timestamp 1569139307
transform 1 0 3880 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3365
timestamp 1569139307
transform 1 0 3880 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3366
timestamp 1569139307
transform 1 0 3944 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3367
timestamp 1569139307
transform 1 0 3944 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3368
timestamp 1569139307
transform 1 0 4008 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3369
timestamp 1569139307
transform 1 0 3816 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3370
timestamp 1569139307
transform 1 0 4008 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3371
timestamp 1569139307
transform 1 0 3880 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3372
timestamp 1569139307
transform 1 0 3944 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3373
timestamp 1569139307
transform 1 0 3816 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3374
timestamp 1569139307
transform 1 0 3816 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3375
timestamp 1569139307
transform 1 0 3816 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3376
timestamp 1569139307
transform 1 0 3752 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3377
timestamp 1569139307
transform 1 0 3752 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3378
timestamp 1569139307
transform 1 0 3944 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3379
timestamp 1569139307
transform 1 0 4072 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3380
timestamp 1569139307
transform 1 0 4264 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3381
timestamp 1569139307
transform 1 0 4264 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3382
timestamp 1569139307
transform 1 0 4200 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3383
timestamp 1569139307
transform 1 0 4072 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3384
timestamp 1569139307
transform 1 0 4136 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3385
timestamp 1569139307
transform 1 0 4328 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3386
timestamp 1569139307
transform 1 0 4072 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3387
timestamp 1569139307
transform 1 0 4200 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3388
timestamp 1569139307
transform 1 0 4136 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3389
timestamp 1569139307
transform 1 0 4328 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3390
timestamp 1569139307
transform 1 0 4328 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3391
timestamp 1569139307
transform 1 0 4264 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3392
timestamp 1569139307
transform 1 0 4328 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3393
timestamp 1569139307
transform 1 0 4200 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3394
timestamp 1569139307
transform 1 0 4136 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3395
timestamp 1569139307
transform 1 0 4200 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3396
timestamp 1569139307
transform 1 0 4072 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3397
timestamp 1569139307
transform 1 0 4264 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3398
timestamp 1569139307
transform 1 0 4136 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3399
timestamp 1569139307
transform 1 0 4264 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3400
timestamp 1569139307
transform 1 0 4072 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3401
timestamp 1569139307
transform 1 0 4328 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3402
timestamp 1569139307
transform 1 0 3944 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3403
timestamp 1569139307
transform 1 0 4200 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3404
timestamp 1569139307
transform 1 0 4136 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3405
timestamp 1569139307
transform 1 0 3752 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3406
timestamp 1569139307
transform 1 0 4008 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3407
timestamp 1569139307
transform 1 0 3816 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3408
timestamp 1569139307
transform 1 0 3880 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3409
timestamp 1569139307
transform 1 0 4776 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3410
timestamp 1569139307
transform 1 0 4840 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3411
timestamp 1569139307
transform 1 0 4712 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3412
timestamp 1569139307
transform 1 0 4840 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3413
timestamp 1569139307
transform 1 0 4712 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3414
timestamp 1569139307
transform 1 0 4776 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3415
timestamp 1569139307
transform 1 0 4904 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3416
timestamp 1569139307
transform 1 0 4776 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3417
timestamp 1569139307
transform 1 0 4904 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3418
timestamp 1569139307
transform 1 0 4840 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3419
timestamp 1569139307
transform 1 0 4840 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3420
timestamp 1569139307
transform 1 0 4712 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3421
timestamp 1569139307
transform 1 0 4904 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3422
timestamp 1569139307
transform 1 0 4776 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3423
timestamp 1569139307
transform 1 0 4712 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3424
timestamp 1569139307
transform 1 0 4904 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3425
timestamp 1569139307
transform 1 0 4648 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3426
timestamp 1569139307
transform 1 0 4584 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3427
timestamp 1569139307
transform 1 0 4456 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3428
timestamp 1569139307
transform 1 0 4456 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3429
timestamp 1569139307
transform 1 0 4648 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3430
timestamp 1569139307
transform 1 0 4456 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3431
timestamp 1569139307
transform 1 0 4456 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3432
timestamp 1569139307
transform 1 0 4584 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3433
timestamp 1569139307
transform 1 0 4584 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3434
timestamp 1569139307
transform 1 0 4520 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3435
timestamp 1569139307
transform 1 0 4520 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3436
timestamp 1569139307
transform 1 0 4392 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3437
timestamp 1569139307
transform 1 0 4520 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3438
timestamp 1569139307
transform 1 0 4520 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3439
timestamp 1569139307
transform 1 0 4392 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3440
timestamp 1569139307
transform 1 0 4392 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3441
timestamp 1569139307
transform 1 0 4392 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3442
timestamp 1569139307
transform 1 0 4584 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3443
timestamp 1569139307
transform 1 0 4648 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3444
timestamp 1569139307
transform 1 0 4648 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3445
timestamp 1569139307
transform 1 0 4392 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3446
timestamp 1569139307
transform 1 0 4392 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3447
timestamp 1569139307
transform 1 0 4648 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3448
timestamp 1569139307
transform 1 0 4520 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3449
timestamp 1569139307
transform 1 0 4584 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3450
timestamp 1569139307
transform 1 0 4520 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3451
timestamp 1569139307
transform 1 0 4392 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3452
timestamp 1569139307
transform 1 0 4456 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3453
timestamp 1569139307
transform 1 0 4520 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3454
timestamp 1569139307
transform 1 0 4392 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3455
timestamp 1569139307
transform 1 0 4456 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3456
timestamp 1569139307
transform 1 0 4648 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3457
timestamp 1569139307
transform 1 0 4456 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3458
timestamp 1569139307
transform 1 0 4584 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3459
timestamp 1569139307
transform 1 0 4648 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3460
timestamp 1569139307
transform 1 0 4584 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3461
timestamp 1569139307
transform 1 0 4456 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3462
timestamp 1569139307
transform 1 0 4648 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3463
timestamp 1569139307
transform 1 0 4584 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3464
timestamp 1569139307
transform 1 0 4520 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3465
timestamp 1569139307
transform 1 0 4712 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3466
timestamp 1569139307
transform 1 0 4904 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3467
timestamp 1569139307
transform 1 0 4776 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3468
timestamp 1569139307
transform 1 0 4840 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3469
timestamp 1569139307
transform 1 0 4712 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3470
timestamp 1569139307
transform 1 0 4840 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3471
timestamp 1569139307
transform 1 0 4712 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3472
timestamp 1569139307
transform 1 0 4904 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3473
timestamp 1569139307
transform 1 0 4712 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3474
timestamp 1569139307
transform 1 0 4904 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3475
timestamp 1569139307
transform 1 0 4904 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3476
timestamp 1569139307
transform 1 0 4840 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3477
timestamp 1569139307
transform 1 0 4776 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3478
timestamp 1569139307
transform 1 0 4840 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3479
timestamp 1569139307
transform 1 0 4776 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3480
timestamp 1569139307
transform 1 0 4776 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3481
timestamp 1569139307
transform 1 0 4840 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3482
timestamp 1569139307
transform 1 0 4712 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3483
timestamp 1569139307
transform 1 0 4392 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3484
timestamp 1569139307
transform 1 0 4776 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3485
timestamp 1569139307
transform 1 0 4456 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3486
timestamp 1569139307
transform 1 0 4520 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3487
timestamp 1569139307
transform 1 0 4904 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3488
timestamp 1569139307
transform 1 0 4584 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3489
timestamp 1569139307
transform 1 0 4648 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3490
timestamp 1569139307
transform 1 0 3624 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3491
timestamp 1569139307
transform 1 0 3496 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3492
timestamp 1569139307
transform 1 0 3496 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3493
timestamp 1569139307
transform 1 0 3496 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3494
timestamp 1569139307
transform 1 0 3624 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3495
timestamp 1569139307
transform 1 0 3560 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3496
timestamp 1569139307
transform 1 0 3560 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3497
timestamp 1569139307
transform 1 0 3624 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3498
timestamp 1569139307
transform 1 0 3624 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3499
timestamp 1569139307
transform 1 0 3560 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3500
timestamp 1569139307
transform 1 0 3688 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3501
timestamp 1569139307
transform 1 0 3688 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3502
timestamp 1569139307
transform 1 0 3688 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3503
timestamp 1569139307
transform 1 0 3560 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3504
timestamp 1569139307
transform 1 0 3688 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3505
timestamp 1569139307
transform 1 0 3688 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3506
timestamp 1569139307
transform 1 0 3560 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3507
timestamp 1569139307
transform 1 0 3496 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3508
timestamp 1569139307
transform 1 0 3624 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3509
timestamp 1569139307
transform 1 0 3496 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3510
timestamp 1569139307
transform 1 0 3368 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3511
timestamp 1569139307
transform 1 0 3368 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3512
timestamp 1569139307
transform 1 0 3304 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3513
timestamp 1569139307
transform 1 0 3176 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3514
timestamp 1569139307
transform 1 0 3176 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3515
timestamp 1569139307
transform 1 0 3176 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3516
timestamp 1569139307
transform 1 0 3176 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3517
timestamp 1569139307
transform 1 0 3176 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3518
timestamp 1569139307
transform 1 0 3304 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3519
timestamp 1569139307
transform 1 0 3240 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3520
timestamp 1569139307
transform 1 0 3240 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3521
timestamp 1569139307
transform 1 0 3240 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3522
timestamp 1569139307
transform 1 0 3240 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3523
timestamp 1569139307
transform 1 0 3240 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3524
timestamp 1569139307
transform 1 0 3304 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3525
timestamp 1569139307
transform 1 0 3304 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3526
timestamp 1569139307
transform 1 0 3304 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3527
timestamp 1569139307
transform 1 0 3368 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3528
timestamp 1569139307
transform 1 0 3368 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3529
timestamp 1569139307
transform 1 0 3368 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3530
timestamp 1569139307
transform 1 0 3176 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3531
timestamp 1569139307
transform 1 0 3240 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3532
timestamp 1569139307
transform 1 0 3304 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3533
timestamp 1569139307
transform 1 0 3368 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3534
timestamp 1569139307
transform 1 0 3304 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3535
timestamp 1569139307
transform 1 0 3304 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3536
timestamp 1569139307
transform 1 0 3176 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3537
timestamp 1569139307
transform 1 0 3368 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3538
timestamp 1569139307
transform 1 0 3368 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3539
timestamp 1569139307
transform 1 0 3368 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3540
timestamp 1569139307
transform 1 0 3176 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3541
timestamp 1569139307
transform 1 0 3368 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3542
timestamp 1569139307
transform 1 0 3304 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3543
timestamp 1569139307
transform 1 0 3240 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3544
timestamp 1569139307
transform 1 0 3240 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3545
timestamp 1569139307
transform 1 0 3240 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3546
timestamp 1569139307
transform 1 0 3240 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3547
timestamp 1569139307
transform 1 0 3304 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3548
timestamp 1569139307
transform 1 0 3176 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3549
timestamp 1569139307
transform 1 0 3176 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3550
timestamp 1569139307
transform 1 0 3688 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3551
timestamp 1569139307
transform 1 0 3624 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3552
timestamp 1569139307
transform 1 0 3688 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3553
timestamp 1569139307
transform 1 0 3496 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3554
timestamp 1569139307
transform 1 0 3496 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3555
timestamp 1569139307
transform 1 0 3688 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3556
timestamp 1569139307
transform 1 0 3496 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3557
timestamp 1569139307
transform 1 0 3496 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3558
timestamp 1569139307
transform 1 0 3688 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3559
timestamp 1569139307
transform 1 0 3688 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3560
timestamp 1569139307
transform 1 0 3560 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3561
timestamp 1569139307
transform 1 0 3496 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3562
timestamp 1569139307
transform 1 0 3560 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3563
timestamp 1569139307
transform 1 0 3560 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3564
timestamp 1569139307
transform 1 0 3560 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3565
timestamp 1569139307
transform 1 0 3560 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3566
timestamp 1569139307
transform 1 0 3624 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3567
timestamp 1569139307
transform 1 0 3624 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3568
timestamp 1569139307
transform 1 0 3624 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3569
timestamp 1569139307
transform 1 0 3624 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3570
timestamp 1569139307
transform 1 0 3432 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3571
timestamp 1569139307
transform 1 0 3432 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3572
timestamp 1569139307
transform 1 0 3432 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3573
timestamp 1569139307
transform 1 0 3432 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3574
timestamp 1569139307
transform 1 0 3432 0 1 2536
box -8 -8 8 8
use VIA2  VIA2_3575
timestamp 1569139307
transform 1 0 3432 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3576
timestamp 1569139307
transform 1 0 3432 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3577
timestamp 1569139307
transform 1 0 3432 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3578
timestamp 1569139307
transform 1 0 3432 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3579
timestamp 1569139307
transform 1 0 3432 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3580
timestamp 1569139307
transform 1 0 3048 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3581
timestamp 1569139307
transform 1 0 3048 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3582
timestamp 1569139307
transform 1 0 3112 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3583
timestamp 1569139307
transform 1 0 2600 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3584
timestamp 1569139307
transform 1 0 2856 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3585
timestamp 1569139307
transform 1 0 2856 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3586
timestamp 1569139307
transform 1 0 2856 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3587
timestamp 1569139307
transform 1 0 2856 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3588
timestamp 1569139307
transform 1 0 2792 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3589
timestamp 1569139307
transform 1 0 2792 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3590
timestamp 1569139307
transform 1 0 2792 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3591
timestamp 1569139307
transform 1 0 2792 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3592
timestamp 1569139307
transform 1 0 3112 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3593
timestamp 1569139307
transform 1 0 3112 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3594
timestamp 1569139307
transform 1 0 2920 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3595
timestamp 1569139307
transform 1 0 2920 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3596
timestamp 1569139307
transform 1 0 2920 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3597
timestamp 1569139307
transform 1 0 2920 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3598
timestamp 1569139307
transform 1 0 3112 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3599
timestamp 1569139307
transform 1 0 3048 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3600
timestamp 1569139307
transform 1 0 3048 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3601
timestamp 1569139307
transform 1 0 3048 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3602
timestamp 1569139307
transform 1 0 3048 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3603
timestamp 1569139307
transform 1 0 3112 0 1 2600
box -8 -8 8 8
use VIA2  VIA2_3604
timestamp 1569139307
transform 1 0 2664 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3605
timestamp 1569139307
transform 1 0 2664 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3606
timestamp 1569139307
transform 1 0 3112 0 1 2664
box -8 -8 8 8
use VIA2  VIA2_3607
timestamp 1569139307
transform 1 0 3112 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3608
timestamp 1569139307
transform 1 0 3112 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3609
timestamp 1569139307
transform 1 0 3112 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3610
timestamp 1569139307
transform 1 0 2856 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3611
timestamp 1569139307
transform 1 0 2920 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3612
timestamp 1569139307
transform 1 0 2920 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3613
timestamp 1569139307
transform 1 0 2984 0 1 2728
box -8 -8 8 8
use VIA2  VIA2_3614
timestamp 1569139307
transform 1 0 2984 0 1 2792
box -8 -8 8 8
use VIA2  VIA2_3615
timestamp 1569139307
transform 1 0 2984 0 1 2856
box -8 -8 8 8
use VIA2  VIA2_3616
timestamp 1569139307
transform 1 0 2728 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3617
timestamp 1569139307
transform 1 0 2728 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3618
timestamp 1569139307
transform 1 0 2984 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3619
timestamp 1569139307
transform 1 0 2984 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3620
timestamp 1569139307
transform 1 0 2984 0 1 3048
box -8 -8 8 8
use VIA2  VIA2_3621
timestamp 1569139307
transform 1 0 2984 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3622
timestamp 1569139307
transform 1 0 2728 0 1 3112
box -8 -8 8 8
use VIA2  VIA2_3623
timestamp 1569139307
transform 1 0 3048 0 1 2920
box -8 -8 8 8
use VIA2  VIA2_3624
timestamp 1569139307
transform 1 0 3048 0 1 2984
box -8 -8 8 8
use VIA2  VIA2_3625
timestamp 1569139307
transform 1 0 2984 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3626
timestamp 1569139307
transform 1 0 2984 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3627
timestamp 1569139307
transform 1 0 2920 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3628
timestamp 1569139307
transform 1 0 3112 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3629
timestamp 1569139307
transform 1 0 3048 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3630
timestamp 1569139307
transform 1 0 3112 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3631
timestamp 1569139307
transform 1 0 2920 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3632
timestamp 1569139307
transform 1 0 2920 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3633
timestamp 1569139307
transform 1 0 3048 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3634
timestamp 1569139307
transform 1 0 2856 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3635
timestamp 1569139307
transform 1 0 3112 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3636
timestamp 1569139307
transform 1 0 2920 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3637
timestamp 1569139307
transform 1 0 3048 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3638
timestamp 1569139307
transform 1 0 2856 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3639
timestamp 1569139307
transform 1 0 2856 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3640
timestamp 1569139307
transform 1 0 2856 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3641
timestamp 1569139307
transform 1 0 2984 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3642
timestamp 1569139307
transform 1 0 3048 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3643
timestamp 1569139307
transform 1 0 3112 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3644
timestamp 1569139307
transform 1 0 2984 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3645
timestamp 1569139307
transform 1 0 2600 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3646
timestamp 1569139307
transform 1 0 2600 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3647
timestamp 1569139307
transform 1 0 2792 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3648
timestamp 1569139307
transform 1 0 2600 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3649
timestamp 1569139307
transform 1 0 2536 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3650
timestamp 1569139307
transform 1 0 2536 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3651
timestamp 1569139307
transform 1 0 2728 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3652
timestamp 1569139307
transform 1 0 2792 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3653
timestamp 1569139307
transform 1 0 2728 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3654
timestamp 1569139307
transform 1 0 2600 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3655
timestamp 1569139307
transform 1 0 2536 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3656
timestamp 1569139307
transform 1 0 2728 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3657
timestamp 1569139307
transform 1 0 2664 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3658
timestamp 1569139307
transform 1 0 2792 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3659
timestamp 1569139307
transform 1 0 2664 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3660
timestamp 1569139307
transform 1 0 2536 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3661
timestamp 1569139307
transform 1 0 2728 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3662
timestamp 1569139307
transform 1 0 2664 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3663
timestamp 1569139307
transform 1 0 2792 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3664
timestamp 1569139307
transform 1 0 2664 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3665
timestamp 1569139307
transform 1 0 2600 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3666
timestamp 1569139307
transform 1 0 2536 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3667
timestamp 1569139307
transform 1 0 2728 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3668
timestamp 1569139307
transform 1 0 2728 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3669
timestamp 1569139307
transform 1 0 2792 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3670
timestamp 1569139307
transform 1 0 2536 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3671
timestamp 1569139307
transform 1 0 2728 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3672
timestamp 1569139307
transform 1 0 2792 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3673
timestamp 1569139307
transform 1 0 2728 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3674
timestamp 1569139307
transform 1 0 2792 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3675
timestamp 1569139307
transform 1 0 2792 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3676
timestamp 1569139307
transform 1 0 2600 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3677
timestamp 1569139307
transform 1 0 2664 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3678
timestamp 1569139307
transform 1 0 2664 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3679
timestamp 1569139307
transform 1 0 2664 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3680
timestamp 1569139307
transform 1 0 2536 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3681
timestamp 1569139307
transform 1 0 2600 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3682
timestamp 1569139307
transform 1 0 2664 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3683
timestamp 1569139307
transform 1 0 2536 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3684
timestamp 1569139307
transform 1 0 2600 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3685
timestamp 1569139307
transform 1 0 2856 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3686
timestamp 1569139307
transform 1 0 2984 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3687
timestamp 1569139307
transform 1 0 2984 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3688
timestamp 1569139307
transform 1 0 2984 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3689
timestamp 1569139307
transform 1 0 2856 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3690
timestamp 1569139307
transform 1 0 2856 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3691
timestamp 1569139307
transform 1 0 3048 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3692
timestamp 1569139307
transform 1 0 2984 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3693
timestamp 1569139307
transform 1 0 3048 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3694
timestamp 1569139307
transform 1 0 2920 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3695
timestamp 1569139307
transform 1 0 2920 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3696
timestamp 1569139307
transform 1 0 3112 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3697
timestamp 1569139307
transform 1 0 2920 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3698
timestamp 1569139307
transform 1 0 3048 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3699
timestamp 1569139307
transform 1 0 3048 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3700
timestamp 1569139307
transform 1 0 3112 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3701
timestamp 1569139307
transform 1 0 3112 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3702
timestamp 1569139307
transform 1 0 2920 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3703
timestamp 1569139307
transform 1 0 3112 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3704
timestamp 1569139307
transform 1 0 2856 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3705
timestamp 1569139307
transform 1 0 2984 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3706
timestamp 1569139307
transform 1 0 3048 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3707
timestamp 1569139307
transform 1 0 2728 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3708
timestamp 1569139307
transform 1 0 2600 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3709
timestamp 1569139307
transform 1 0 2792 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3710
timestamp 1569139307
transform 1 0 2664 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3711
timestamp 1569139307
transform 1 0 3112 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3712
timestamp 1569139307
transform 1 0 2856 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3713
timestamp 1569139307
transform 1 0 2920 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3714
timestamp 1569139307
transform 1 0 2536 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3715
timestamp 1569139307
transform 1 0 3688 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3716
timestamp 1569139307
transform 1 0 3496 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3717
timestamp 1569139307
transform 1 0 3496 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3718
timestamp 1569139307
transform 1 0 3496 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3719
timestamp 1569139307
transform 1 0 3496 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3720
timestamp 1569139307
transform 1 0 3688 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3721
timestamp 1569139307
transform 1 0 3560 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3722
timestamp 1569139307
transform 1 0 3560 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3723
timestamp 1569139307
transform 1 0 3560 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3724
timestamp 1569139307
transform 1 0 3560 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3725
timestamp 1569139307
transform 1 0 3688 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3726
timestamp 1569139307
transform 1 0 3624 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3727
timestamp 1569139307
transform 1 0 3624 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3728
timestamp 1569139307
transform 1 0 3688 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3729
timestamp 1569139307
transform 1 0 3624 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3730
timestamp 1569139307
transform 1 0 3624 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3731
timestamp 1569139307
transform 1 0 3304 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3732
timestamp 1569139307
transform 1 0 3176 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3733
timestamp 1569139307
transform 1 0 3176 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3734
timestamp 1569139307
transform 1 0 3304 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3735
timestamp 1569139307
transform 1 0 3304 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3736
timestamp 1569139307
transform 1 0 3304 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3737
timestamp 1569139307
transform 1 0 3176 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3738
timestamp 1569139307
transform 1 0 3176 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3739
timestamp 1569139307
transform 1 0 3240 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3740
timestamp 1569139307
transform 1 0 3240 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3741
timestamp 1569139307
transform 1 0 3240 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3742
timestamp 1569139307
transform 1 0 3240 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3743
timestamp 1569139307
transform 1 0 3368 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3744
timestamp 1569139307
transform 1 0 3368 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3745
timestamp 1569139307
transform 1 0 3368 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3746
timestamp 1569139307
transform 1 0 3368 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3747
timestamp 1569139307
transform 1 0 3176 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3748
timestamp 1569139307
transform 1 0 3176 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3749
timestamp 1569139307
transform 1 0 3368 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3750
timestamp 1569139307
transform 1 0 3240 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3751
timestamp 1569139307
transform 1 0 3240 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3752
timestamp 1569139307
transform 1 0 3240 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3753
timestamp 1569139307
transform 1 0 3240 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3754
timestamp 1569139307
transform 1 0 3368 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3755
timestamp 1569139307
transform 1 0 3368 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3756
timestamp 1569139307
transform 1 0 3176 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3757
timestamp 1569139307
transform 1 0 3176 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3758
timestamp 1569139307
transform 1 0 3304 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3759
timestamp 1569139307
transform 1 0 3304 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3760
timestamp 1569139307
transform 1 0 3304 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3761
timestamp 1569139307
transform 1 0 3304 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3762
timestamp 1569139307
transform 1 0 3368 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3763
timestamp 1569139307
transform 1 0 3688 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3764
timestamp 1569139307
transform 1 0 3688 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3765
timestamp 1569139307
transform 1 0 3688 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3766
timestamp 1569139307
transform 1 0 3688 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3767
timestamp 1569139307
transform 1 0 3496 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3768
timestamp 1569139307
transform 1 0 3496 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3769
timestamp 1569139307
transform 1 0 3560 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3770
timestamp 1569139307
transform 1 0 3560 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3771
timestamp 1569139307
transform 1 0 3624 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3772
timestamp 1569139307
transform 1 0 3624 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3773
timestamp 1569139307
transform 1 0 3496 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3774
timestamp 1569139307
transform 1 0 3496 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3775
timestamp 1569139307
transform 1 0 3624 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3776
timestamp 1569139307
transform 1 0 3624 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3777
timestamp 1569139307
transform 1 0 3560 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3778
timestamp 1569139307
transform 1 0 3560 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3779
timestamp 1569139307
transform 1 0 3240 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3780
timestamp 1569139307
transform 1 0 3304 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3781
timestamp 1569139307
transform 1 0 3432 0 1 3560
box -8 -8 8 8
use VIA2  VIA2_3782
timestamp 1569139307
transform 1 0 3496 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3783
timestamp 1569139307
transform 1 0 3560 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3784
timestamp 1569139307
transform 1 0 3624 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3785
timestamp 1569139307
transform 1 0 3432 0 1 3624
box -8 -8 8 8
use VIA2  VIA2_3786
timestamp 1569139307
transform 1 0 3432 0 1 3688
box -8 -8 8 8
use VIA2  VIA2_3787
timestamp 1569139307
transform 1 0 3368 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3788
timestamp 1569139307
transform 1 0 3432 0 1 3176
box -8 -8 8 8
use VIA2  VIA2_3789
timestamp 1569139307
transform 1 0 3432 0 1 3240
box -8 -8 8 8
use VIA2  VIA2_3790
timestamp 1569139307
transform 1 0 3432 0 1 3304
box -8 -8 8 8
use VIA2  VIA2_3791
timestamp 1569139307
transform 1 0 3432 0 1 3368
box -8 -8 8 8
use VIA2  VIA2_3792
timestamp 1569139307
transform 1 0 3432 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3793
timestamp 1569139307
transform 1 0 3432 0 1 3496
box -8 -8 8 8
use VIA2  VIA2_3794
timestamp 1569139307
transform 1 0 3688 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3795
timestamp 1569139307
transform 1 0 3176 0 1 3432
box -8 -8 8 8
use VIA2  VIA2_3796
timestamp 1569139307
transform 1 0 3688 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3797
timestamp 1569139307
transform 1 0 3624 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3798
timestamp 1569139307
transform 1 0 3560 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3799
timestamp 1569139307
transform 1 0 3496 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3800
timestamp 1569139307
transform 1 0 3688 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3801
timestamp 1569139307
transform 1 0 3624 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3802
timestamp 1569139307
transform 1 0 3688 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3803
timestamp 1569139307
transform 1 0 3624 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3804
timestamp 1569139307
transform 1 0 3496 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3805
timestamp 1569139307
transform 1 0 3560 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3806
timestamp 1569139307
transform 1 0 3496 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3807
timestamp 1569139307
transform 1 0 3560 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3808
timestamp 1569139307
transform 1 0 3624 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3809
timestamp 1569139307
transform 1 0 3560 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3810
timestamp 1569139307
transform 1 0 3688 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3811
timestamp 1569139307
transform 1 0 3560 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3812
timestamp 1569139307
transform 1 0 3688 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3813
timestamp 1569139307
transform 1 0 3624 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3814
timestamp 1569139307
transform 1 0 3496 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3815
timestamp 1569139307
transform 1 0 3496 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3816
timestamp 1569139307
transform 1 0 3368 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3817
timestamp 1569139307
transform 1 0 3368 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3818
timestamp 1569139307
transform 1 0 3240 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3819
timestamp 1569139307
transform 1 0 3176 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3820
timestamp 1569139307
transform 1 0 3240 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3821
timestamp 1569139307
transform 1 0 3240 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3822
timestamp 1569139307
transform 1 0 3304 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3823
timestamp 1569139307
transform 1 0 3176 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3824
timestamp 1569139307
transform 1 0 3368 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3825
timestamp 1569139307
transform 1 0 3304 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3826
timestamp 1569139307
transform 1 0 3304 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3827
timestamp 1569139307
transform 1 0 3304 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3828
timestamp 1569139307
transform 1 0 3240 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3829
timestamp 1569139307
transform 1 0 3176 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3830
timestamp 1569139307
transform 1 0 3176 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3831
timestamp 1569139307
transform 1 0 3368 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3832
timestamp 1569139307
transform 1 0 3304 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3833
timestamp 1569139307
transform 1 0 3368 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3834
timestamp 1569139307
transform 1 0 3176 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3835
timestamp 1569139307
transform 1 0 3240 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3836
timestamp 1569139307
transform 1 0 3304 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3837
timestamp 1569139307
transform 1 0 3240 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3838
timestamp 1569139307
transform 1 0 3176 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3839
timestamp 1569139307
transform 1 0 3240 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3840
timestamp 1569139307
transform 1 0 3176 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3841
timestamp 1569139307
transform 1 0 3176 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3842
timestamp 1569139307
transform 1 0 3368 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3843
timestamp 1569139307
transform 1 0 3304 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3844
timestamp 1569139307
transform 1 0 3240 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3845
timestamp 1569139307
transform 1 0 3240 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3846
timestamp 1569139307
transform 1 0 3368 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3847
timestamp 1569139307
transform 1 0 3176 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3848
timestamp 1569139307
transform 1 0 3304 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3849
timestamp 1569139307
transform 1 0 3368 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3850
timestamp 1569139307
transform 1 0 3304 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3851
timestamp 1569139307
transform 1 0 3304 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3852
timestamp 1569139307
transform 1 0 3240 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3853
timestamp 1569139307
transform 1 0 3368 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3854
timestamp 1569139307
transform 1 0 3176 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3855
timestamp 1569139307
transform 1 0 3368 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3856
timestamp 1569139307
transform 1 0 3624 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3857
timestamp 1569139307
transform 1 0 3624 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3858
timestamp 1569139307
transform 1 0 3688 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3859
timestamp 1569139307
transform 1 0 3496 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3860
timestamp 1569139307
transform 1 0 3624 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3861
timestamp 1569139307
transform 1 0 3688 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3862
timestamp 1569139307
transform 1 0 3560 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3863
timestamp 1569139307
transform 1 0 3688 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3864
timestamp 1569139307
transform 1 0 3688 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3865
timestamp 1569139307
transform 1 0 3496 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3866
timestamp 1569139307
transform 1 0 3688 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3867
timestamp 1569139307
transform 1 0 3624 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3868
timestamp 1569139307
transform 1 0 3496 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3869
timestamp 1569139307
transform 1 0 3496 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3870
timestamp 1569139307
transform 1 0 3560 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3871
timestamp 1569139307
transform 1 0 3560 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3872
timestamp 1569139307
transform 1 0 3496 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3873
timestamp 1569139307
transform 1 0 3560 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3874
timestamp 1569139307
transform 1 0 3560 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3875
timestamp 1569139307
transform 1 0 3624 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3876
timestamp 1569139307
transform 1 0 3432 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3877
timestamp 1569139307
transform 1 0 3432 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3878
timestamp 1569139307
transform 1 0 3432 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3879
timestamp 1569139307
transform 1 0 3432 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3880
timestamp 1569139307
transform 1 0 3432 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3881
timestamp 1569139307
transform 1 0 3432 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3882
timestamp 1569139307
transform 1 0 3432 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3883
timestamp 1569139307
transform 1 0 3432 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3884
timestamp 1569139307
transform 1 0 3432 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3885
timestamp 1569139307
transform 1 0 3432 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3886
timestamp 1569139307
transform 1 0 2984 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3887
timestamp 1569139307
transform 1 0 3112 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3888
timestamp 1569139307
transform 1 0 2984 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3889
timestamp 1569139307
transform 1 0 2920 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3890
timestamp 1569139307
transform 1 0 3112 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3891
timestamp 1569139307
transform 1 0 2920 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3892
timestamp 1569139307
transform 1 0 2856 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3893
timestamp 1569139307
transform 1 0 2984 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3894
timestamp 1569139307
transform 1 0 2984 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3895
timestamp 1569139307
transform 1 0 2984 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3896
timestamp 1569139307
transform 1 0 3112 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3897
timestamp 1569139307
transform 1 0 2856 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3898
timestamp 1569139307
transform 1 0 3048 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3899
timestamp 1569139307
transform 1 0 2856 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3900
timestamp 1569139307
transform 1 0 2920 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3901
timestamp 1569139307
transform 1 0 2920 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3902
timestamp 1569139307
transform 1 0 3048 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3903
timestamp 1569139307
transform 1 0 3112 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3904
timestamp 1569139307
transform 1 0 2856 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3905
timestamp 1569139307
transform 1 0 3048 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3906
timestamp 1569139307
transform 1 0 3048 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3907
timestamp 1569139307
transform 1 0 3112 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3908
timestamp 1569139307
transform 1 0 3048 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3909
timestamp 1569139307
transform 1 0 2920 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3910
timestamp 1569139307
transform 1 0 2856 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3911
timestamp 1569139307
transform 1 0 2664 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3912
timestamp 1569139307
transform 1 0 2536 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3913
timestamp 1569139307
transform 1 0 2728 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3914
timestamp 1569139307
transform 1 0 2536 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3915
timestamp 1569139307
transform 1 0 2728 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3916
timestamp 1569139307
transform 1 0 2536 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3917
timestamp 1569139307
transform 1 0 2728 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3918
timestamp 1569139307
transform 1 0 2600 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3919
timestamp 1569139307
transform 1 0 2600 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3920
timestamp 1569139307
transform 1 0 2664 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3921
timestamp 1569139307
transform 1 0 2600 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3922
timestamp 1569139307
transform 1 0 2664 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3923
timestamp 1569139307
transform 1 0 2728 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3924
timestamp 1569139307
transform 1 0 2728 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3925
timestamp 1569139307
transform 1 0 2600 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3926
timestamp 1569139307
transform 1 0 2664 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3927
timestamp 1569139307
transform 1 0 2792 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3928
timestamp 1569139307
transform 1 0 2600 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3929
timestamp 1569139307
transform 1 0 2792 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3930
timestamp 1569139307
transform 1 0 2536 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3931
timestamp 1569139307
transform 1 0 2792 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_3932
timestamp 1569139307
transform 1 0 2664 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_3933
timestamp 1569139307
transform 1 0 2536 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_3934
timestamp 1569139307
transform 1 0 2792 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_3935
timestamp 1569139307
transform 1 0 2792 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_3936
timestamp 1569139307
transform 1 0 2792 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3937
timestamp 1569139307
transform 1 0 2664 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3938
timestamp 1569139307
transform 1 0 2536 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3939
timestamp 1569139307
transform 1 0 2536 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3940
timestamp 1569139307
transform 1 0 2600 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3941
timestamp 1569139307
transform 1 0 2600 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3942
timestamp 1569139307
transform 1 0 2728 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3943
timestamp 1569139307
transform 1 0 2600 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3944
timestamp 1569139307
transform 1 0 2664 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3945
timestamp 1569139307
transform 1 0 2728 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3946
timestamp 1569139307
transform 1 0 2792 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3947
timestamp 1569139307
transform 1 0 2792 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3948
timestamp 1569139307
transform 1 0 2728 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3949
timestamp 1569139307
transform 1 0 2664 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3950
timestamp 1569139307
transform 1 0 2792 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3951
timestamp 1569139307
transform 1 0 2536 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3952
timestamp 1569139307
transform 1 0 2792 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3953
timestamp 1569139307
transform 1 0 2536 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3954
timestamp 1569139307
transform 1 0 2536 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3955
timestamp 1569139307
transform 1 0 2728 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3956
timestamp 1569139307
transform 1 0 2600 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3957
timestamp 1569139307
transform 1 0 2664 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3958
timestamp 1569139307
transform 1 0 2664 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3959
timestamp 1569139307
transform 1 0 2728 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3960
timestamp 1569139307
transform 1 0 2600 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3961
timestamp 1569139307
transform 1 0 2856 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3962
timestamp 1569139307
transform 1 0 2984 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3963
timestamp 1569139307
transform 1 0 2984 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3964
timestamp 1569139307
transform 1 0 3112 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3965
timestamp 1569139307
transform 1 0 3112 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3966
timestamp 1569139307
transform 1 0 2984 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3967
timestamp 1569139307
transform 1 0 2920 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3968
timestamp 1569139307
transform 1 0 2920 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3969
timestamp 1569139307
transform 1 0 3048 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3970
timestamp 1569139307
transform 1 0 3048 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3971
timestamp 1569139307
transform 1 0 2920 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3972
timestamp 1569139307
transform 1 0 2920 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3973
timestamp 1569139307
transform 1 0 2920 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3974
timestamp 1569139307
transform 1 0 2984 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3975
timestamp 1569139307
transform 1 0 2984 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_3976
timestamp 1569139307
transform 1 0 3048 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3977
timestamp 1569139307
transform 1 0 3048 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3978
timestamp 1569139307
transform 1 0 3048 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3979
timestamp 1569139307
transform 1 0 3112 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3980
timestamp 1569139307
transform 1 0 3112 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3981
timestamp 1569139307
transform 1 0 3112 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3982
timestamp 1569139307
transform 1 0 2856 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_3983
timestamp 1569139307
transform 1 0 2856 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_3984
timestamp 1569139307
transform 1 0 2856 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_3985
timestamp 1569139307
transform 1 0 2856 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_3986
timestamp 1569139307
transform 1 0 2856 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3987
timestamp 1569139307
transform 1 0 3112 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3988
timestamp 1569139307
transform 1 0 2920 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3989
timestamp 1569139307
transform 1 0 3048 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3990
timestamp 1569139307
transform 1 0 2920 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_3991
timestamp 1569139307
transform 1 0 3048 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3992
timestamp 1569139307
transform 1 0 3112 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3993
timestamp 1569139307
transform 1 0 3048 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_3994
timestamp 1569139307
transform 1 0 2856 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_3995
timestamp 1569139307
transform 1 0 2920 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3996
timestamp 1569139307
transform 1 0 2984 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_3997
timestamp 1569139307
transform 1 0 2856 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3998
timestamp 1569139307
transform 1 0 3112 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_3999
timestamp 1569139307
transform 1 0 2984 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4000
timestamp 1569139307
transform 1 0 2920 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4001
timestamp 1569139307
transform 1 0 3048 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4002
timestamp 1569139307
transform 1 0 2920 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4003
timestamp 1569139307
transform 1 0 2984 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4004
timestamp 1569139307
transform 1 0 2856 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4005
timestamp 1569139307
transform 1 0 3048 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4006
timestamp 1569139307
transform 1 0 2984 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4007
timestamp 1569139307
transform 1 0 2856 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4008
timestamp 1569139307
transform 1 0 3112 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4009
timestamp 1569139307
transform 1 0 2984 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4010
timestamp 1569139307
transform 1 0 3112 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4011
timestamp 1569139307
transform 1 0 2536 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4012
timestamp 1569139307
transform 1 0 2600 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4013
timestamp 1569139307
transform 1 0 2664 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4014
timestamp 1569139307
transform 1 0 2664 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4015
timestamp 1569139307
transform 1 0 2536 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4016
timestamp 1569139307
transform 1 0 2728 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4017
timestamp 1569139307
transform 1 0 2664 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4018
timestamp 1569139307
transform 1 0 2536 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4019
timestamp 1569139307
transform 1 0 2728 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4020
timestamp 1569139307
transform 1 0 2664 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4021
timestamp 1569139307
transform 1 0 2536 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4022
timestamp 1569139307
transform 1 0 2664 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4023
timestamp 1569139307
transform 1 0 2536 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4024
timestamp 1569139307
transform 1 0 2792 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4025
timestamp 1569139307
transform 1 0 2600 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4026
timestamp 1569139307
transform 1 0 2728 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4027
timestamp 1569139307
transform 1 0 2728 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4028
timestamp 1569139307
transform 1 0 2600 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4029
timestamp 1569139307
transform 1 0 2792 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4030
timestamp 1569139307
transform 1 0 2792 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4031
timestamp 1569139307
transform 1 0 2728 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4032
timestamp 1569139307
transform 1 0 2600 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4033
timestamp 1569139307
transform 1 0 2792 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4034
timestamp 1569139307
transform 1 0 2600 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4035
timestamp 1569139307
transform 1 0 2792 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4036
timestamp 1569139307
transform 1 0 2536 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4037
timestamp 1569139307
transform 1 0 2792 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4038
timestamp 1569139307
transform 1 0 2664 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4039
timestamp 1569139307
transform 1 0 2664 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4040
timestamp 1569139307
transform 1 0 2728 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4041
timestamp 1569139307
transform 1 0 2664 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4042
timestamp 1569139307
transform 1 0 2728 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4043
timestamp 1569139307
transform 1 0 2600 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4044
timestamp 1569139307
transform 1 0 2536 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4045
timestamp 1569139307
transform 1 0 2600 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4046
timestamp 1569139307
transform 1 0 2664 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4047
timestamp 1569139307
transform 1 0 2792 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4048
timestamp 1569139307
transform 1 0 2536 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4049
timestamp 1569139307
transform 1 0 2728 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4050
timestamp 1569139307
transform 1 0 2536 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4051
timestamp 1569139307
transform 1 0 2728 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4052
timestamp 1569139307
transform 1 0 2792 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4053
timestamp 1569139307
transform 1 0 2600 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4054
timestamp 1569139307
transform 1 0 2600 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4055
timestamp 1569139307
transform 1 0 2792 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4056
timestamp 1569139307
transform 1 0 3112 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4057
timestamp 1569139307
transform 1 0 2920 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4058
timestamp 1569139307
transform 1 0 2920 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4059
timestamp 1569139307
transform 1 0 2984 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4060
timestamp 1569139307
transform 1 0 2984 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4061
timestamp 1569139307
transform 1 0 2984 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4062
timestamp 1569139307
transform 1 0 3048 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4063
timestamp 1569139307
transform 1 0 3112 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4064
timestamp 1569139307
transform 1 0 3112 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4065
timestamp 1569139307
transform 1 0 3048 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4066
timestamp 1569139307
transform 1 0 2856 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4067
timestamp 1569139307
transform 1 0 2920 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4068
timestamp 1569139307
transform 1 0 3048 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4069
timestamp 1569139307
transform 1 0 2984 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4070
timestamp 1569139307
transform 1 0 3112 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4071
timestamp 1569139307
transform 1 0 3048 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4072
timestamp 1569139307
transform 1 0 2856 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4073
timestamp 1569139307
transform 1 0 2856 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4074
timestamp 1569139307
transform 1 0 2856 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4075
timestamp 1569139307
transform 1 0 2920 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4076
timestamp 1569139307
transform 1 0 3496 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4077
timestamp 1569139307
transform 1 0 3496 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4078
timestamp 1569139307
transform 1 0 3496 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4079
timestamp 1569139307
transform 1 0 3688 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4080
timestamp 1569139307
transform 1 0 3688 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4081
timestamp 1569139307
transform 1 0 3688 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4082
timestamp 1569139307
transform 1 0 3560 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4083
timestamp 1569139307
transform 1 0 3560 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4084
timestamp 1569139307
transform 1 0 3560 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4085
timestamp 1569139307
transform 1 0 3560 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4086
timestamp 1569139307
transform 1 0 3560 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4087
timestamp 1569139307
transform 1 0 3688 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4088
timestamp 1569139307
transform 1 0 3688 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4089
timestamp 1569139307
transform 1 0 3624 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4090
timestamp 1569139307
transform 1 0 3624 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4091
timestamp 1569139307
transform 1 0 3624 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4092
timestamp 1569139307
transform 1 0 3624 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4093
timestamp 1569139307
transform 1 0 3496 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4094
timestamp 1569139307
transform 1 0 3624 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4095
timestamp 1569139307
transform 1 0 3496 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4096
timestamp 1569139307
transform 1 0 3304 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4097
timestamp 1569139307
transform 1 0 3240 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4098
timestamp 1569139307
transform 1 0 3176 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4099
timestamp 1569139307
transform 1 0 3304 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4100
timestamp 1569139307
transform 1 0 3176 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4101
timestamp 1569139307
transform 1 0 3240 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4102
timestamp 1569139307
transform 1 0 3176 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4103
timestamp 1569139307
transform 1 0 3176 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4104
timestamp 1569139307
transform 1 0 3176 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4105
timestamp 1569139307
transform 1 0 3240 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4106
timestamp 1569139307
transform 1 0 3368 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4107
timestamp 1569139307
transform 1 0 3368 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4108
timestamp 1569139307
transform 1 0 3368 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4109
timestamp 1569139307
transform 1 0 3304 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4110
timestamp 1569139307
transform 1 0 3240 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4111
timestamp 1569139307
transform 1 0 3304 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4112
timestamp 1569139307
transform 1 0 3240 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4113
timestamp 1569139307
transform 1 0 3368 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4114
timestamp 1569139307
transform 1 0 3368 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4115
timestamp 1569139307
transform 1 0 3304 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4116
timestamp 1569139307
transform 1 0 3368 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4117
timestamp 1569139307
transform 1 0 3240 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4118
timestamp 1569139307
transform 1 0 3240 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4119
timestamp 1569139307
transform 1 0 3368 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4120
timestamp 1569139307
transform 1 0 3240 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4121
timestamp 1569139307
transform 1 0 3176 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4122
timestamp 1569139307
transform 1 0 3304 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4123
timestamp 1569139307
transform 1 0 3304 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4124
timestamp 1569139307
transform 1 0 3176 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4125
timestamp 1569139307
transform 1 0 3304 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4126
timestamp 1569139307
transform 1 0 3176 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4127
timestamp 1569139307
transform 1 0 3176 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4128
timestamp 1569139307
transform 1 0 3240 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4129
timestamp 1569139307
transform 1 0 3304 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4130
timestamp 1569139307
transform 1 0 3368 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4131
timestamp 1569139307
transform 1 0 3368 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4132
timestamp 1569139307
transform 1 0 3624 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4133
timestamp 1569139307
transform 1 0 3624 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4134
timestamp 1569139307
transform 1 0 3496 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4135
timestamp 1569139307
transform 1 0 3560 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4136
timestamp 1569139307
transform 1 0 3624 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4137
timestamp 1569139307
transform 1 0 3624 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4138
timestamp 1569139307
transform 1 0 3496 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4139
timestamp 1569139307
transform 1 0 3496 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4140
timestamp 1569139307
transform 1 0 3496 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4141
timestamp 1569139307
transform 1 0 3560 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4142
timestamp 1569139307
transform 1 0 3560 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4143
timestamp 1569139307
transform 1 0 3560 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4144
timestamp 1569139307
transform 1 0 3688 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4145
timestamp 1569139307
transform 1 0 3688 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4146
timestamp 1569139307
transform 1 0 3688 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4147
timestamp 1569139307
transform 1 0 3688 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4148
timestamp 1569139307
transform 1 0 3432 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4149
timestamp 1569139307
transform 1 0 3432 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4150
timestamp 1569139307
transform 1 0 3432 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4151
timestamp 1569139307
transform 1 0 3432 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4152
timestamp 1569139307
transform 1 0 3432 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4153
timestamp 1569139307
transform 1 0 3432 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4154
timestamp 1569139307
transform 1 0 3432 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4155
timestamp 1569139307
transform 1 0 3432 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4156
timestamp 1569139307
transform 1 0 3432 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4157
timestamp 1569139307
transform 1 0 4712 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4158
timestamp 1569139307
transform 1 0 4520 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4159
timestamp 1569139307
transform 1 0 4520 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4160
timestamp 1569139307
transform 1 0 4712 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4161
timestamp 1569139307
transform 1 0 4904 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4162
timestamp 1569139307
transform 1 0 4584 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4163
timestamp 1569139307
transform 1 0 4840 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4164
timestamp 1569139307
transform 1 0 4840 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4165
timestamp 1569139307
transform 1 0 4648 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4166
timestamp 1569139307
transform 1 0 4456 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4167
timestamp 1569139307
transform 1 0 4456 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4168
timestamp 1569139307
transform 1 0 4648 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4169
timestamp 1569139307
transform 1 0 4584 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4170
timestamp 1569139307
transform 1 0 4584 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4171
timestamp 1569139307
transform 1 0 4904 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4172
timestamp 1569139307
transform 1 0 4776 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4173
timestamp 1569139307
transform 1 0 4904 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4174
timestamp 1569139307
transform 1 0 4648 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4175
timestamp 1569139307
transform 1 0 4712 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4176
timestamp 1569139307
transform 1 0 4520 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4177
timestamp 1569139307
transform 1 0 4392 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4178
timestamp 1569139307
transform 1 0 4840 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4179
timestamp 1569139307
transform 1 0 4776 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4180
timestamp 1569139307
transform 1 0 4776 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4181
timestamp 1569139307
transform 1 0 4328 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4182
timestamp 1569139307
transform 1 0 3752 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4183
timestamp 1569139307
transform 1 0 3752 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_4184
timestamp 1569139307
transform 1 0 3752 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_4185
timestamp 1569139307
transform 1 0 3752 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_4186
timestamp 1569139307
transform 1 0 3752 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_4187
timestamp 1569139307
transform 1 0 3752 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_4188
timestamp 1569139307
transform 1 0 3752 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_4189
timestamp 1569139307
transform 1 0 3752 0 1 4200
box -8 -8 8 8
use VIA2  VIA2_4190
timestamp 1569139307
transform 1 0 3816 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4191
timestamp 1569139307
transform 1 0 3816 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_4192
timestamp 1569139307
transform 1 0 3816 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_4193
timestamp 1569139307
transform 1 0 3816 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_4194
timestamp 1569139307
transform 1 0 3816 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_4195
timestamp 1569139307
transform 1 0 3816 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_4196
timestamp 1569139307
transform 1 0 3816 0 1 4136
box -8 -8 8 8
use VIA2  VIA2_4197
timestamp 1569139307
transform 1 0 3880 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4198
timestamp 1569139307
transform 1 0 3880 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_4199
timestamp 1569139307
transform 1 0 3880 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_4200
timestamp 1569139307
transform 1 0 3880 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_4201
timestamp 1569139307
transform 1 0 3880 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_4202
timestamp 1569139307
transform 1 0 3880 0 1 4072
box -8 -8 8 8
use VIA2  VIA2_4203
timestamp 1569139307
transform 1 0 3944 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4204
timestamp 1569139307
transform 1 0 3944 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_4205
timestamp 1569139307
transform 1 0 3944 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_4206
timestamp 1569139307
transform 1 0 3944 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_4207
timestamp 1569139307
transform 1 0 3944 0 1 4008
box -8 -8 8 8
use VIA2  VIA2_4208
timestamp 1569139307
transform 1 0 4008 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_4209
timestamp 1569139307
transform 1 0 4008 0 1 3944
box -8 -8 8 8
use VIA2  VIA2_4210
timestamp 1569139307
transform 1 0 4072 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4211
timestamp 1569139307
transform 1 0 4072 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_4212
timestamp 1569139307
transform 1 0 4072 0 1 3880
box -8 -8 8 8
use VIA2  VIA2_4213
timestamp 1569139307
transform 1 0 4136 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4214
timestamp 1569139307
transform 1 0 4136 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_4215
timestamp 1569139307
transform 1 0 3752 0 1 4264
box -8 -8 8 8
use VIA2  VIA2_4216
timestamp 1569139307
transform 1 0 3752 0 1 4328
box -8 -8 8 8
use VIA2  VIA2_4217
timestamp 1569139307
transform 1 0 4200 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4218
timestamp 1569139307
transform 1 0 4264 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4219
timestamp 1569139307
transform 1 0 4008 0 1 3752
box -8 -8 8 8
use VIA2  VIA2_4220
timestamp 1569139307
transform 1 0 4008 0 1 3816
box -8 -8 8 8
use VIA2  VIA2_4221
timestamp 1569139307
transform 1 0 4264 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4222
timestamp 1569139307
transform 1 0 4328 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4223
timestamp 1569139307
transform 1 0 4264 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4224
timestamp 1569139307
transform 1 0 3752 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4225
timestamp 1569139307
transform 1 0 3752 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4226
timestamp 1569139307
transform 1 0 3752 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4227
timestamp 1569139307
transform 1 0 3752 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4228
timestamp 1569139307
transform 1 0 3752 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4229
timestamp 1569139307
transform 1 0 4264 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4230
timestamp 1569139307
transform 1 0 3752 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4231
timestamp 1569139307
transform 1 0 4328 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4232
timestamp 1569139307
transform 1 0 4328 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4233
timestamp 1569139307
transform 1 0 4328 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4234
timestamp 1569139307
transform 1 0 4328 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4235
timestamp 1569139307
transform 1 0 4328 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4236
timestamp 1569139307
transform 1 0 4328 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4237
timestamp 1569139307
transform 1 0 4328 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4238
timestamp 1569139307
transform 1 0 3752 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4239
timestamp 1569139307
transform 1 0 4264 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4240
timestamp 1569139307
transform 1 0 4264 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4241
timestamp 1569139307
transform 1 0 3752 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4242
timestamp 1569139307
transform 1 0 4264 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4243
timestamp 1569139307
transform 1 0 3752 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4244
timestamp 1569139307
transform 1 0 4264 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4245
timestamp 1569139307
transform 1 0 4456 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4246
timestamp 1569139307
transform 1 0 4520 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4247
timestamp 1569139307
transform 1 0 4520 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4248
timestamp 1569139307
transform 1 0 4520 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4249
timestamp 1569139307
transform 1 0 4520 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4250
timestamp 1569139307
transform 1 0 4584 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4251
timestamp 1569139307
transform 1 0 4584 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4252
timestamp 1569139307
transform 1 0 4584 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4253
timestamp 1569139307
transform 1 0 4392 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4254
timestamp 1569139307
transform 1 0 4456 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4255
timestamp 1569139307
transform 1 0 4648 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4256
timestamp 1569139307
transform 1 0 4776 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4257
timestamp 1569139307
transform 1 0 4776 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4258
timestamp 1569139307
transform 1 0 4648 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4259
timestamp 1569139307
transform 1 0 4776 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4260
timestamp 1569139307
transform 1 0 4776 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4261
timestamp 1569139307
transform 1 0 4776 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4262
timestamp 1569139307
transform 1 0 4840 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4263
timestamp 1569139307
transform 1 0 4840 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4264
timestamp 1569139307
transform 1 0 4840 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4265
timestamp 1569139307
transform 1 0 4840 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4266
timestamp 1569139307
transform 1 0 4840 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4267
timestamp 1569139307
transform 1 0 4840 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4268
timestamp 1569139307
transform 1 0 4904 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4269
timestamp 1569139307
transform 1 0 4904 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4270
timestamp 1569139307
transform 1 0 4904 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4271
timestamp 1569139307
transform 1 0 4904 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4272
timestamp 1569139307
transform 1 0 4712 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4273
timestamp 1569139307
transform 1 0 4904 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4274
timestamp 1569139307
transform 1 0 4904 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4275
timestamp 1569139307
transform 1 0 4712 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4276
timestamp 1569139307
transform 1 0 4712 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4277
timestamp 1569139307
transform 1 0 4712 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4278
timestamp 1569139307
transform 1 0 4968 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4279
timestamp 1569139307
transform 1 0 4968 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4280
timestamp 1569139307
transform 1 0 4968 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4281
timestamp 1569139307
transform 1 0 4968 0 1 4904
box -8 -8 8 8
use VIA2  VIA2_4282
timestamp 1569139307
transform 1 0 4712 0 1 4968
box -8 -8 8 8
use VIA2  VIA2_4283
timestamp 1569139307
transform 1 0 4776 0 1 4968
box -8 -8 8 8
use VIA2  VIA2_4284
timestamp 1569139307
transform 1 0 4840 0 1 4968
box -8 -8 8 8
use VIA2  VIA2_4285
timestamp 1569139307
transform 1 0 4904 0 1 4968
box -8 -8 8 8
use VIA2  VIA2_4286
timestamp 1569139307
transform 1 0 4968 0 1 4968
box -8 -8 8 8
use VIA2  VIA2_4287
timestamp 1569139307
transform 1 0 4392 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4288
timestamp 1569139307
transform 1 0 4392 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4289
timestamp 1569139307
transform 1 0 4392 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4290
timestamp 1569139307
transform 1 0 4392 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4291
timestamp 1569139307
transform 1 0 4392 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4292
timestamp 1569139307
transform 1 0 4392 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4293
timestamp 1569139307
transform 1 0 4392 0 1 4776
box -8 -8 8 8
use VIA2  VIA2_4294
timestamp 1569139307
transform 1 0 4392 0 1 4840
box -8 -8 8 8
use VIA2  VIA2_4295
timestamp 1569139307
transform 1 0 4456 0 1 4392
box -8 -8 8 8
use VIA2  VIA2_4296
timestamp 1569139307
transform 1 0 4456 0 1 4456
box -8 -8 8 8
use VIA2  VIA2_4297
timestamp 1569139307
transform 1 0 4456 0 1 4520
box -8 -8 8 8
use VIA2  VIA2_4298
timestamp 1569139307
transform 1 0 4456 0 1 4584
box -8 -8 8 8
use VIA2  VIA2_4299
timestamp 1569139307
transform 1 0 4456 0 1 4648
box -8 -8 8 8
use VIA2  VIA2_4300
timestamp 1569139307
transform 1 0 4456 0 1 4712
box -8 -8 8 8
use VIA2  VIA2_4301
timestamp 1569139307
transform 1 0 4456 0 1 4776
box -8 -8 8 8
<< end >>
