/* Verilog module written by vlog2Verilog (qflow) */

module ALU8_Mult(
    input [7:0] ABCmd_i,
    output [7:0] ACC_o,
    input Flag_i,
    input LoadA_i,
    input LoadB_i,
    input LoadCmd_i,
    input MulH_i,
    input MulL_i,
    input clk,
    input reset
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire [7:0] ABCmd_i ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire LoadA_i ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _899_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire BCD ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _893_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire HC ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire [3:0] alu_op ;
wire _902_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _878_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire MUL ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [7:0] ACC_o ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire [7:0] _919_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _898_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _895_ ;
wire _475_ ;
wire _284_ ;
wire [7:0] _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire _913_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire MulH_i ;
wire _719_ ;
wire _892_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _889_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _904_ ;
wire _713_ ;
wire [6:0] ACC ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire Flag_i ;
wire [6:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire LoadB_i ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire MUL_bF$buf0 ;
wire MUL_bF$buf1 ;
wire MUL_bF$buf2 ;
wire MUL_bF$buf3 ;
wire MUL_bF$buf4 ;
wire MUL_bF$buf5 ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire LoadCmd_i ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _897_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire shr ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _894_ ;
wire _474_ ;
wire _283_ ;
wire MulL_i ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _912_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _891_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _903_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire CI ;
wire CO ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire reset ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire alu_op_2_bF$buf0 ;
wire alu_op_2_bF$buf1 ;
wire alu_op_2_bF$buf2 ;
wire alu_op_2_bF$buf3 ;
wire _779_ ;
wire _359_ ;

FILL FILL_0__1241_ (
);

FILL FILL_2__1259_ (
);

FILL FILL_1__1822_ (
);

FILL FILL_1__1402_ (
);

DFFPOSX1 _1677_ (
    .D(_18_),
    .CLK(clk_bF$buf2),
    .Q(BI[0])
);

NAND3X1 _1257_ (
    .A(_343_),
    .B(_344_),
    .C(_345_),
    .Y(_349_)
);

FILL FILL_0__1717_ (
);

FILL FILL_0__1890_ (
);

FILL FILL_0__1470_ (
);

FILL FILL_0__1050_ (
);

FILL FILL_1__1631_ (
);

FILL FILL_1__1211_ (
);

OAI21X1 _1486_ (
    .A(_574_),
    .B(_571_),
    .C(_712_),
    .Y(_575_)
);

NAND2X1 _1066_ (
    .A(MUL_bF$buf5),
    .B(AI[6]),
    .Y(_158_)
);

FILL FILL_0__1526_ (
);

FILL FILL_0__1106_ (
);

FILL FILL_1__1860_ (
);

FILL FILL_1__1440_ (
);

FILL FILL_1__1020_ (
);

NAND3X1 _1295_ (
    .A(_384_),
    .B(_134_),
    .C(_385_),
    .Y(_386_)
);

FILL FILL_0__1755_ (
);

FILL FILL_0__1335_ (
);

FILL FILL_0__1564_ (
);

FILL FILL_0__1144_ (
);

FILL FILL_1__1725_ (
);

FILL FILL_1__1305_ (
);

FILL FILL_0__1793_ (
);

FILL FILL_0__1373_ (
);

FILL FILL_1__1534_ (
);

FILL FILL_1__1114_ (
);

OR2X2 _1389_ (
    .A(_477_),
    .B(_478_),
    .Y(_479_)
);

FILL FILL_0__1849_ (
);

FILL FILL_0__1429_ (
);

FILL FILL_0__1009_ (
);

FILL FILL_0__1182_ (
);

NAND2X1 _1601_ (
    .A(LoadCmd_i),
    .B(ABCmd_i[1]),
    .Y(_683_)
);

NAND3X1 _932_ (
    .A(MUL_bF$buf4),
    .B(BI[2]),
    .C(AI[1]),
    .Y(_724_)
);

FILL FILL_1__1763_ (
);

FILL FILL_1__1343_ (
);

NAND2X1 _1198_ (
    .A(AI[1]),
    .B(_289_),
    .Y(_290_)
);

FILL FILL_0__1238_ (
);

FILL FILL_1__1819_ (
);

FILL FILL86850x39750 (
);

NAND2X1 _1830_ (
    .A(_801_),
    .B(_790_),
    .Y(_802_)
);

OAI21X1 _1410_ (
    .A(_316_),
    .B(_499_),
    .C(_486_),
    .Y(_500_)
);

FILL FILL_1__1572_ (
);

FILL FILL_1__1152_ (
);

FILL FILL_0__1887_ (
);

FILL FILL_0__1467_ (
);

FILL FILL_0__1047_ (
);

FILL FILL_1__1628_ (
);

FILL FILL_1__1208_ (
);

NAND3X1 _970_ (
    .A(_58_),
    .B(_61_),
    .C(_49_),
    .Y(_62_)
);

FILL FILL_1__1381_ (
);

FILL FILL_2__1030_ (
);

FILL FILL_0__1696_ (
);

FILL FILL_0__1276_ (
);

FILL FILL_1__1857_ (
);

FILL FILL_1__1437_ (
);

FILL FILL_1__1017_ (
);

FILL FILL_1__1190_ (
);

FILL FILL_0__1085_ (
);

NAND3X1 _1504_ (
    .A(_586_),
    .B(_591_),
    .C(_585_),
    .Y(_592_)
);

FILL FILL_1__1246_ (
);

FILL FILL_2__1735_ (
);

NAND3X1 _1733_ (
    .A(_873_),
    .B(_898_),
    .C(_903_),
    .Y(_904_)
);

NAND3X1 _1313_ (
    .A(AI[5]),
    .B(_399_),
    .C(_713_),
    .Y(_404_)
);

FILL FILL_1__1895_ (
);

FILL FILL_1__1475_ (
);

FILL FILL_1__1055_ (
);

OAI21X1 _1542_ (
    .A(_628_),
    .B(_626_),
    .C(_712_),
    .Y(_629_)
);

NAND3X1 _1122_ (
    .A(_146_),
    .B(_213_),
    .C(_209_),
    .Y(_214_)
);

FILL FILL_1__1284_ (
);

FILL FILL_0__1599_ (
);

FILL FILL_0__1179_ (
);

FILL FILL_0__926_ (
);

NAND3X1 _929_ (
    .A(MUL_bF$buf4),
    .B(BI[1]),
    .C(AI[2]),
    .Y(_721_)
);

OAI21X1 _1771_ (
    .A(_743_),
    .B(_745_),
    .C(_746_),
    .Y(_747_)
);

OAI21X1 _1351_ (
    .A(_438_),
    .B(_441_),
    .C(_377_),
    .Y(_442_)
);

FILL FILL_1__1093_ (
);

FILL FILL_0__1811_ (
);

FILL FILL_2__1409_ (
);

FILL FILL_2__920_ (
);

OAI21X1 _1827_ (
    .A(_877_),
    .B(_798_),
    .C(_796_),
    .Y(_799_)
);

INVX1 _1407_ (
    .A(_486_),
    .Y(_497_)
);

FILL FILL_1__1569_ (
);

FILL FILL_1__1149_ (
);

NAND2X1 _1580_ (
    .A(_665_),
    .B(_664_),
    .Y(_666_)
);

INVX1 _1160_ (
    .A(_251_),
    .Y(_252_)
);

FILL FILL_1__942_ (
);

FILL FILL_2__1638_ (
);

FILL FILL_0__1620_ (
);

FILL FILL_0__1200_ (
);

NAND2X1 _1636_ (
    .A(ABCmd_i[0]),
    .B(LoadB_i),
    .Y(_703_)
);

OR2X2 _1216_ (
    .A(_168_),
    .B(_303_),
    .Y(_308_)
);

FILL FILL_0__964_ (
);

NOR2X1 _967_ (
    .A(_50_),
    .B(_51_),
    .Y(_59_)
);

FILL FILL_1__1798_ (
);

FILL FILL_1__1378_ (
);

INVX1 _1865_ (
    .A(_830_),
    .Y(_834_)
);

OAI21X1 _1445_ (
    .A(_401_),
    .B(_135_),
    .C(_533_),
    .Y(_534_)
);

NAND2X1 _1025_ (
    .A(_115_),
    .B(_116_),
    .Y(_117_)
);

FILL FILL_1__1187_ (
);

FILL FILL_1__980_ (
);

DFFPOSX1 _1674_ (
    .D(_15_),
    .CLK(clk_bF$buf1),
    .Q(AI[5])
);

AOI21X1 _1254_ (
    .A(_345_),
    .B(_344_),
    .C(_343_),
    .Y(_346_)
);

FILL FILL_0__1714_ (
);

INVX1 _1483_ (
    .A(AV),
    .Y(_572_)
);

INVX1 _1063_ (
    .A(_154_),
    .Y(_155_)
);

FILL FILL_0__1523_ (
);

FILL FILL_0__1103_ (
);

AOI21X1 _1539_ (
    .A(_617_),
    .B(_624_),
    .C(_625_),
    .Y(_626_)
);

NAND3X1 _1119_ (
    .A(_203_),
    .B(_205_),
    .C(_206_),
    .Y(_211_)
);

INVX1 _1292_ (
    .A(_382_),
    .Y(_383_)
);

FILL FILL_0__1752_ (
);

FILL FILL_0__1332_ (
);

OAI21X1 _1768_ (
    .A(alu_op_2_bF$buf3),
    .B(BI[3]),
    .C(_858_),
    .Y(_744_)
);

NAND3X1 _1348_ (
    .A(_429_),
    .B(_422_),
    .C(_432_),
    .Y(_439_)
);

FILL FILL_0__1808_ (
);

FILL FILL_0__1561_ (
);

FILL FILL_2__1579_ (
);

FILL FILL_0__1141_ (
);

FILL FILL_1__1722_ (
);

FILL FILL_1__1302_ (
);

AOI21X1 _1577_ (
    .A(_405_),
    .B(_134_),
    .C(_634_),
    .Y(_663_)
);

OAI21X1 _1157_ (
    .A(_247_),
    .B(_248_),
    .C(_246_),
    .Y(_249_)
);

FILL FILL_1__939_ (
);

FILL FILL86550x50550 (
);

FILL FILL_0__1617_ (
);

FILL FILL_0__1790_ (
);

FILL FILL_0__1370_ (
);

FILL FILL_1__1531_ (
);

FILL FILL_1__1111_ (
);

INVX1 _1386_ (
    .A(_475_),
    .Y(_476_)
);

FILL FILL_0__1846_ (
);

FILL FILL_0__1426_ (
);

FILL FILL_0__1006_ (
);

FILL FILL_1__1760_ (
);

FILL FILL_1__1340_ (
);

OAI21X1 _1195_ (
    .A(_207_),
    .B(_186_),
    .C(_206_),
    .Y(_287_)
);

FILL FILL_1__977_ (
);

FILL FILL_0__1235_ (
);

FILL FILL_1__1816_ (
);

FILL FILL_0__999_ (
);

FILL FILL_0__1884_ (
);

FILL FILL_0__1464_ (
);

FILL FILL_0__1044_ (
);

FILL FILL_1__1625_ (
);

FILL FILL_1__1205_ (
);

FILL FILL_0__1693_ (
);

FILL FILL_0__1273_ (
);

FILL FILL_1__1854_ (
);

FILL FILL_1__1434_ (
);

FILL FILL_1__1014_ (
);

NOR3X1 _1289_ (
    .A(_329_),
    .B(_330_),
    .C(_301_),
    .Y(_380_)
);

FILL FILL_0__1749_ (
);

FILL FILL_0__1329_ (
);

FILL FILL_0__1082_ (
);

INVX1 _1501_ (
    .A(_182_),
    .Y(_589_)
);

FILL FILL_1__1243_ (
);

AOI21X1 _1098_ (
    .A(_188_),
    .B(_189_),
    .C(_187_),
    .Y(_190_)
);

FILL FILL_0__1558_ (
);

FILL FILL_0__1138_ (
);

FILL FILL_1__1719_ (
);

OAI21X1 _1730_ (
    .A(_870_),
    .B(_862_),
    .C(BI[0]),
    .Y(_901_)
);

INVX1 _1310_ (
    .A(AI[5]),
    .Y(_401_)
);

FILL FILL_1__1892_ (
);

FILL FILL_1__1472_ (
);

FILL FILL_1__1052_ (
);

FILL FILL_0__1787_ (
);

FILL FILL_0__1367_ (
);

FILL FILL_1__1528_ (
);

FILL FILL_1__1108_ (
);

FILL FILL_1__1281_ (
);

FILL FILL86850x25350 (
);

FILL FILL_2__1350_ (
);

FILL FILL_0__1596_ (
);

FILL FILL_0__1176_ (
);

FILL FILL_0__923_ (
);

NAND2X1 _926_ (
    .A(BI[3]),
    .B(_717_),
    .Y(_718_)
);

FILL FILL_1__1757_ (
);

FILL FILL_1__1337_ (
);

FILL FILL_1__1090_ (
);

FILL FILL_2__1826_ (
);

OAI22X1 _1824_ (
    .A(_868_),
    .B(_791_),
    .C(_795_),
    .D(_794_),
    .Y(_796_)
);

NAND3X1 _1404_ (
    .A(_490_),
    .B(_493_),
    .C(_459_),
    .Y(_494_)
);

FILL FILL_1__1566_ (
);

FILL FILL_1__1146_ (
);

OAI21X1 _1633_ (
    .A(LoadA_i),
    .B(_480_),
    .C(_701_),
    .Y(_16_)
);

AND2X2 _1213_ (
    .A(_168_),
    .B(_303_),
    .Y(_305_)
);

FILL FILL_0__961_ (
);

NAND3X1 _964_ (
    .A(MUL_bF$buf4),
    .B(BI[2]),
    .C(AI[3]),
    .Y(_56_)
);

FILL FILL_1__1795_ (
);

FILL FILL_1__1375_ (
);

FILL FILL_2__1024_ (
);

NAND2X1 _1862_ (
    .A(_830_),
    .B(_790_),
    .Y(_831_)
);

OAI21X1 _1442_ (
    .A(_475_),
    .B(_484_),
    .C(_479_),
    .Y(_531_)
);

OAI21X1 _1022_ (
    .A(_111_),
    .B(_113_),
    .C(_108_),
    .Y(_114_)
);

FILL FILL_1__1184_ (
);

FILL FILL_0__1499_ (
);

FILL FILL_0__1079_ (
);

DFFPOSX1 _1671_ (
    .D(_12_),
    .CLK(clk_bF$buf3),
    .Q(AI[2])
);

INVX1 _1251_ (
    .A(_286_),
    .Y(_343_)
);

FILL FILL_0__1711_ (
);

INVX1 _1727_ (
    .A(_876_),
    .Y(_898_)
);

NAND3X1 _1307_ (
    .A(MUL_bF$buf3),
    .B(AI[5]),
    .C(BI[4]),
    .Y(_398_)
);

FILL FILL_1__1889_ (
);

FILL FILL_1__1469_ (
);

FILL FILL_1__1049_ (
);

NAND2X1 _1480_ (
    .A(_262_),
    .B(_273_),
    .Y(_569_)
);

NOR2X1 _1060_ (
    .A(_150_),
    .B(_151_),
    .Y(_152_)
);

FILL FILL_0__1520_ (
);

FILL FILL_0__1100_ (
);

FILL FILL_2__1291_ (
);

OAI21X1 _1536_ (
    .A(_712_),
    .B(_616_),
    .C(_623_),
    .Y(_0_[4])
);

NAND3X1 _1116_ (
    .A(_205_),
    .B(_206_),
    .C(_207_),
    .Y(_208_)
);

FILL FILL_1__1698_ (
);

FILL FILL_1__1278_ (
);

FILL FILL85950x10950 (
);

AOI22X1 _1765_ (
    .A(_862_),
    .B(BI[3]),
    .C(_740_),
    .D(_863_),
    .Y(_741_)
);

AOI21X1 _1345_ (
    .A(_434_),
    .B(_435_),
    .C(_395_),
    .Y(_436_)
);

FILL FILL_1__1087_ (
);

FILL FILL_0__1805_ (
);

AOI21X1 _1574_ (
    .A(_613_),
    .B(_614_),
    .C(_659_),
    .Y(_660_)
);

NAND3X1 _1154_ (
    .A(_244_),
    .B(_245_),
    .C(_235_),
    .Y(_246_)
);

FILL FILL_1__936_ (
);

FILL FILL_0__1614_ (
);

FILL FILL_0__958_ (
);

OAI21X1 _1383_ (
    .A(_471_),
    .B(_472_),
    .C(_460_),
    .Y(_473_)
);

FILL FILL_0__1843_ (
);

FILL FILL_0__1423_ (
);

FILL FILL_0__1003_ (
);

OAI21X1 _1859_ (
    .A(_799_),
    .B(_816_),
    .C(_815_),
    .Y(_828_)
);

AOI21X1 _1439_ (
    .A(_491_),
    .B(_488_),
    .C(_487_),
    .Y(_528_)
);

NOR2X1 _1019_ (
    .A(_109_),
    .B(_110_),
    .Y(_111_)
);

AOI21X1 _1192_ (
    .A(_209_),
    .B(_146_),
    .C(_216_),
    .Y(_284_)
);

FILL FILL_1__974_ (
);

FILL FILL_0__1652_ (
);

FILL FILL_0__1232_ (
);

FILL FILL_1__1813_ (
);

DFFSR _1668_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[7]),
    .CLK(clk_bF$buf4),
    .Q(_919_[7])
);

AOI21X1 _1248_ (
    .A(_327_),
    .B(_331_),
    .C(_300_),
    .Y(_340_)
);

FILL FILL_0__996_ (
);

AOI21X1 _999_ (
    .A(_55_),
    .B(_57_),
    .C(_59_),
    .Y(_91_)
);

FILL FILL_0__1708_ (
);

FILL FILL_0__1881_ (
);

FILL FILL_0__1461_ (
);

FILL FILL_0__1041_ (
);

FILL FILL_1__1622_ (
);

FILL FILL_1__1202_ (
);

BUFX2 _1897_ (
    .A(_919_[7]),
    .Y(ACC_o[7])
);

INVX1 _1477_ (
    .A(_560_),
    .Y(_566_)
);

AOI21X1 _1057_ (
    .A(_100_),
    .B(_97_),
    .C(_94_),
    .Y(_149_)
);

FILL FILL_0__1517_ (
);

FILL FILL_0__1690_ (
);

FILL FILL_0__1270_ (
);

FILL FILL_1__1851_ (
);

FILL FILL_1__1431_ (
);

FILL FILL_1__1011_ (
);

AOI21X1 _1286_ (
    .A(_286_),
    .B(_341_),
    .C(_376_),
    .Y(_377_)
);

FILL FILL86850x7350 (
);

FILL FILL_2__1500_ (
);

FILL FILL_0__1746_ (
);

FILL FILL_0__1326_ (
);

FILL FILL_1__1240_ (
);

AOI21X1 _1095_ (
    .A(_119_),
    .B(_102_),
    .C(_122_),
    .Y(_187_)
);

FILL FILL_0__1555_ (
);

FILL FILL_0__1135_ (
);

FILL FILL_1__1716_ (
);

FILL FILL_0__1784_ (
);

FILL FILL_0__1364_ (
);

FILL FILL_1__1525_ (
);

FILL FILL_1__1105_ (
);

FILL FILL_0__1593_ (
);

FILL FILL_0__1173_ (
);

FILL FILL_0__920_ (
);

INVX1 _923_ (
    .A(MUL_bF$buf3),
    .Y(_715_)
);

FILL FILL_1__1754_ (
);

FILL FILL_1__1334_ (
);

FILL FILL86850x46950 (
);

INVX1 _1189_ (
    .A(_280_),
    .Y(_281_)
);

FILL FILL_0__1649_ (
);

FILL FILL_0__1229_ (
);

NAND2X1 _1821_ (
    .A(AI[6]),
    .B(_792_),
    .Y(_793_)
);

AND2X2 _1401_ (
    .A(_473_),
    .B(_470_),
    .Y(_491_)
);

FILL FILL_1__1563_ (
);

FILL FILL_1__1143_ (
);

FILL FILL_0__1878_ (
);

FILL FILL_0__1458_ (
);

FILL FILL_0__1038_ (
);

FILL FILL_1__1619_ (
);

NAND2X1 _1630_ (
    .A(ABCmd_i[5]),
    .B(LoadA_i),
    .Y(_700_)
);

NAND3X1 _1210_ (
    .A(MUL_bF$buf2),
    .B(AI[3]),
    .C(BI[5]),
    .Y(_302_)
);

INVX1 _961_ (
    .A(BI[0]),
    .Y(_53_)
);

FILL FILL_1__1792_ (
);

FILL FILL_1__1372_ (
);

FILL FILL_0__1687_ (
);

FILL FILL_0__1267_ (
);

FILL FILL_1__1848_ (
);

FILL FILL_1__1428_ (
);

FILL FILL_1__1008_ (
);

FILL FILL_1__1181_ (
);

FILL FILL_0__1496_ (
);

FILL FILL_0__1076_ (
);

FILL FILL_1_BUFX2_insert5 (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

FILL FILL_1__1237_ (
);

OAI21X1 _1724_ (
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_894_),
    .Y(_895_)
);

NAND2X1 _1304_ (
    .A(_390_),
    .B(_394_),
    .Y(_395_)
);

FILL FILL_1__1886_ (
);

FILL FILL_1__1466_ (
);

FILL FILL_1__1046_ (
);

FILL FILL_2__1115_ (
);

OAI21X1 _1533_ (
    .A(CO),
    .B(_364_),
    .C(_365_),
    .Y(_621_)
);

NAND3X1 _1113_ (
    .A(_189_),
    .B(_187_),
    .C(_188_),
    .Y(_205_)
);

FILL FILL_1__1695_ (
);

FILL FILL_1__1275_ (
);

FILL FILL_2__1344_ (
);

NAND2X1 _1762_ (
    .A(shr),
    .B(AI[4]),
    .Y(_738_)
);

AOI21X1 _1342_ (
    .A(_426_),
    .B(_428_),
    .C(_423_),
    .Y(_433_)
);

FILL FILL_1__1084_ (
);

FILL FILL_0__1802_ (
);

FILL FILL_0__1399_ (
);

OAI21X1 _1818_ (
    .A(_784_),
    .B(_787_),
    .C(_783_),
    .Y(_790_)
);

OAI21X1 _1571_ (
    .A(_655_),
    .B(_654_),
    .C(_656_),
    .Y(_657_)
);

INVX1 _1151_ (
    .A(_242_),
    .Y(_243_)
);

FILL FILL_1__933_ (
);

FILL FILL_0__1611_ (
);

OAI21X1 _1627_ (
    .A(LoadA_i),
    .B(_387_),
    .C(_698_),
    .Y(_13_)
);

OAI21X1 _1207_ (
    .A(_297_),
    .B(_298_),
    .C(_290_),
    .Y(_299_)
);

FILL FILL_0__955_ (
);

NAND3X1 _958_ (
    .A(MUL_bF$buf4),
    .B(BI[1]),
    .C(AI[4]),
    .Y(_50_)
);

FILL FILL_1__1789_ (
);

FILL FILL_1__1369_ (
);

NAND3X1 _1380_ (
    .A(_461_),
    .B(_469_),
    .C(_467_),
    .Y(_470_)
);

FILL FILL_0__1840_ (
);

FILL FILL_0__1420_ (
);

FILL FILL_0__1000_ (
);

AND2X2 _1856_ (
    .A(_825_),
    .B(_822_),
    .Y(AZ)
);

AOI21X1 _1436_ (
    .A(_457_),
    .B(_505_),
    .C(_524_),
    .Y(_525_)
);

INVX1 _1016_ (
    .A(_107_),
    .Y(_108_)
);

FILL FILL_1__1598_ (
);

FILL FILL_1__1178_ (
);

FILL FILL_1__971_ (
);

FILL FILL_1__1810_ (
);

DFFSR _1665_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[4]),
    .CLK(clk_bF$buf4),
    .Q(_919_[4])
);

NAND3X1 _1245_ (
    .A(_332_),
    .B(_336_),
    .C(_287_),
    .Y(_337_)
);

FILL FILL_0__993_ (
);

AOI21X1 _996_ (
    .A(_86_),
    .B(_80_),
    .C(_48_),
    .Y(_88_)
);

FILL FILL_0__1705_ (
);

FILL FILL_2__1056_ (
);

BUFX2 _1894_ (
    .A(_919_[4]),
    .Y(ACC_o[4])
);

NOR2X1 _1474_ (
    .A(_360_),
    .B(_448_),
    .Y(_563_)
);

INVX1 _1054_ (
    .A(_132_),
    .Y(_146_)
);

FILL FILL_0__1514_ (
);

FILL FILL_2__1285_ (
);

NAND2X1 _1283_ (
    .A(_373_),
    .B(_371_),
    .Y(_374_)
);

FILL FILL_0__1743_ (
);

FILL FILL_0__1323_ (
);

INVX1 _1759_ (
    .A(_735_),
    .Y(ACC[2])
);

NAND3X1 _1339_ (
    .A(_422_),
    .B(_429_),
    .C(_381_),
    .Y(_430_)
);

NAND2X1 _1092_ (
    .A(_181_),
    .B(_183_),
    .Y(_184_)
);

FILL FILL_0__1552_ (
);

FILL FILL_0__1132_ (
);

FILL FILL_1__1713_ (
);

AOI21X1 _1568_ (
    .A(_653_),
    .B(_357_),
    .C(_281_),
    .Y(_654_)
);

NAND2X1 _1148_ (
    .A(_237_),
    .B(_239_),
    .Y(_240_)
);

FILL FILL_0__1608_ (
);

FILL FILL_0__1781_ (
);

FILL FILL_0__1361_ (
);

FILL FILL_1__1522_ (
);

FILL FILL_1__1102_ (
);

OAI21X1 _1797_ (
    .A(_751_),
    .B(_771_),
    .C(_757_),
    .Y(HC)
);

OAI21X1 _1377_ (
    .A(_462_),
    .B(_407_),
    .C(_466_),
    .Y(_467_)
);

FILL FILL_0__1837_ (
);

FILL FILL_0__1417_ (
);

FILL FILL_2__946_ (
);

FILL FILL_0__1590_ (
);

FILL FILL_0__1170_ (
);

INVX2 _920_ (
    .A(MulH_i),
    .Y(_712_)
);

FILL FILL_1__1751_ (
);

FILL FILL_1__1331_ (
);

NAND3X1 _1186_ (
    .A(_719_),
    .B(_87_),
    .C(_232_),
    .Y(_278_)
);

FILL FILL_1__968_ (
);

FILL FILL_2__1820_ (
);

FILL FILL85950x18150 (
);

FILL FILL_0__1646_ (
);

FILL FILL_0__1226_ (
);

FILL FILL_1__1807_ (
);

FILL FILL_1__1560_ (
);

FILL FILL_1__1140_ (
);

FILL FILL_0__1875_ (
);

FILL FILL_0__1455_ (
);

FILL FILL_0__1035_ (
);

FILL FILL_1__1616_ (
);

FILL FILL_0__1264_ (
);

FILL FILL_1__1845_ (
);

FILL FILL_1__1425_ (
);

FILL FILL_1__1005_ (
);

FILL FILL_0__1493_ (
);

FILL FILL_0__1073_ (
);

FILL FILL_1__1234_ (
);

NAND3X1 _1089_ (
    .A(_167_),
    .B(_171_),
    .C(_175_),
    .Y(_181_)
);

FILL FILL_0__1549_ (
);

FILL FILL_0__1129_ (
);

OAI21X1 _1721_ (
    .A(alu_op_2_bF$buf0),
    .B(BI[1]),
    .C(_858_),
    .Y(_892_)
);

NOR2X1 _1301_ (
    .A(_391_),
    .B(_388_),
    .Y(_392_)
);

FILL FILL_1__1883_ (
);

FILL FILL_1__1463_ (
);

FILL FILL_1__1043_ (
);

FILL FILL_0__1778_ (
);

FILL FILL_0__1358_ (
);

FILL FILL_1__1519_ (
);

FILL FILL86850x32550 (
);

OAI21X1 _1530_ (
    .A(_275_),
    .B(_252_),
    .C(_274_),
    .Y(_618_)
);

NAND3X1 _1110_ (
    .A(_191_),
    .B(_201_),
    .C(_200_),
    .Y(_202_)
);

FILL FILL_1__1692_ (
);

FILL FILL_1__1272_ (
);

FILL FILL_2__1761_ (
);

FILL FILL_0__1587_ (
);

FILL FILL_0__1167_ (
);

FILL FILL_1__1748_ (
);

FILL FILL_1__1328_ (
);

FILL FILL_1__1081_ (
);

FILL FILL_0__1396_ (
);

NAND2X1 _1815_ (
    .A(_784_),
    .B(_787_),
    .Y(_788_)
);

FILL FILL_1__1557_ (
);

FILL FILL_1__1137_ (
);

FILL FILL_1__930_ (
);

NAND2X1 _1624_ (
    .A(ABCmd_i[2]),
    .B(LoadA_i),
    .Y(_697_)
);

NAND3X1 _1204_ (
    .A(_291_),
    .B(_295_),
    .C(_294_),
    .Y(_296_)
);

FILL FILL_0__952_ (
);

AOI21X1 _955_ (
    .A(_39_),
    .B(_41_),
    .C(_29_),
    .Y(_47_)
);

FILL FILL_1__1786_ (
);

FILL FILL_1__1366_ (
);

FILL FILL_2__1435_ (
);

NOR2X1 _1853_ (
    .A(_801_),
    .B(_790_),
    .Y(_823_)
);

NAND2X1 _1433_ (
    .A(_712_),
    .B(_522_),
    .Y(_523_)
);

OAI21X1 _1013_ (
    .A(_94_),
    .B(_95_),
    .C(_96_),
    .Y(_105_)
);

FILL FILL_1__1595_ (
);

FILL FILL_1__1175_ (
);

DFFSR _1662_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[1]),
    .CLK(clk_bF$buf4),
    .Q(_919_[1])
);

NAND3X1 _1242_ (
    .A(_322_),
    .B(_326_),
    .C(_328_),
    .Y(_334_)
);

FILL FILL_0__990_ (
);

NAND2X1 _993_ (
    .A(_84_),
    .B(_83_),
    .Y(_85_)
);

FILL FILL_0__1702_ (
);

FILL FILL_0__1299_ (
);

NOR2X1 _1718_ (
    .A(alu_op[0]),
    .B(_888_),
    .Y(_889_)
);

BUFX2 _1891_ (
    .A(_919_[1]),
    .Y(ACC_o[1])
);

NAND2X1 _1471_ (
    .A(_559_),
    .B(_556_),
    .Y(_560_)
);

NAND2X1 _1051_ (
    .A(_142_),
    .B(_139_),
    .Y(_143_)
);

FILL FILL_0__1511_ (
);

FILL FILL_2__1109_ (
);

NAND3X1 _1527_ (
    .A(_603_),
    .B(_614_),
    .C(_613_),
    .Y(_615_)
);

NAND3X1 _1107_ (
    .A(_192_),
    .B(_198_),
    .C(_195_),
    .Y(_199_)
);

FILL FILL_1__1689_ (
);

FILL FILL_1__1269_ (
);

OAI21X1 _1280_ (
    .A(_267_),
    .B(_370_),
    .C(MulL_i),
    .Y(_371_)
);

FILL FILL_0__1740_ (
);

FILL FILL_0__1320_ (
);

OAI21X1 _1756_ (
    .A(_918_),
    .B(_727_),
    .C(_732_),
    .Y(_733_)
);

AOI21X1 _1336_ (
    .A(_323_),
    .B(_325_),
    .C(_424_),
    .Y(_427_)
);

FILL FILL_1__1498_ (
);

FILL FILL_1__1078_ (
);

FILL FILL_1__1710_ (
);

NAND3X1 _1565_ (
    .A(MulH_i),
    .B(_647_),
    .C(_651_),
    .Y(_652_)
);

INVX1 _1145_ (
    .A(_236_),
    .Y(_237_)
);

FILL FILL_1__927_ (
);

FILL FILL_0__1605_ (
);

FILL FILL_2__1376_ (
);

FILL FILL_0__949_ (
);

NOR2X1 _1794_ (
    .A(_730_),
    .B(_911_),
    .Y(_769_)
);

NOR2X1 _1374_ (
    .A(_715_),
    .B(_463_),
    .Y(_464_)
);

FILL FILL_0__1834_ (
);

FILL FILL_0__1414_ (
);

AOI21X1 _1183_ (
    .A(_250_),
    .B(_234_),
    .C(_249_),
    .Y(_275_)
);

FILL FILL_1__965_ (
);

FILL FILL_0__1643_ (
);

FILL FILL_0__1223_ (
);

FILL FILL_1__1804_ (
);

DFFPOSX1 _1659_ (
    .D(_8_),
    .CLK(clk_bF$buf2),
    .Q(BCD)
);

OAI21X1 _1239_ (
    .A(_329_),
    .B(_330_),
    .C(_328_),
    .Y(_331_)
);

FILL FILL_0__987_ (
);

FILL FILL85950x39750 (
);

FILL FILL_0__1872_ (
);

FILL FILL_0__1452_ (
);

FILL FILL_0__1032_ (
);

FILL FILL_1__1613_ (
);

NAND2X1 _1888_ (
    .A(CO),
    .B(_855_),
    .Y(_856_)
);

AOI21X1 _1468_ (
    .A(_490_),
    .B(_493_),
    .C(_495_),
    .Y(_557_)
);

NAND3X1 _1048_ (
    .A(_128_),
    .B(_127_),
    .C(_126_),
    .Y(_140_)
);

FILL FILL_0__1508_ (
);

FILL FILL_0__1261_ (
);

FILL FILL_1__1842_ (
);

FILL FILL_1__1422_ (
);

FILL FILL_1__1002_ (
);

INVX1 _1697_ (
    .A(BI[0]),
    .Y(_869_)
);

NAND2X1 _1277_ (
    .A(_712_),
    .B(_368_),
    .Y(_369_)
);

FILL FILL_0__1737_ (
);

FILL FILL_0__1317_ (
);

FILL FILL86550x10950 (
);

FILL FILL_0__1490_ (
);

FILL FILL_0__1070_ (
);

FILL FILL_1__1651_ (
);

FILL FILL_1__1231_ (
);

NAND3X1 _1086_ (
    .A(_161_),
    .B(_177_),
    .C(_165_),
    .Y(_178_)
);

FILL FILL_0__1546_ (
);

FILL FILL_0__1126_ (
);

FILL FILL_1__1707_ (
);

FILL FILL_1__1880_ (
);

FILL FILL_1__1460_ (
);

FILL FILL_1__1040_ (
);

FILL FILL_0__1775_ (
);

FILL FILL_0__1355_ (
);

FILL FILL_1__1516_ (
);

FILL FILL_0__1584_ (
);

FILL FILL_0__1164_ (
);

FILL FILL_1__1745_ (
);

FILL FILL_1__1325_ (
);

FILL FILL_0__1393_ (
);

INVX1 _1812_ (
    .A(_784_),
    .Y(_785_)
);

FILL FILL_1__1554_ (
);

FILL FILL_1__1134_ (
);

FILL FILL_0__1869_ (
);

FILL FILL_0__1449_ (
);

FILL FILL_0__1029_ (
);

OAI21X1 _1621_ (
    .A(LoadA_i),
    .B(_43_),
    .C(_695_),
    .Y(_10_)
);

AOI22X1 _1201_ (
    .A(_116_),
    .B(_174_),
    .C(_171_),
    .D(_167_),
    .Y(_293_)
);

NAND2X1 _952_ (
    .A(MUL_bF$buf0),
    .B(BI[4]),
    .Y(_44_)
);

FILL FILL_1__1783_ (
);

FILL FILL_1__1363_ (
);

FILL FILL_2__1852_ (
);

FILL FILL_0__1258_ (
);

FILL FILL_1__1839_ (
);

FILL FILL_1__1419_ (
);

NOR2X1 _1850_ (
    .A(ACC[0]),
    .B(_770_),
    .Y(_820_)
);

NOR2X1 _1430_ (
    .A(Flag_i),
    .B(ACC[2]),
    .Y(_520_)
);

NAND3X1 _1010_ (
    .A(_91_),
    .B(_98_),
    .C(_101_),
    .Y(_102_)
);

FILL FILL_1__1592_ (
);

FILL FILL_1__1172_ (
);

FILL FILL_0__1487_ (
);

FILL FILL_0__1067_ (
);

FILL FILL_1__1648_ (
);

FILL FILL_1__1228_ (
);

AOI21X1 _990_ (
    .A(_58_),
    .B(_61_),
    .C(_49_),
    .Y(_82_)
);

FILL FILL_2__1050_ (
);

FILL FILL_0__1296_ (
);

NAND3X1 _1715_ (
    .A(AI[1]),
    .B(BI[1]),
    .C(_864_),
    .Y(_886_)
);

FILL FILL_1__1877_ (
);

FILL FILL_1__1457_ (
);

FILL FILL_1__1037_ (
);

FILL FILL86250x7350 (
);

NOR2X1 _1524_ (
    .A(_560_),
    .B(_512_),
    .Y(_612_)
);

NAND2X1 _1104_ (
    .A(AI[1]),
    .B(_134_),
    .Y(_196_)
);

FILL FILL_1__1686_ (
);

FILL FILL_1__1266_ (
);

FILL FILL_2__1755_ (
);

MUX2X1 _1753_ (
    .A(_729_),
    .B(_728_),
    .S(_918_),
    .Y(_730_)
);

AND2X2 _1333_ (
    .A(_318_),
    .B(_320_),
    .Y(_424_)
);

FILL FILL_1__1495_ (
);

FILL FILL_1__1075_ (
);

AOI21X1 _1809_ (
    .A(alu_op_2_bF$buf3),
    .B(BI[5]),
    .C(_781_),
    .Y(_782_)
);

AOI21X1 _1562_ (
    .A(_613_),
    .B(_614_),
    .C(_603_),
    .Y(_649_)
);

NAND3X1 _1142_ (
    .A(_42_),
    .B(_228_),
    .C(_227_),
    .Y(_234_)
);

FILL FILL_1__924_ (
);

FILL FILL_0__1602_ (
);

FILL FILL_0__1199_ (
);

NAND2X1 _1618_ (
    .A(LoadCmd_i),
    .B(ABCmd_i[7]),
    .Y(_694_)
);

FILL FILL_0__946_ (
);

OAI21X1 _949_ (
    .A(_34_),
    .B(_40_),
    .C(_30_),
    .Y(_41_)
);

OAI21X1 _1791_ (
    .A(_877_),
    .B(_765_),
    .C(_763_),
    .Y(_766_)
);

INVX1 _1371_ (
    .A(_460_),
    .Y(_461_)
);

FILL FILL_0__1831_ (
);

FILL FILL_0__1411_ (
);

FILL FILL_2__1429_ (
);

FILL FILL_2__940_ (
);

OAI21X1 _1847_ (
    .A(_805_),
    .B(_806_),
    .C(_817_),
    .Y(_818_)
);

AND2X2 _1427_ (
    .A(_264_),
    .B(_269_),
    .Y(_517_)
);

OR2X2 _1007_ (
    .A(_92_),
    .B(_93_),
    .Y(_99_)
);

FILL FILL_1__1589_ (
);

FILL FILL_1__1169_ (
);

INVX1 _1180_ (
    .A(_246_),
    .Y(_272_)
);

FILL FILL_1__962_ (
);

FILL FILL_0__1640_ (
);

FILL FILL_0__1220_ (
);

FILL FILL_1__1801_ (
);

DFFPOSX1 _1656_ (
    .D(_5_),
    .CLK(clk_bF$buf3),
    .Q(alu_op[3])
);

OAI21X1 _1236_ (
    .A(_184_),
    .B(_179_),
    .C(_165_),
    .Y(_328_)
);

FILL FILL_0__984_ (
);

NAND2X1 _987_ (
    .A(_78_),
    .B(_76_),
    .Y(_79_)
);

FILL FILL_1__1398_ (
);

FILL FILL_1__1610_ (
);

NAND3X1 _1885_ (
    .A(_850_),
    .B(_819_),
    .C(_818_),
    .Y(_853_)
);

NAND3X1 _1465_ (
    .A(_526_),
    .B(_552_),
    .C(_553_),
    .Y(_554_)
);

NAND2X1 _1045_ (
    .A(_136_),
    .B(_132_),
    .Y(_137_)
);

FILL FILL_0__1505_ (
);

FILL FILL_2__1696_ (
);

NAND2X1 _1694_ (
    .A(AI[0]),
    .B(alu_op[1]),
    .Y(_866_)
);

OAI21X1 _1274_ (
    .A(HC),
    .B(_364_),
    .C(_365_),
    .Y(_366_)
);

FILL FILL_0__1734_ (
);

FILL FILL_0__1314_ (
);

NAND2X1 _1083_ (
    .A(_116_),
    .B(_174_),
    .Y(_175_)
);

FILL FILL_0__1543_ (
);

FILL FILL_0__1123_ (
);

FILL FILL_1__1704_ (
);

NAND2X1 _1559_ (
    .A(_644_),
    .B(_645_),
    .Y(_646_)
);

NAND3X1 _1139_ (
    .A(_66_),
    .B(_62_),
    .C(_85_),
    .Y(_231_)
);

FILL FILL_0__1772_ (
);

FILL FILL_0__1352_ (
);

FILL FILL_1__1513_ (
);

OAI21X1 _1788_ (
    .A(_762_),
    .B(_761_),
    .C(_758_),
    .Y(_763_)
);

INVX1 _1368_ (
    .A(_457_),
    .Y(_458_)
);

FILL FILL_0__1828_ (
);

FILL FILL_0__1408_ (
);

FILL FILL_0__1581_ (
);

FILL FILL_0__1161_ (
);

FILL FILL85950x25350 (
);

FILL FILL_1__1742_ (
);

FILL FILL_1__1322_ (
);

INVX1 _1597_ (
    .A(alu_op[0]),
    .Y(_680_)
);

OAI21X1 _1177_ (
    .A(_268_),
    .B(_67_),
    .C(_263_),
    .Y(_269_)
);

FILL FILL_1__959_ (
);

FILL FILL_0__1637_ (
);

FILL FILL_0__1217_ (
);

FILL FILL_0__1390_ (
);

FILL FILL_1__1551_ (
);

FILL FILL_1__1131_ (
);

FILL FILL_2__1200_ (
);

FILL FILL_0__1866_ (
);

FILL FILL_0__1446_ (
);

FILL FILL_0__1026_ (
);

FILL FILL_1__1607_ (
);

FILL FILL_1__1780_ (
);

FILL FILL_1__1360_ (
);

FILL FILL_1__997_ (
);

FILL FILL_0__1255_ (
);

FILL FILL_1__1836_ (
);

FILL FILL_1__1416_ (
);

FILL FILL_0__1484_ (
);

FILL FILL_0__1064_ (
);

FILL FILL_1__1645_ (
);

FILL FILL_1__1225_ (
);

FILL FILL_0__1293_ (
);

NOR2X1 _1712_ (
    .A(_876_),
    .B(_874_),
    .Y(_883_)
);

FILL FILL_1__1874_ (
);

FILL FILL_1__1454_ (
);

FILL FILL_1__1034_ (
);

FILL FILL_0__1769_ (
);

FILL FILL_0__1349_ (
);

OAI21X1 _1521_ (
    .A(_453_),
    .B(_359_),
    .C(_608_),
    .Y(_609_)
);

AOI21X1 _1101_ (
    .A(_108_),
    .B(_112_),
    .C(_111_),
    .Y(_193_)
);

FILL FILL_1__1263_ (
);

FILL FILL_0__1578_ (
);

FILL FILL_0__1158_ (
);

FILL FILL_1__1739_ (
);

FILL FILL_1__1319_ (
);

AOI21X1 _1750_ (
    .A(alu_op_2_bF$buf1),
    .B(BI[2]),
    .C(_726_),
    .Y(_727_)
);

AOI21X1 _1330_ (
    .A(_409_),
    .B(_413_),
    .C(_420_),
    .Y(_421_)
);

FILL FILL86550x18150 (
);

FILL FILL_1__1492_ (
);

FILL FILL_1__1072_ (
);

FILL FILL_2__1141_ (
);

FILL FILL_0__1387_ (
);

OAI21X1 _1806_ (
    .A(AI[5]),
    .B(_776_),
    .C(_868_),
    .Y(_779_)
);

FILL FILL_1__1548_ (
);

FILL FILL_1__1128_ (
);

FILL FILL_1__921_ (
);

FILL FILL_2__1370_ (
);

FILL FILL_0__1196_ (
);

INVX1 _1615_ (
    .A(BCD),
    .Y(_692_)
);

FILL FILL_0__943_ (
);

OAI21X1 _946_ (
    .A(_36_),
    .B(_37_),
    .C(_32_),
    .Y(_38_)
);

FILL FILL_1__1777_ (
);

FILL FILL_1__1357_ (
);

FILL FILL_2__1846_ (
);

OAI21X1 _1844_ (
    .A(_877_),
    .B(_814_),
    .C(_812_),
    .Y(_815_)
);

NAND2X1 _1424_ (
    .A(_513_),
    .B(_456_),
    .Y(_514_)
);

NAND3X1 _1004_ (
    .A(MUL_bF$buf1),
    .B(BI[2]),
    .C(AI[4]),
    .Y(_96_)
);

FILL FILL_1__1586_ (
);

FILL FILL_1__1166_ (
);

DFFPOSX1 _1653_ (
    .D(_2_),
    .CLK(clk_bF$buf3),
    .Q(alu_op[0])
);

OAI21X1 _1233_ (
    .A(_316_),
    .B(_317_),
    .C(_313_),
    .Y(_325_)
);

FILL FILL_0__981_ (
);

OAI21X1 _984_ (
    .A(_73_),
    .B(_75_),
    .C(_70_),
    .Y(_76_)
);

FILL FILL_1__1395_ (
);

OAI21X1 _1709_ (
    .A(shr),
    .B(_859_),
    .C(_879_),
    .Y(_881_)
);

NAND2X1 _1882_ (
    .A(_848_),
    .B(_849_),
    .Y(_850_)
);

OAI21X1 _1462_ (
    .A(_489_),
    .B(_474_),
    .C(_492_),
    .Y(_551_)
);

NOR2X1 _1042_ (
    .A(_715_),
    .B(_133_),
    .Y(_134_)
);

FILL FILL_0__1502_ (
);

FILL FILL_0__1099_ (
);

OAI21X1 _1518_ (
    .A(_525_),
    .B(_555_),
    .C(_605_),
    .Y(_606_)
);

NAND2X1 _1691_ (
    .A(alu_op[0]),
    .B(_862_),
    .Y(_863_)
);

NOR2X1 _1271_ (
    .A(ACC[0]),
    .B(Flag_i),
    .Y(_363_)
);

FILL FILL_0__1731_ (
);

FILL FILL_0__1311_ (
);

FILL FILL_2__1082_ (
);

OAI21X1 _1747_ (
    .A(AI[2]),
    .B(_914_),
    .C(_868_),
    .Y(_917_)
);

OAI21X1 _1327_ (
    .A(_417_),
    .B(_26_),
    .C(_314_),
    .Y(_418_)
);

FILL FILL_1__1489_ (
);

FILL FILL_1__1069_ (
);

OAI21X1 _1080_ (
    .A(_110_),
    .B(_168_),
    .C(_171_),
    .Y(_172_)
);

FILL FILL_0__1540_ (
);

FILL FILL_0__1120_ (
);

FILL FILL_1__1701_ (
);

NAND2X1 _1556_ (
    .A(_642_),
    .B(_640_),
    .Y(_643_)
);

NAND3X1 _1136_ (
    .A(_222_),
    .B(_223_),
    .C(_224_),
    .Y(_228_)
);

FILL FILL_1__1298_ (
);

FILL FILL_2__1787_ (
);

FILL FILL_1__1510_ (
);

NAND2X1 _1785_ (
    .A(AI[4]),
    .B(_759_),
    .Y(_760_)
);

NAND2X1 _1365_ (
    .A(_442_),
    .B(_454_),
    .Y(_455_)
);

FILL FILL_0__1825_ (
);

FILL FILL_0__1405_ (
);

FILL FILL86250x64950 (
);

AOI21X1 _1594_ (
    .A(_627_),
    .B(AN),
    .C(MulH_i),
    .Y(_679_)
);

NAND2X1 _1174_ (
    .A(BI[0]),
    .B(_717_),
    .Y(_266_)
);

FILL FILL_1__956_ (
);

FILL FILL85950x46950 (
);

FILL FILL_0__1634_ (
);

FILL FILL_0__1214_ (
);

FILL FILL_0__978_ (
);

FILL FILL_0__1863_ (
);

FILL FILL_0__1443_ (
);

FILL FILL_0__1023_ (
);

FILL FILL_2__972_ (
);

FILL FILL_1__1604_ (
);

NAND2X1 _1879_ (
    .A(_845_),
    .B(_846_),
    .Y(_847_)
);

NAND2X1 _1459_ (
    .A(_543_),
    .B(_546_),
    .Y(_548_)
);

AOI21X1 _1039_ (
    .A(_70_),
    .B(_74_),
    .C(_73_),
    .Y(_131_)
);

FILL FILL_1__994_ (
);

FILL FILL_0__1252_ (
);

FILL FILL_1__1833_ (
);

FILL FILL_1__1413_ (
);

NOR2X1 _1688_ (
    .A(shr),
    .B(_859_),
    .Y(_860_)
);

NAND2X1 _1268_ (
    .A(_351_),
    .B(_347_),
    .Y(_360_)
);

FILL FILL_0__1728_ (
);

FILL FILL_0__1308_ (
);

FILL FILL_0__1481_ (
);

FILL FILL_0__1061_ (
);

FILL FILL_1__1642_ (
);

FILL FILL_1__1222_ (
);

OR2X2 _1497_ (
    .A(_584_),
    .B(_581_),
    .Y(_585_)
);

INVX1 _1077_ (
    .A(BI[4]),
    .Y(_169_)
);

FILL FILL_0__1537_ (
);

FILL FILL_0__1117_ (
);

FILL FILL_0__1290_ (
);

FILL FILL_1__1871_ (
);

FILL FILL_1__1451_ (
);

FILL FILL_1__1031_ (
);

FILL FILL_2__1520_ (
);

FILL FILL_0__1766_ (
);

FILL FILL_0__1346_ (
);

FILL FILL_1__1507_ (
);

FILL FILL_1__1260_ (
);

FILL FILL_0__1575_ (
);

FILL FILL_0__1155_ (
);

FILL FILL_1__1736_ (
);

FILL FILL_1__1316_ (
);

FILL FILL_0__1384_ (
);

FILL FILL86550x39750 (
);

AND2X2 _1803_ (
    .A(_864_),
    .B(BI[5]),
    .Y(_776_)
);

FILL FILL_1__1545_ (
);

FILL FILL_1__1125_ (
);

FILL FILL_0__1193_ (
);

INVX1 _1612_ (
    .A(shr),
    .Y(_690_)
);

FILL FILL_0__940_ (
);

INVX1 _943_ (
    .A(_34_),
    .Y(_35_)
);

FILL FILL_1__1774_ (
);

FILL FILL_1__1354_ (
);

FILL FILL_0__1249_ (
);

OAI21X1 _1841_ (
    .A(_811_),
    .B(_810_),
    .C(_807_),
    .Y(_812_)
);

NAND3X1 _1421_ (
    .A(_503_),
    .B(_506_),
    .C(_510_),
    .Y(_511_)
);

NAND3X1 _1001_ (
    .A(MUL_bF$buf1),
    .B(BI[0]),
    .C(AI[6]),
    .Y(_93_)
);

FILL FILL_1__1583_ (
);

FILL FILL_1__1163_ (
);

FILL FILL_0__1478_ (
);

FILL FILL_0__1058_ (
);

FILL FILL_1__1639_ (
);

FILL FILL_1__1219_ (
);

OAI21X1 _1650_ (
    .A(LoadB_i),
    .B(_133_),
    .C(_710_),
    .Y(_24_)
);

NAND3X1 _1230_ (
    .A(_319_),
    .B(_312_),
    .C(_321_),
    .Y(_322_)
);

NOR2X1 _981_ (
    .A(_71_),
    .B(_72_),
    .Y(_73_)
);

FILL FILL_1__1392_ (
);

FILL FILL_2__1461_ (
);

FILL FILL_0__1287_ (
);

OAI21X1 _1706_ (
    .A(_877_),
    .B(_876_),
    .C(_874_),
    .Y(_878_)
);

FILL FILL_1__1868_ (
);

FILL FILL_1__1448_ (
);

FILL FILL_1__1028_ (
);

FILL FILL_0__1096_ (
);

NAND2X1 _1515_ (
    .A(_602_),
    .B(_601_),
    .Y(_603_)
);

FILL FILL_1__1257_ (
);

NOR2X1 _1744_ (
    .A(alu_op[0]),
    .B(_913_),
    .Y(_914_)
);

AOI21X1 _1324_ (
    .A(_326_),
    .B(_324_),
    .C(_414_),
    .Y(_415_)
);

FILL FILL_1__1486_ (
);

FILL FILL_1__1066_ (
);

FILL FILL_2__1135_ (
);

NAND2X1 _1553_ (
    .A(_633_),
    .B(_639_),
    .Y(_640_)
);

AOI21X1 _1133_ (
    .A(_224_),
    .B(_223_),
    .C(_222_),
    .Y(_225_)
);

FILL FILL_1__1295_ (
);

FILL FILL_1_CLKBUF1_insert0 (
);

FILL FILL_1_CLKBUF1_insert1 (
);

FILL FILL_1_CLKBUF1_insert2 (
);

FILL FILL_1_CLKBUF1_insert3 (
);

FILL FILL_1_CLKBUF1_insert4 (
);

INVX1 _1609_ (
    .A(CI),
    .Y(_688_)
);

FILL FILL_0__937_ (
);

AOI21X1 _1782_ (
    .A(_755_),
    .B(_748_),
    .C(_756_),
    .Y(_757_)
);

OAI21X1 _1362_ (
    .A(_449_),
    .B(_452_),
    .C(_374_),
    .Y(_0_[1])
);

FILL FILL_0__1822_ (
);

FILL FILL_0__1402_ (
);

NAND2X1 _1838_ (
    .A(\u_ALU8.AI7 ),
    .B(_808_),
    .Y(_809_)
);

NAND3X1 _1418_ (
    .A(_439_),
    .B(_445_),
    .C(_507_),
    .Y(_508_)
);

NOR2X1 _1591_ (
    .A(_219_),
    .B(_354_),
    .Y(_676_)
);

NAND2X1 _1171_ (
    .A(_242_),
    .B(_240_),
    .Y(_263_)
);

FILL FILL_1__953_ (
);

FILL FILL_0__1631_ (
);

FILL FILL_0__1211_ (
);

NAND2X1 _1647_ (
    .A(ABCmd_i[5]),
    .B(LoadB_i),
    .Y(_709_)
);

NAND2X1 _1227_ (
    .A(_313_),
    .B(_318_),
    .Y(_319_)
);

FILL FILL_0__975_ (
);

INVX1 _978_ (
    .A(_69_),
    .Y(_70_)
);

FILL FILL_1__1389_ (
);

FILL FILL_0__1860_ (
);

FILL FILL_0__1440_ (
);

FILL FILL_0__1020_ (
);

FILL FILL_1__1601_ (
);

AND2X2 _1876_ (
    .A(_842_),
    .B(_816_),
    .Y(_844_)
);

INVX1 _1456_ (
    .A(_542_),
    .Y(_545_)
);

NAND3X1 _1036_ (
    .A(_102_),
    .B(_106_),
    .C(_123_),
    .Y(_128_)
);

FILL FILL_1__1198_ (
);

FILL FILL_1__991_ (
);

FILL FILL_1__1830_ (
);

FILL FILL_1__1410_ (
);

INVX1 _1685_ (
    .A(alu_op_2_bF$buf1),
    .Y(_857_)
);

NAND3X1 _1265_ (
    .A(_144_),
    .B(_258_),
    .C(_256_),
    .Y(_357_)
);

FILL FILL_0__1725_ (
);

FILL FILL_0__1305_ (
);

FILL FILL_2__1076_ (
);

NAND2X1 _1494_ (
    .A(BI[6]),
    .B(_405_),
    .Y(_582_)
);

NAND3X1 _1074_ (
    .A(MUL_bF$buf5),
    .B(BI[5]),
    .C(AI[2]),
    .Y(_166_)
);

FILL FILL_0__1534_ (
);

FILL FILL_0__1114_ (
);

FILL FILL86250x50550 (
);

BUFX2 BUFX2_insert5 (
    .A(MUL),
    .Y(MUL_bF$buf5)
);

BUFX2 BUFX2_insert6 (
    .A(MUL),
    .Y(MUL_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .A(MUL),
    .Y(MUL_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .A(MUL),
    .Y(MUL_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .A(MUL),
    .Y(MUL_bF$buf1)
);

FILL FILL_0__1763_ (
);

FILL FILL_0__1343_ (
);

FILL FILL_1__1504_ (
);

NAND3X1 _1779_ (
    .A(_749_),
    .B(_750_),
    .C(_753_),
    .Y(_754_)
);

OAI21X1 _1359_ (
    .A(_360_),
    .B(_359_),
    .C(_351_),
    .Y(_450_)
);

FILL FILL_0__1819_ (
);

FILL FILL_0__1572_ (
);

FILL FILL_0__1152_ (
);

FILL FILL_1__1733_ (
);

FILL FILL_1__1313_ (
);

NAND2X1 _1588_ (
    .A(_658_),
    .B(_673_),
    .Y(_0_[6])
);

INVX1 _1168_ (
    .A(_247_),
    .Y(_260_)
);

FILL FILL_0__1628_ (
);

FILL FILL_0__1208_ (
);

FILL FILL_0__1381_ (
);

NOR2X1 _1800_ (
    .A(_768_),
    .B(_773_),
    .Y(ACC[4])
);

FILL FILL_1__1542_ (
);

FILL FILL_1__1122_ (
);

AOI21X1 _1397_ (
    .A(_413_),
    .B(_416_),
    .C(_486_),
    .Y(_487_)
);

FILL FILL_2__1611_ (
);

FILL FILL_0__1857_ (
);

FILL FILL_0__1437_ (
);

FILL FILL_0__1017_ (
);

FILL FILL_2__966_ (
);

FILL FILL_0__1190_ (
);

NAND3X1 _940_ (
    .A(MUL_bF$buf0),
    .B(BI[0]),
    .C(AI[4]),
    .Y(_32_)
);

FILL FILL_1__1771_ (
);

FILL FILL_1__1351_ (
);

FILL FILL_1__988_ (
);

FILL FILL_0__1246_ (
);

FILL FILL_1__1827_ (
);

FILL FILL_1__1407_ (
);

FILL FILL_1__1580_ (
);

FILL FILL_1__1160_ (
);

FILL FILL_0__1895_ (
);

FILL FILL_0__1475_ (
);

FILL FILL_0__1055_ (
);

FILL FILL_1__1636_ (
);

FILL FILL_1__1216_ (
);

FILL FILL_0__1284_ (
);

OAI21X1 _1703_ (
    .A(BI[0]),
    .B(alu_op_2_bF$buf1),
    .C(_858_),
    .Y(_875_)
);

FILL FILL_1__1865_ (
);

FILL FILL_1__1445_ (
);

FILL FILL_1__1025_ (
);

FILL FILL_2__1514_ (
);

FILL FILL_0__1093_ (
);

NAND2X1 _1512_ (
    .A(_596_),
    .B(_599_),
    .Y(_600_)
);

FILL FILL_1__1254_ (
);

FILL FILL86550x25350 (
);

FILL FILL_0__1569_ (
);

FILL FILL_0__1149_ (
);

OAI21X1 _1741_ (
    .A(_910_),
    .B(_905_),
    .C(_906_),
    .Y(_911_)
);

NOR2X1 _1321_ (
    .A(_408_),
    .B(_316_),
    .Y(_412_)
);

FILL FILL_1__1483_ (
);

FILL FILL_1__1063_ (
);

FILL FILL_0__1798_ (
);

FILL FILL_0__1378_ (
);

FILL FILL_1__1539_ (
);

FILL FILL_1__1119_ (
);

OR2X2 _1550_ (
    .A(_592_),
    .B(_636_),
    .Y(_637_)
);

AOI21X1 _1130_ (
    .A(_221_),
    .B(_27_),
    .C(_722_),
    .Y(_222_)
);

FILL FILL_1__1292_ (
);

FILL FILL_2__1781_ (
);

FILL FILL_0__1187_ (
);

INVX1 _1606_ (
    .A(alu_op[3]),
    .Y(_686_)
);

FILL FILL_0__934_ (
);

OAI21X1 _937_ (
    .A(_724_),
    .B(_28_),
    .C(_723_),
    .Y(_29_)
);

FILL FILL_1__1768_ (
);

FILL FILL_1__1348_ (
);

FILL FILL86850x68550 (
);

AOI21X1 _1835_ (
    .A(_786_),
    .B(_783_),
    .C(_800_),
    .Y(_806_)
);

OAI21X1 _1415_ (
    .A(_496_),
    .B(_501_),
    .C(_459_),
    .Y(_505_)
);

FILL FILL_1__1577_ (
);

FILL FILL_1__1157_ (
);

FILL FILL_1__950_ (
);

FILL FILL_2__1226_ (
);

NAND2X1 _1644_ (
    .A(ABCmd_i[4]),
    .B(LoadB_i),
    .Y(_707_)
);

NOR2X1 _1224_ (
    .A(_314_),
    .B(_315_),
    .Y(_316_)
);

FILL FILL_0__972_ (
);

NAND2X1 _975_ (
    .A(MUL_bF$buf5),
    .B(AI[0]),
    .Y(_67_)
);

FILL FILL_1__1386_ (
);

FILL FILL_2__1455_ (
);

AOI21X1 _1873_ (
    .A(AN),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

NAND2X1 _1453_ (
    .A(_541_),
    .B(_540_),
    .Y(_542_)
);

AOI21X1 _1033_ (
    .A(_120_),
    .B(_124_),
    .C(_90_),
    .Y(_125_)
);

FILL FILL_1__1195_ (
);

OR2X2 _1509_ (
    .A(_593_),
    .B(_546_),
    .Y(_597_)
);

DFFPOSX1 _1682_ (
    .D(_23_),
    .CLK(clk_bF$buf1),
    .Q(BI[5])
);

INVX1 _1262_ (
    .A(_218_),
    .Y(_354_)
);

FILL FILL_0__1722_ (
);

FILL FILL_0__1302_ (
);

NAND2X1 _1738_ (
    .A(_908_),
    .B(_897_),
    .Y(_909_)
);

OAI22X1 _1318_ (
    .A(_316_),
    .B(_408_),
    .C(_407_),
    .D(_403_),
    .Y(_409_)
);

OAI21X1 _1491_ (
    .A(_529_),
    .B(_578_),
    .C(_532_),
    .Y(_579_)
);

NAND3X1 _1071_ (
    .A(_159_),
    .B(_155_),
    .C(_157_),
    .Y(_163_)
);

FILL FILL_0__1531_ (
);

FILL FILL_0__1111_ (
);

NAND2X1 _1547_ (
    .A(\u_ALU8.AI7 ),
    .B(_289_),
    .Y(_634_)
);

AOI21X1 _1127_ (
    .A(_217_),
    .B(_214_),
    .C(_145_),
    .Y(_219_)
);

FILL FILL_1__1289_ (
);

FILL FILL_0__1760_ (
);

FILL FILL_0__1340_ (
);

FILL FILL_1__1501_ (
);

INVX1 _1776_ (
    .A(_751_),
    .Y(ACC[3])
);

NAND3X1 _1356_ (
    .A(_445_),
    .B(_446_),
    .C(_444_),
    .Y(_447_)
);

FILL FILL_1__1098_ (
);

FILL FILL_0__1816_ (
);

FILL FILL_2__1167_ (
);

FILL FILL_1__1730_ (
);

FILL FILL_1__1310_ (
);

INVX1 _1585_ (
    .A(_661_),
    .Y(_671_)
);

INVX1 _1165_ (
    .A(_89_),
    .Y(_257_)
);

FILL FILL_1__947_ (
);

FILL FILL_0__1625_ (
);

FILL FILL_0__1205_ (
);

FILL FILL_2__1396_ (
);

FILL FILL_0__969_ (
);

AND2X2 _1394_ (
    .A(_477_),
    .B(_478_),
    .Y(_484_)
);

FILL FILL_0__1854_ (
);

FILL FILL_0__1434_ (
);

FILL FILL_0__1014_ (
);

FILL FILL_1__985_ (
);

FILL FILL_0__1243_ (
);

FILL FILL_1__1824_ (
);

FILL FILL_1__1404_ (
);

DFFPOSX1 _1679_ (
    .D(_20_),
    .CLK(clk_bF$buf3),
    .Q(BI[2])
);

NAND3X1 _1259_ (
    .A(_349_),
    .B(_350_),
    .C(_348_),
    .Y(_351_)
);

FILL FILL_0__1719_ (
);

FILL FILL_0__1892_ (
);

FILL FILL_0__1472_ (
);

FILL FILL_0__1052_ (
);

FILL FILL_1__1633_ (
);

FILL FILL_1__1213_ (
);

OAI21X1 _1488_ (
    .A(_528_),
    .B(_548_),
    .C(_554_),
    .Y(_576_)
);

NAND3X1 _1068_ (
    .A(_159_),
    .B(_154_),
    .C(_157_),
    .Y(_160_)
);

FILL FILL_2__1702_ (
);

FILL FILL_0__1528_ (
);

FILL FILL_0__1108_ (
);

FILL FILL_0__1281_ (
);

NAND2X1 _1700_ (
    .A(_868_),
    .B(_871_),
    .Y(_872_)
);

FILL FILL_1__1862_ (
);

FILL FILL_1__1442_ (
);

FILL FILL_1__1022_ (
);

AOI21X1 _1297_ (
    .A(_307_),
    .B(_310_),
    .C(_304_),
    .Y(_388_)
);

FILL FILL_0__1757_ (
);

FILL FILL_0__1337_ (
);

FILL FILL_0__1090_ (
);

FILL FILL_1__1251_ (
);

FILL FILL_0__1566_ (
);

FILL FILL_0__1146_ (
);

FILL FILL_1__1727_ (
);

FILL FILL_1__1307_ (
);

FILL FILL86550x46950 (
);

FILL FILL_1__1480_ (
);

FILL FILL_1__1060_ (
);

FILL FILL_0__1795_ (
);

FILL FILL_0__1375_ (
);

FILL FILL_1__1536_ (
);

FILL FILL_1__1116_ (
);

FILL FILL_2__1605_ (
);

FILL FILL_0__1184_ (
);

INVX1 _1603_ (
    .A(alu_op_2_bF$buf2),
    .Y(_684_)
);

FILL FILL_0__931_ (
);

NAND2X1 _934_ (
    .A(MUL_bF$buf2),
    .B(BI[1]),
    .Y(_26_)
);

FILL FILL_1__1765_ (
);

FILL FILL_1__1345_ (
);

NAND2X1 _1832_ (
    .A(_803_),
    .B(_802_),
    .Y(_804_)
);

OAI21X1 _1412_ (
    .A(_496_),
    .B(_501_),
    .C(_495_),
    .Y(_502_)
);

FILL FILL_1__1574_ (
);

FILL FILL_1__1154_ (
);

FILL FILL_0__1889_ (
);

FILL FILL_0__1469_ (
);

FILL FILL_0__1049_ (
);

OAI21X1 _1641_ (
    .A(LoadB_i),
    .B(_268_),
    .C(_705_),
    .Y(_20_)
);

AOI21X1 _1221_ (
    .A(_159_),
    .B(_155_),
    .C(_152_),
    .Y(_313_)
);

OAI21X1 _972_ (
    .A(_59_),
    .B(_60_),
    .C(_57_),
    .Y(_64_)
);

FILL FILL_1__1383_ (
);

FILL FILL_2__1872_ (
);

FILL FILL_0__1698_ (
);

FILL FILL_0__1278_ (
);

FILL FILL_1__1859_ (
);

FILL FILL_1__1439_ (
);

FILL FILL_1__1019_ (
);

OAI21X1 _1870_ (
    .A(_826_),
    .B(_827_),
    .C(_838_),
    .Y(CO)
);

NAND2X1 _1450_ (
    .A(\u_ALU8.AI7 ),
    .B(_713_),
    .Y(_539_)
);

AOI21X1 _1030_ (
    .A(_101_),
    .B(_98_),
    .C(_91_),
    .Y(_122_)
);

FILL FILL_1__1192_ (
);

FILL FILL_0__1087_ (
);

NOR2X1 _1506_ (
    .A(_546_),
    .B(_593_),
    .Y(_594_)
);

FILL FILL_1__1248_ (
);

OAI21X1 _1735_ (
    .A(_877_),
    .B(_893_),
    .C(_891_),
    .Y(_906_)
);

NAND3X1 _1315_ (
    .A(BI[3]),
    .B(_398_),
    .C(_405_),
    .Y(_406_)
);

FILL FILL_1__1897_ (
);

FILL FILL_1__1477_ (
);

FILL FILL_1__1057_ (
);

FILL FILL_2__1546_ (
);

INVX1 _1544_ (
    .A(_581_),
    .Y(_631_)
);

AOI21X1 _1124_ (
    .A(_204_),
    .B(_208_),
    .C(_147_),
    .Y(_216_)
);

FILL FILL86850x54150 (
);

FILL FILL_1__1286_ (
);

FILL FILL_0__928_ (
);

OAI21X1 _1773_ (
    .A(_736_),
    .B(_737_),
    .C(_748_),
    .Y(_749_)
);

OAI21X1 _1353_ (
    .A(_343_),
    .B(_443_),
    .C(_337_),
    .Y(_444_)
);

FILL FILL_1__1095_ (
);

FILL FILL_0__1813_ (
);

INVX1 _1829_ (
    .A(_800_),
    .Y(_801_)
);

INVX1 _1409_ (
    .A(_413_),
    .Y(_499_)
);

OAI21X1 _1582_ (
    .A(_661_),
    .B(_660_),
    .C(_667_),
    .Y(_668_)
);

OAI21X1 _1162_ (
    .A(_88_),
    .B(_253_),
    .C(_719_),
    .Y(_254_)
);

FILL FILL_1__944_ (
);

FILL FILL_0__1622_ (
);

FILL FILL_0__1202_ (
);

NAND2X1 _1638_ (
    .A(ABCmd_i[1]),
    .B(LoadB_i),
    .Y(_704_)
);

OAI21X1 _1218_ (
    .A(_309_),
    .B(_54_),
    .C(_168_),
    .Y(_310_)
);

FILL FILL_0__966_ (
);

OAI21X1 _969_ (
    .A(_59_),
    .B(_60_),
    .C(_56_),
    .Y(_61_)
);

OAI21X1 _1391_ (
    .A(_480_),
    .B(_44_),
    .C(_478_),
    .Y(_481_)
);

FILL FILL_0__1851_ (
);

FILL FILL_0__1431_ (
);

FILL FILL_0__1011_ (
);

INVX1 _1867_ (
    .A(_832_),
    .Y(_836_)
);

INVX1 _1447_ (
    .A(_535_),
    .Y(_536_)
);

NAND2X1 _1027_ (
    .A(_118_),
    .B(_114_),
    .Y(_119_)
);

FILL FILL_1__1189_ (
);

FILL FILL_1__982_ (
);

FILL FILL_0__1240_ (
);

FILL FILL_1__1821_ (
);

FILL FILL_1__1401_ (
);

DFFPOSX1 _1676_ (
    .D(_17_),
    .CLK(clk_bF$buf1),
    .Q(\u_ALU8.AI7 )
);

OAI21X1 _1256_ (
    .A(_132_),
    .B(_215_),
    .C(_213_),
    .Y(_348_)
);

FILL FILL_0__1716_ (
);

FILL FILL_2__1487_ (
);

FILL FILL_1__1630_ (
);

FILL FILL_1__1210_ (
);

AOI21X1 _1485_ (
    .A(Flag_i),
    .B(_572_),
    .C(_573_),
    .Y(_574_)
);

OR2X2 _1065_ (
    .A(_150_),
    .B(_151_),
    .Y(_157_)
);

FILL FILL_0__1525_ (
);

FILL FILL_0__1105_ (
);

OAI21X1 _1294_ (
    .A(_302_),
    .B(_305_),
    .C(_308_),
    .Y(_385_)
);

FILL FILL_0__1754_ (
);

FILL FILL_0__1334_ (
);

FILL FILL_0__1563_ (
);

FILL FILL_0__1143_ (
);

FILL FILL_1__1724_ (
);

FILL FILL_1__1304_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

FILL FILL_0_BUFX2_insert12 (
);

FILL FILL_0_BUFX2_insert13 (
);

NAND2X1 _1579_ (
    .A(_663_),
    .B(_662_),
    .Y(_665_)
);

FILL FILL_0_BUFX2_insert14 (
);

NAND3X1 _1159_ (
    .A(_234_),
    .B(_249_),
    .C(_250_),
    .Y(_251_)
);

FILL FILL_0__1619_ (
);

FILL FILL_0__1792_ (
);

FILL FILL_0__1372_ (
);

FILL FILL_1__1533_ (
);

FILL FILL_1__1113_ (
);

NAND3X1 _1388_ (
    .A(MUL_bF$buf3),
    .B(\u_ALU8.AI7 ),
    .C(BI[3]),
    .Y(_478_)
);

FILL FILL_0__1848_ (
);

FILL FILL_0__1428_ (
);

FILL FILL_0__1008_ (
);

FILL FILL_0__1181_ (
);

INVX1 _1600_ (
    .A(alu_op[1]),
    .Y(_682_)
);

INVX1 _931_ (
    .A(_722_),
    .Y(_723_)
);

FILL FILL_1__1762_ (
);

FILL FILL_1__1342_ (
);

NOR2X1 _1197_ (
    .A(_715_),
    .B(_288_),
    .Y(_289_)
);

FILL FILL_1__979_ (
);

FILL FILL_0__1237_ (
);

FILL FILL_1__1818_ (
);

FILL FILL_1__1571_ (
);

FILL FILL_1__1151_ (
);

FILL FILL_2__1220_ (
);

FILL FILL_0__1886_ (
);

FILL FILL_0__1466_ (
);

FILL FILL_0__1046_ (
);

FILL FILL_1__1627_ (
);

FILL FILL_1__1207_ (
);

FILL FILL_1__1380_ (
);

FILL FILL_0__1695_ (
);

FILL FILL_0__1275_ (
);

FILL FILL_1__1856_ (
);

FILL FILL_1__1436_ (
);

FILL FILL_1__1016_ (
);

FILL FILL_0__1084_ (
);

FILL FILL86550x32550 (
);

INVX1 _1503_ (
    .A(_590_),
    .Y(_591_)
);

FILL FILL_1__1245_ (
);

NAND3X1 _1732_ (
    .A(_868_),
    .B(_871_),
    .C(_902_),
    .Y(_903_)
);

AOI21X1 _1312_ (
    .A(_400_),
    .B(_402_),
    .C(_397_),
    .Y(_403_)
);

FILL FILL_1__1894_ (
);

FILL FILL_1__1474_ (
);

FILL FILL_1__1054_ (
);

FILL FILL_0__1789_ (
);

FILL FILL_0__1369_ (
);

AND2X2 _1541_ (
    .A(_627_),
    .B(ACC[5]),
    .Y(_628_)
);

NAND3X1 _1121_ (
    .A(_211_),
    .B(_210_),
    .C(_212_),
    .Y(_213_)
);

FILL FILL_1__1283_ (
);

FILL FILL_0__1598_ (
);

FILL FILL_0__1178_ (
);

FILL FILL86850x75750 (
);

FILL FILL_0__925_ (
);

NAND3X1 _928_ (
    .A(MUL_bF$buf2),
    .B(BI[0]),
    .C(AI[3]),
    .Y(_720_)
);

FILL FILL_1__1759_ (
);

FILL FILL_1__1339_ (
);

OAI21X1 _1770_ (
    .A(_877_),
    .B(_745_),
    .C(_743_),
    .Y(_746_)
);

AOI21X1 _1350_ (
    .A(_440_),
    .B(_439_),
    .C(_378_),
    .Y(_441_)
);

FILL FILL_1__1092_ (
);

FILL FILL_0__1810_ (
);

FILL FILL_2__1161_ (
);

AOI21X1 _1826_ (
    .A(alu_op_2_bF$buf2),
    .B(BI[6]),
    .C(_797_),
    .Y(_798_)
);

AOI22X1 _1406_ (
    .A(_470_),
    .B(_473_),
    .C(_492_),
    .D(_488_),
    .Y(_496_)
);

FILL FILL_1__1568_ (
);

FILL FILL_1__1148_ (
);

FILL FILL_1__941_ (
);

OAI21X1 _1635_ (
    .A(LoadA_i),
    .B(_417_),
    .C(_702_),
    .Y(_17_)
);

INVX1 _1215_ (
    .A(_302_),
    .Y(_307_)
);

FILL FILL_0__963_ (
);

NAND3X1 _966_ (
    .A(_55_),
    .B(_57_),
    .C(_52_),
    .Y(_58_)
);

FILL FILL_1__1797_ (
);

FILL FILL_1__1377_ (
);

FILL FILL_2__1866_ (
);

NAND3X1 _1864_ (
    .A(_829_),
    .B(_832_),
    .C(_831_),
    .Y(_833_)
);

AOI21X1 _1444_ (
    .A(_476_),
    .B(_481_),
    .C(_483_),
    .Y(_533_)
);

INVX1 _1024_ (
    .A(_110_),
    .Y(_116_)
);

FILL FILL_1__1186_ (
);

DFFPOSX1 _1673_ (
    .D(_14_),
    .CLK(clk_bF$buf2),
    .Q(AI[4])
);

OAI21X1 _1253_ (
    .A(_339_),
    .B(_340_),
    .C(_287_),
    .Y(_345_)
);

FILL FILL86250x150 (
);

FILL FILL_0__1713_ (
);

MUX2X1 _1729_ (
    .A(alu_op[1]),
    .B(_869_),
    .S(alu_op[0]),
    .Y(_900_)
);

OR2X2 _1309_ (
    .A(_398_),
    .B(_399_),
    .Y(_400_)
);

AOI21X1 _1482_ (
    .A(_270_),
    .B(_569_),
    .C(_570_),
    .Y(_571_)
);

NAND3X1 _1062_ (
    .A(MUL_bF$buf1),
    .B(BI[2]),
    .C(AI[5]),
    .Y(_154_)
);

FILL FILL_0__1522_ (
);

FILL FILL_0__1102_ (
);

OAI21X1 _1538_ (
    .A(_617_),
    .B(_624_),
    .C(MulL_i),
    .Y(_625_)
);

OAI21X1 _1118_ (
    .A(_137_),
    .B(_125_),
    .C(_141_),
    .Y(_210_)
);

NAND2X1 _1291_ (
    .A(AI[2]),
    .B(_289_),
    .Y(_382_)
);

FILL FILL_0__1751_ (
);

FILL FILL_0__1331_ (
);

OAI21X1 _1767_ (
    .A(_742_),
    .B(_741_),
    .C(_738_),
    .Y(_743_)
);

AOI21X1 _1347_ (
    .A(_430_),
    .B(_437_),
    .C(_379_),
    .Y(_438_)
);

FILL FILL_1__1089_ (
);

FILL FILL_0__1807_ (
);

FILL FILL_0__1560_ (
);

FILL FILL_0__1140_ (
);

FILL FILL_1__1721_ (
);

FILL FILL_1__1301_ (
);

OAI21X1 _1576_ (
    .A(_592_),
    .B(_636_),
    .C(_642_),
    .Y(_662_)
);

AOI21X1 _1156_ (
    .A(_235_),
    .B(_245_),
    .C(_244_),
    .Y(_248_)
);

FILL FILL_1__938_ (
);

FILL FILL_0__1616_ (
);

FILL FILL_1__1530_ (
);

FILL FILL85650x39750 (
);

FILL FILL_1__1110_ (
);

NAND3X1 _1385_ (
    .A(MUL_bF$buf3),
    .B(AI[5]),
    .C(BI[5]),
    .Y(_475_)
);

FILL FILL_0__1845_ (
);

FILL FILL_0__1425_ (
);

FILL FILL_0__1005_ (
);

OAI21X1 _1194_ (
    .A(_191_),
    .B(_285_),
    .C(_200_),
    .Y(_286_)
);

FILL FILL_1__976_ (
);

FILL FILL_0__1234_ (
);

FILL FILL_1__1815_ (
);

FILL FILL_0__998_ (
);

FILL FILL86250x10950 (
);

FILL FILL_0__1883_ (
);

FILL FILL_0__1463_ (
);

FILL FILL_0__1043_ (
);

FILL FILL_2__992_ (
);

FILL FILL_1__1624_ (
);

FILL FILL_1__1204_ (
);

NAND2X1 _1479_ (
    .A(_561_),
    .B(_567_),
    .Y(_568_)
);

NAND3X1 _1059_ (
    .A(MUL_bF$buf5),
    .B(BI[0]),
    .C(\u_ALU8.AI7 ),
    .Y(_151_)
);

FILL FILL_0__1519_ (
);

FILL FILL_0__1692_ (
);

FILL FILL_0__1272_ (
);

FILL FILL_1__1853_ (
);

FILL FILL_1__1433_ (
);

FILL FILL_1__1013_ (
);

INVX1 _1288_ (
    .A(_378_),
    .Y(_379_)
);

FILL FILL_0__1748_ (
);

FILL FILL_0__1328_ (
);

FILL FILL_0__1081_ (
);

OAI21X1 _1500_ (
    .A(_417_),
    .B(_182_),
    .C(_587_),
    .Y(_588_)
);

FILL FILL_1__1242_ (
);

NAND3X1 _1097_ (
    .A(_161_),
    .B(_165_),
    .C(_184_),
    .Y(_189_)
);

FILL FILL_2__1311_ (
);

FILL FILL_0__1557_ (
);

FILL FILL_0__1137_ (
);

FILL FILL_1__1718_ (
);

FILL FILL_1__1891_ (
);

FILL FILL_1__1471_ (
);

FILL FILL_1__1051_ (
);

FILL FILL_2__1540_ (
);

FILL FILL_0__1786_ (
);

FILL FILL_0__1366_ (
);

FILL FILL_1__1527_ (
);

FILL FILL_1__1107_ (
);

FILL FILL_1__1280_ (
);

FILL FILL_0__1595_ (
);

FILL FILL_0__1175_ (
);

FILL FILL_0__922_ (
);

NOR2X1 _925_ (
    .A(_715_),
    .B(_716_),
    .Y(_717_)
);

FILL FILL_1__1756_ (
);

FILL FILL_1__1336_ (
);

OAI21X1 _1823_ (
    .A(AI[6]),
    .B(_792_),
    .C(_868_),
    .Y(_795_)
);

NAND3X1 _1403_ (
    .A(_492_),
    .B(_488_),
    .C(_491_),
    .Y(_493_)
);

FILL FILL_1__1565_ (
);

FILL FILL_1__1145_ (
);

NAND2X1 _1632_ (
    .A(ABCmd_i[6]),
    .B(LoadA_i),
    .Y(_701_)
);

NOR2X1 _1212_ (
    .A(_168_),
    .B(_303_),
    .Y(_304_)
);

FILL FILL_0__960_ (
);

OAI21X1 _963_ (
    .A(_53_),
    .B(_54_),
    .C(_50_),
    .Y(_55_)
);

FILL FILL_1__1794_ (
);

FILL FILL_1__1374_ (
);

FILL FILL_0__1689_ (
);

FILL FILL_0__1269_ (
);

NOR2X1 _1861_ (
    .A(_816_),
    .B(_800_),
    .Y(_830_)
);

INVX1 _1441_ (
    .A(_529_),
    .Y(_530_)
);

INVX1 _1021_ (
    .A(_112_),
    .Y(_113_)
);

FILL FILL_1__1183_ (
);

FILL FILL_2__1252_ (
);

FILL FILL_0__1498_ (
);

FILL FILL_0__1078_ (
);

FILL FILL_1__1239_ (
);

DFFPOSX1 _1670_ (
    .D(_11_),
    .CLK(clk_bF$buf0),
    .Q(AI[1])
);

AOI21X1 _1250_ (
    .A(_337_),
    .B(_341_),
    .C(_286_),
    .Y(_342_)
);

FILL FILL_0__1710_ (
);

FILL FILL_2__1728_ (
);

FILL FILL_2__1481_ (
);

NAND2X1 _1726_ (
    .A(_896_),
    .B(_884_),
    .Y(_897_)
);

INVX1 _1306_ (
    .A(_396_),
    .Y(_397_)
);

FILL FILL_1__1888_ (
);

FILL FILL_1__1468_ (
);

FILL FILL_1__1048_ (
);

FILL FILL86850x28950 (
);

NAND2X1 _1535_ (
    .A(_712_),
    .B(_622_),
    .Y(_623_)
);

AND2X2 _1115_ (
    .A(_199_),
    .B(_202_),
    .Y(_207_)
);

FILL FILL_1__1697_ (
);

FILL FILL_1__1277_ (
);

NAND2X1 _1764_ (
    .A(AI[3]),
    .B(_739_),
    .Y(_740_)
);

OAI21X1 _1344_ (
    .A(_424_),
    .B(_330_),
    .C(_414_),
    .Y(_435_)
);

FILL FILL_1__1086_ (
);

FILL FILL_0__1804_ (
);

NAND3X1 _1573_ (
    .A(_601_),
    .B(_602_),
    .C(_650_),
    .Y(_659_)
);

OAI21X1 _1153_ (
    .A(_722_),
    .B(_28_),
    .C(_724_),
    .Y(_245_)
);

FILL FILL_1__935_ (
);

FILL FILL_0__1613_ (
);

OAI21X1 _1629_ (
    .A(LoadA_i),
    .B(_463_),
    .C(_699_),
    .Y(_14_)
);

AOI21X1 _1209_ (
    .A(_161_),
    .B(_177_),
    .C(_180_),
    .Y(_301_)
);

FILL FILL_0__957_ (
);

AND2X2 _1382_ (
    .A(_468_),
    .B(_465_),
    .Y(_472_)
);

FILL FILL_0__1842_ (
);

FILL FILL_0__1422_ (
);

FILL FILL_0__1002_ (
);

FILL FILL_2__1193_ (
);

NAND2X1 _1858_ (
    .A(BCD),
    .B(_824_),
    .Y(_827_)
);

INVX1 _1438_ (
    .A(_526_),
    .Y(_527_)
);

NAND3X1 _1018_ (
    .A(MUL_bF$buf1),
    .B(BI[3]),
    .C(AI[3]),
    .Y(_110_)
);

OAI21X1 _1191_ (
    .A(_219_),
    .B(_282_),
    .C(_218_),
    .Y(_283_)
);

FILL FILL_1__973_ (
);

FILL FILL_0__1651_ (
);

FILL FILL_0__1231_ (
);

FILL FILL_1__1812_ (
);

DFFSR _1667_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[6]),
    .CLK(clk_bF$buf4),
    .Q(_919_[6])
);

AOI21X1 _1247_ (
    .A(_334_),
    .B(_335_),
    .C(_333_),
    .Y(_339_)
);

FILL FILL_0__995_ (
);

OAI21X1 _998_ (
    .A(_85_),
    .B(_82_),
    .C(_62_),
    .Y(_90_)
);

FILL FILL_0__1707_ (
);

FILL FILL_0__1880_ (
);

FILL FILL_0__1460_ (
);

FILL FILL_0__1040_ (
);

FILL FILL_1__1621_ (
);

FILL FILL_1__1201_ (
);

BUFX2 _1896_ (
    .A(_919_[6]),
    .Y(ACC_o[6])
);

AOI21X1 _1476_ (
    .A(_564_),
    .B(_455_),
    .C(_512_),
    .Y(_565_)
);

OAI21X1 _1056_ (
    .A(_121_),
    .B(_123_),
    .C(_106_),
    .Y(_148_)
);

FILL FILL_0__1516_ (
);

FILL FILL_1__1850_ (
);

FILL FILL_1__1430_ (
);

FILL FILL_1__1010_ (
);

NOR2X1 _1285_ (
    .A(_338_),
    .B(_375_),
    .Y(_376_)
);

FILL FILL_0__1745_ (
);

FILL FILL_0__1325_ (
);

FILL FILL_2__1096_ (
);

AOI21X1 _1094_ (
    .A(_178_),
    .B(_185_),
    .C(_148_),
    .Y(_186_)
);

FILL FILL_0__1554_ (
);

FILL FILL_0__1134_ (
);

FILL FILL_1__1715_ (
);

FILL FILL_0__1783_ (
);

FILL FILL_0__1363_ (
);

FILL FILL_1__1524_ (
);

FILL FILL_1__1104_ (
);

NOR2X1 _1799_ (
    .A(_772_),
    .B(HC),
    .Y(_773_)
);

OAI21X1 _1379_ (
    .A(_463_),
    .B(_135_),
    .C(_468_),
    .Y(_469_)
);

FILL FILL_0__1839_ (
);

FILL FILL_0__1419_ (
);

FILL FILL_0__1592_ (
);

FILL FILL_0__1172_ (
);

NAND2X1 _922_ (
    .A(AI[0]),
    .B(_713_),
    .Y(_714_)
);

FILL FILL_1__1753_ (
);

FILL FILL_1__1333_ (
);

NAND3X1 _1188_ (
    .A(_276_),
    .B(_255_),
    .C(_279_),
    .Y(_280_)
);

FILL FILL_2__1402_ (
);

FILL FILL_0__1648_ (
);

FILL FILL_0__1228_ (
);

FILL FILL_1__1809_ (
);

AND2X2 _1820_ (
    .A(_864_),
    .B(BI[6]),
    .Y(_792_)
);

OAI21X1 _1400_ (
    .A(_487_),
    .B(_489_),
    .C(_474_),
    .Y(_490_)
);

FILL FILL_1__1562_ (
);

FILL FILL_1__1142_ (
);

FILL FILL_2__1631_ (
);

FILL FILL_0__1877_ (
);

FILL FILL_0__1457_ (
);

FILL FILL_0__1037_ (
);

FILL FILL_2__986_ (
);

FILL FILL_1__1618_ (
);

OR2X2 _960_ (
    .A(_50_),
    .B(_51_),
    .Y(_52_)
);

FILL FILL_1__1791_ (
);

FILL FILL_1__1371_ (
);

FILL FILL_0__1686_ (
);

FILL FILL_0__1266_ (
);

FILL FILL_1__1847_ (
);

FILL FILL_1__1427_ (
);

FILL FILL_1__1007_ (
);

FILL FILL_1__1180_ (
);

FILL FILL_0__1495_ (
);

FILL FILL_0__1075_ (
);

FILL FILL_1__1236_ (
);

FILL FILL_2__1305_ (
);

INVX1 _1723_ (
    .A(_893_),
    .Y(_894_)
);

OAI21X1 _1303_ (
    .A(_392_),
    .B(_393_),
    .C(_382_),
    .Y(_394_)
);

FILL FILL86250x18150 (
);

FILL FILL_1__1885_ (
);

FILL FILL_1__1465_ (
);

FILL FILL_1__1045_ (
);

NOR2X1 _1532_ (
    .A(Flag_i),
    .B(ACC[4]),
    .Y(_620_)
);

OAI21X1 _1112_ (
    .A(_190_),
    .B(_186_),
    .C(_203_),
    .Y(_204_)
);

FILL FILL86850x82950 (
);

FILL FILL_1__1694_ (
);

FILL FILL_1__1274_ (
);

FILL FILL_0__1589_ (
);

FILL FILL_0__1169_ (
);

AND2X2 _1761_ (
    .A(_911_),
    .B(_730_),
    .Y(_737_)
);

OAI21X1 _1341_ (
    .A(_300_),
    .B(_431_),
    .C(_334_),
    .Y(_432_)
);

FILL FILL_1__1083_ (
);

FILL FILL_0__1801_ (
);

FILL FILL_2__1572_ (
);

FILL FILL_0__1398_ (
);

INVX1 _1817_ (
    .A(_789_),
    .Y(ACC[5])
);

FILL FILL_1__1559_ (
);

FILL FILL_1__1139_ (
);

NAND2X1 _1570_ (
    .A(ACC[6]),
    .B(_627_),
    .Y(_656_)
);

OAI21X1 _1150_ (
    .A(_716_),
    .B(_26_),
    .C(_236_),
    .Y(_242_)
);

FILL FILL_1__932_ (
);

FILL FILL_0__1610_ (
);

NAND2X1 _1626_ (
    .A(ABCmd_i[3]),
    .B(LoadA_i),
    .Y(_698_)
);

AND2X2 _1206_ (
    .A(_293_),
    .B(_292_),
    .Y(_298_)
);

FILL FILL_0__954_ (
);

OAI21X1 _957_ (
    .A(_30_),
    .B(_40_),
    .C(_35_),
    .Y(_49_)
);

FILL FILL_1__1788_ (
);

FILL FILL_1__1368_ (
);

FILL FILL_2__1017_ (
);

NOR2X1 _1855_ (
    .A(_824_),
    .B(AN),
    .Y(_825_)
);

NOR3X1 _1435_ (
    .A(_496_),
    .B(_501_),
    .C(_459_),
    .Y(_524_)
);

NAND3X1 _1015_ (
    .A(MUL_bF$buf1),
    .B(BI[5]),
    .C(AI[1]),
    .Y(_107_)
);

FILL FILL_1__1597_ (
);

FILL FILL_1__1177_ (
);

FILL FILL_1__970_ (
);

FILL FILL_2__1246_ (
);

DFFSR _1664_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[3]),
    .CLK(clk_bF$buf4),
    .Q(_919_[3])
);

NAND3X1 _1244_ (
    .A(_333_),
    .B(_335_),
    .C(_334_),
    .Y(_336_)
);

FILL FILL_0__992_ (
);

NAND3X1 _995_ (
    .A(_80_),
    .B(_86_),
    .C(_48_),
    .Y(_87_)
);

FILL FILL_0__1704_ (
);

FILL FILL86850x14550 (
);

BUFX2 _1893_ (
    .A(_919_[3]),
    .Y(ACC_o[3])
);

INVX1 _1473_ (
    .A(_511_),
    .Y(_562_)
);

INVX1 _1053_ (
    .A(_144_),
    .Y(_145_)
);

FILL FILL_0__1513_ (
);

INVX1 _1529_ (
    .A(_276_),
    .Y(_617_)
);

OAI21X1 _1109_ (
    .A(_716_),
    .B(_135_),
    .C(_193_),
    .Y(_201_)
);

AOI21X1 _1282_ (
    .A(_372_),
    .B(_365_),
    .C(MulH_i),
    .Y(_373_)
);

FILL FILL_0__1742_ (
);

FILL FILL_0__1322_ (
);

NAND2X1 _1758_ (
    .A(_731_),
    .B(_734_),
    .Y(_735_)
);

NAND3X1 _1338_ (
    .A(_428_),
    .B(_423_),
    .C(_426_),
    .Y(_429_)
);

OAI21X1 _1091_ (
    .A(_725_),
    .B(_182_),
    .C(_172_),
    .Y(_183_)
);

FILL FILL_0__1551_ (
);

FILL FILL_0__1131_ (
);

FILL FILL_1__1712_ (
);

NAND2X1 _1567_ (
    .A(_255_),
    .B(_356_),
    .Y(_653_)
);

INVX1 _1147_ (
    .A(_238_),
    .Y(_239_)
);

FILL FILL_1__929_ (
);

FILL FILL_0__1607_ (
);

FILL FILL85650x46950 (
);

FILL FILL_0__1780_ (
);

FILL FILL_0__1360_ (
);

FILL FILL_1__1521_ (
);

FILL FILL_1__1101_ (
);

NAND2X1 _1796_ (
    .A(BCD),
    .B(_770_),
    .Y(_771_)
);

INVX1 _1376_ (
    .A(_465_),
    .Y(_466_)
);

FILL FILL_0__1836_ (
);

FILL FILL_0__1416_ (
);

FILL FILL_2__1187_ (
);

FILL FILL_1__1750_ (
);

FILL FILL_1__1330_ (
);

OAI21X1 _1185_ (
    .A(_88_),
    .B(_253_),
    .C(_220_),
    .Y(_277_)
);

FILL FILL_1__967_ (
);

FILL FILL_0__1645_ (
);

FILL FILL_0__1225_ (
);

FILL FILL_1__1806_ (
);

FILL FILL_0__989_ (
);

FILL FILL_0__1874_ (
);

FILL FILL_0__1454_ (
);

FILL FILL_0__1034_ (
);

FILL FILL_1__1615_ (
);

FILL FILL_0__1263_ (
);

FILL FILL_1__1844_ (
);

FILL FILL_1__1424_ (
);

FILL FILL_1__1004_ (
);

OAI21X1 _1699_ (
    .A(alu_op[0]),
    .B(_869_),
    .C(_870_),
    .Y(_871_)
);

AND2X2 _1279_ (
    .A(_266_),
    .B(_265_),
    .Y(_370_)
);

FILL FILL_0__1739_ (
);

FILL FILL_0__1319_ (
);

FILL FILL_0__1492_ (
);

FILL FILL_0__1072_ (
);

FILL FILL_1__1233_ (
);

AOI21X1 _1088_ (
    .A(_160_),
    .B(_156_),
    .C(_149_),
    .Y(_180_)
);

FILL FILL_2__1722_ (
);

FILL FILL_0__1548_ (
);

FILL FILL_0__1128_ (
);

FILL FILL_1__1709_ (
);

OAI21X1 _1720_ (
    .A(_887_),
    .B(_890_),
    .C(_885_),
    .Y(_891_)
);

NAND2X1 _1300_ (
    .A(BI[6]),
    .B(_384_),
    .Y(_391_)
);

FILL FILL_1__1882_ (
);

FILL FILL_1__1462_ (
);

FILL FILL_1__1042_ (
);

FILL FILL_0__1777_ (
);

FILL FILL_0__1357_ (
);

FILL FILL86250x39750 (
);

FILL FILL_1__1518_ (
);

FILL FILL_1__1691_ (
);

FILL FILL_1__1271_ (
);

FILL FILL86550x150 (
);

FILL FILL_0__1586_ (
);

FILL FILL_0__1166_ (
);

FILL FILL_1__1747_ (
);

FILL FILL_1__1327_ (
);

FILL FILL_1__1080_ (
);

FILL FILL_0__1395_ (
);

AOI21X1 _1814_ (
    .A(HC),
    .B(_772_),
    .C(_774_),
    .Y(_787_)
);

FILL FILL_1__1556_ (
);

FILL FILL_1__1136_ (
);

FILL FILL_2__1625_ (
);

OAI21X1 _1623_ (
    .A(LoadA_i),
    .B(_716_),
    .C(_696_),
    .Y(_11_)
);

OAI21X1 _1203_ (
    .A(_725_),
    .B(_135_),
    .C(_293_),
    .Y(_295_)
);

FILL FILL_0__951_ (
);

NAND2X1 _954_ (
    .A(_45_),
    .B(_719_),
    .Y(_46_)
);

FILL FILL_1__1785_ (
);

FILL FILL_1__1365_ (
);

NOR2X1 _1852_ (
    .A(_821_),
    .B(ACC[4]),
    .Y(_822_)
);

OAI21X1 _1432_ (
    .A(_520_),
    .B(_521_),
    .C(_519_),
    .Y(_522_)
);

NAND3X1 _1012_ (
    .A(_100_),
    .B(_97_),
    .C(_99_),
    .Y(_104_)
);

FILL FILL_1__1594_ (
);

FILL FILL_1__1174_ (
);

FILL FILL_0__1489_ (
);

FILL FILL_0__1069_ (
);

DFFSR _1661_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[0]),
    .CLK(clk_bF$buf4),
    .Q(_919_[0])
);

AND2X2 _1241_ (
    .A(_296_),
    .B(_299_),
    .Y(_333_)
);

OAI21X1 _992_ (
    .A(_73_),
    .B(_75_),
    .C(_69_),
    .Y(_84_)
);

FILL FILL_0__1701_ (
);

FILL FILL_2__1892_ (
);

FILL FILL_0__1298_ (
);

INVX1 _1717_ (
    .A(BI[1]),
    .Y(_888_)
);

FILL FILL_1__1879_ (
);

FILL FILL_1__1459_ (
);

FILL FILL_1__1039_ (
);

BUFX2 _1890_ (
    .A(_919_[0]),
    .Y(ACC_o[0])
);

NAND3X1 _1470_ (
    .A(_550_),
    .B(_554_),
    .C(_558_),
    .Y(_559_)
);

NAND3X1 _1050_ (
    .A(_137_),
    .B(_141_),
    .C(_140_),
    .Y(_142_)
);

FILL FILL_0__1510_ (
);

NAND3X1 _1526_ (
    .A(_283_),
    .B(_612_),
    .C(_563_),
    .Y(_614_)
);

NAND2X1 _1106_ (
    .A(_193_),
    .B(_197_),
    .Y(_198_)
);

FILL FILL_1__1688_ (
);

FILL FILL_1__1268_ (
);

FILL FILL_2__1337_ (
);

OAI21X1 _1755_ (
    .A(_877_),
    .B(_727_),
    .C(_918_),
    .Y(_732_)
);

OAI21X1 _1335_ (
    .A(_424_),
    .B(_330_),
    .C(_425_),
    .Y(_426_)
);

FILL FILL_1__1497_ (
);

FILL FILL_1__1077_ (
);

FILL FILL_2__1566_ (
);

OAI21X1 _1564_ (
    .A(_648_),
    .B(_649_),
    .C(_650_),
    .Y(_651_)
);

NAND3X1 _1144_ (
    .A(MUL_bF$buf0),
    .B(BI[0]),
    .C(AI[2]),
    .Y(_236_)
);

FILL FILL_1__926_ (
);

FILL FILL_0__1604_ (
);

FILL FILL_0__948_ (
);

FILL FILL_2_BUFX2_insert14 (
);

AOI21X1 _1793_ (
    .A(_754_),
    .B(_757_),
    .C(_767_),
    .Y(_768_)
);

INVX1 _1373_ (
    .A(AI[4]),
    .Y(_463_)
);

FILL FILL_0__1833_ (
);

FILL FILL_0__1413_ (
);

AND2X2 _1849_ (
    .A(_818_),
    .B(_819_),
    .Y(AN)
);

OAI21X1 _1429_ (
    .A(_267_),
    .B(_517_),
    .C(_518_),
    .Y(_519_)
);

NAND3X1 _1009_ (
    .A(_100_),
    .B(_96_),
    .C(_99_),
    .Y(_101_)
);

NAND3X1 _1182_ (
    .A(_271_),
    .B(_262_),
    .C(_273_),
    .Y(_274_)
);

FILL FILL_1__964_ (
);

FILL FILL_0__1642_ (
);

FILL FILL_0__1222_ (
);

FILL FILL_1__1803_ (
);

DFFPOSX1 _1658_ (
    .D(_7_),
    .CLK(clk_bF$buf2),
    .Q(shr)
);

AOI21X1 _1238_ (
    .A(_321_),
    .B(_319_),
    .C(_312_),
    .Y(_330_)
);

FILL FILL_0__986_ (
);

AOI21X1 _989_ (
    .A(_64_),
    .B(_65_),
    .C(_63_),
    .Y(_81_)
);

FILL FILL_0__1871_ (
);

FILL FILL_0__1451_ (
);

FILL FILL_0__1031_ (
);

FILL FILL_1__1612_ (
);

NAND2X1 _1887_ (
    .A(_853_),
    .B(_852_),
    .Y(_855_)
);

NAND2X1 _1467_ (
    .A(_525_),
    .B(_555_),
    .Y(_556_)
);

OAI21X1 _1047_ (
    .A(_129_),
    .B(_125_),
    .C(_138_),
    .Y(_139_)
);

FILL FILL_0__1507_ (
);

FILL FILL_0__1260_ (
);

FILL FILL_2__1278_ (
);

FILL FILL_1__1841_ (
);

FILL FILL_1__1421_ (
);

FILL FILL_1__1001_ (
);

INVX2 _1696_ (
    .A(shr),
    .Y(_868_)
);

OAI21X1 _1276_ (
    .A(_363_),
    .B(_366_),
    .C(_367_),
    .Y(_368_)
);

FILL FILL_0__1736_ (
);

FILL FILL_0__1316_ (
);

FILL FILL_1__1650_ (
);

FILL FILL_1__1230_ (
);

NAND2X1 _1085_ (
    .A(_176_),
    .B(_173_),
    .Y(_177_)
);

FILL FILL_0__1545_ (
);

FILL FILL_0__1125_ (
);

FILL FILL_1__1706_ (
);

FILL FILL_0__1774_ (
);

FILL FILL_0__1354_ (
);

FILL FILL_1__1515_ (
);

FILL FILL_0__1583_ (
);

FILL FILL_0__1163_ (
);

FILL FILL_1__1744_ (
);

FILL FILL_1__1324_ (
);

OAI21X1 _1599_ (
    .A(LoadCmd_i),
    .B(_680_),
    .C(_681_),
    .Y(_2_)
);

INVX1 _1179_ (
    .A(_270_),
    .Y(_271_)
);

FILL FILL_2__1813_ (
);

FILL FILL_0__1639_ (
);

FILL FILL_0__1219_ (
);

FILL FILL_0__1392_ (
);

OAI21X1 _1811_ (
    .A(_780_),
    .B(_782_),
    .C(_783_),
    .Y(_784_)
);

FILL FILL_1__1553_ (
);

FILL FILL_1__1133_ (
);

FILL FILL_0__1868_ (
);

FILL FILL_0__1448_ (
);

FILL FILL_0__1028_ (
);

FILL FILL_1__1609_ (
);

NAND2X1 _1620_ (
    .A(ABCmd_i[0]),
    .B(LoadA_i),
    .Y(_695_)
);

NAND2X1 _1200_ (
    .A(AI[2]),
    .B(_134_),
    .Y(_292_)
);

INVX1 _951_ (
    .A(AI[0]),
    .Y(_43_)
);

FILL FILL_1__1782_ (
);

FILL FILL_1__1362_ (
);

FILL FILL_1__999_ (
);

FILL FILL_2__1011_ (
);

FILL FILL_0__1257_ (
);

FILL FILL_1__1838_ (
);

FILL FILL_1__1418_ (
);

FILL FILL_1__1591_ (
);

FILL FILL_1__1171_ (
);

FILL FILL_0__1486_ (
);

FILL FILL_0__1066_ (
);

FILL FILL_1__1647_ (
);

FILL FILL_1__1227_ (
);

FILL FILL86250x25350 (
);

FILL FILL_0__1295_ (
);

NAND2X1 _1714_ (
    .A(shr),
    .B(AI[2]),
    .Y(_885_)
);

FILL FILL_1__1876_ (
);

FILL FILL_1__1456_ (
);

FILL FILL_1__1036_ (
);

OAI21X1 _1523_ (
    .A(_351_),
    .B(_448_),
    .C(_447_),
    .Y(_611_)
);

OAI21X1 _1103_ (
    .A(_716_),
    .B(_135_),
    .C(_194_),
    .Y(_195_)
);

FILL FILL_1__1685_ (
);

FILL FILL_1__1265_ (
);

OAI21X1 _1752_ (
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_728_),
    .Y(_729_)
);

AND2X2 _1332_ (
    .A(_394_),
    .B(_390_),
    .Y(_423_)
);

FILL FILL_1__1494_ (
);

FILL FILL_1__1074_ (
);

FILL FILL86550x68550 (
);

FILL FILL_0__1389_ (
);

OAI21X1 _1808_ (
    .A(alu_op_2_bF$buf3),
    .B(BI[5]),
    .C(_858_),
    .Y(_781_)
);

INVX1 _1561_ (
    .A(_602_),
    .Y(_648_)
);

NAND3X1 _1141_ (
    .A(_220_),
    .B(_87_),
    .C(_232_),
    .Y(_233_)
);

FILL FILL_1__923_ (
);

FILL FILL_0__1601_ (
);

FILL FILL_0__1198_ (
);

OAI21X1 _1617_ (
    .A(LoadCmd_i),
    .B(_692_),
    .C(_693_),
    .Y(_8_)
);

FILL FILL_0__945_ (
);

INVX1 _948_ (
    .A(_38_),
    .Y(_40_)
);

FILL FILL_1__1779_ (
);

FILL FILL_1__1359_ (
);

AOI21X1 _1790_ (
    .A(alu_op_2_bF$buf2),
    .B(BI[4]),
    .C(_764_),
    .Y(_765_)
);

NAND2X1 _1370_ (
    .A(BI[7]),
    .B(_384_),
    .Y(_460_)
);

FILL FILL_0__1830_ (
);

FILL FILL_0__1410_ (
);

INVX1 _1846_ (
    .A(_816_),
    .Y(_817_)
);

NAND2X1 _1426_ (
    .A(_514_),
    .B(_515_),
    .Y(_516_)
);

OAI21X1 _1006_ (
    .A(_94_),
    .B(_95_),
    .C(_97_),
    .Y(_98_)
);

FILL FILL_1__1588_ (
);

FILL FILL_1__1168_ (
);

FILL FILL_1__961_ (
);

FILL FILL86850x21750 (
);

FILL FILL_1__1800_ (
);

DFFPOSX1 _1655_ (
    .D(_4_),
    .CLK(clk_bF$buf3),
    .Q(alu_op[2])
);

NAND3X1 _1235_ (
    .A(_322_),
    .B(_326_),
    .C(_301_),
    .Y(_327_)
);

FILL FILL_0__983_ (
);

NAND3X1 _986_ (
    .A(_69_),
    .B(_74_),
    .C(_77_),
    .Y(_78_)
);

FILL FILL_1__1397_ (
);

OAI21X1 _1884_ (
    .A(_843_),
    .B(_844_),
    .C(_851_),
    .Y(_852_)
);

NAND2X1 _1464_ (
    .A(_548_),
    .B(_528_),
    .Y(_553_)
);

OAI21X1 _1044_ (
    .A(_43_),
    .B(_135_),
    .C(_131_),
    .Y(_136_)
);

FILL FILL_0__1504_ (
);

NAND2X1 _1693_ (
    .A(BI[0]),
    .B(_864_),
    .Y(_865_)
);

INVX2 _1273_ (
    .A(MulL_i),
    .Y(_365_)
);

FILL FILL_0__1733_ (
);

FILL FILL_0__1313_ (
);

OAI21X1 _1749_ (
    .A(alu_op_2_bF$buf1),
    .B(BI[2]),
    .C(_858_),
    .Y(_726_)
);

OAI21X1 _1329_ (
    .A(_312_),
    .B(_419_),
    .C(_324_),
    .Y(_420_)
);

INVX1 _1082_ (
    .A(_168_),
    .Y(_174_)
);

FILL FILL_0__1542_ (
);

FILL FILL_0__1122_ (
);

FILL FILL_1__1703_ (
);

OR2X2 _1558_ (
    .A(_643_),
    .B(_630_),
    .Y(_645_)
);

OAI21X1 _1138_ (
    .A(_81_),
    .B(_82_),
    .C(_79_),
    .Y(_230_)
);

FILL FILL_0__1771_ (
);

FILL FILL_0__1351_ (
);

FILL FILL_1__1512_ (
);

OAI21X1 _1787_ (
    .A(AI[4]),
    .B(_759_),
    .C(_868_),
    .Y(_762_)
);

OAI21X1 _1367_ (
    .A(_382_),
    .B(_393_),
    .C(_386_),
    .Y(_457_)
);

FILL FILL_0__1827_ (
);

FILL FILL_0__1407_ (
);

FILL FILL_0__1580_ (
);

FILL FILL_2__1598_ (
);

FILL FILL_0__1160_ (
);

FILL FILL_1__1741_ (
);

FILL FILL_1__1321_ (
);

INVX4 _1596_ (
    .A(reset),
    .Y(_1_)
);

INVX1 _1176_ (
    .A(BI[2]),
    .Y(_268_)
);

FILL FILL_1__958_ (
);

FILL FILL_0__1636_ (
);

FILL FILL_0__1216_ (
);

FILL FILL_1__1550_ (
);

FILL FILL_1__1130_ (
);

FILL FILL_0__1865_ (
);

FILL FILL_0__1445_ (
);

FILL FILL_0__1025_ (
);

FILL FILL_1__1606_ (
);

FILL FILL_1__996_ (
);

FILL FILL_0__1254_ (
);

FILL FILL_1__1835_ (
);

FILL FILL_1__1415_ (
);

FILL FILL_0__1483_ (
);

FILL FILL_0__1063_ (
);

FILL FILL_1__1644_ (
);

FILL FILL_1__1224_ (
);

NAND2X1 _1499_ (
    .A(_586_),
    .B(_585_),
    .Y(_587_)
);

OAI21X1 _1079_ (
    .A(_169_),
    .B(_37_),
    .C(_170_),
    .Y(_171_)
);

FILL FILL_0__1539_ (
);

FILL FILL_0__1119_ (
);

FILL FILL_0__1292_ (
);

INVX1 _1711_ (
    .A(_882_),
    .Y(ACC[0])
);

FILL FILL86250x46950 (
);

FILL FILL_1__1873_ (
);

FILL FILL_1__1453_ (
);

FILL FILL_1__1033_ (
);

FILL FILL_2__1102_ (
);

FILL FILL_0__1768_ (
);

FILL FILL_0__1348_ (
);

FILL FILL_1__1509_ (
);

AOI22X1 _1520_ (
    .A(_556_),
    .B(_607_),
    .C(_454_),
    .D(_442_),
    .Y(_608_)
);

INVX1 _1100_ (
    .A(_191_),
    .Y(_192_)
);

FILL FILL_1__1262_ (
);

FILL FILL_2__1331_ (
);

FILL FILL_0__1577_ (
);

FILL FILL_0__1157_ (
);

FILL FILL_1__1738_ (
);

FILL FILL_1__1318_ (
);

FILL FILL_1__1491_ (
);

FILL FILL_1__1071_ (
);

FILL FILL_2__1807_ (
);

FILL FILL86850x3750 (
);

FILL FILL_0__1386_ (
);

AOI22X1 _1805_ (
    .A(_862_),
    .B(BI[5]),
    .C(_777_),
    .D(_863_),
    .Y(_778_)
);

FILL FILL_1__1547_ (
);

FILL FILL_1__1127_ (
);

FILL FILL_1__920_ (
);

FILL FILL_0__1195_ (
);

OAI21X1 _1614_ (
    .A(LoadCmd_i),
    .B(_690_),
    .C(_691_),
    .Y(_7_)
);

FILL FILL_0__942_ (
);

NAND2X1 _945_ (
    .A(MUL_bF$buf2),
    .B(AI[3]),
    .Y(_37_)
);

FILL FILL_1__1776_ (
);

FILL FILL_1__1356_ (
);

AOI21X1 _1843_ (
    .A(alu_op_2_bF$buf2),
    .B(BI[7]),
    .C(_813_),
    .Y(_814_)
);

INVX1 _1423_ (
    .A(_512_),
    .Y(_513_)
);

AND2X2 _1003_ (
    .A(_92_),
    .B(_93_),
    .Y(_95_)
);

FILL FILL_1__1585_ (
);

FILL FILL_1__1165_ (
);

OAI21X1 _1652_ (
    .A(LoadB_i),
    .B(_288_),
    .C(_711_),
    .Y(_25_)
);

NAND2X1 _1232_ (
    .A(_320_),
    .B(_318_),
    .Y(_324_)
);

FILL FILL_0__980_ (
);

INVX1 _983_ (
    .A(_74_),
    .Y(_75_)
);

FILL FILL_1__1394_ (
);

FILL FILL_2__1043_ (
);

FILL FILL_0__1289_ (
);

OR2X2 _1708_ (
    .A(_879_),
    .B(_861_),
    .Y(_880_)
);

OR2X2 _1881_ (
    .A(_847_),
    .B(\u_ALU8.AI7 ),
    .Y(_849_)
);

NAND3X1 _1461_ (
    .A(_527_),
    .B(_549_),
    .C(_547_),
    .Y(_550_)
);

INVX1 _1041_ (
    .A(BI[6]),
    .Y(_133_)
);

FILL FILL_0__1501_ (
);

FILL FILL_2__1272_ (
);

FILL FILL_0__1098_ (
);

NAND2X1 _1517_ (
    .A(_556_),
    .B(_508_),
    .Y(_605_)
);

FILL FILL86550x54150 (
);

FILL FILL_1__1259_ (
);

INVX2 _1690_ (
    .A(alu_op[1]),
    .Y(_862_)
);

NAND2X1 _1270_ (
    .A(_353_),
    .B(_361_),
    .Y(_362_)
);

FILL FILL_0__1730_ (
);

FILL FILL_2__1748_ (
);

FILL FILL_0__1310_ (
);

AOI22X1 _1746_ (
    .A(_862_),
    .B(BI[2]),
    .C(_915_),
    .D(_863_),
    .Y(_916_)
);

INVX2 _1326_ (
    .A(\u_ALU8.AI7 ),
    .Y(_417_)
);

FILL FILL_1__1488_ (
);

FILL FILL_1__1068_ (
);

FILL FILL_1__1700_ (
);

NAND3X1 _1555_ (
    .A(_641_),
    .B(_638_),
    .C(_637_),
    .Y(_642_)
);

NOR2X1 _1135_ (
    .A(_220_),
    .B(_226_),
    .Y(_227_)
);

FILL FILL_1__1297_ (
);

FILL FILL_2_CLKBUF1_insert1 (
);

FILL FILL_0__939_ (
);

AND2X2 _1784_ (
    .A(_864_),
    .B(BI[4]),
    .Y(_759_)
);

NAND2X1 _1364_ (
    .A(_447_),
    .B(_351_),
    .Y(_454_)
);

FILL FILL_0__1824_ (
);

FILL FILL_0__1404_ (
);

FILL FILL_2__933_ (
);

OAI21X1 _1593_ (
    .A(_676_),
    .B(_358_),
    .C(_677_),
    .Y(_678_)
);

NAND2X1 _1173_ (
    .A(BI[1]),
    .B(_68_),
    .Y(_265_)
);

FILL FILL_1__955_ (
);

FILL FILL_0__1633_ (
);

FILL FILL_0__1213_ (
);

NAND2X1 _1649_ (
    .A(ABCmd_i[6]),
    .B(LoadB_i),
    .Y(_710_)
);

OAI21X1 _1229_ (
    .A(_316_),
    .B(_317_),
    .C(_320_),
    .Y(_321_)
);

FILL FILL_0__977_ (
);

FILL FILL86850x150 (
);

FILL FILL_0__1862_ (
);

FILL FILL_0__1442_ (
);

FILL FILL_0__1022_ (
);

FILL FILL_1__1603_ (
);

NAND2X1 _1878_ (
    .A(_877_),
    .B(_812_),
    .Y(_846_)
);

NAND3X1 _1458_ (
    .A(_543_),
    .B(_546_),
    .C(_528_),
    .Y(_547_)
);

NAND2X1 _1038_ (
    .A(BI[6]),
    .B(_68_),
    .Y(_130_)
);

FILL FILL_1__993_ (
);

FILL FILL_2__1689_ (
);

FILL FILL_0__1251_ (
);

FILL FILL_1__1832_ (
);

FILL FILL_1__1412_ (
);

OAI21X1 _1687_ (
    .A(_857_),
    .B(_858_),
    .C(CI),
    .Y(_859_)
);

AOI21X1 _1267_ (
    .A(_355_),
    .B(_358_),
    .C(_354_),
    .Y(_359_)
);

FILL FILL_0__1727_ (
);

FILL FILL_0__1307_ (
);

FILL FILL_0__1480_ (
);

FILL FILL_0__1060_ (
);

FILL FILL_1__1641_ (
);

FILL FILL_1__1221_ (
);

OAI21X1 _1496_ (
    .A(_135_),
    .B(_540_),
    .C(_583_),
    .Y(_584_)
);

NAND3X1 _1076_ (
    .A(MUL_bF$buf5),
    .B(AI[4]),
    .C(BI[4]),
    .Y(_168_)
);

FILL FILL_0__1536_ (
);

FILL FILL_0__1116_ (
);

FILL FILL_1__1870_ (
);

FILL FILL_1__1450_ (
);

FILL FILL_1__1030_ (
);

FILL FILL_0__1765_ (
);

FILL FILL_0__1345_ (
);

FILL FILL_1__1506_ (
);

FILL FILL85950x82950 (
);

FILL FILL_0__1574_ (
);

FILL FILL_0__1154_ (
);

FILL FILL_1__1735_ (
);

FILL FILL_1__1315_ (
);

FILL FILL_0__1383_ (
);

NAND2X1 _1802_ (
    .A(shr),
    .B(AI[6]),
    .Y(_775_)
);

FILL FILL_1__1544_ (
);

FILL FILL_1__1124_ (
);

INVX1 _1399_ (
    .A(_488_),
    .Y(_489_)
);

FILL FILL_0__1859_ (
);

FILL FILL_0__1439_ (
);

FILL FILL_0__1019_ (
);

FILL FILL_0__1192_ (
);

OAI21X1 _1611_ (
    .A(LoadCmd_i),
    .B(_688_),
    .C(_689_),
    .Y(_6_)
);

NOR2X1 _942_ (
    .A(_32_),
    .B(_33_),
    .Y(_34_)
);

FILL FILL_1__1773_ (
);

FILL FILL_1__1353_ (
);

FILL FILL_2__1422_ (
);

FILL FILL_0__1248_ (
);

FILL FILL_1__1829_ (
);

FILL FILL_1__1409_ (
);

OAI21X1 _1840_ (
    .A(\u_ALU8.AI7 ),
    .B(_808_),
    .C(_868_),
    .Y(_811_)
);

OAI21X1 _1420_ (
    .A(_379_),
    .B(_509_),
    .C(_439_),
    .Y(_510_)
);

NAND3X1 _1000_ (
    .A(MUL_bF$buf1),
    .B(BI[1]),
    .C(AI[5]),
    .Y(_92_)
);

FILL FILL_1__1582_ (
);

FILL FILL_1__1162_ (
);

FILL FILL_2__1651_ (
);

FILL FILL_0__1897_ (
);

FILL FILL_0__1477_ (
);

FILL FILL_0__1057_ (
);

FILL FILL86250x32550 (
);

FILL FILL_1__1638_ (
);

FILL FILL_1__1218_ (
);

NAND3X1 _980_ (
    .A(MUL_bF$buf4),
    .B(BI[3]),
    .C(AI[2]),
    .Y(_72_)
);

FILL FILL_1__1391_ (
);

FILL FILL_0__1286_ (
);

NOR2X1 _1705_ (
    .A(alu_op_2_bF$buf3),
    .B(_858_),
    .Y(_877_)
);

FILL FILL_1__1867_ (
);

FILL FILL_1__1447_ (
);

FILL FILL_1__1027_ (
);

FILL FILL_0__1095_ (
);

NAND3X1 _1514_ (
    .A(_576_),
    .B(_596_),
    .C(_599_),
    .Y(_602_)
);

FILL FILL_1__1256_ (
);

FILL FILL86550x75750 (
);

INVX1 _1743_ (
    .A(BI[2]),
    .Y(_913_)
);

NAND2X1 _1323_ (
    .A(_413_),
    .B(_409_),
    .Y(_414_)
);

FILL FILL_1__1485_ (
);

FILL FILL_1__1065_ (
);

NAND2X1 _1552_ (
    .A(_638_),
    .B(_637_),
    .Y(_639_)
);

NAND3X1 _1132_ (
    .A(_30_),
    .B(_38_),
    .C(_35_),
    .Y(_224_)
);

FILL FILL_1__1294_ (
);

FILL FILL_2__1363_ (
);

FILL FILL_0__1189_ (
);

OAI21X1 _1608_ (
    .A(LoadCmd_i),
    .B(_686_),
    .C(_687_),
    .Y(_5_)
);

FILL FILL_0__936_ (
);

INVX1 _939_ (
    .A(_30_),
    .Y(_31_)
);

INVX1 _1781_ (
    .A(_746_),
    .Y(_756_)
);

OAI21X1 _1361_ (
    .A(_451_),
    .B(_450_),
    .C(MulH_i),
    .Y(_452_)
);

FILL FILL_0__1821_ (
);

FILL FILL_2__1839_ (
);

FILL FILL_0__1401_ (
);

FILL FILL_2__1592_ (
);

AND2X2 _1837_ (
    .A(_864_),
    .B(BI[7]),
    .Y(_808_)
);

NAND2X1 _1417_ (
    .A(_503_),
    .B(_506_),
    .Y(_507_)
);

FILL FILL_1__1579_ (
);

FILL FILL_1__1159_ (
);

NOR2X1 _1590_ (
    .A(_712_),
    .B(_674_),
    .Y(_675_)
);

NAND3X1 _1170_ (
    .A(_246_),
    .B(_260_),
    .C(_261_),
    .Y(_262_)
);

FILL FILL_1__952_ (
);

FILL FILL_0__1630_ (
);

FILL FILL_0__1210_ (
);

INVX1 _1646_ (
    .A(BI[5]),
    .Y(_708_)
);

NOR2X1 _1226_ (
    .A(_316_),
    .B(_317_),
    .Y(_318_)
);

FILL FILL_0__974_ (
);

NAND2X1 _977_ (
    .A(BI[5]),
    .B(_68_),
    .Y(_69_)
);

FILL FILL_1__1388_ (
);

FILL FILL_2__1037_ (
);

FILL FILL_1__1600_ (
);

NOR2X1 _1875_ (
    .A(_816_),
    .B(_842_),
    .Y(_843_)
);

INVX1 _1455_ (
    .A(_537_),
    .Y(_544_)
);

OAI21X1 _1035_ (
    .A(_122_),
    .B(_121_),
    .C(_119_),
    .Y(_127_)
);

FILL FILL_1__1197_ (
);

FILL FILL_1__990_ (
);

DFFPOSX1 _1684_ (
    .D(_25_),
    .CLK(clk_bF$buf2),
    .Q(BI[7])
);

NAND2X1 _1264_ (
    .A(_144_),
    .B(_258_),
    .Y(_356_)
);

FILL FILL_0__1724_ (
);

FILL FILL_0__1304_ (
);

NAND2X1 _1493_ (
    .A(AI[5]),
    .B(_289_),
    .Y(_581_)
);

NAND3X1 _1073_ (
    .A(_164_),
    .B(_162_),
    .C(_163_),
    .Y(_165_)
);

FILL FILL_0__1533_ (
);

FILL FILL_0__1113_ (
);

OAI21X1 _1549_ (
    .A(_582_),
    .B(_634_),
    .C(_635_),
    .Y(_636_)
);

INVX1 _1129_ (
    .A(_724_),
    .Y(_221_)
);

FILL FILL_0__1762_ (
);

FILL FILL_0__1342_ (
);

FILL FILL_1__1503_ (
);

AOI21X1 _1778_ (
    .A(_735_),
    .B(_909_),
    .C(_752_),
    .Y(_753_)
);

AOI21X1 _1358_ (
    .A(_353_),
    .B(_351_),
    .C(_448_),
    .Y(_449_)
);

FILL FILL_0__1818_ (
);

FILL FILL_2__927_ (
);

FILL FILL_0__1571_ (
);

FILL FILL_0__1151_ (
);

FILL FILL_1__1732_ (
);

FILL FILL_1__1312_ (
);

NAND3X1 _1587_ (
    .A(MulH_i),
    .B(_672_),
    .C(_668_),
    .Y(_673_)
);

AND2X2 _1167_ (
    .A(_258_),
    .B(_144_),
    .Y(_259_)
);

FILL FILL_1__949_ (
);

FILL FILL_0__1627_ (
);

FILL FILL_0__1207_ (
);

FILL FILL_0__1380_ (
);

FILL FILL_1__1541_ (
);

FILL FILL_1__1121_ (
);

NAND2X1 _1396_ (
    .A(_485_),
    .B(_482_),
    .Y(_486_)
);

FILL FILL_0__1856_ (
);

FILL FILL_0__1436_ (
);

FILL FILL_0__1016_ (
);

FILL FILL_1__1770_ (
);

FILL FILL_1__1350_ (
);

FILL FILL_1__987_ (
);

FILL FILL_0__1245_ (
);

FILL FILL_1__1826_ (
);

FILL FILL_1__1406_ (
);

FILL FILL_0__1894_ (
);

FILL FILL_0__1474_ (
);

FILL FILL_0__1054_ (
);

FILL FILL_1__1635_ (
);

FILL FILL_1__1215_ (
);

FILL FILL_0__1283_ (
);

OAI21X1 _1702_ (
    .A(_867_),
    .B(_872_),
    .C(_873_),
    .Y(_874_)
);

FILL FILL_1__1864_ (
);

FILL FILL_1__1444_ (
);

FILL FILL_1__1024_ (
);

NAND3X1 _1299_ (
    .A(_383_),
    .B(_389_),
    .C(_386_),
    .Y(_390_)
);

FILL FILL_0__1759_ (
);

FILL FILL_0__1339_ (
);

FILL FILL_0__1092_ (
);

NAND3X1 _1511_ (
    .A(_579_),
    .B(_598_),
    .C(_597_),
    .Y(_599_)
);

FILL FILL_1__1253_ (
);

FILL FILL_0__1568_ (
);

FILL FILL_0__1148_ (
);

FILL FILL_1__1729_ (
);

FILL FILL_1__1309_ (
);

NOR2X1 _1740_ (
    .A(_893_),
    .B(_891_),
    .Y(_910_)
);

NAND3X1 _1320_ (
    .A(_397_),
    .B(_402_),
    .C(_400_),
    .Y(_411_)
);

FILL FILL_1__1482_ (
);

FILL FILL_1__1062_ (
);

FILL FILL_0__1797_ (
);

FILL FILL_0__1377_ (
);

FILL FILL_1__1538_ (
);

FILL FILL_1__1118_ (
);

FILL FILL_1__1291_ (
);

FILL FILL_0__1186_ (
);

OAI21X1 _1605_ (
    .A(LoadCmd_i),
    .B(_684_),
    .C(_685_),
    .Y(_4_)
);

FILL FILL_0__933_ (
);

INVX1 _936_ (
    .A(_27_),
    .Y(_28_)
);

FILL FILL_1__1767_ (
);

FILL FILL_1__1347_ (
);

FILL FILL_2__1416_ (
);

INVX1 _1834_ (
    .A(_799_),
    .Y(_805_)
);

NAND3X1 _1414_ (
    .A(_490_),
    .B(_493_),
    .C(_495_),
    .Y(_504_)
);

FILL FILL_1__1576_ (
);

FILL FILL_1__1156_ (
);

OAI21X1 _1643_ (
    .A(LoadB_i),
    .B(_309_),
    .C(_706_),
    .Y(_21_)
);

NAND3X1 _1223_ (
    .A(MUL_bF$buf5),
    .B(\u_ALU8.AI7 ),
    .C(BI[1]),
    .Y(_315_)
);

FILL FILL_0__971_ (
);

NAND3X1 _974_ (
    .A(_63_),
    .B(_65_),
    .C(_64_),
    .Y(_66_)
);

FILL FILL_1__1385_ (
);

NAND2X1 _1872_ (
    .A(_833_),
    .B(_837_),
    .Y(_840_)
);

OAI21X1 _1452_ (
    .A(_417_),
    .B(_44_),
    .C(_538_),
    .Y(_541_)
);

OAI21X1 _1032_ (
    .A(_122_),
    .B(_121_),
    .C(_123_),
    .Y(_124_)
);

FILL FILL_0_CLKBUF1_insert0 (
);

FILL FILL_0_CLKBUF1_insert1 (
);

FILL FILL_0_CLKBUF1_insert2 (
);

FILL FILL_0_CLKBUF1_insert3 (
);

FILL FILL_0_CLKBUF1_insert4 (
);

FILL FILL_1__1194_ (
);

FILL FILL_0__1089_ (
);

OAI21X1 _1508_ (
    .A(_594_),
    .B(_595_),
    .C(_580_),
    .Y(_596_)
);

DFFPOSX1 _1681_ (
    .D(_22_),
    .CLK(clk_bF$buf0),
    .Q(BI[4])
);

NAND2X1 _1261_ (
    .A(_352_),
    .B(_283_),
    .Y(_353_)
);

FILL FILL_0__1721_ (
);

FILL FILL_0__1301_ (
);

NAND2X1 _1737_ (
    .A(_905_),
    .B(_907_),
    .Y(_908_)
);

NAND3X1 _1317_ (
    .A(MUL_bF$buf0),
    .B(\u_ALU8.AI7 ),
    .C(BI[2]),
    .Y(_408_)
);

FILL FILL_1__1479_ (
);

FILL FILL_1__1059_ (
);

NAND2X1 _1490_ (
    .A(_534_),
    .B(_532_),
    .Y(_578_)
);

OAI21X1 _1070_ (
    .A(_96_),
    .B(_95_),
    .C(_99_),
    .Y(_162_)
);

FILL FILL_0__1530_ (
);

FILL FILL_2__1128_ (
);

FILL FILL_0__1110_ (
);

AOI21X1 _1546_ (
    .A(_631_),
    .B(_583_),
    .C(_632_),
    .Y(_633_)
);

NAND3X1 _1126_ (
    .A(_145_),
    .B(_214_),
    .C(_217_),
    .Y(_218_)
);

FILL FILL_1__1288_ (
);

FILL FILL_2__1357_ (
);

FILL FILL_1__1500_ (
);

NAND2X1 _1775_ (
    .A(_750_),
    .B(_749_),
    .Y(_751_)
);

NAND3X1 _1355_ (
    .A(_379_),
    .B(_437_),
    .C(_430_),
    .Y(_446_)
);

FILL FILL_1__1097_ (
);

FILL FILL_0__1815_ (
);

NAND3X1 _1584_ (
    .A(_606_),
    .B(_669_),
    .C(_609_),
    .Y(_670_)
);

INVX1 _1164_ (
    .A(_255_),
    .Y(_256_)
);

FILL FILL_1__946_ (
);

FILL FILL_0__1624_ (
);

FILL FILL_0__1204_ (
);

FILL FILL_0__968_ (
);

NOR2X1 _1393_ (
    .A(_477_),
    .B(_478_),
    .Y(_483_)
);

FILL FILL_0__1853_ (
);

FILL FILL_0__1433_ (
);

FILL FILL_0__1013_ (
);

AND2X2 _1869_ (
    .A(_837_),
    .B(_833_),
    .Y(_838_)
);

NAND2X1 _1449_ (
    .A(BI[5]),
    .B(_405_),
    .Y(_538_)
);

AOI21X1 _1029_ (
    .A(_104_),
    .B(_105_),
    .C(_103_),
    .Y(_121_)
);

FILL FILL_1__984_ (
);

FILL FILL_0__1242_ (
);

FILL FILL_1__1823_ (
);

FILL FILL_1__1403_ (
);

DFFPOSX1 _1678_ (
    .D(_19_),
    .CLK(clk_bF$buf0),
    .Q(BI[1])
);

NAND3X1 _1258_ (
    .A(_286_),
    .B(_341_),
    .C(_337_),
    .Y(_350_)
);

FILL FILL_0__1718_ (
);

FILL FILL_0__1891_ (
);

FILL FILL_0__1471_ (
);

FILL FILL_0__1051_ (
);

FILL FILL_2__1069_ (
);

FILL FILL86850x36150 (
);

FILL FILL_1__1632_ (
);

FILL FILL_1__1212_ (
);

OAI21X1 _1487_ (
    .A(_712_),
    .B(_568_),
    .C(_575_),
    .Y(_0_[3])
);

OAI21X1 _1067_ (
    .A(_36_),
    .B(_158_),
    .C(_151_),
    .Y(_159_)
);

FILL FILL_0__1527_ (
);

FILL FILL_0__1107_ (
);

FILL FILL_2__1298_ (
);

FILL FILL_0__1280_ (
);

FILL FILL_1__1861_ (
);

FILL FILL_1__1441_ (
);

FILL FILL_1__1021_ (
);

INVX1 _1296_ (
    .A(AI[3]),
    .Y(_387_)
);

FILL FILL_0__1756_ (
);

FILL FILL_0__1336_ (
);

FILL FILL_1__1250_ (
);

FILL FILL_0__1565_ (
);

FILL FILL_0__1145_ (
);

FILL FILL_1__1726_ (
);

FILL FILL_1__1306_ (
);

FILL FILL_0__1794_ (
);

FILL FILL_0__1374_ (
);

FILL FILL_1__1535_ (
);

FILL FILL_1__1115_ (
);

FILL FILL_2__959_ (
);

FILL FILL_0__1183_ (
);

OAI21X1 _1602_ (
    .A(LoadCmd_i),
    .B(_682_),
    .C(_683_),
    .Y(_3_)
);

FILL FILL_0__930_ (
);

INVX2 _933_ (
    .A(AI[2]),
    .Y(_725_)
);

FILL FILL_1__1764_ (
);

FILL FILL_1__1344_ (
);

INVX1 _1199_ (
    .A(_290_),
    .Y(_291_)
);

FILL FILL_2__1833_ (
);

FILL FILL_0__1239_ (
);

NAND3X1 _1831_ (
    .A(_783_),
    .B(_800_),
    .C(_786_),
    .Y(_803_)
);

AOI21X1 _1411_ (
    .A(_498_),
    .B(_500_),
    .C(_474_),
    .Y(_501_)
);

FILL FILL_1__1573_ (
);

FILL FILL_1__1153_ (
);

FILL FILL_0__1888_ (
);

FILL FILL_0__1468_ (
);

FILL FILL_0__1048_ (
);

FILL FILL_1__1629_ (
);

FILL FILL_1__1209_ (
);

NAND2X1 _1640_ (
    .A(ABCmd_i[2]),
    .B(LoadB_i),
    .Y(_705_)
);

NAND2X1 _1220_ (
    .A(_306_),
    .B(_311_),
    .Y(_312_)
);

AOI21X1 _971_ (
    .A(_31_),
    .B(_38_),
    .C(_34_),
    .Y(_63_)
);

FILL FILL_1__1382_ (
);

FILL FILL_0__1697_ (
);

FILL FILL_0__1277_ (
);

FILL FILL_1__1858_ (
);

FILL FILL_1__1438_ (
);

FILL FILL_1__1018_ (
);

FILL FILL_1__1191_ (
);

FILL FILL_2__1507_ (
);

FILL FILL_0__1086_ (
);

NAND2X1 _1505_ (
    .A(_592_),
    .B(_588_),
    .Y(_593_)
);

FILL FILL_1__1247_ (
);

FILL FILL86550x82950 (
);

AOI22X1 _1734_ (
    .A(_874_),
    .B(_899_),
    .C(_904_),
    .D(_860_),
    .Y(_905_)
);

AND2X2 _1314_ (
    .A(MUL_bF$buf3),
    .B(AI[6]),
    .Y(_405_)
);

FILL FILL_1__1896_ (
);

FILL FILL_1__1476_ (
);

FILL FILL_1__1056_ (
);

AOI21X1 _1543_ (
    .A(_579_),
    .B(_598_),
    .C(_594_),
    .Y(_630_)
);

AOI21X1 _1123_ (
    .A(_212_),
    .B(_211_),
    .C(_210_),
    .Y(_215_)
);

FILL FILL_1__1285_ (
);

FILL FILL_2__1774_ (
);

FILL FILL_0__927_ (
);

INVX1 _1772_ (
    .A(_747_),
    .Y(_748_)
);

AOI21X1 _1352_ (
    .A(_332_),
    .B(_336_),
    .C(_287_),
    .Y(_443_)
);

FILL FILL_1__1094_ (
);

FILL FILL_0__1812_ (
);

OAI21X1 _1828_ (
    .A(_796_),
    .B(_798_),
    .C(_799_),
    .Y(_800_)
);

NAND3X1 _1408_ (
    .A(_416_),
    .B(_413_),
    .C(_497_),
    .Y(_498_)
);

INVX1 _1581_ (
    .A(_666_),
    .Y(_667_)
);

AOI21X1 _1161_ (
    .A(_230_),
    .B(_231_),
    .C(_229_),
    .Y(_253_)
);

FILL FILL_1__943_ (
);

FILL FILL_0__1621_ (
);

FILL FILL_0__1201_ (
);

OAI21X1 _1637_ (
    .A(LoadB_i),
    .B(_53_),
    .C(_703_),
    .Y(_18_)
);

INVX1 _1217_ (
    .A(BI[3]),
    .Y(_309_)
);

FILL FILL_0__965_ (
);

INVX1 _968_ (
    .A(_55_),
    .Y(_60_)
);

FILL FILL_1__1799_ (
);

FILL FILL_1__1379_ (
);

INVX1 _1390_ (
    .A(AI[6]),
    .Y(_480_)
);

FILL FILL_0__1850_ (
);

FILL FILL_2__1448_ (
);

FILL FILL_0__1430_ (
);

FILL FILL_0__1010_ (
);

AOI21X1 _1866_ (
    .A(_786_),
    .B(_783_),
    .C(_834_),
    .Y(_835_)
);

NAND3X1 _1446_ (
    .A(_530_),
    .B(_534_),
    .C(_532_),
    .Y(_535_)
);

NAND3X1 _1026_ (
    .A(_107_),
    .B(_112_),
    .C(_117_),
    .Y(_118_)
);

FILL FILL_1__1188_ (
);

FILL FILL_1__981_ (
);

FILL FILL_1__1820_ (
);

FILL FILL_1__1400_ (
);

DFFPOSX1 _1675_ (
    .D(_16_),
    .CLK(clk_bF$buf1),
    .Q(AI[6])
);

OAI21X1 _1255_ (
    .A(_346_),
    .B(_342_),
    .C(_284_),
    .Y(_347_)
);

FILL FILL_0__1715_ (
);

OAI21X1 _1484_ (
    .A(Flag_i),
    .B(ACC[3]),
    .C(_365_),
    .Y(_573_)
);

OAI21X1 _1064_ (
    .A(_152_),
    .B(_153_),
    .C(_155_),
    .Y(_156_)
);

FILL FILL86850x57750 (
);

FILL FILL_0__1524_ (
);

FILL FILL_0__1104_ (
);

INVX1 _1293_ (
    .A(_37_),
    .Y(_384_)
);

FILL FILL_0__1753_ (
);

FILL FILL_0__1333_ (
);

AOI21X1 _1769_ (
    .A(alu_op_2_bF$buf3),
    .B(BI[3]),
    .C(_744_),
    .Y(_745_)
);

OAI21X1 _1349_ (
    .A(_433_),
    .B(_436_),
    .C(_381_),
    .Y(_440_)
);

FILL FILL_0__1809_ (
);

FILL FILL_0__1562_ (
);

FILL FILL_0__1142_ (
);

FILL FILL_1__1723_ (
);

FILL FILL_1__1303_ (
);

OR2X2 _1578_ (
    .A(_662_),
    .B(_663_),
    .Y(_664_)
);

OAI21X1 _1158_ (
    .A(_225_),
    .B(_47_),
    .C(_46_),
    .Y(_250_)
);

FILL FILL_0__1618_ (
);

FILL FILL_0__1791_ (
);

FILL FILL_2__1389_ (
);

FILL FILL_0__1371_ (
);

FILL FILL_1__1532_ (
);

FILL FILL_1__1112_ (
);

NAND3X1 _1387_ (
    .A(MUL_bF$buf3),
    .B(AI[6]),
    .C(BI[4]),
    .Y(_477_)
);

FILL FILL_0__1847_ (
);

FILL FILL_0__1427_ (
);

FILL FILL_0__1007_ (
);

FILL FILL_0__1180_ (
);

NOR2X1 _930_ (
    .A(_720_),
    .B(_721_),
    .Y(_722_)
);

FILL FILL_1__1761_ (
);

FILL FILL_1__1341_ (
);

INVX1 _1196_ (
    .A(BI[7]),
    .Y(_288_)
);

FILL FILL_1__978_ (
);

FILL FILL_0__1236_ (
);

FILL FILL_1__1817_ (
);

FILL FILL_1__1570_ (
);

FILL FILL_1__1150_ (
);

BUFX2 BUFX2_insert10 (
    .A(MUL),
    .Y(MUL_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf3)
);

BUFX2 BUFX2_insert12 (
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf0)
);

FILL FILL_0__1885_ (
);

FILL FILL_0__1465_ (
);

FILL FILL_0__1045_ (
);

FILL FILL_1__1626_ (
);

FILL FILL_1__1206_ (
);

FILL FILL_0__1694_ (
);

FILL FILL_0__1274_ (
);

FILL FILL_1__1855_ (
);

FILL FILL_1__1435_ (
);

FILL FILL_1__1015_ (
);

FILL FILL_0__1083_ (
);

NAND2X1 _1502_ (
    .A(\u_ALU8.AI7 ),
    .B(_589_),
    .Y(_590_)
);

FILL FILL_1__1244_ (
);

NAND2X1 _1099_ (
    .A(BI[7]),
    .B(_68_),
    .Y(_191_)
);

FILL FILL_0__1559_ (
);

FILL FILL_0__1139_ (
);

NAND2X1 _1731_ (
    .A(_901_),
    .B(_900_),
    .Y(_902_)
);

OAI21X1 _1311_ (
    .A(_401_),
    .B(_44_),
    .C(_399_),
    .Y(_402_)
);

FILL FILL_1__1893_ (
);

FILL FILL_1__1473_ (
);

FILL FILL_1__1053_ (
);

FILL FILL_2__1122_ (
);

FILL FILL_0__1788_ (
);

FILL FILL_0__1368_ (
);

FILL FILL_1__1529_ (
);

FILL FILL_1__1109_ (
);

NOR2X1 _1540_ (
    .A(Flag_i),
    .B(MulL_i),
    .Y(_627_)
);

OAI21X1 _1120_ (
    .A(_190_),
    .B(_186_),
    .C(_207_),
    .Y(_212_)
);

FILL FILL_1__1282_ (
);

FILL FILL_0__1597_ (
);

FILL FILL_0__1177_ (
);

FILL FILL_0__924_ (
);

OR2X2 _927_ (
    .A(_718_),
    .B(_714_),
    .Y(_719_)
);

FILL FILL_1__1758_ (
);

FILL FILL_1__1338_ (
);

FILL FILL_1__1091_ (
);

OAI21X1 _1825_ (
    .A(alu_op_2_bF$buf2),
    .B(BI[6]),
    .C(_858_),
    .Y(_797_)
);

OAI21X1 _1405_ (
    .A(_395_),
    .B(_421_),
    .C(_426_),
    .Y(_495_)
);

FILL FILL_1__1567_ (
);

FILL FILL_1__1147_ (
);

FILL FILL_1__940_ (
);

NAND2X1 _1634_ (
    .A(ABCmd_i[7]),
    .B(LoadA_i),
    .Y(_702_)
);

OAI21X1 _1214_ (
    .A(_304_),
    .B(_305_),
    .C(_302_),
    .Y(_306_)
);

FILL FILL_0__962_ (
);

INVX1 _965_ (
    .A(_56_),
    .Y(_57_)
);

FILL FILL_1__1796_ (
);

FILL FILL_1__1376_ (
);

NOR2X1 _1863_ (
    .A(_870_),
    .B(_868_),
    .Y(_832_)
);

NAND3X1 _1443_ (
    .A(AI[5]),
    .B(_134_),
    .C(_531_),
    .Y(_532_)
);

INVX1 _1023_ (
    .A(_109_),
    .Y(_115_)
);

FILL FILL_1__1185_ (
);

DFFPOSX1 _1672_ (
    .D(_13_),
    .CLK(clk_bF$buf0),
    .Q(AI[3])
);

NAND3X1 _1252_ (
    .A(_332_),
    .B(_336_),
    .C(_338_),
    .Y(_344_)
);

FILL FILL_0__1712_ (
);

FILL FILL_2__1063_ (
);

OAI21X1 _1728_ (
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_898_),
    .Y(_899_)
);

NAND3X1 _1308_ (
    .A(MUL_bF$buf0),
    .B(AI[6]),
    .C(BI[3]),
    .Y(_399_)
);

OAI21X1 _1481_ (
    .A(_270_),
    .B(_569_),
    .C(MulL_i),
    .Y(_570_)
);

AND2X2 _1061_ (
    .A(_150_),
    .B(_151_),
    .Y(_153_)
);

FILL FILL_0__1521_ (
);

FILL FILL_0__1101_ (
);

NAND2X1 _1537_ (
    .A(_255_),
    .B(_279_),
    .Y(_624_)
);

NAND3X1 _1117_ (
    .A(_208_),
    .B(_204_),
    .C(_147_),
    .Y(_209_)
);

FILL FILL_1__1699_ (
);

FILL FILL_1__1279_ (
);

AOI21X1 _1290_ (
    .A(_333_),
    .B(_335_),
    .C(_380_),
    .Y(_381_)
);

FILL FILL_2__1768_ (
);

FILL FILL_0__1750_ (
);

FILL FILL_0__1330_ (
);

OAI21X1 _1766_ (
    .A(AI[3]),
    .B(_739_),
    .C(_868_),
    .Y(_742_)
);

OAI21X1 _1346_ (
    .A(_436_),
    .B(_433_),
    .C(_432_),
    .Y(_437_)
);

FILL FILL_1__1088_ (
);

FILL FILL_0__1806_ (
);

FILL FILL_1__1720_ (
);

FILL FILL_1__1300_ (
);

OAI21X1 _1575_ (
    .A(_602_),
    .B(_646_),
    .C(_645_),
    .Y(_661_)
);

NAND2X1 _1155_ (
    .A(BI[3]),
    .B(_68_),
    .Y(_247_)
);

FILL FILL_1__937_ (
);

FILL FILL_0__1615_ (
);

FILL FILL_0__959_ (
);

NAND2X1 _1384_ (
    .A(_470_),
    .B(_473_),
    .Y(_474_)
);

FILL FILL_0__1844_ (
);

FILL FILL_0__1424_ (
);

FILL FILL_0__1004_ (
);

FILL FILL_2__953_ (
);

NOR2X1 _1193_ (
    .A(_197_),
    .B(_194_),
    .Y(_285_)
);

FILL FILL_1__975_ (
);

FILL FILL_0__1233_ (
);

FILL FILL_1__1814_ (
);

FILL FILL86850x43350 (
);

DFFPOSX1 _1669_ (
    .D(_10_),
    .CLK(clk_bF$buf0),
    .Q(AI[0])
);

OAI21X1 _1249_ (
    .A(_339_),
    .B(_340_),
    .C(_338_),
    .Y(_341_)
);

FILL FILL_0__997_ (
);

FILL FILL_0__1709_ (
);

FILL FILL_0__1882_ (
);

FILL FILL_0__1462_ (
);

FILL FILL_0__1042_ (
);

FILL FILL_1__1623_ (
);

FILL FILL_1__1203_ (
);

OAI21X1 _1478_ (
    .A(_562_),
    .B(_565_),
    .C(_566_),
    .Y(_567_)
);

NAND3X1 _1058_ (
    .A(MUL_bF$buf5),
    .B(BI[1]),
    .C(AI[6]),
    .Y(_150_)
);

FILL FILL_0__1518_ (
);

FILL FILL_0__1691_ (
);

FILL FILL_0__1271_ (
);

FILL FILL_1__1852_ (
);

FILL FILL_1__1432_ (
);

FILL FILL_1__1012_ (
);

OAI21X1 _1287_ (
    .A(_290_),
    .B(_298_),
    .C(_294_),
    .Y(_378_)
);

FILL FILL_0__1747_ (
);

FILL FILL_0__1327_ (
);

FILL FILL_0__1080_ (
);

FILL FILL_1__1241_ (
);

OAI21X1 _1096_ (
    .A(_180_),
    .B(_179_),
    .C(_177_),
    .Y(_188_)
);

FILL FILL_0__1556_ (
);

FILL FILL_0__1136_ (
);

FILL FILL_1__1717_ (
);

FILL FILL_1__1890_ (
);

FILL FILL_1__1470_ (
);

FILL FILL_1__1050_ (
);

FILL FILL_0__1785_ (
);

FILL FILL_0__1365_ (
);

FILL FILL_1__1526_ (
);

FILL FILL_1__1106_ (
);

FILL FILL_0__1594_ (
);

FILL FILL_0__1174_ (
);

FILL FILL_0__921_ (
);

INVX2 _924_ (
    .A(AI[1]),
    .Y(_716_)
);

FILL FILL_1__1755_ (
);

FILL FILL_1__1335_ (
);

AOI22X1 _1822_ (
    .A(_862_),
    .B(BI[6]),
    .C(_793_),
    .D(_863_),
    .Y(_794_)
);

INVX1 _1402_ (
    .A(_487_),
    .Y(_492_)
);

FILL FILL_1__1564_ (
);

FILL FILL_1__1144_ (
);

FILL FILL_2__1213_ (
);

FILL FILL_0__1879_ (
);

FILL FILL_0__1459_ (
);

FILL FILL_0__1039_ (
);

OAI21X1 _1631_ (
    .A(LoadA_i),
    .B(_401_),
    .C(_700_),
    .Y(_15_)
);

NAND3X1 _1211_ (
    .A(MUL_bF$buf5),
    .B(AI[5]),
    .C(BI[3]),
    .Y(_303_)
);

NAND2X1 _962_ (
    .A(MUL_bF$buf2),
    .B(AI[5]),
    .Y(_54_)
);

FILL FILL_1__1793_ (
);

FILL FILL_1__1373_ (
);

FILL FILL_2__1442_ (
);

FILL FILL_0__1688_ (
);

FILL FILL_0__1268_ (
);

FILL FILL_1__1849_ (
);

FILL FILL_1__1429_ (
);

FILL FILL_1__1009_ (
);

INVX1 _1860_ (
    .A(_828_),
    .Y(_829_)
);

NAND2X1 _1440_ (
    .A(BI[7]),
    .B(_464_),
    .Y(_529_)
);

OAI21X1 _1020_ (
    .A(_725_),
    .B(_44_),
    .C(_110_),
    .Y(_112_)
);

FILL FILL_1__1182_ (
);

FILL FILL_0__1497_ (
);

FILL FILL_0__1077_ (
);

FILL FILL_1__1238_ (
);

MUX2X1 _1725_ (
    .A(_895_),
    .B(_894_),
    .S(_891_),
    .Y(_896_)
);

NAND3X1 _1305_ (
    .A(MUL_bF$buf3),
    .B(AI[4]),
    .C(BI[5]),
    .Y(_396_)
);

FILL FILL_1__1887_ (
);

FILL FILL_1__1467_ (
);

FILL FILL_1__1047_ (
);

FILL FILL86250x68550 (
);

OAI21X1 _1534_ (
    .A(_620_),
    .B(_621_),
    .C(_619_),
    .Y(_622_)
);

NAND3X1 _1114_ (
    .A(_178_),
    .B(_185_),
    .C(_148_),
    .Y(_206_)
);

FILL FILL_1__1696_ (
);

FILL FILL_1__1276_ (
);

AND2X2 _1763_ (
    .A(_864_),
    .B(BI[3]),
    .Y(_739_)
);

NAND2X1 _1343_ (
    .A(_427_),
    .B(_425_),
    .Y(_434_)
);

FILL FILL_1__1085_ (
);

FILL FILL_0__1803_ (
);

FILL FILL_2__1154_ (
);

INVX1 _1819_ (
    .A(\u_ALU8.AI7 ),
    .Y(_791_)
);

NAND2X1 _1572_ (
    .A(_712_),
    .B(_657_),
    .Y(_658_)
);

OAI21X1 _1152_ (
    .A(_241_),
    .B(_243_),
    .C(_240_),
    .Y(_244_)
);

FILL FILL_1__934_ (
);

FILL FILL_0__1612_ (
);

FILL FILL_2__1383_ (
);

NAND2X1 _1628_ (
    .A(ABCmd_i[4]),
    .B(LoadA_i),
    .Y(_699_)
);

NAND2X1 _1208_ (
    .A(_299_),
    .B(_296_),
    .Y(_300_)
);

FILL FILL_0__956_ (
);

NAND3X1 _959_ (
    .A(MUL_bF$buf2),
    .B(BI[0]),
    .C(AI[5]),
    .Y(_51_)
);

NOR2X1 _1381_ (
    .A(_465_),
    .B(_468_),
    .Y(_471_)
);

FILL FILL_0__1841_ (
);

FILL FILL_2__1859_ (
);

FILL FILL_0__1421_ (
);

FILL FILL_0__1001_ (
);

NAND2X1 _1857_ (
    .A(_819_),
    .B(_818_),
    .Y(_826_)
);

OAI21X1 _1437_ (
    .A(_460_),
    .B(_472_),
    .C(_467_),
    .Y(_526_)
);

NAND3X1 _1017_ (
    .A(MUL_bF$buf1),
    .B(BI[4]),
    .C(AI[2]),
    .Y(_109_)
);

FILL FILL_1__1599_ (
);

FILL FILL_1__1179_ (
);

OAI21X1 _1190_ (
    .A(_256_),
    .B(_281_),
    .C(_259_),
    .Y(_282_)
);

FILL FILL_1__972_ (
);

FILL FILL_0__1650_ (
);

FILL FILL_0__1230_ (
);

FILL FILL_1__1811_ (
);

DFFSR _1666_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[5]),
    .CLK(clk_bF$buf3),
    .Q(_919_[5])
);

AOI21X1 _1246_ (
    .A(_203_),
    .B(_205_),
    .C(_190_),
    .Y(_338_)
);

FILL FILL_0__994_ (
);

OAI21X1 _997_ (
    .A(_719_),
    .B(_88_),
    .C(_87_),
    .Y(_89_)
);

FILL FILL_0__1706_ (
);

FILL FILL86850x64950 (
);

FILL FILL_1__1620_ (
);

FILL FILL_1__1200_ (
);

BUFX2 _1895_ (
    .A(_919_[5]),
    .Y(ACC_o[5])
);

NAND2X1 _1475_ (
    .A(_283_),
    .B(_563_),
    .Y(_564_)
);

AOI21X1 _1055_ (
    .A(_138_),
    .B(_140_),
    .C(_129_),
    .Y(_147_)
);

FILL FILL_0__1515_ (
);

NAND2X1 _1284_ (
    .A(_332_),
    .B(_336_),
    .Y(_375_)
);

FILL FILL_0__1744_ (
);

FILL FILL_0__1324_ (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

FILL FILL_1_BUFX2_insert12 (
);

FILL FILL_1_BUFX2_insert13 (
);

FILL FILL_1_BUFX2_insert14 (
);

OAI21X1 _1093_ (
    .A(_180_),
    .B(_179_),
    .C(_184_),
    .Y(_185_)
);

FILL FILL_0__1553_ (
);

FILL FILL_0__1133_ (
);

FILL FILL_1__1714_ (
);

OAI21X1 _1569_ (
    .A(_280_),
    .B(_356_),
    .C(MulL_i),
    .Y(_655_)
);

NAND2X1 _1149_ (
    .A(BI[2]),
    .B(_68_),
    .Y(_241_)
);

FILL FILL_0__1609_ (
);

FILL FILL_0__1782_ (
);

FILL FILL_0__1362_ (
);

FILL FILL_1__1523_ (
);

FILL FILL_1__1103_ (
);

INVX1 _1798_ (
    .A(_767_),
    .Y(_772_)
);

AOI21X1 _1378_ (
    .A(_397_),
    .B(_402_),
    .C(_462_),
    .Y(_468_)
);

FILL FILL_0__1838_ (
);

FILL FILL_0__1418_ (
);

FILL FILL_0__1591_ (
);

FILL FILL_0__1171_ (
);

AND2X2 _921_ (
    .A(MUL_bF$buf3),
    .B(BI[4]),
    .Y(_713_)
);

FILL FILL_1__1752_ (
);

FILL FILL_1__1332_ (
);

NAND3X1 _1187_ (
    .A(_251_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

FILL FILL_1__969_ (
);

FILL FILL_0__1647_ (
);

FILL FILL_0__1227_ (
);

FILL FILL_1__1808_ (
);

FILL FILL_1__1561_ (
);

FILL FILL_1__1141_ (
);

FILL FILL_0__1876_ (
);

FILL FILL_0__1456_ (
);

FILL FILL_0__1036_ (
);

FILL FILL_1__1617_ (
);

FILL FILL_1__1790_ (
);

FILL FILL_1__1370_ (
);

FILL FILL_0__1685_ (
);

FILL FILL_0__1265_ (
);

FILL FILL86550x7350 (
);

FILL FILL_1__1846_ (
);

FILL FILL_1__1426_ (
);

FILL FILL_1__1006_ (
);

FILL FILL_0__1494_ (
);

FILL FILL_0__1074_ (
);

FILL FILL_1__1235_ (
);

AOI21X1 _1722_ (
    .A(alu_op_2_bF$buf0),
    .B(BI[1]),
    .C(_892_),
    .Y(_893_)
);

AND2X2 _1302_ (
    .A(_388_),
    .B(_391_),
    .Y(_393_)
);

FILL FILL_1__1884_ (
);

FILL FILL_1__1464_ (
);

FILL FILL_1__1044_ (
);

FILL FILL_2__1533_ (
);

FILL FILL_0__1779_ (
);

FILL FILL_0__1359_ (
);

NAND3X1 _1531_ (
    .A(MulL_i),
    .B(_618_),
    .C(_617_),
    .Y(_619_)
);

NAND2X1 _1111_ (
    .A(_202_),
    .B(_199_),
    .Y(_203_)
);

FILL FILL_1__1693_ (
);

FILL FILL_1__1273_ (
);

FILL FILL_0__1588_ (
);

FILL FILL_0__1168_ (
);

FILL FILL_1__1749_ (
);

FILL FILL_1__1329_ (
);

INVX1 _1760_ (
    .A(_732_),
    .Y(_736_)
);

AOI21X1 _1340_ (
    .A(_322_),
    .B(_326_),
    .C(_328_),
    .Y(_431_)
);

FILL FILL_1__1082_ (
);

FILL FILL_0__1800_ (
);

FILL FILL_0__1397_ (
);

NAND2X1 _1816_ (
    .A(_786_),
    .B(_788_),
    .Y(_789_)
);

FILL FILL_1__1558_ (
);

FILL FILL_1__1138_ (
);

FILL FILL_1__931_ (
);

FILL FILL_2__1207_ (
);

OAI21X1 _1625_ (
    .A(LoadA_i),
    .B(_725_),
    .C(_697_),
    .Y(_12_)
);

NOR2X1 _1205_ (
    .A(_292_),
    .B(_293_),
    .Y(_297_)
);

FILL FILL_0__953_ (
);

OAI21X1 _956_ (
    .A(_46_),
    .B(_47_),
    .C(_42_),
    .Y(_48_)
);

FILL FILL_1__1787_ (
);

FILL FILL_1__1367_ (
);

OAI21X1 _1854_ (
    .A(_806_),
    .B(_823_),
    .C(_789_),
    .Y(_824_)
);

OAI21X1 _1434_ (
    .A(_712_),
    .B(_516_),
    .C(_523_),
    .Y(_0_[2])
);

NAND3X1 _1014_ (
    .A(_104_),
    .B(_105_),
    .C(_103_),
    .Y(_106_)
);

FILL FILL_1__1596_ (
);

FILL FILL_1__1176_ (
);

DFFSR _1663_ (
    .R(_1_),
    .S(vdd),
    .D(_0_[2]),
    .CLK(clk_bF$buf4),
    .Q(_919_[2])
);

OAI21X1 _1243_ (
    .A(_329_),
    .B(_330_),
    .C(_301_),
    .Y(_335_)
);

FILL FILL_0__991_ (
);

OAI21X1 _994_ (
    .A(_81_),
    .B(_82_),
    .C(_85_),
    .Y(_86_)
);

FILL FILL_0__1703_ (
);

FILL FILL_2__1474_ (
);

OAI21X1 _1719_ (
    .A(AI[1]),
    .B(_889_),
    .C(_868_),
    .Y(_890_)
);

BUFX2 _1892_ (
    .A(_919_[2]),
    .Y(ACC_o[2])
);

NAND3X1 _1472_ (
    .A(_511_),
    .B(_560_),
    .C(_514_),
    .Y(_561_)
);

NAND2X1 _1052_ (
    .A(_89_),
    .B(_143_),
    .Y(_144_)
);

FILL FILL_0__1512_ (
);

NAND2X1 _1528_ (
    .A(_615_),
    .B(_610_),
    .Y(_616_)
);

NAND2X1 _1108_ (
    .A(_197_),
    .B(_194_),
    .Y(_200_)
);

MUX2X1 _1281_ (
    .A(AN),
    .B(ACC[1]),
    .S(Flag_i),
    .Y(_372_)
);

FILL FILL_0__1741_ (
);

FILL FILL_0__1321_ (
);

NAND3X1 _1757_ (
    .A(_906_),
    .B(_733_),
    .C(_897_),
    .Y(_734_)
);

NAND2X1 _1337_ (
    .A(_414_),
    .B(_427_),
    .Y(_428_)
);

FILL FILL_1__1499_ (
);

FILL FILL_1__1079_ (
);

NAND2X1 _1090_ (
    .A(MUL_bF$buf0),
    .B(BI[5]),
    .Y(_182_)
);

FILL FILL_0__1550_ (
);

FILL FILL_0__1130_ (
);

FILL FILL_2__1148_ (
);

FILL FILL_1__1711_ (
);

NAND2X1 _1566_ (
    .A(_629_),
    .B(_652_),
    .Y(_0_[5])
);

NAND3X1 _1146_ (
    .A(MUL_bF$buf0),
    .B(BI[1]),
    .C(AI[1]),
    .Y(_238_)
);

FILL FILL_1__928_ (
);

FILL FILL_0__1606_ (
);

FILL FILL_1__1520_ (
);

FILL FILL_1__1100_ (
);

OAI21X1 _1795_ (
    .A(_769_),
    .B(_737_),
    .C(_909_),
    .Y(_770_)
);

NAND2X1 _1375_ (
    .A(BI[6]),
    .B(_464_),
    .Y(_465_)
);

FILL FILL_0__1835_ (
);

FILL FILL_0__1415_ (
);

NOR3X1 _1184_ (
    .A(_275_),
    .B(_274_),
    .C(_252_),
    .Y(_276_)
);

FILL FILL_1__966_ (
);

FILL FILL86850x50550 (
);

FILL FILL_0__1644_ (
);

FILL FILL_0__1224_ (
);

FILL FILL_1__1805_ (
);

FILL FILL_0__988_ (
);

FILL FILL_0__1873_ (
);

FILL FILL_0__1453_ (
);

FILL FILL_0__1033_ (
);

FILL FILL_1__1614_ (
);

AND2X2 _1889_ (
    .A(_854_),
    .B(_856_),
    .Y(AV)
);

OAI21X1 _1469_ (
    .A(_458_),
    .B(_557_),
    .C(_504_),
    .Y(_558_)
);

NAND3X1 _1049_ (
    .A(_120_),
    .B(_124_),
    .C(_90_),
    .Y(_141_)
);

FILL FILL_0__1509_ (
);

FILL FILL_0__1262_ (
);

FILL FILL_1__1843_ (
);

FILL FILL_1__1423_ (
);

FILL FILL_1__1003_ (
);

INVX1 _1698_ (
    .A(AI[0]),
    .Y(_870_)
);

OAI21X1 _1278_ (
    .A(_712_),
    .B(_362_),
    .C(_369_),
    .Y(_0_[0])
);

FILL FILL_0__1738_ (
);

FILL FILL_0__1318_ (
);

FILL FILL_0__1491_ (
);

FILL FILL_2__1089_ (
);

FILL FILL_0__1071_ (
);

FILL FILL_1__1652_ (
);

FILL FILL_1__1232_ (
);

AOI21X1 _1087_ (
    .A(_163_),
    .B(_164_),
    .C(_162_),
    .Y(_179_)
);

FILL FILL85650x82950 (
);

FILL FILL_0__1547_ (
);

FILL FILL_0__1127_ (
);

FILL FILL_1__1708_ (
);

FILL FILL_1__1881_ (
);

FILL FILL_1__1461_ (
);

FILL FILL_1__1041_ (
);

FILL FILL_0__1776_ (
);

FILL FILL_0__1356_ (
);

FILL FILL_1__1517_ (
);

FILL FILL_1__1690_ (
);

FILL FILL_1__1270_ (
);

FILL FILL_0__1585_ (
);

FILL FILL_0__1165_ (
);

FILL FILL_1__1746_ (
);

FILL FILL_1__1326_ (
);

FILL FILL_0__1394_ (
);

OAI21X1 _1813_ (
    .A(_774_),
    .B(_768_),
    .C(_785_),
    .Y(_786_)
);

FILL FILL_1__1555_ (
);

FILL FILL_1__1135_ (
);

FILL FILL_2__979_ (
);

NAND2X1 _1622_ (
    .A(ABCmd_i[1]),
    .B(LoadA_i),
    .Y(_696_)
);

OR2X2 _1202_ (
    .A(_293_),
    .B(_292_),
    .Y(_294_)
);

FILL FILL_0__950_ (
);

OAI21X1 _953_ (
    .A(_43_),
    .B(_44_),
    .C(_718_),
    .Y(_45_)
);

FILL FILL_1__1784_ (
);

FILL FILL_1__1364_ (
);

FILL FILL_0__1259_ (
);

NAND2X1 _1851_ (
    .A(_751_),
    .B(_820_),
    .Y(_821_)
);

OAI21X1 _1431_ (
    .A(AZ),
    .B(_364_),
    .C(_365_),
    .Y(_521_)
);

OAI21X1 _1011_ (
    .A(_56_),
    .B(_60_),
    .C(_52_),
    .Y(_103_)
);

FILL FILL_1__1593_ (
);

FILL FILL_1__1173_ (
);

FILL FILL_0__1488_ (
);

FILL FILL_0__1068_ (
);

FILL FILL_1__1649_ (
);

FILL FILL_1__1229_ (
);

DFFPOSX1 _1660_ (
    .D(_9_),
    .CLK(clk_bF$buf1),
    .Q(MUL)
);

NAND3X1 _1240_ (
    .A(_300_),
    .B(_331_),
    .C(_327_),
    .Y(_332_)
);

NAND3X1 _991_ (
    .A(_74_),
    .B(_77_),
    .C(_70_),
    .Y(_83_)
);

FILL FILL_0__1700_ (
);

FILL FILL_0__1297_ (
);

AOI22X1 _1716_ (
    .A(_862_),
    .B(BI[1]),
    .C(_886_),
    .D(_863_),
    .Y(_887_)
);

FILL FILL_1__1878_ (
);

FILL FILL_1__1458_ (
);

FILL FILL_1__1038_ (
);

FILL FILL_2__1527_ (
);

AOI22X1 _1525_ (
    .A(_556_),
    .B(_607_),
    .C(_612_),
    .D(_611_),
    .Y(_613_)
);

INVX1 _1105_ (
    .A(_196_),
    .Y(_197_)
);

FILL FILL_1__1687_ (
);

FILL FILL_1__1267_ (
);

NAND2X1 _1754_ (
    .A(_730_),
    .B(_911_),
    .Y(_731_)
);

AND2X2 _1334_ (
    .A(_409_),
    .B(_413_),
    .Y(_425_)
);

FILL FILL_1__1496_ (
);

FILL FILL_1__1076_ (
);

AND2X2 _1563_ (
    .A(_645_),
    .B(_644_),
    .Y(_650_)
);

NAND3X1 _1143_ (
    .A(_221_),
    .B(_27_),
    .C(_723_),
    .Y(_235_)
);

FILL FILL_1__925_ (
);

FILL FILL_0__1603_ (
);

FILL FILL_2__1794_ (
);

OAI21X1 _1619_ (
    .A(LoadCmd_i),
    .B(_715_),
    .C(_694_),
    .Y(_9_)
);

FILL FILL_0__947_ (
);

OAI21X1 _1792_ (
    .A(_763_),
    .B(_765_),
    .C(_766_),
    .Y(_767_)
);

NOR2X1 _1372_ (
    .A(_398_),
    .B(_399_),
    .Y(_462_)
);

FILL FILL_0__1832_ (
);

FILL FILL_0__1412_ (
);

NAND3X1 _1848_ (
    .A(_799_),
    .B(_816_),
    .C(_802_),
    .Y(_819_)
);

NOR2X1 _1428_ (
    .A(_365_),
    .B(_271_),
    .Y(_518_)
);

OAI21X1 _1008_ (
    .A(_36_),
    .B(_54_),
    .C(_93_),
    .Y(_100_)
);

OAI21X1 _1181_ (
    .A(_248_),
    .B(_272_),
    .C(_247_),
    .Y(_273_)
);

FILL FILL_1__963_ (
);

FILL FILL_0__1641_ (
);

FILL FILL_2__1239_ (
);

FILL FILL_0__1221_ (
);

FILL FILL_1__1802_ (
);

DFFPOSX1 _1657_ (
    .D(_6_),
    .CLK(clk_bF$buf3),
    .Q(CI)
);

AOI22X1 _1237_ (
    .A(_306_),
    .B(_311_),
    .C(_324_),
    .D(_325_),
    .Y(_329_)
);

FILL FILL_0__985_ (
);

NAND3X1 _988_ (
    .A(_66_),
    .B(_62_),
    .C(_79_),
    .Y(_80_)
);

FILL FILL_1__1399_ (
);

FILL FILL_0__1870_ (
);

FILL FILL_2__1468_ (
);

FILL FILL_0__1450_ (
);

FILL FILL_0__1030_ (
);

FILL FILL_1__1611_ (
);

NAND3X1 _1886_ (
    .A(_852_),
    .B(_853_),
    .C(_841_),
    .Y(_854_)
);

NAND2X1 _1466_ (
    .A(_554_),
    .B(_550_),
    .Y(_555_)
);

INVX1 _1046_ (
    .A(_137_),
    .Y(_138_)
);

FILL FILL_0__1506_ (
);

FILL FILL_1__1840_ (
);

FILL FILL_1__1420_ (
);

FILL FILL_1__1000_ (
);

AOI22X1 _1695_ (
    .A(BI[0]),
    .B(_866_),
    .C(_863_),
    .D(_865_),
    .Y(_867_)
);

NAND3X1 _1275_ (
    .A(BI[0]),
    .B(MulL_i),
    .C(_68_),
    .Y(_367_)
);

FILL FILL_0__1735_ (
);

FILL FILL_0__1315_ (
);

NAND3X1 _1084_ (
    .A(_166_),
    .B(_171_),
    .C(_175_),
    .Y(_176_)
);

FILL FILL_0__1544_ (
);

FILL FILL_0__1124_ (
);

FILL FILL_1__1705_ (
);

FILL FILL_0__1773_ (
);

FILL FILL_0__1353_ (
);

FILL FILL_1__1514_ (
);

OAI21X1 _1789_ (
    .A(alu_op_2_bF$buf3),
    .B(BI[4]),
    .C(_858_),
    .Y(_764_)
);

AOI21X1 _1369_ (
    .A(_423_),
    .B(_428_),
    .C(_415_),
    .Y(_459_)
);

FILL FILL_0__1829_ (
);

FILL FILL_0__1409_ (
);

FILL FILL_0__1582_ (
);

FILL FILL_0__1162_ (
);

FILL FILL_1__1743_ (
);

FILL FILL_1__1323_ (
);

NAND2X1 _1598_ (
    .A(ABCmd_i[0]),
    .B(LoadCmd_i),
    .Y(_681_)
);

NAND3X1 _1178_ (
    .A(_267_),
    .B(_269_),
    .C(_264_),
    .Y(_270_)
);

FILL FILL_0__1638_ (
);

FILL FILL_0__1218_ (
);

FILL FILL_0__1391_ (
);

OAI21X1 _1810_ (
    .A(_877_),
    .B(_782_),
    .C(_780_),
    .Y(_783_)
);

FILL FILL_1__1552_ (
);

FILL FILL_1__1132_ (
);

FILL FILL_0__1867_ (
);

FILL FILL_0__1447_ (
);

FILL FILL_0__1027_ (
);

FILL FILL_1__1608_ (
);

NAND3X1 _950_ (
    .A(_41_),
    .B(_29_),
    .C(_39_),
    .Y(_42_)
);

FILL FILL_1__1781_ (
);

FILL FILL_1__1361_ (
);

FILL FILL_1__998_ (
);

FILL FILL_0__1256_ (
);

FILL FILL_1__1837_ (
);

FILL FILL_1__1417_ (
);

FILL FILL_1__1590_ (
);

FILL FILL_1__1170_ (
);

FILL FILL_0__1485_ (
);

FILL FILL_0__1065_ (
);

FILL FILL_1__1646_ (
);

FILL FILL_1__1226_ (
);

FILL FILL_2__1715_ (
);

FILL FILL_0__1294_ (
);

OAI21X1 _1713_ (
    .A(_861_),
    .B(_883_),
    .C(_878_),
    .Y(_884_)
);

FILL FILL_1__1875_ (
);

FILL FILL_1__1455_ (
);

FILL FILL_1__1035_ (
);

NAND3X1 _1522_ (
    .A(_604_),
    .B(_606_),
    .C(_609_),
    .Y(_610_)
);

INVX1 _1102_ (
    .A(_193_),
    .Y(_194_)
);

FILL FILL_1__1264_ (
);

FILL FILL_0__1579_ (
);

FILL FILL_0__1159_ (
);

INVX1 _1751_ (
    .A(_727_),
    .Y(_728_)
);

OAI21X1 _1331_ (
    .A(_415_),
    .B(_421_),
    .C(_395_),
    .Y(_422_)
);

FILL FILL_1__1493_ (
);

FILL FILL_1__1073_ (
);

FILL FILL_0__1388_ (
);

OAI21X1 _1807_ (
    .A(_779_),
    .B(_778_),
    .C(_775_),
    .Y(_780_)
);

FILL FILL_1__1549_ (
);

FILL FILL_1__1129_ (
);

NAND3X1 _1560_ (
    .A(_602_),
    .B(_646_),
    .C(_610_),
    .Y(_647_)
);

NAND3X1 _1140_ (
    .A(_231_),
    .B(_230_),
    .C(_229_),
    .Y(_232_)
);

FILL FILL_1__922_ (
);

FILL FILL_2__1618_ (
);

FILL FILL_0__1600_ (
);

FILL FILL_0__1197_ (
);

NAND2X1 _1616_ (
    .A(LoadCmd_i),
    .B(ABCmd_i[6]),
    .Y(_693_)
);

FILL FILL_0__944_ (
);

NAND3X1 _947_ (
    .A(_31_),
    .B(_38_),
    .C(_35_),
    .Y(_39_)
);

FILL FILL_1__1778_ (
);

FILL FILL_1__1358_ (
);

FILL FILL_2__1180_ (
);

OAI21X1 _1845_ (
    .A(_812_),
    .B(_814_),
    .C(_815_),
    .Y(_816_)
);

OR2X2 _1425_ (
    .A(_456_),
    .B(_513_),
    .Y(_515_)
);

INVX1 _1005_ (
    .A(_96_),
    .Y(_97_)
);

FILL FILL_1__1587_ (
);

FILL FILL_1__1167_ (
);

FILL FILL_1__960_ (
);

DFFPOSX1 _1654_ (
    .D(_3_),
    .CLK(clk_bF$buf2),
    .Q(alu_op[1])
);

NAND3X1 _1234_ (
    .A(_324_),
    .B(_325_),
    .C(_323_),
    .Y(_326_)
);

FILL FILL_0__982_ (
);

INVX1 _985_ (
    .A(_73_),
    .Y(_77_)
);

FILL FILL_1__1396_ (
);

FILL FILL_2__1885_ (
);

INVX1 _1883_ (
    .A(_850_),
    .Y(_851_)
);

NAND3X1 _1463_ (
    .A(_543_),
    .B(_546_),
    .C(_551_),
    .Y(_552_)
);

INVX4 _1043_ (
    .A(_134_),
    .Y(_135_)
);

FILL FILL_0__1503_ (
);

OAI21X1 _1519_ (
    .A(_525_),
    .B(_555_),
    .C(_511_),
    .Y(_607_)
);

INVX2 _1692_ (
    .A(alu_op[0]),
    .Y(_864_)
);

INVX1 _1272_ (
    .A(Flag_i),
    .Y(_364_)
);

FILL FILL_0__1732_ (
);

FILL FILL_0__1312_ (
);

OAI21X1 _1748_ (
    .A(_917_),
    .B(_916_),
    .C(_912_),
    .Y(_918_)
);

AOI21X1 _1328_ (
    .A(_416_),
    .B(_418_),
    .C(_320_),
    .Y(_419_)
);

NAND2X1 _1081_ (
    .A(_167_),
    .B(_172_),
    .Y(_173_)
);

FILL FILL_2__1559_ (
);

FILL FILL_0__1541_ (
);

FILL FILL_0__1121_ (
);

FILL FILL_1__1702_ (
);

NAND2X1 _1557_ (
    .A(_630_),
    .B(_643_),
    .Y(_644_)
);

AOI21X1 _1137_ (
    .A(_227_),
    .B(_228_),
    .C(_225_),
    .Y(_229_)
);

FILL FILL_1__1299_ (
);

FILL FILL_0__1770_ (
);

FILL FILL_0__1350_ (
);

FILL FILL_1__1511_ (
);

AOI22X1 _1786_ (
    .A(_862_),
    .B(BI[4]),
    .C(_760_),
    .D(_863_),
    .Y(_761_)
);

OAI21X1 _1366_ (
    .A(_453_),
    .B(_359_),
    .C(_455_),
    .Y(_456_)
);

FILL FILL_0__1826_ (
);

FILL FILL_0__1406_ (
);

FILL FILL_1__1740_ (
);

FILL FILL_1__1320_ (
);

AOI22X1 _1595_ (
    .A(_678_),
    .B(_679_),
    .C(_668_),
    .D(_675_),
    .Y(_0_[7])
);

NOR2X1 _1175_ (
    .A(_265_),
    .B(_266_),
    .Y(_267_)
);

FILL FILL_1__957_ (
);

FILL FILL_0__1635_ (
);

FILL FILL_0__1215_ (
);

FILL FILL_0__979_ (
);

FILL FILL_0__1864_ (
);

FILL FILL_0__1444_ (
);

FILL FILL_0__1024_ (
);

FILL FILL86550x36150 (
);

FILL FILL_1__1605_ (
);

FILL FILL_1__995_ (
);

FILL FILL_0__1253_ (
);

FILL FILL_1__1834_ (
);

FILL FILL_1__1414_ (
);

INVX1 _1689_ (
    .A(_860_),
    .Y(_861_)
);

NAND2X1 _1269_ (
    .A(_360_),
    .B(_359_),
    .Y(_361_)
);

FILL FILL_0__1729_ (
);

FILL FILL_0__1309_ (
);

FILL FILL_0__1482_ (
);

FILL FILL_0__1062_ (
);

FILL FILL_1__1643_ (
);

FILL FILL_1__1223_ (
);

OAI21X1 _1498_ (
    .A(_288_),
    .B(_54_),
    .C(_584_),
    .Y(_586_)
);

NAND3X1 _1078_ (
    .A(MUL_bF$buf2),
    .B(BI[3]),
    .C(AI[4]),
    .Y(_170_)
);

FILL FILL_0__1538_ (
);

FILL FILL_0__1118_ (
);

FILL FILL86850x79350 (
);

FILL FILL_0__1291_ (
);

NAND2X1 _1710_ (
    .A(_881_),
    .B(_880_),
    .Y(_882_)
);

FILL FILL_1__1872_ (
);

FILL FILL_1__1452_ (
);

FILL FILL_1__1032_ (
);

FILL FILL_0__1767_ (
);

FILL FILL_0__1347_ (
);

FILL FILL_1__1508_ (
);

FILL FILL_1__1261_ (
);

FILL FILL_0__1576_ (
);

FILL FILL_0__1156_ (
);

FILL FILL_1__1737_ (
);

FILL FILL_1__1317_ (
);

FILL FILL_1__1490_ (
);

FILL FILL_1__1070_ (
);

FILL FILL_0__1385_ (
);

NAND2X1 _1804_ (
    .A(AI[5]),
    .B(_776_),
    .Y(_777_)
);

FILL FILL_1__1546_ (
);

FILL FILL_1__1126_ (
);

FILL FILL_0__1194_ (
);

NAND2X1 _1613_ (
    .A(LoadCmd_i),
    .B(ABCmd_i[5]),
    .Y(_691_)
);

FILL FILL_0__941_ (
);

INVX1 _944_ (
    .A(BI[1]),
    .Y(_36_)
);

FILL FILL_1__1775_ (
);

FILL FILL_1__1355_ (
);

FILL FILL_2__1004_ (
);

OAI21X1 _1842_ (
    .A(alu_op_2_bF$buf2),
    .B(BI[7]),
    .C(_858_),
    .Y(_813_)
);

NAND2X1 _1422_ (
    .A(_511_),
    .B(_508_),
    .Y(_512_)
);

NOR2X1 _1002_ (
    .A(_92_),
    .B(_93_),
    .Y(_94_)
);

FILL FILL_1__1584_ (
);

FILL FILL_1__1164_ (
);

FILL FILL_2__1233_ (
);

FILL FILL_0__1479_ (
);

FILL FILL_0__1059_ (
);

FILL FILL86250x82950 (
);

NAND2X1 _1651_ (
    .A(ABCmd_i[7]),
    .B(LoadB_i),
    .Y(_711_)
);

AND2X2 _1231_ (
    .A(_311_),
    .B(_306_),
    .Y(_323_)
);

OAI21X1 _982_ (
    .A(_716_),
    .B(_44_),
    .C(_72_),
    .Y(_74_)
);

FILL FILL_1__1393_ (
);

FILL FILL_2__1709_ (
);

FILL FILL_0__1288_ (
);

OAI21X1 _1707_ (
    .A(_874_),
    .B(_876_),
    .C(_878_),
    .Y(_879_)
);

FILL FILL85950x64950 (
);

FILL FILL_1__1869_ (
);

FILL FILL_1__1449_ (
);

FILL FILL_1__1029_ (
);

NAND2X1 _1880_ (
    .A(\u_ALU8.AI7 ),
    .B(_847_),
    .Y(_848_)
);

OAI21X1 _1460_ (
    .A(_487_),
    .B(_501_),
    .C(_548_),
    .Y(_549_)
);

OR2X2 _1040_ (
    .A(_131_),
    .B(_130_),
    .Y(_132_)
);

FILL FILL_0__1500_ (
);

FILL FILL_0__1097_ (
);

INVX1 _1516_ (
    .A(_603_),
    .Y(_604_)
);

FILL FILL_1__1258_ (
);

NAND2X1 _1745_ (
    .A(AI[2]),
    .B(_914_),
    .Y(_915_)
);

OR2X2 _1325_ (
    .A(_314_),
    .B(_315_),
    .Y(_416_)
);

FILL FILL_1__1487_ (
);

FILL FILL_1__1067_ (
);

INVX1 _1554_ (
    .A(_633_),
    .Y(_641_)
);

AND2X2 _1134_ (
    .A(_718_),
    .B(_714_),
    .Y(_226_)
);

FILL FILL_1__1296_ (
);

FILL FILL_0__938_ (
);

NAND2X1 _1783_ (
    .A(shr),
    .B(AI[5]),
    .Y(_758_)
);

NAND2X1 _1363_ (
    .A(_352_),
    .B(_451_),
    .Y(_453_)
);

FILL FILL_0__1823_ (
);

FILL FILL_0__1403_ (
);

FILL FILL_2__1174_ (
);

AOI22X1 _1839_ (
    .A(_862_),
    .B(BI[7]),
    .C(_809_),
    .D(_863_),
    .Y(_810_)
);

AOI21X1 _1419_ (
    .A(_422_),
    .B(_429_),
    .C(_432_),
    .Y(_509_)
);

AOI21X1 _1592_ (
    .A(_676_),
    .B(_358_),
    .C(_365_),
    .Y(_677_)
);

OR2X2 _1172_ (
    .A(_263_),
    .B(_241_),
    .Y(_264_)
);

FILL FILL_1__954_ (
);

FILL FILL_0__1632_ (
);

FILL FILL_0__1212_ (
);

OAI21X1 _1648_ (
    .A(LoadB_i),
    .B(_708_),
    .C(_709_),
    .Y(_23_)
);

OAI21X1 _1228_ (
    .A(_153_),
    .B(_154_),
    .C(_157_),
    .Y(_320_)
);

FILL FILL_0__976_ (
);

NAND3X1 _979_ (
    .A(MUL_bF$buf4),
    .B(BI[4]),
    .C(AI[1]),
    .Y(_71_)
);

FILL FILL_2__1879_ (
);

FILL FILL_0__1861_ (
);

FILL FILL_0__1441_ (
);

FILL FILL_0__1021_ (
);

FILL FILL_1__1602_ (
);

INVX1 _1877_ (
    .A(_814_),
    .Y(_845_)
);

NAND3X1 _1457_ (
    .A(_535_),
    .B(_545_),
    .C(_544_),
    .Y(_546_)
);

AOI21X1 _1037_ (
    .A(_127_),
    .B(_128_),
    .C(_126_),
    .Y(_129_)
);

FILL FILL_1__1199_ (
);

FILL FILL_1__992_ (
);

FILL FILL_0__1250_ (
);

FILL FILL_1__1831_ (
);

FILL FILL_1__1411_ (
);

INVX4 _1686_ (
    .A(alu_op[3]),
    .Y(_858_)
);

OAI21X1 _1266_ (
    .A(_280_),
    .B(_356_),
    .C(_357_),
    .Y(_358_)
);

FILL FILL_0__1726_ (
);

FILL FILL_0__1306_ (
);

FILL FILL_1__1640_ (
);

FILL FILL_1__1220_ (
);

FILL FILL85950x7350 (
);

OAI21X1 _1495_ (
    .A(_538_),
    .B(_539_),
    .C(_582_),
    .Y(_583_)
);

INVX1 _1075_ (
    .A(_166_),
    .Y(_167_)
);

FILL FILL_0__1535_ (
);

FILL FILL_0__1115_ (
);

FILL FILL_0__1764_ (
);

FILL FILL_0__1344_ (
);

FILL FILL86850x10950 (
);

FILL FILL_1__1505_ (
);

FILL FILL_0__1573_ (
);

FILL FILL_0__1153_ (
);

FILL FILL_1__1734_ (
);

FILL FILL_1__1314_ (
);

OAI21X1 _1589_ (
    .A(_582_),
    .B(_634_),
    .C(_665_),
    .Y(_674_)
);

INVX1 _1169_ (
    .A(_248_),
    .Y(_261_)
);

FILL FILL_0__1629_ (
);

FILL FILL_0__1209_ (
);

FILL FILL_0__1382_ (
);

INVX1 _1801_ (
    .A(_766_),
    .Y(_774_)
);

FILL FILL_1__1543_ (
);

FILL FILL_1__1123_ (
);

NAND3X1 _1398_ (
    .A(_416_),
    .B(_486_),
    .C(_413_),
    .Y(_488_)
);

FILL FILL_0__1858_ (
);

FILL FILL_0__1438_ (
);

FILL FILL_0__1018_ (
);

FILL FILL_0__1191_ (
);

NAND2X1 _1610_ (
    .A(LoadCmd_i),
    .B(ABCmd_i[4]),
    .Y(_689_)
);

NAND3X1 _941_ (
    .A(MUL_bF$buf4),
    .B(BI[1]),
    .C(AI[3]),
    .Y(_33_)
);

FILL FILL_1__1772_ (
);

FILL FILL_1__1352_ (
);

FILL FILL_1__989_ (
);

FILL FILL_0__1247_ (
);

FILL FILL_1__1828_ (
);

FILL FILL_1__1408_ (
);

FILL FILL_1__1581_ (
);

FILL FILL_1__1161_ (
);

FILL FILL_0__1896_ (
);

FILL FILL_0__1476_ (
);

FILL FILL_0__1056_ (
);

FILL FILL_1__1637_ (
);

FILL FILL_1__1217_ (
);

FILL FILL_1__1390_ (
);

FILL FILL_0_BUFX2_insert5 (
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_0__1285_ (
);

AOI21X1 _1704_ (
    .A(BI[0]),
    .B(alu_op_2_bF$buf1),
    .C(_875_),
    .Y(_876_)
);

FILL FILL_1__1866_ (
);

FILL FILL_1__1446_ (
);

FILL FILL_1__1026_ (
);

FILL FILL_0__1094_ (
);

NAND2X1 _1513_ (
    .A(_577_),
    .B(_600_),
    .Y(_601_)
);

FILL FILL_1__1255_ (
);

FILL FILL_2__1324_ (
);

NAND2X1 _1742_ (
    .A(shr),
    .B(AI[3]),
    .Y(_912_)
);

NAND3X1 _1322_ (
    .A(_410_),
    .B(_412_),
    .C(_411_),
    .Y(_413_)
);

FILL FILL_1__1484_ (
);

FILL FILL_1__1064_ (
);

FILL FILL_2__1553_ (
);

FILL FILL_0__1799_ (
);

FILL FILL_0__1379_ (
);

OAI21X1 _1551_ (
    .A(_590_),
    .B(_587_),
    .C(_636_),
    .Y(_638_)
);

OAI21X1 _1131_ (
    .A(_34_),
    .B(_40_),
    .C(_31_),
    .Y(_223_)
);

FILL FILL_1__1293_ (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_0__1188_ (
);

NAND2X1 _1607_ (
    .A(LoadCmd_i),
    .B(ABCmd_i[3]),
    .Y(_687_)
);

FILL FILL_0__935_ (
);

NAND3X1 _938_ (
    .A(MUL_bF$buf4),
    .B(BI[2]),
    .C(AI[2]),
    .Y(_30_)
);

FILL FILL_1__1769_ (
);

FILL FILL_1__1349_ (
);

NAND2X1 _1780_ (
    .A(_732_),
    .B(_731_),
    .Y(_755_)
);

AND2X2 _1360_ (
    .A(_442_),
    .B(_447_),
    .Y(_451_)
);

FILL FILL_0__1820_ (
);

FILL FILL_0__1400_ (
);

NAND2X1 _1836_ (
    .A(shr),
    .B(CI),
    .Y(_807_)
);

NAND3X1 _1416_ (
    .A(_457_),
    .B(_504_),
    .C(_505_),
    .Y(_506_)
);

FILL FILL_1__1578_ (
);

FILL FILL_1__1158_ (
);

FILL FILL_1__951_ (
);

FILL FILL85950x50550 (
);

OAI21X1 _1645_ (
    .A(LoadB_i),
    .B(_169_),
    .C(_707_),
    .Y(_22_)
);

AND2X2 _1225_ (
    .A(_314_),
    .B(_315_),
    .Y(_317_)
);

FILL FILL_0__973_ (
);

INVX2 _976_ (
    .A(_67_),
    .Y(_68_)
);

FILL FILL_1__1387_ (
);

AOI21X1 _1874_ (
    .A(_790_),
    .B(_801_),
    .C(_805_),
    .Y(_842_)
);

OAI21X1 _1454_ (
    .A(_537_),
    .B(_536_),
    .C(_542_),
    .Y(_543_)
);

AOI21X1 _1034_ (
    .A(_79_),
    .B(_66_),
    .C(_81_),
    .Y(_126_)
);

FILL FILL_1__1196_ (
);

FILL FILL_2__1265_ (
);

DFFPOSX1 _1683_ (
    .D(_24_),
    .CLK(clk_bF$buf1),
    .Q(BI[6])
);

INVX1 _1263_ (
    .A(_219_),
    .Y(_355_)
);

FILL FILL_0__1723_ (
);

FILL FILL_0__1303_ (
);

FILL FILL_2__1494_ (
);

INVX1 _1739_ (
    .A(_909_),
    .Y(ACC[1])
);

NAND3X1 _1319_ (
    .A(_396_),
    .B(_404_),
    .C(_406_),
    .Y(_410_)
);

INVX1 _1492_ (
    .A(_579_),
    .Y(_580_)
);

OAI21X1 _1072_ (
    .A(_152_),
    .B(_153_),
    .C(_154_),
    .Y(_164_)
);

FILL FILL_0__1532_ (
);

FILL FILL_0__1112_ (
);

OAI22X1 _1548_ (
    .A(_288_),
    .B(_158_),
    .C(_417_),
    .D(_135_),
    .Y(_635_)
);

NOR2X1 _1128_ (
    .A(_714_),
    .B(_718_),
    .Y(_220_)
);

FILL FILL_0__1761_ (
);

FILL FILL_0__1341_ (
);

FILL FILL_1__1502_ (
);

INVX1 _1777_ (
    .A(BCD),
    .Y(_752_)
);

NAND2X1 _1357_ (
    .A(_447_),
    .B(_442_),
    .Y(_448_)
);

FILL FILL_1__1099_ (
);

FILL FILL_0__1817_ (
);

FILL FILL_0__1570_ (
);

FILL FILL_0__1150_ (
);

FILL FILL_1__1731_ (
);

FILL FILL_1__1311_ (
);

NAND3X1 _1586_ (
    .A(_671_),
    .B(_666_),
    .C(_670_),
    .Y(_672_)
);

NAND3X1 _1166_ (
    .A(_139_),
    .B(_142_),
    .C(_257_),
    .Y(_258_)
);

FILL FILL_1__948_ (
);

FILL FILL_2__1800_ (
);

FILL FILL_0__1626_ (
);

FILL FILL_0__1206_ (
);

FILL FILL86550x43350 (
);

FILL FILL_1__1540_ (
);

FILL FILL_1__1120_ (
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf0)
);

OAI21X1 _1395_ (
    .A(_483_),
    .B(_484_),
    .C(_475_),
    .Y(_485_)
);

FILL FILL_0__1855_ (
);

FILL FILL_0__1435_ (
);

FILL FILL_0__1015_ (
);

FILL FILL_1__986_ (
);

FILL FILL_0__1244_ (
);

FILL FILL_1__1825_ (
);

FILL FILL_1__1405_ (
);

FILL FILL_0__1893_ (
);

FILL FILL_0__1473_ (
);

FILL FILL_0__1053_ (
);

FILL FILL_1__1634_ (
);

FILL FILL_1__1214_ (
);

INVX1 _1489_ (
    .A(_576_),
    .Y(_577_)
);

NAND3X1 _1069_ (
    .A(_149_),
    .B(_156_),
    .C(_160_),
    .Y(_161_)
);

FILL FILL_0__1529_ (
);

FILL FILL_0__1109_ (
);

FILL FILL_0__1282_ (
);

NAND2X1 _1701_ (
    .A(AI[1]),
    .B(shr),
    .Y(_873_)
);

FILL FILL_1__1863_ (
);

FILL FILL_1__1443_ (
);

FILL FILL_1__1023_ (
);

OAI21X1 _1298_ (
    .A(_387_),
    .B(_135_),
    .C(_388_),
    .Y(_389_)
);

FILL FILL_0__1758_ (
);

FILL FILL_0__1338_ (
);

FILL FILL_0__1091_ (
);

NAND2X1 _1510_ (
    .A(_546_),
    .B(_593_),
    .Y(_598_)
);

FILL FILL_1__1252_ (
);

FILL FILL_2__1741_ (
);

FILL FILL_0__1567_ (
);

FILL FILL_0__1147_ (
);

FILL FILL_1__1728_ (
);

FILL FILL_1__1308_ (
);

FILL FILL_1__1481_ (
);

FILL FILL_1__1061_ (
);

FILL FILL_0__1796_ (
);

FILL FILL_0__1376_ (
);

FILL FILL_1__1537_ (
);

FILL FILL_1__1117_ (
);

FILL FILL_1__1290_ (
);

FILL FILL_0__1185_ (
);

NAND2X1 _1604_ (
    .A(LoadCmd_i),
    .B(ABCmd_i[2]),
    .Y(_685_)
);

FILL FILL_0__932_ (
);

OAI21X1 _935_ (
    .A(_725_),
    .B(_26_),
    .C(_720_),
    .Y(_27_)
);

FILL FILL_1__1766_ (
);

FILL FILL_1__1346_ (
);

FILL FILL86850x18150 (
);

INVX1 _1833_ (
    .A(_804_),
    .Y(ACC[6])
);

NAND3X1 _1413_ (
    .A(_458_),
    .B(_502_),
    .C(_494_),
    .Y(_503_)
);

FILL FILL_1__1575_ (
);

FILL FILL_1__1155_ (
);

FILL FILL_2__1644_ (
);

FILL FILL_2__999_ (
);

NAND2X1 _1642_ (
    .A(ABCmd_i[3]),
    .B(LoadB_i),
    .Y(_706_)
);

NAND3X1 _1222_ (
    .A(MUL_bF$buf2),
    .B(AI[6]),
    .C(BI[2]),
    .Y(_314_)
);

FILL FILL_0__970_ (
);

NAND3X1 _973_ (
    .A(_55_),
    .B(_56_),
    .C(_52_),
    .Y(_65_)
);

FILL FILL_1__1384_ (
);

FILL FILL_0__1699_ (
);

FILL FILL_0__1279_ (
);

AOI21X1 _1871_ (
    .A(_804_),
    .B(_789_),
    .C(_752_),
    .Y(_839_)
);

OR2X2 _1451_ (
    .A(_538_),
    .B(_539_),
    .Y(_540_)
);

AND2X2 _1031_ (
    .A(_114_),
    .B(_118_),
    .Y(_123_)
);

FILL FILL_1__1193_ (
);

FILL FILL_0__1088_ (
);

AND2X2 _1507_ (
    .A(_593_),
    .B(_546_),
    .Y(_595_)
);

FILL FILL_1__1249_ (
);

DFFPOSX1 _1680_ (
    .D(_21_),
    .CLK(clk_bF$buf0),
    .Q(BI[3])
);

AND2X2 _1260_ (
    .A(_347_),
    .B(_351_),
    .Y(_352_)
);

FILL FILL_0__1720_ (
);

FILL FILL_2__1318_ (
);

FILL FILL_0__1300_ (
);

OAI21X1 _1736_ (
    .A(_891_),
    .B(_893_),
    .C(_906_),
    .Y(_907_)
);

AOI21X1 _1316_ (
    .A(_404_),
    .B(_406_),
    .C(_396_),
    .Y(_407_)
);

FILL FILL_1__1478_ (
);

FILL FILL_1__1058_ (
);

NOR2X1 _1545_ (
    .A(_135_),
    .B(_540_),
    .Y(_632_)
);

OAI21X1 _1125_ (
    .A(_215_),
    .B(_216_),
    .C(_132_),
    .Y(_217_)
);

FILL FILL_1__1287_ (
);

FILL FILL_0__929_ (
);

NAND3X1 _1774_ (
    .A(_732_),
    .B(_747_),
    .C(_731_),
    .Y(_750_)
);

NAND3X1 _1354_ (
    .A(_378_),
    .B(_439_),
    .C(_440_),
    .Y(_445_)
);

FILL FILL_1__1096_ (
);

FILL FILL_0__1814_ (
);

FILL FILL_2__1585_ (
);

NOR2X1 _1583_ (
    .A(_646_),
    .B(_603_),
    .Y(_669_)
);

NAND3X1 _1163_ (
    .A(_233_),
    .B(_252_),
    .C(_254_),
    .Y(_255_)
);

FILL FILL_1__945_ (
);

FILL FILL_0__1623_ (
);

FILL FILL_0__1203_ (
);

OAI21X1 _1639_ (
    .A(LoadB_i),
    .B(_36_),
    .C(_704_),
    .Y(_19_)
);

NAND3X1 _1219_ (
    .A(_307_),
    .B(_310_),
    .C(_308_),
    .Y(_311_)
);

FILL FILL_0__967_ (
);

NAND3X1 _1392_ (
    .A(_476_),
    .B(_481_),
    .C(_479_),
    .Y(_482_)
);

FILL FILL_0__1852_ (
);

FILL FILL_0__1432_ (
);

FILL FILL_0__1012_ (
);

FILL FILL86550x64950 (
);

OAI21X1 _1868_ (
    .A(_828_),
    .B(_835_),
    .C(_836_),
    .Y(_837_)
);

AOI21X1 _1448_ (
    .A(_532_),
    .B(_534_),
    .C(_530_),
    .Y(_537_)
);

NAND3X1 _1028_ (
    .A(_102_),
    .B(_119_),
    .C(_106_),
    .Y(_120_)
);

FILL FILL_1__983_ (
);

endmodule
