magic
tech scmos
magscale 1 2
timestamp 1726836556
<< nwell >>
rect -12 154 132 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
<< ptransistor >>
rect 20 166 24 246
rect 30 166 34 246
rect 60 166 64 246
rect 70 166 74 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 44 40 54
rect 24 14 26 44
rect 38 14 40 44
rect 44 14 46 54
rect 58 14 60 54
rect 64 26 66 54
rect 78 26 80 54
rect 64 14 80 26
rect 84 14 86 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 30 246
rect 34 166 36 246
rect 58 166 60 246
rect 64 166 70 246
rect 74 166 76 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 44
rect 46 14 58 54
rect 66 26 78 54
rect 86 14 98 54
<< pdcontact >>
rect 6 166 18 246
rect 36 166 58 246
rect 76 166 88 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 126 266
<< polysilicon >>
rect 20 246 24 250
rect 30 246 34 250
rect 60 246 64 250
rect 70 246 74 250
rect 20 162 24 166
rect 10 158 24 162
rect 30 162 34 166
rect 30 158 44 162
rect 10 129 16 158
rect 10 82 16 117
rect 40 103 44 158
rect 36 91 44 103
rect 10 76 24 82
rect 20 54 24 76
rect 40 54 44 91
rect 60 54 64 166
rect 70 162 74 166
rect 70 158 88 162
rect 84 129 88 158
rect 84 82 88 117
rect 80 76 88 82
rect 80 54 84 76
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 4 117 16 129
rect 24 91 36 103
rect 84 117 96 129
rect 64 91 76 103
<< metal1 >>
rect -6 266 126 268
rect -6 252 126 254
rect 6 246 18 252
rect 76 246 88 252
rect 44 117 52 166
rect 43 72 52 103
rect 43 64 74 72
rect 6 54 58 56
rect 68 54 74 64
rect 18 50 46 54
rect 58 14 86 20
rect 26 8 38 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 3 103 17 117
rect 23 103 37 117
rect 43 103 57 117
rect 63 103 77 117
rect 83 103 97 117
<< metal2 >>
rect 26 117 34 135
rect 66 117 74 135
rect 6 87 14 103
rect 46 87 54 103
rect 86 87 94 103
<< m1p >>
rect -6 252 126 268
rect -6 -8 126 8
<< m2p >>
rect 26 119 34 135
rect 66 119 74 135
rect 6 87 14 101
rect 46 87 54 101
rect 86 87 94 101
<< labels >>
rlabel metal1 -6 252 106 268 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 7 nsew ground bidirectional abutment
rlabel metal2 10 91 10 91 1 A
port 1 n signal input
rlabel metal2 30 131 30 131 1 B
port 2 n signal input
rlabel metal2 50 89 50 89 5 Y
port 5 n signal output
rlabel metal2 70 131 70 131 1 D
port 4 n signal input
rlabel metal2 90 91 90 91 1 C
port 3 n signal input
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
