magic
tech scmos
magscale 1 30
timestamp 1724567886
<< checkpaint >>
rect 9150 149700 181740 180850
rect 9150 136300 182150 149700
rect 9150 9150 181740 136300
<< metal1 >>
rect 138300 103900 144500 113100
rect 44600 78200 49600 84800
<< m2contact >>
rect 144500 103900 145500 113100
rect 44100 78200 44600 84800
<< metal2 >>
rect 44100 140600 47600 141000
rect 47200 139900 47600 140600
rect 48900 140800 49400 145900
rect 62500 141500 62900 145900
rect 76000 142600 76400 145900
rect 76000 142200 95800 142600
rect 62500 141100 90400 141500
rect 48900 140400 83300 140800
rect 47200 139500 81100 139900
rect 48200 138300 66100 138700
rect 44100 116400 46000 116800
rect 48200 103200 48600 138300
rect 65700 137300 66100 138300
rect 80700 137300 81100 139500
rect 82900 137300 83300 140400
rect 90000 137300 90400 141100
rect 95400 137300 95800 142200
rect 100300 137700 100700 145900
rect 113700 144500 114200 145900
rect 127300 144900 127700 145900
rect 119800 144500 127700 144900
rect 113700 144100 118600 144500
rect 99700 137300 100700 137700
rect 102300 137300 102700 144000
rect 118200 137300 118600 144100
rect 119800 137300 120200 144500
rect 140800 143600 141200 145900
rect 142200 140800 145900 141200
rect 143600 127300 145900 127700
rect 145500 103900 145900 113100
rect 44100 102800 48600 103200
rect 44100 89300 45000 89700
rect 144900 89500 145900 89900
rect 142700 76000 145900 76400
rect 141800 73300 145900 73700
rect 44100 62300 46500 62700
rect 140400 59700 145900 60200
rect 87000 53000 87400 54300
rect 48900 52600 87400 53000
rect 48900 44100 49400 52600
rect 88200 52100 88600 54300
rect 73200 51700 88600 52100
rect 73200 44100 73700 51700
rect 88900 49200 89300 54300
rect 75900 48800 89300 49200
rect 75900 44100 76400 48800
rect 90400 45900 90800 54300
rect 93100 47700 93500 54300
rect 95200 49300 95600 54300
rect 107500 52200 107900 54300
rect 107500 51800 141200 52200
rect 95200 48900 113700 49300
rect 93100 47300 127700 47700
rect 90400 45500 100800 45900
rect 100300 44100 100800 45500
rect 113700 44100 114200 45100
rect 127200 44100 127700 47300
rect 140700 44100 141200 51800
<< m3contact >>
rect 46000 116400 46400 117200
rect 101900 144000 102700 144400
rect 140200 143200 141200 143600
rect 141500 140800 142200 141200
rect 142900 127300 143600 127700
rect 45000 89300 45400 90000
rect 144200 89500 144900 89900
rect 142000 76000 142700 76400
rect 141100 73300 141800 73700
rect 46500 62300 46900 63100
rect 139800 59700 140400 60200
rect 113700 48500 114200 49300
rect 113700 45100 114200 45900
<< metal3 >>
rect 46000 144000 101900 144400
rect 46000 117200 46400 144000
rect 45000 99400 48800 99800
rect 45000 90000 45400 99400
rect 46500 95100 48600 95500
rect 46500 63100 46900 95100
rect 140200 94700 140600 143200
rect 139400 94300 140600 94700
rect 141500 92000 141900 140800
rect 139400 91600 141900 92000
rect 142900 89600 143300 127300
rect 139400 89200 143300 89600
rect 144200 88100 144600 89500
rect 139400 87700 144600 88100
rect 139300 87000 142400 87400
rect 139400 83700 141500 84100
rect 139400 76500 140200 76900
rect 139800 60200 140200 76500
rect 141100 73700 141500 83700
rect 142000 76400 142400 87000
rect 113700 45900 114200 48500
use PIC  CIN_0
timestamp 1537935238
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_1
timestamp 1537935238
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_2
timestamp 1537935238
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_3
timestamp 1537935238
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use PIC  CIN_4
timestamp 1537935238
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC  CIN_5
timestamp 1537935238
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC  CLK
timestamp 1537935238
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use fir_pe_Core  fir_pe_Core_0
timestamp 1724553464
transform 1 0 50345 0 1 54560
box -1920 -375 89280 82845
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1719894731
transform 0 -1 171100 -1 0 75646
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_1
timestamp 1719894731
transform 0 -1 171100 -1 0 62146
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_2
timestamp 1719894731
transform 0 -1 171100 -1 0 102646
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_3
timestamp 1719894731
transform 0 -1 171100 -1 0 89146
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_4
timestamp 1719894731
transform 0 -1 171100 -1 0 129646
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_5
timestamp 1719894731
transform 0 -1 171100 -1 0 116146
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_6
timestamp 1719894731
transform 1 0 73845 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_7
timestamp 1719894731
transform 1 0 60345 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_8
timestamp 1719894731
transform 1 0 100845 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_9
timestamp 1719894731
transform 1 0 87345 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_10
timestamp 1719894731
transform 1 0 127845 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_11
timestamp 1719894731
transform 1 0 114345 0 1 18900
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_12
timestamp 1719894731
transform 0 1 18900 -1 0 75655
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_13
timestamp 1719894731
transform 0 1 18900 -1 0 62155
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_14
timestamp 1719894731
transform 0 1 18900 -1 0 102655
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_15
timestamp 1719894731
transform 0 1 18900 -1 0 89155
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_16
timestamp 1719894731
transform 1 0 73845 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_17
timestamp 1719894731
transform 0 1 18900 -1 0 116155
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_18
timestamp 1719894731
transform 0 1 18900 -1 0 129655
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_19
timestamp 1719894731
transform 1 0 60345 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_20
timestamp 1719894731
transform 1 0 100845 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_21
timestamp 1719894731
transform 1 0 87345 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_22
timestamp 1719894731
transform 1 0 127845 0 -1 171099
box 0 0 1800 25050
use IOFILLER18  IOFILLER18_23
timestamp 1719894731
transform 1 0 114345 0 -1 171099
box 0 0 1800 25050
use IOFILLER50  IOFILLER50_0
timestamp 1537935238
transform 1 0 43585 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 141465 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1537935238
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1537935238
transform 1 0 43585 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1537935238
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1537935238
transform 0 1 18900 -1 0 146415
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1537935238
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1537935238
transform 0 -1 171100 -1 0 146415
box -35 0 5035 25060
use MY_LOGO  MY_LOGO_0
timestamp 1724157349
transform 1 0 149430 0 1 12135
box 60 75 7170 3015
use PIC  PAD_27
timestamp 1537935238
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PCORNER  PCORNER_0
timestamp 1537935238
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1537935238
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1537935238
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1537935238
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  RDY
timestamp 1537935238
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PVDD  VDD_0
timestamp 1537935238
transform 0 1 18900 -1 0 87500
box 0 -9150 12000 25300
use PIC  VLD
timestamp 1537935238
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PVSS  VSS_0
timestamp 1537935238
transform 0 -1 171100 1 0 102500
box 0 -9150 12000 25300
use PIC  XIN_0
timestamp 1537935238
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  XIN_1
timestamp 1537935238
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  XIN_2
timestamp 1537935238
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use PIC  XIN_3
timestamp 1537935238
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use POB8  XOUT_0
timestamp 1537935238
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use POB8  XOUT_1
timestamp 1537935238
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  XOUT_2
timestamp 1537935238
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use POB8  XOUT_3
timestamp 1537935238
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use PIC  YIN_0
timestamp 1537935238
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  YIN_1
timestamp 1537935238
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  YIN_2
timestamp 1537935238
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  YIN_3
timestamp 1537935238
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT_0
timestamp 1537935238
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use POB8  YOUT_1
timestamp 1537935238
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT_2
timestamp 1537935238
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT_3
timestamp 1537935238
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
<< end >>
