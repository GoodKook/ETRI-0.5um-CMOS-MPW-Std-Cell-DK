magic
tech scmos
magscale 1 2
timestamp 1727572430
<< nwell >>
rect -12 152 252 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 34
rect 52 14 56 34
rect 72 14 76 34
rect 82 14 86 34
rect 104 14 108 34
rect 148 14 152 34
rect 158 14 162 34
rect 178 14 182 34
rect 188 14 192 34
rect 208 14 212 54
<< ptransistor >>
rect 20 166 24 246
rect 40 206 44 246
rect 52 206 56 246
rect 72 206 76 246
rect 84 206 88 246
rect 104 206 108 246
rect 148 206 152 246
rect 158 206 162 246
rect 178 226 182 246
rect 188 226 192 246
rect 208 166 212 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 34 35 54
rect 197 34 208 54
rect 24 14 26 34
rect 38 14 40 34
rect 44 14 52 34
rect 56 14 58 34
rect 70 14 72 34
rect 76 14 82 34
rect 86 14 88 34
rect 100 14 104 34
rect 108 14 110 34
rect 146 14 148 34
rect 152 14 158 34
rect 162 14 164 34
rect 176 14 178 34
rect 182 14 188 34
rect 192 14 194 34
rect 206 14 208 34
rect 212 14 214 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 206 52 246
rect 56 206 58 246
rect 70 206 72 246
rect 76 206 84 246
rect 88 206 90 246
rect 102 206 104 246
rect 108 206 110 246
rect 146 206 148 246
rect 152 206 158 246
rect 162 226 164 246
rect 176 226 178 246
rect 182 226 188 246
rect 192 226 194 246
rect 206 226 208 246
rect 162 206 172 226
rect 24 166 35 206
rect 197 166 208 226
rect 212 166 214 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 34
rect 58 14 70 34
rect 88 14 100 34
rect 110 14 122 34
rect 134 14 146 34
rect 164 14 176 34
rect 194 14 206 34
rect 214 14 226 54
<< pdcontact >>
rect 6 166 18 246
rect 26 206 38 246
rect 58 206 70 246
rect 90 206 102 246
rect 110 206 122 246
rect 134 206 146 246
rect 164 226 176 246
rect 194 226 206 246
rect 214 166 226 246
<< psubstratepcontact >>
rect -6 -6 246 6
<< nsubstratencontact >>
rect -6 254 246 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 52 246 56 250
rect 72 246 76 250
rect 84 246 88 250
rect 104 246 108 250
rect 148 246 152 250
rect 158 246 162 250
rect 178 246 182 250
rect 188 246 192 250
rect 208 246 212 250
rect 20 146 24 166
rect 12 140 24 146
rect 12 76 16 140
rect 40 129 44 206
rect 52 162 56 206
rect 72 200 76 206
rect 84 200 88 206
rect 64 150 76 154
rect 36 117 44 129
rect 12 64 19 76
rect 20 54 24 64
rect 40 34 44 117
rect 52 34 56 60
rect 72 34 76 150
rect 84 54 88 188
rect 104 148 108 206
rect 148 202 152 206
rect 82 52 88 54
rect 82 40 84 52
rect 82 34 86 40
rect 104 34 108 136
rect 116 200 152 202
rect 128 198 152 200
rect 158 197 162 206
rect 156 192 162 197
rect 116 42 120 188
rect 134 50 138 168
rect 156 76 160 192
rect 178 184 182 226
rect 180 172 182 184
rect 188 163 192 226
rect 158 69 160 76
rect 180 159 192 163
rect 180 115 184 159
rect 180 69 184 103
rect 158 64 172 69
rect 180 64 192 69
rect 168 50 172 64
rect 134 46 162 50
rect 168 46 182 50
rect 116 38 152 42
rect 148 34 152 38
rect 158 34 162 46
rect 178 34 182 46
rect 188 34 192 64
rect 208 54 212 166
rect 20 10 24 14
rect 40 10 44 14
rect 52 10 56 14
rect 72 10 76 14
rect 82 10 86 14
rect 104 10 108 14
rect 148 10 152 14
rect 158 10 162 14
rect 178 10 182 14
rect 188 10 192 14
rect 208 10 212 14
<< polycontact >>
rect 64 188 76 200
rect 84 188 96 200
rect 52 150 64 162
rect 24 117 36 129
rect 19 64 31 76
rect 52 60 64 72
rect 96 136 108 148
rect 84 40 96 52
rect 116 188 128 200
rect 134 168 146 180
rect 168 172 180 184
rect 146 64 158 76
rect 196 132 208 144
rect 180 103 192 115
<< metal1 >>
rect -6 266 246 268
rect -6 252 246 254
rect 26 246 38 252
rect 90 246 102 252
rect 134 246 146 252
rect 194 246 206 252
rect 46 206 58 214
rect 164 206 176 226
rect 46 202 57 206
rect 110 200 122 206
rect 96 192 116 200
rect 64 182 76 188
rect 146 172 168 180
rect 6 162 18 166
rect 134 162 140 168
rect 6 154 52 162
rect 6 54 12 154
rect 64 154 140 162
rect 57 136 96 144
rect 176 132 196 140
rect 214 117 222 166
rect 192 103 203 115
rect 217 103 222 117
rect 31 74 63 76
rect 103 76 117 83
rect 77 74 146 76
rect 31 72 146 74
rect 31 68 52 72
rect 64 68 146 72
rect 214 54 222 103
rect 96 40 118 48
rect 46 34 57 40
rect 110 34 118 40
rect 46 27 58 34
rect 162 28 164 34
rect 26 8 38 14
rect 88 8 100 14
rect 134 8 146 14
rect 194 8 206 14
rect -6 6 246 8
rect -6 -8 246 -6
<< m2contact >>
rect 43 188 57 202
rect 162 192 176 206
rect 63 168 77 182
rect 43 130 57 144
rect 162 130 176 144
rect 23 103 37 117
rect 203 103 217 117
rect 63 74 77 88
rect 103 83 117 97
rect 43 40 57 54
rect 162 34 176 48
<< metal2 >>
rect 47 144 54 188
rect 23 83 37 103
rect 47 54 54 130
rect 67 88 76 168
rect 162 144 170 192
rect 103 97 117 117
rect 162 48 170 130
rect 203 83 217 103
<< m2p >>
rect 103 103 117 117
rect 23 83 37 97
rect 203 83 217 97
<< labels >>
rlabel metal2 23 83 37 97 0 D
port 0 nsew signal input
rlabel metal2 103 103 117 117 0 CLK
port 1 nsew clock input
rlabel metal2 203 83 217 97 0 Q
port 2 nsew signal output
rlabel metal1 -6 252 246 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 246 8 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 240 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
