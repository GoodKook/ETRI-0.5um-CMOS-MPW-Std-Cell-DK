magic
tech scmos
magscale 1 2
timestamp 1727487319
<< nwell >>
rect -6 154 106 272
<< ntransistor >>
rect 24 14 28 54
rect 34 14 38 54
rect 56 14 60 34
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
<< ndiffusion >>
rect 22 14 24 54
rect 28 14 34 54
rect 38 14 40 54
rect 52 14 56 34
rect 60 14 62 34
<< pdiffusion >>
rect 18 174 20 246
rect 6 166 20 174
rect 24 178 26 246
rect 38 178 40 246
rect 24 166 40 178
rect 44 166 46 246
rect 58 166 60 246
rect 64 166 66 246
<< ndcontact >>
rect 10 14 22 54
rect 40 14 52 54
rect 62 14 74 34
<< pdcontact >>
rect 6 174 18 246
rect 26 178 38 246
rect 46 166 58 246
rect 66 166 78 246
<< psubstratepcontact >>
rect 0 -6 100 6
<< nsubstratencontact >>
rect 0 254 100 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 20 152 24 166
rect 40 152 44 166
rect 9 146 24 152
rect 30 146 44 152
rect 9 123 15 146
rect 30 129 36 146
rect 60 123 64 166
rect 10 64 16 111
rect 30 82 36 117
rect 56 111 64 123
rect 30 72 38 82
rect 10 58 28 64
rect 24 54 28 58
rect 34 54 38 72
rect 56 34 60 111
rect 24 10 28 14
rect 34 10 38 14
rect 56 10 60 14
<< polycontact >>
rect 4 111 16 123
rect 24 117 36 129
rect 44 111 56 123
<< metal1 >>
rect 0 266 100 268
rect 0 252 100 254
rect 26 246 38 252
rect 6 172 18 174
rect 6 166 46 172
rect 66 117 74 166
rect 66 54 74 103
rect 52 46 74 54
rect 10 8 22 14
rect 62 8 74 14
rect 0 6 100 8
rect 0 -8 100 -6
<< m2contact >>
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect 63 103 77 117
<< metal2 >>
rect 3 137 17 157
rect 43 137 57 157
rect 23 83 37 103
rect 63 83 77 103
<< m2p >>
rect 3 143 17 157
rect 43 143 57 157
rect 23 83 37 97
rect 63 83 77 97
<< labels >>
rlabel metal2 3 143 17 157 0 A
port 0 nsew signal input
rlabel metal2 23 83 37 97 0 B
port 1 nsew signal input
rlabel metal2 63 83 77 97 0 Y
port 3 nsew signal output
rlabel metal2 43 143 57 157 0 C
port 2 nsew signal input
rlabel metal1 0 252 100 254 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 0 -8 100 -6 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 0 266 100 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 0 254 100 266 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 0 6 100 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 0 -6 100 6 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
