magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -60 -60 148 202
use pmos4_CDNS_7230122529110  pmos4_CDNS_7230122529110_0
timestamp 1555596690
transform 1 0 8 0 1 8
box -8 -8 80 134
<< end >>
