#--------------------------------------------------
# LEF file for Route & Via Rile
#  Ported from osu050 by GoodKook@gmail.com
#

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.15 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.6 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH	    0.9 ;   # ETRI050 Rule: WIDTH=0.8
  SPACING	1.05 ;  # ETRI050 Rule: SPACING=0.8(1.0)
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 3.2e-05 ;
END metal1

LAYER via1
  TYPE	CUT ;
  SPACING	0.9 ;
END via1

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.05 ;  # ETRI050 Rule: WIDTH=1.0
  SPACING	1.2 ;   # ETRI050 Rule: SPACING=1.0(1.2)
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 1.6e-05 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.9 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.2 ;   # ETRI050 Rule: WIDTH=1.2
  SPACING	1.2 ;   # ETRI050 Rule: SPACING=1.0(1.2)
  RESISTANCE	RPERSQ 0.05 ;
  CAPACITANCE	CPERSQDIST 1e-05 ;
END metal3

SPACING
  SAMENET cc   via1	0.900 ;
  SAMENET via1 via2	0.900 ;
END SPACING

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via1 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via2 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal3 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M3_M2


VIARULE viagen21 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via1 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen32

VIARULE TURN1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END TURN3

SITE  corner
    CLASS	PAD ;
    SYMMETRY	R90 Y ;
    SIZE	300.000 BY 300.000 ;
END  corner

SITE  IO
    CLASS	PAD ;
    SYMMETRY	Y ;
    SIZE	90.000 BY 300.000 ;
END  IO

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	3.000 BY 30.000 ;
END  core

# =====================================================================
#  Core MACROS
# =====================================================================
