magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -15 -15 505 505
use pnp10_CDNS_723012252910  pnp10_CDNS_723012252910_0
timestamp 1554524574
transform 1 0 0 0 1 0
box 45 45 445 445
<< end >>
