magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -56 -56 84 324
<< genericcontact >>
rect 11 243 17 249
rect 11 215 17 221
rect 11 187 17 193
rect 11 159 17 165
rect 11 131 17 137
rect 11 103 17 109
rect 11 75 17 81
rect 11 47 17 53
rect 11 19 17 25
<< metal1 >>
rect 4 4 24 264
<< end >>
