magic
tech scmos
magscale 1 2
timestamp 1756350801
<< error_s >>
rect 4 6244 7916 6256
rect 4 6004 7916 6016
rect 4 5764 7916 5776
rect 4 5524 7916 5536
rect 4 5284 7916 5296
rect 4 5044 7916 5056
rect 4 4804 7916 4816
rect 4 4564 7916 4576
rect 4 4324 7916 4336
rect 4 4084 7916 4096
rect 4 3844 7916 3856
rect 4 3604 7916 3616
rect 4 3364 7916 3376
rect 4 3124 7916 3136
rect 4 2884 7916 2896
rect 4 2644 7916 2656
rect 4 2404 7916 2416
rect 4 2164 7916 2176
rect 4 1924 7916 1936
rect 4 1684 7916 1696
rect 4 1444 7916 1456
rect 4 1204 7916 1216
rect 4 964 7916 976
rect 4 724 7916 736
rect 4 484 7916 496
rect 4 244 7916 256
rect 4 4 7916 16
<< metal1 >>
rect -62 6242 30 6258
rect -62 5778 -2 6242
rect 7657 6107 7663 6173
rect 7922 6018 7982 6258
rect 7890 6002 7982 6018
rect 4207 5937 4233 5943
rect 6767 5917 6813 5923
rect 7037 5843 7043 5913
rect 7027 5837 7043 5843
rect -62 5762 30 5778
rect -62 5298 -2 5762
rect 5617 5603 5623 5673
rect 5607 5597 5623 5603
rect 7357 5583 7363 5673
rect 7347 5577 7363 5583
rect 7922 5538 7982 6002
rect 7890 5522 7982 5538
rect 6847 5437 6863 5443
rect 2407 5377 2433 5383
rect 6857 5383 6863 5437
rect 6857 5377 6873 5383
rect -62 5282 30 5298
rect -62 4818 -2 5282
rect 7922 5058 7982 5522
rect 7890 5042 7982 5058
rect 6917 4957 6933 4963
rect 6917 4927 6923 4957
rect 7227 4957 7243 4963
rect 7237 4923 7243 4957
rect 7237 4917 7273 4923
rect 7537 4907 7543 4973
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 6317 4647 6323 4713
rect 7147 4697 7213 4703
rect 7922 4578 7982 5042
rect 7890 4562 7982 4578
rect 7577 4523 7583 4533
rect 7427 4517 7443 4523
rect 7577 4517 7603 4523
rect 127 4497 153 4503
rect 5397 4497 5413 4503
rect 767 4477 783 4483
rect 777 4403 783 4477
rect 2477 4447 2483 4493
rect 5397 4427 5403 4497
rect 7307 4477 7333 4483
rect 3327 4417 3353 4423
rect 7437 4407 7443 4517
rect 7567 4497 7583 4503
rect 767 4397 783 4403
rect 7557 4403 7563 4473
rect 7547 4397 7563 4403
rect 7577 4383 7583 4497
rect 7597 4427 7603 4517
rect 7567 4377 7583 4383
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 2707 4257 2733 4263
rect 497 4163 503 4253
rect 5087 4237 5103 4243
rect 1267 4197 1283 4203
rect 487 4157 503 4163
rect 1277 4163 1283 4197
rect 1277 4157 1293 4163
rect 1537 4163 1543 4213
rect 1537 4157 1573 4163
rect 1637 4163 1643 4213
rect 1637 4157 1653 4163
rect 1857 4163 1863 4233
rect 1857 4157 1873 4163
rect 2257 4163 2263 4213
rect 2707 4177 2773 4183
rect 3357 4183 3363 4233
rect 3357 4177 3373 4183
rect 2257 4157 2273 4163
rect 4877 4143 4883 4193
rect 5097 4163 5103 4237
rect 7687 4237 7743 4243
rect 7387 4217 7403 4223
rect 5087 4157 5103 4163
rect 7397 4163 7403 4217
rect 7737 4183 7743 4237
rect 7737 4177 7753 4183
rect 7397 4157 7433 4163
rect 4867 4137 4883 4143
rect 7922 4098 7982 4562
rect 7890 4082 7982 4098
rect 297 4017 313 4023
rect 297 3947 303 4017
rect 547 3997 563 4003
rect 557 3987 563 3997
rect 1257 3967 1263 4033
rect 1957 4023 1963 4033
rect 1937 4017 1963 4023
rect 2117 4017 2133 4023
rect 1937 3923 1943 4017
rect 2117 3947 2123 4017
rect 2227 4017 2273 4023
rect 2657 4017 2673 4023
rect 2497 3943 2503 3973
rect 2497 3937 2553 3943
rect 2657 3943 2663 4017
rect 7757 4017 7813 4023
rect 2737 3977 2753 3983
rect 2627 3937 2673 3943
rect 2737 3943 2743 3977
rect 2717 3937 2743 3943
rect 5077 3943 5083 4013
rect 5387 3997 5403 4003
rect 5397 3947 5403 3997
rect 7627 3997 7643 4003
rect 5077 3937 5093 3943
rect 2717 3927 2723 3937
rect 5187 3937 5213 3943
rect 7537 3927 7543 3993
rect 1927 3917 1943 3923
rect 7637 3923 7643 3997
rect 7757 3967 7763 4017
rect 7707 3957 7753 3963
rect 7627 3917 7643 3923
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 2767 3777 2783 3783
rect 1357 3683 1363 3753
rect 1527 3737 1543 3743
rect 1357 3677 1373 3683
rect 1537 3663 1543 3737
rect 2567 3737 2583 3743
rect 1797 3683 1803 3713
rect 1787 3677 1803 3683
rect 2197 3683 2203 3713
rect 2187 3677 2203 3683
rect 2297 3683 2303 3733
rect 2297 3677 2333 3683
rect 1527 3657 1543 3663
rect 2577 3663 2583 3737
rect 2777 3703 2783 3777
rect 7587 3777 7603 3783
rect 2777 3697 2793 3703
rect 7597 3703 7603 3777
rect 7567 3697 7603 3703
rect 2577 3657 2593 3663
rect 7922 3618 7982 4082
rect 7890 3602 7982 3618
rect 2657 3557 2713 3563
rect 1947 3537 2013 3543
rect 1787 3517 1803 3523
rect 1797 3467 1803 3517
rect 1977 3497 1993 3503
rect 1977 3427 1983 3497
rect 2557 3443 2563 3533
rect 2657 3483 2663 3557
rect 3707 3537 3753 3543
rect 3447 3517 3463 3523
rect 2647 3477 2663 3483
rect 2547 3437 2563 3443
rect 2817 3443 2823 3513
rect 2817 3437 2833 3443
rect 3457 3443 3463 3517
rect 7757 3517 7773 3523
rect 7757 3487 7763 3517
rect 3447 3437 3463 3443
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 1427 3257 1453 3263
rect 647 3217 693 3223
rect 2337 3223 2343 3293
rect 2337 3217 2353 3223
rect 3497 3203 3503 3233
rect 6207 3217 6253 3223
rect 3497 3197 3513 3203
rect 7922 3138 7982 3602
rect 7890 3122 7982 3138
rect 3047 3077 3093 3083
rect 2887 3057 2933 3063
rect 3317 3063 3323 3073
rect 3307 3057 3323 3063
rect 3527 3057 3553 3063
rect 7607 3057 7633 3063
rect 987 3037 1003 3043
rect 997 2983 1003 3037
rect 3407 3037 3423 3043
rect 997 2977 1023 2983
rect 1017 2967 1023 2977
rect 3417 2963 3423 3037
rect 7507 3037 7523 3043
rect 7517 3003 7523 3037
rect 7517 2997 7543 3003
rect 7537 2983 7543 2997
rect 7537 2977 7553 2983
rect 3407 2957 3423 2963
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 1847 2797 1873 2803
rect 1237 2777 1253 2783
rect 1237 2703 1243 2777
rect 1237 2697 1253 2703
rect 7922 2658 7982 3122
rect 7890 2642 7982 2658
rect 7447 2597 7463 2603
rect 2467 2577 2513 2583
rect 2687 2577 2713 2583
rect 4817 2577 4833 2583
rect 3307 2557 3343 2563
rect 3337 2523 3343 2557
rect 3337 2517 3373 2523
rect 4817 2507 4823 2577
rect 4907 2557 4933 2563
rect 7457 2507 7463 2597
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 737 2243 743 2273
rect 2057 2257 2093 2263
rect 737 2237 753 2243
rect 2057 2223 2063 2257
rect 2157 2263 2163 2333
rect 3297 2317 3313 2323
rect 2157 2257 2173 2263
rect 3297 2247 3303 2317
rect 6757 2263 6763 2273
rect 6757 2257 6813 2263
rect 2047 2217 2063 2223
rect 2147 2197 2193 2203
rect 7922 2178 7982 2642
rect 7890 2162 7982 2178
rect 307 2097 323 2103
rect 317 2027 323 2097
rect 487 2097 553 2103
rect 2457 2097 2473 2103
rect 2457 2047 2463 2097
rect 2817 2007 2823 2113
rect 3967 2097 3983 2103
rect 3977 2043 3983 2097
rect 4097 2083 4103 2113
rect 4087 2077 4103 2083
rect 3977 2037 3993 2043
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 707 1857 723 1863
rect 657 1763 663 1813
rect 647 1757 663 1763
rect 717 1763 723 1857
rect 717 1757 733 1763
rect 797 1763 803 1833
rect 787 1757 803 1763
rect 1197 1817 1213 1823
rect 1197 1743 1203 1817
rect 3797 1817 3813 1823
rect 3797 1767 3803 1817
rect 2587 1757 2613 1763
rect 1187 1737 1203 1743
rect 5747 1737 5773 1743
rect 7287 1737 7313 1743
rect 7787 1737 7833 1743
rect 7922 1698 7982 2162
rect 7890 1682 7982 1698
rect 2337 1617 2353 1623
rect 1397 1597 1413 1603
rect 1397 1543 1403 1597
rect 2337 1603 2343 1617
rect 2527 1617 2543 1623
rect 2297 1597 2343 1603
rect 2297 1587 2303 1597
rect 2537 1587 2543 1617
rect 7887 1617 7903 1623
rect 3337 1567 3343 1613
rect 7897 1587 7903 1617
rect 1387 1537 1403 1543
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 1707 1297 1773 1303
rect 1007 1277 1033 1283
rect 7922 1218 7982 1682
rect 7890 1202 7982 1218
rect 2727 1157 2753 1163
rect 1977 1137 1993 1143
rect 327 1097 353 1103
rect 1977 1063 1983 1137
rect 2307 1137 2333 1143
rect 1977 1057 1993 1063
rect 2437 1063 2443 1153
rect 2437 1057 2453 1063
rect -62 962 30 978
rect -62 498 -2 962
rect 7922 738 7982 1202
rect 7890 722 7982 738
rect 647 637 663 643
rect 657 607 663 637
rect 1667 637 1683 643
rect 1677 587 1683 637
rect 6747 597 6793 603
rect 7657 587 7663 633
rect -62 482 30 498
rect -62 18 -2 482
rect 287 377 413 383
rect 527 317 553 323
rect 7922 258 7982 722
rect 7890 242 7982 258
rect 6147 177 6173 183
rect -62 2 30 18
rect 7922 2 7982 242
<< m2contact >>
rect 1433 6253 1447 6267
rect 3153 6253 3167 6267
rect 7653 6173 7667 6187
rect 7653 6093 7667 6107
rect 4193 5933 4207 5947
rect 4233 5933 4247 5947
rect 6753 5913 6767 5927
rect 6813 5913 6827 5927
rect 7033 5913 7047 5927
rect 7013 5833 7027 5847
rect 4073 5773 4087 5787
rect 4213 5773 4227 5787
rect 1113 5753 1127 5767
rect 3693 5753 3707 5767
rect 5053 5753 5067 5767
rect 5613 5673 5627 5687
rect 7353 5673 7367 5687
rect 5593 5593 5607 5607
rect 7333 5573 7347 5587
rect 6833 5433 6847 5447
rect 2393 5373 2407 5387
rect 2433 5373 2447 5387
rect 6873 5373 6887 5387
rect 3313 5273 3327 5287
rect 3733 5273 3747 5287
rect 4193 5273 4207 5287
rect 4353 5273 4367 5287
rect 4813 5273 4827 5287
rect 7533 4973 7547 4987
rect 6933 4953 6947 4967
rect 7213 4953 7227 4967
rect 6913 4913 6927 4927
rect 7273 4913 7287 4927
rect 7533 4893 7547 4907
rect 4373 4813 4387 4827
rect 3813 4793 3827 4807
rect 4293 4793 4307 4807
rect 6313 4713 6327 4727
rect 7133 4693 7147 4707
rect 7213 4693 7227 4707
rect 6313 4633 6327 4647
rect 7573 4533 7587 4547
rect 7413 4513 7427 4527
rect 113 4493 127 4507
rect 153 4493 167 4507
rect 2473 4493 2487 4507
rect 753 4473 767 4487
rect 753 4393 767 4407
rect 2473 4433 2487 4447
rect 5413 4493 5427 4507
rect 7293 4473 7307 4487
rect 7333 4473 7347 4487
rect 3313 4413 3327 4427
rect 3353 4413 3367 4427
rect 5393 4413 5407 4427
rect 7553 4493 7567 4507
rect 7553 4473 7567 4487
rect 7433 4393 7447 4407
rect 7533 4393 7547 4407
rect 7553 4373 7567 4387
rect 7593 4413 7607 4427
rect 4193 4313 4207 4327
rect 493 4253 507 4267
rect 2693 4253 2707 4267
rect 2733 4253 2747 4267
rect 473 4153 487 4167
rect 1853 4233 1867 4247
rect 3353 4233 3367 4247
rect 5073 4233 5087 4247
rect 1533 4213 1547 4227
rect 1633 4213 1647 4227
rect 1253 4193 1267 4207
rect 1293 4153 1307 4167
rect 1573 4153 1587 4167
rect 1653 4153 1667 4167
rect 2253 4213 2267 4227
rect 1873 4153 1887 4167
rect 2693 4173 2707 4187
rect 2773 4173 2787 4187
rect 4873 4193 4887 4207
rect 3373 4173 3387 4187
rect 2273 4153 2287 4167
rect 4853 4133 4867 4147
rect 5073 4153 5087 4167
rect 7673 4233 7687 4247
rect 7373 4213 7387 4227
rect 7753 4173 7767 4187
rect 7433 4153 7447 4167
rect 1253 4033 1267 4047
rect 1953 4033 1967 4047
rect 313 4013 327 4027
rect 533 3993 547 4007
rect 553 3973 567 3987
rect 1253 3953 1267 3967
rect 293 3933 307 3947
rect 1913 3913 1927 3927
rect 2133 4013 2147 4027
rect 2213 4013 2227 4027
rect 2273 4013 2287 4027
rect 2493 3973 2507 3987
rect 2113 3933 2127 3947
rect 2553 3933 2567 3947
rect 2613 3933 2627 3947
rect 2673 4013 2687 4027
rect 5073 4013 5087 4027
rect 2673 3933 2687 3947
rect 2753 3973 2767 3987
rect 5373 3993 5387 4007
rect 7533 3993 7547 4007
rect 7613 3993 7627 4007
rect 5093 3933 5107 3947
rect 5173 3933 5187 3947
rect 5213 3933 5227 3947
rect 5393 3933 5407 3947
rect 2713 3913 2727 3927
rect 7533 3913 7547 3927
rect 7613 3913 7627 3927
rect 7813 4013 7827 4027
rect 7693 3953 7707 3967
rect 7753 3953 7767 3967
rect 3913 3853 3927 3867
rect 4233 3833 4247 3847
rect 4653 3833 4667 3847
rect 4773 3833 4787 3847
rect 7593 3833 7607 3847
rect 2753 3773 2767 3787
rect 1353 3753 1367 3767
rect 1513 3733 1527 3747
rect 1373 3673 1387 3687
rect 1513 3653 1527 3667
rect 2293 3733 2307 3747
rect 2553 3733 2567 3747
rect 1793 3713 1807 3727
rect 2193 3713 2207 3727
rect 1773 3673 1787 3687
rect 2173 3673 2187 3687
rect 2333 3673 2347 3687
rect 7573 3773 7587 3787
rect 2793 3693 2807 3707
rect 7553 3693 7567 3707
rect 2593 3653 2607 3667
rect 1933 3533 1947 3547
rect 2013 3533 2027 3547
rect 2553 3533 2567 3547
rect 1773 3513 1787 3527
rect 1793 3453 1807 3467
rect 1993 3493 2007 3507
rect 2533 3433 2547 3447
rect 2633 3473 2647 3487
rect 2713 3553 2727 3567
rect 3693 3533 3707 3547
rect 3753 3533 3767 3547
rect 2813 3513 2827 3527
rect 3433 3513 3447 3527
rect 2833 3433 2847 3447
rect 3433 3433 3447 3447
rect 7773 3513 7787 3527
rect 7753 3473 7767 3487
rect 1973 3413 1987 3427
rect 4153 3373 4167 3387
rect 4533 3373 4547 3387
rect 4733 3353 4747 3367
rect 5433 3353 5447 3367
rect 7133 3353 7147 3367
rect 7813 3353 7827 3367
rect 2333 3293 2347 3307
rect 1413 3253 1427 3267
rect 1453 3253 1467 3267
rect 633 3213 647 3227
rect 693 3213 707 3227
rect 3493 3233 3507 3247
rect 2353 3213 2367 3227
rect 6193 3213 6207 3227
rect 6253 3213 6267 3227
rect 3513 3193 3527 3207
rect 3033 3073 3047 3087
rect 3093 3073 3107 3087
rect 3313 3073 3327 3087
rect 2873 3053 2887 3067
rect 2933 3053 2947 3067
rect 3293 3053 3307 3067
rect 3513 3053 3527 3067
rect 3553 3053 3567 3067
rect 7593 3053 7607 3067
rect 7633 3053 7647 3067
rect 973 3033 987 3047
rect 3393 3033 3407 3047
rect 1013 2953 1027 2967
rect 3393 2953 3407 2967
rect 7493 3033 7507 3047
rect 7553 2973 7567 2987
rect 3973 2873 3987 2887
rect 4853 2873 4867 2887
rect 4953 2873 4967 2887
rect 5533 2873 5547 2887
rect 5933 2873 5947 2887
rect 6233 2873 6247 2887
rect 6573 2873 6587 2887
rect 7433 2873 7447 2887
rect 7753 2873 7767 2887
rect 1833 2793 1847 2807
rect 1873 2793 1887 2807
rect 1253 2773 1267 2787
rect 1253 2693 1267 2707
rect 7433 2593 7447 2607
rect 2453 2573 2467 2587
rect 2513 2573 2527 2587
rect 2673 2573 2687 2587
rect 2713 2573 2727 2587
rect 3293 2553 3307 2567
rect 3373 2513 3387 2527
rect 4833 2573 4847 2587
rect 4893 2553 4907 2567
rect 4933 2553 4947 2567
rect 4813 2493 4827 2507
rect 7453 2493 7467 2507
rect 4353 2413 4367 2427
rect 4613 2413 4627 2427
rect 5933 2413 5947 2427
rect 6473 2413 6487 2427
rect 7473 2393 7487 2407
rect 2153 2333 2167 2347
rect 733 2273 747 2287
rect 753 2233 767 2247
rect 2033 2213 2047 2227
rect 2093 2253 2107 2267
rect 2173 2253 2187 2267
rect 3313 2313 3327 2327
rect 6753 2273 6767 2287
rect 6813 2253 6827 2267
rect 3293 2233 3307 2247
rect 2133 2193 2147 2207
rect 2193 2193 2207 2207
rect 2813 2113 2827 2127
rect 4093 2113 4107 2127
rect 293 2093 307 2107
rect 473 2093 487 2107
rect 553 2093 567 2107
rect 2473 2093 2487 2107
rect 2453 2033 2467 2047
rect 313 2013 327 2027
rect 3953 2093 3967 2107
rect 4073 2073 4087 2087
rect 3993 2033 4007 2047
rect 2813 1993 2827 2007
rect 6133 1933 6147 1947
rect 5393 1913 5407 1927
rect 7893 1913 7907 1927
rect 693 1853 707 1867
rect 653 1813 667 1827
rect 633 1753 647 1767
rect 793 1833 807 1847
rect 733 1753 747 1767
rect 773 1753 787 1767
rect 1173 1733 1187 1747
rect 1213 1813 1227 1827
rect 3813 1813 3827 1827
rect 2573 1753 2587 1767
rect 2613 1753 2627 1767
rect 3793 1753 3807 1767
rect 5733 1733 5747 1747
rect 5773 1733 5787 1747
rect 7273 1733 7287 1747
rect 7313 1733 7327 1747
rect 7773 1733 7787 1747
rect 7833 1733 7847 1747
rect 1373 1533 1387 1547
rect 1413 1593 1427 1607
rect 2353 1613 2367 1627
rect 2513 1613 2527 1627
rect 3333 1613 3347 1627
rect 7873 1613 7887 1627
rect 2293 1573 2307 1587
rect 2533 1573 2547 1587
rect 7893 1573 7907 1587
rect 3333 1553 3347 1567
rect 1693 1293 1707 1307
rect 1773 1293 1787 1307
rect 993 1273 1007 1287
rect 1033 1273 1047 1287
rect 2433 1153 2447 1167
rect 2713 1153 2727 1167
rect 2753 1153 2767 1167
rect 313 1093 327 1107
rect 353 1093 367 1107
rect 1993 1133 2007 1147
rect 2293 1133 2307 1147
rect 2333 1133 2347 1147
rect 1993 1053 2007 1067
rect 2453 1053 2467 1067
rect 6313 973 6327 987
rect 6453 953 6467 967
rect 7773 953 7787 967
rect 633 633 647 647
rect 1653 633 1667 647
rect 653 593 667 607
rect 7653 633 7667 647
rect 6733 593 6747 607
rect 6793 593 6807 607
rect 1673 573 1687 587
rect 7653 573 7667 587
rect 5693 473 5707 487
rect 7893 473 7907 487
rect 273 373 287 387
rect 413 373 427 387
rect 513 313 527 327
rect 553 313 567 327
rect 6133 173 6147 187
rect 6173 173 6187 187
<< metal2 >>
rect 16 5887 23 6153
rect 176 6136 183 6303
rect 276 6136 283 6303
rect 356 6136 363 6303
rect 456 6136 463 6303
rect 536 6136 543 6303
rect 36 5923 43 6133
rect 96 6067 103 6103
rect 36 5916 63 5923
rect 56 5667 63 5916
rect 156 5916 163 5973
rect 76 5656 83 5873
rect 196 5687 203 6123
rect 256 5967 263 6123
rect 316 5987 323 6133
rect 216 5683 223 5953
rect 216 5676 243 5683
rect 36 4936 43 5473
rect 56 5423 63 5633
rect 96 5487 103 5643
rect 136 5623 143 5653
rect 236 5643 243 5676
rect 216 5636 243 5643
rect 136 5616 163 5623
rect 56 5416 83 5423
rect 136 5143 143 5473
rect 196 5436 203 5623
rect 276 5487 283 5913
rect 296 5667 303 5933
rect 316 5916 323 5973
rect 436 5683 443 6123
rect 516 5907 523 6123
rect 556 6103 563 6133
rect 656 6123 663 6133
rect 636 6116 663 6123
rect 1316 6116 1343 6123
rect 556 6096 583 6103
rect 736 6096 763 6103
rect 816 6096 843 6103
rect 736 6087 743 6096
rect 536 5916 543 5933
rect 436 5676 463 5683
rect 236 5436 263 5443
rect 176 5387 183 5413
rect 256 5167 263 5436
rect 316 5267 323 5433
rect 76 4983 83 5143
rect 116 5136 143 5143
rect 256 5143 263 5153
rect 236 5136 263 5143
rect 76 4976 103 4983
rect 96 4963 103 4976
rect 96 4956 123 4963
rect 76 4656 103 4663
rect 16 4476 43 4483
rect 76 4476 83 4656
rect 116 4507 123 4956
rect 276 4956 303 4963
rect 136 4647 143 4663
rect 16 4443 23 4476
rect 16 4436 43 4443
rect 16 4167 23 4333
rect 36 4227 43 4436
rect 56 4347 63 4463
rect 96 4267 103 4463
rect 56 4207 63 4233
rect 96 4207 103 4253
rect 116 4187 123 4293
rect 36 4107 43 4183
rect 76 4167 83 4183
rect 56 4083 63 4113
rect 36 4076 63 4083
rect 16 3467 23 4053
rect 16 2507 23 3433
rect 36 3427 43 4076
rect 76 3787 83 4153
rect 96 4023 103 4173
rect 136 4027 143 4613
rect 196 4496 203 4573
rect 156 4247 163 4493
rect 216 4223 223 4533
rect 236 4247 243 4773
rect 256 4587 263 4653
rect 276 4647 283 4956
rect 336 4703 343 5653
rect 356 5463 363 5673
rect 456 5643 463 5676
rect 436 5636 463 5643
rect 376 5547 383 5623
rect 356 5456 383 5463
rect 356 5147 363 5433
rect 376 5416 383 5456
rect 436 5447 443 5533
rect 516 5436 523 5473
rect 416 5403 423 5423
rect 396 5396 423 5403
rect 396 5156 403 5396
rect 376 4927 383 4953
rect 316 4696 343 4703
rect 316 4547 323 4696
rect 336 4607 343 4663
rect 376 4647 383 4663
rect 276 4476 283 4513
rect 376 4503 383 4593
rect 396 4527 403 5113
rect 376 4496 403 4503
rect 316 4476 343 4483
rect 216 4216 243 4223
rect 196 4196 203 4213
rect 96 4016 123 4023
rect 96 3647 103 3703
rect 116 3607 123 4016
rect 156 3987 163 4193
rect 176 4147 183 4183
rect 236 4127 243 4216
rect 256 4127 263 4453
rect 316 4227 323 4333
rect 336 4283 343 4476
rect 396 4476 403 4496
rect 416 4487 423 5253
rect 476 4627 483 4933
rect 556 4787 563 5593
rect 576 5447 583 5873
rect 596 5587 603 5623
rect 616 5436 623 5533
rect 616 5163 623 5353
rect 596 5156 623 5163
rect 596 4947 603 5156
rect 616 4807 623 4943
rect 616 4703 623 4793
rect 596 4696 623 4703
rect 596 4663 603 4696
rect 456 4563 463 4593
rect 496 4567 503 4653
rect 436 4556 463 4563
rect 336 4276 363 4283
rect 316 4207 323 4213
rect 276 4087 283 4173
rect 296 4147 303 4183
rect 156 3707 163 3953
rect 36 3047 43 3393
rect 76 3127 83 3553
rect 96 3516 103 3573
rect 136 3523 143 3693
rect 156 3547 163 3653
rect 136 3516 163 3523
rect 116 3447 123 3493
rect 96 3207 103 3223
rect 36 2607 43 2773
rect 76 2567 83 2833
rect 96 2787 103 3033
rect 116 2827 123 3413
rect 156 3387 163 3516
rect 136 3267 143 3373
rect 156 3107 163 3313
rect 176 3087 183 4013
rect 236 4003 243 4033
rect 256 4016 263 4033
rect 216 3996 243 4003
rect 216 3696 223 3773
rect 236 3503 243 3973
rect 296 3963 303 4113
rect 316 4027 323 4073
rect 336 4067 343 4173
rect 356 4167 363 4276
rect 376 4027 383 4273
rect 396 4227 403 4433
rect 416 4196 423 4233
rect 436 4227 443 4556
rect 456 4307 463 4513
rect 496 4456 503 4513
rect 516 4447 523 4493
rect 536 4456 543 4553
rect 507 4256 513 4263
rect 456 4196 463 4253
rect 396 4147 403 4183
rect 476 4167 483 4183
rect 496 4163 503 4233
rect 536 4207 543 4413
rect 556 4287 563 4613
rect 576 4607 583 4663
rect 596 4656 623 4663
rect 596 4647 603 4656
rect 636 4627 643 6073
rect 656 5967 663 6053
rect 656 5936 663 5953
rect 716 5923 723 5953
rect 796 5923 803 5933
rect 816 5923 823 6096
rect 836 6087 843 6096
rect 1096 6087 1103 6103
rect 1336 6087 1343 6116
rect 1436 6107 1443 6253
rect 1456 6087 1463 6103
rect 1476 6087 1483 6133
rect 1676 6103 1683 6153
rect 1656 6096 1683 6103
rect 1696 6136 1723 6143
rect 716 5916 743 5923
rect 796 5916 823 5923
rect 856 5916 863 5973
rect 676 5867 683 5903
rect 676 5647 683 5853
rect 696 5487 703 5613
rect 716 5507 723 5633
rect 796 5587 803 5916
rect 816 5587 823 5623
rect 716 5416 723 5493
rect 736 5396 743 5453
rect 756 5416 763 5453
rect 796 5403 803 5513
rect 776 5396 803 5403
rect 756 5143 763 5153
rect 756 5136 783 5143
rect 776 5127 783 5136
rect 816 5127 823 5573
rect 856 5436 863 5553
rect 896 5447 903 5473
rect 916 5167 923 5953
rect 1236 5936 1243 6033
rect 1256 5967 1263 6083
rect 1456 6067 1463 6073
rect 1516 5967 1523 5993
rect 976 5916 1003 5923
rect 1036 5916 1063 5923
rect 976 5636 983 5916
rect 1056 5887 1063 5916
rect 1196 5916 1223 5923
rect 1136 5763 1143 5883
rect 1127 5756 1143 5763
rect 1156 5727 1163 5893
rect 956 5547 963 5593
rect 996 5427 1003 5653
rect 1036 5547 1043 5643
rect 1156 5643 1163 5713
rect 1196 5667 1203 5916
rect 1296 5876 1303 5913
rect 1316 5896 1323 5933
rect 1256 5663 1263 5873
rect 1336 5687 1343 5873
rect 1256 5656 1283 5663
rect 1156 5636 1183 5643
rect 1216 5636 1223 5653
rect 1256 5623 1263 5656
rect 1236 5616 1263 5623
rect 1016 5436 1023 5453
rect 1056 5436 1063 5573
rect 1276 5456 1283 5553
rect 1296 5507 1303 5643
rect 1316 5567 1323 5653
rect 1356 5643 1363 5953
rect 1456 5907 1463 5933
rect 1476 5916 1483 5933
rect 1516 5916 1523 5953
rect 1396 5703 1403 5903
rect 1376 5696 1403 5703
rect 1376 5667 1383 5696
rect 1396 5656 1403 5673
rect 1436 5656 1463 5663
rect 1336 5636 1363 5643
rect 1356 5487 1363 5636
rect 1176 5383 1183 5403
rect 1296 5387 1303 5413
rect 1176 5376 1203 5383
rect 1196 5156 1203 5376
rect 856 5136 863 5153
rect 996 5127 1003 5143
rect 716 4956 743 4963
rect 776 4956 783 5113
rect 716 4923 723 4956
rect 716 4916 743 4923
rect 576 4407 583 4533
rect 656 4487 663 4833
rect 596 4476 623 4483
rect 596 4447 603 4476
rect 636 4387 643 4453
rect 496 4156 543 4163
rect 356 3996 363 4013
rect 396 3996 403 4073
rect 436 4027 443 4153
rect 276 3956 303 3963
rect 256 3567 263 3833
rect 216 3496 243 3503
rect 216 3247 223 3496
rect 176 3067 183 3073
rect 196 3036 203 3053
rect 96 2627 103 2743
rect 96 2523 103 2573
rect 76 2516 103 2523
rect 16 1103 23 2453
rect 36 2107 43 2493
rect 76 2147 83 2293
rect 96 2247 103 2263
rect 116 2167 123 2773
rect 136 2727 143 2743
rect 136 2307 143 2593
rect 156 2587 163 2993
rect 216 2767 223 3093
rect 236 2947 243 3473
rect 256 3447 263 3533
rect 276 3516 283 3956
rect 296 3867 303 3933
rect 316 3687 323 3893
rect 336 3887 343 3983
rect 356 3703 363 3813
rect 336 3696 363 3703
rect 296 3547 303 3613
rect 316 3536 323 3553
rect 356 3547 363 3673
rect 376 3547 383 3673
rect 396 3667 403 3853
rect 416 3623 423 4013
rect 436 3887 443 3973
rect 456 3967 463 4153
rect 476 3996 483 4053
rect 536 4007 543 4133
rect 556 4003 563 4173
rect 576 4027 583 4313
rect 596 4147 603 4353
rect 616 4196 623 4253
rect 616 4107 623 4153
rect 636 4147 643 4163
rect 596 4016 603 4073
rect 616 4047 623 4093
rect 656 4087 663 4393
rect 676 4167 683 4573
rect 696 4476 703 4493
rect 736 4476 743 4916
rect 756 4487 763 4653
rect 776 4627 783 4643
rect 776 4567 783 4613
rect 816 4567 823 4853
rect 856 4703 863 4953
rect 836 4696 863 4703
rect 836 4647 843 4696
rect 856 4583 863 4663
rect 836 4576 863 4583
rect 836 4527 843 4576
rect 716 4367 723 4463
rect 756 4383 763 4393
rect 736 4376 763 4383
rect 716 4196 723 4233
rect 696 4167 703 4183
rect 736 4147 743 4376
rect 776 4227 783 4473
rect 796 4467 803 4513
rect 836 4487 843 4513
rect 796 4227 803 4453
rect 856 4447 863 4493
rect 876 4456 883 4633
rect 896 4487 903 4573
rect 916 4456 923 4683
rect 936 4487 943 4933
rect 956 4687 963 4753
rect 976 4703 983 5093
rect 996 4723 1003 4943
rect 996 4716 1023 4723
rect 976 4696 1003 4703
rect 816 4387 823 4443
rect 896 4423 903 4433
rect 896 4416 923 4423
rect 836 4347 843 4373
rect 556 3996 583 4003
rect 496 3967 503 3983
rect 456 3727 463 3953
rect 476 3627 483 3873
rect 516 3716 523 3953
rect 556 3947 563 3973
rect 596 3847 603 3973
rect 636 3967 643 4013
rect 496 3687 503 3703
rect 396 3616 423 3623
rect 296 3407 303 3503
rect 336 3367 343 3503
rect 256 3067 263 3253
rect 276 3227 283 3273
rect 296 3256 303 3273
rect 336 3256 343 3293
rect 256 3007 263 3053
rect 316 3007 323 3213
rect 356 3123 363 3493
rect 376 3223 383 3433
rect 396 3327 403 3616
rect 416 3267 423 3593
rect 476 3543 483 3573
rect 496 3567 503 3673
rect 556 3627 563 3713
rect 516 3547 523 3593
rect 476 3536 503 3543
rect 436 3516 463 3523
rect 496 3516 503 3536
rect 536 3516 543 3573
rect 436 3507 443 3516
rect 476 3467 483 3503
rect 476 3247 483 3453
rect 516 3247 523 3313
rect 376 3216 403 3223
rect 396 3127 403 3216
rect 416 3207 423 3223
rect 436 3167 443 3193
rect 456 3147 463 3223
rect 496 3187 503 3223
rect 516 3167 523 3203
rect 356 3116 383 3123
rect 176 2647 183 2753
rect 176 2556 183 2613
rect 216 2556 223 2573
rect 156 2227 163 2433
rect 176 2143 183 2293
rect 216 2267 223 2413
rect 236 2307 243 2793
rect 276 2787 283 2893
rect 336 2847 343 3113
rect 376 2963 383 3116
rect 376 2956 403 2963
rect 276 2756 283 2773
rect 256 2723 263 2733
rect 256 2716 283 2723
rect 276 2627 283 2716
rect 296 2707 303 2713
rect 276 2576 283 2613
rect 296 2547 303 2693
rect 256 2283 263 2513
rect 276 2287 283 2533
rect 236 2276 263 2283
rect 236 2207 243 2276
rect 256 2243 263 2253
rect 256 2236 283 2243
rect 176 2136 203 2143
rect 76 2076 83 2113
rect 116 2076 123 2113
rect 156 2076 163 2133
rect 56 1903 63 2053
rect 96 2047 103 2063
rect 76 1927 83 2033
rect 56 1896 83 1903
rect 36 1596 43 1813
rect 76 1687 83 1896
rect 176 1787 183 2113
rect 196 1907 203 2136
rect 216 1983 223 2173
rect 276 2167 283 2193
rect 236 2087 243 2153
rect 276 2107 283 2153
rect 296 2107 303 2213
rect 256 2076 263 2093
rect 216 1976 243 1983
rect 216 1927 223 1933
rect 136 1767 143 1783
rect 216 1776 223 1913
rect 76 1596 83 1633
rect 136 1623 143 1753
rect 116 1616 143 1623
rect 156 1616 163 1713
rect 96 1547 103 1613
rect 16 1096 43 1103
rect 36 167 43 633
rect 76 387 83 1293
rect 96 1247 103 1303
rect 116 1287 123 1616
rect 216 1596 223 1733
rect 236 1627 243 1976
rect 256 1667 263 2013
rect 276 1987 283 2053
rect 316 2047 323 2753
rect 336 2747 343 2773
rect 336 2227 343 2473
rect 356 2407 363 2813
rect 376 2383 383 2933
rect 396 2827 403 2956
rect 416 2783 423 3073
rect 436 3036 443 3073
rect 456 2807 463 3053
rect 516 2843 523 3033
rect 496 2836 523 2843
rect 496 2807 503 2836
rect 396 2776 423 2783
rect 396 2547 403 2776
rect 436 2756 443 2773
rect 476 2767 483 2773
rect 416 2687 423 2743
rect 456 2727 463 2743
rect 396 2467 403 2533
rect 356 2376 383 2383
rect 356 2243 363 2376
rect 396 2307 403 2373
rect 456 2327 463 2593
rect 496 2407 503 2633
rect 516 2607 523 2813
rect 536 2707 543 3073
rect 556 2867 563 3553
rect 576 3547 583 3793
rect 596 3667 603 3773
rect 616 3707 623 3773
rect 676 3747 683 3983
rect 696 3767 703 4013
rect 716 3807 723 4073
rect 736 3996 743 4073
rect 756 4027 763 4183
rect 816 4167 823 4183
rect 796 4087 803 4153
rect 836 4027 843 4293
rect 856 4196 863 4253
rect 856 4067 863 4153
rect 876 4147 883 4183
rect 796 3996 803 4013
rect 856 3996 863 4053
rect 896 4023 903 4333
rect 916 4207 923 4416
rect 936 4407 943 4443
rect 936 4207 943 4273
rect 916 4167 923 4193
rect 956 4187 963 4553
rect 976 4507 983 4593
rect 996 4503 1003 4696
rect 1016 4647 1023 4716
rect 1036 4507 1043 4773
rect 1056 4727 1063 4953
rect 1076 4847 1083 4963
rect 1156 4956 1163 5113
rect 1216 5107 1223 5123
rect 1296 5087 1303 5373
rect 1336 5127 1343 5143
rect 1336 5047 1343 5113
rect 1196 4956 1223 4963
rect 1216 4887 1223 4956
rect 1356 4907 1363 5473
rect 1376 5427 1383 5633
rect 1416 5627 1423 5643
rect 1456 5527 1463 5656
rect 1536 5647 1543 6093
rect 1556 5643 1563 6013
rect 1636 5987 1643 6083
rect 1696 6047 1703 6136
rect 1796 6136 1803 6153
rect 1736 6027 1743 6123
rect 1816 6047 1823 6123
rect 1836 6087 1843 6133
rect 2096 6127 2103 6153
rect 2116 6136 2143 6143
rect 2176 6136 2183 6153
rect 1576 5907 1583 5923
rect 1656 5916 1663 5953
rect 1556 5636 1583 5643
rect 1516 5587 1523 5623
rect 1596 5607 1603 5633
rect 1616 5616 1623 5633
rect 1676 5623 1683 5953
rect 1696 5916 1703 5933
rect 1716 5887 1723 5913
rect 1716 5707 1723 5873
rect 1676 5616 1703 5623
rect 1476 5467 1483 5553
rect 1556 5527 1563 5603
rect 1676 5567 1683 5616
rect 1756 5603 1763 5673
rect 1736 5596 1763 5603
rect 1436 5436 1463 5443
rect 1476 5436 1483 5453
rect 1456 5427 1463 5436
rect 1496 5147 1503 5433
rect 1376 5107 1383 5143
rect 1576 5143 1583 5553
rect 1676 5436 1683 5473
rect 1716 5456 1723 5473
rect 1696 5436 1703 5453
rect 1736 5436 1743 5596
rect 1656 5387 1663 5423
rect 1676 5143 1683 5393
rect 1756 5163 1763 5473
rect 1776 5387 1783 5413
rect 1796 5407 1803 5973
rect 1816 5367 1823 6013
rect 1856 6007 1863 6123
rect 2056 6116 2083 6123
rect 1956 5923 1963 6103
rect 2076 6087 2083 6116
rect 2036 6067 2043 6083
rect 2096 6047 2103 6113
rect 2116 6087 2123 6136
rect 2996 6136 3023 6143
rect 1876 5916 1903 5923
rect 1956 5916 1983 5923
rect 2016 5916 2023 5953
rect 1896 5887 1903 5916
rect 1876 5656 1903 5663
rect 1976 5656 1983 5873
rect 2056 5667 2063 5893
rect 2096 5887 2103 5923
rect 2156 5896 2163 6033
rect 2236 5987 2243 6113
rect 2256 6067 2263 6103
rect 2236 5936 2243 5973
rect 2256 5887 2263 5903
rect 2276 5887 2283 5913
rect 2296 5847 2303 6093
rect 2356 6087 2363 6123
rect 2896 6123 2903 6133
rect 2736 6116 2763 6123
rect 2876 6116 2903 6123
rect 2436 6103 2443 6113
rect 2736 6107 2743 6116
rect 2416 6096 2443 6103
rect 2336 5936 2343 5973
rect 2396 5727 2403 6033
rect 2416 5927 2423 6096
rect 2636 6096 2663 6103
rect 2556 5967 2563 6093
rect 2656 6083 2663 6096
rect 2656 6076 2683 6083
rect 2456 5867 2463 5883
rect 2516 5867 2523 5893
rect 2556 5847 2563 5903
rect 2596 5887 2603 5933
rect 2736 5923 2743 6093
rect 2876 6027 2883 6116
rect 2976 5967 2983 6103
rect 2996 6087 3003 6136
rect 3156 6103 3163 6253
rect 3096 6007 3103 6103
rect 3136 6096 3163 6103
rect 3276 6067 3283 6103
rect 2976 5936 2983 5953
rect 2716 5916 2743 5923
rect 1896 5587 1903 5656
rect 1896 5436 1903 5553
rect 1916 5547 1923 5573
rect 1916 5367 1923 5533
rect 1956 5456 1963 5513
rect 1976 5487 1983 5593
rect 1996 5587 2003 5643
rect 1976 5456 1983 5473
rect 1736 5156 1763 5163
rect 1776 5156 1803 5163
rect 1836 5156 1843 5353
rect 1576 5136 1603 5143
rect 1676 5136 1703 5143
rect 1416 4956 1423 5033
rect 1596 4987 1603 5136
rect 1696 5067 1703 5136
rect 1736 5123 1743 5156
rect 1736 5116 1763 5123
rect 1796 5047 1803 5156
rect 1856 5087 1863 5123
rect 1796 4987 1803 5013
rect 1956 5007 1963 5143
rect 1996 5027 2003 5143
rect 2016 5127 2023 5553
rect 2036 5347 2043 5633
rect 2056 5623 2063 5653
rect 2096 5636 2103 5693
rect 2156 5643 2163 5713
rect 2136 5636 2163 5643
rect 2216 5636 2223 5673
rect 2256 5636 2283 5643
rect 2056 5616 2083 5623
rect 2076 5436 2083 5473
rect 2116 5436 2123 5453
rect 2156 5436 2163 5533
rect 2196 5527 2203 5623
rect 2276 5607 2283 5636
rect 2376 5636 2383 5673
rect 2236 5587 2243 5603
rect 2316 5567 2323 5633
rect 2336 5607 2343 5623
rect 2396 5587 2403 5613
rect 2176 5427 2183 5453
rect 2136 5407 2143 5423
rect 1736 4956 1763 4963
rect 1796 4956 1803 4973
rect 1056 4696 1063 4713
rect 1076 4643 1083 4683
rect 1136 4676 1143 4733
rect 1076 4636 1103 4643
rect 1096 4627 1103 4636
rect 996 4496 1023 4503
rect 976 4287 983 4453
rect 996 4327 1003 4433
rect 1016 4267 1023 4496
rect 1056 4476 1063 4533
rect 1076 4487 1083 4613
rect 1116 4527 1123 4653
rect 1156 4587 1163 4663
rect 1176 4627 1183 4683
rect 1116 4476 1143 4483
rect 1176 4476 1183 4533
rect 1036 4427 1043 4463
rect 1096 4447 1103 4463
rect 1136 4427 1143 4476
rect 1056 4327 1063 4373
rect 876 4016 903 4023
rect 716 3743 723 3773
rect 696 3736 723 3743
rect 696 3716 703 3736
rect 676 3687 683 3703
rect 716 3687 723 3703
rect 596 3523 603 3653
rect 616 3536 623 3573
rect 636 3567 643 3613
rect 656 3567 663 3673
rect 736 3607 743 3933
rect 756 3847 763 3983
rect 776 3963 783 3973
rect 776 3956 803 3963
rect 756 3747 763 3813
rect 776 3747 783 3913
rect 796 3727 803 3956
rect 816 3947 823 3983
rect 836 3947 843 3983
rect 576 3516 603 3523
rect 636 3516 643 3553
rect 676 3543 683 3573
rect 656 3536 683 3543
rect 576 3327 583 3516
rect 616 3287 623 3493
rect 636 3227 643 3243
rect 576 2923 583 3193
rect 616 3147 623 3223
rect 636 3067 643 3213
rect 576 2916 603 2923
rect 536 2576 543 2673
rect 576 2627 583 2813
rect 596 2787 603 2916
rect 636 2863 643 2993
rect 656 2927 663 3536
rect 716 3516 723 3593
rect 756 3587 763 3713
rect 776 3667 783 3703
rect 756 3523 763 3553
rect 756 3516 783 3523
rect 796 3516 803 3593
rect 816 3547 823 3693
rect 836 3667 843 3853
rect 856 3607 863 3953
rect 676 3487 683 3513
rect 736 3487 743 3503
rect 776 3463 783 3516
rect 756 3456 783 3463
rect 736 3247 743 3413
rect 756 3267 763 3456
rect 696 3227 703 3243
rect 776 3223 783 3433
rect 816 3407 823 3493
rect 856 3407 863 3503
rect 876 3467 883 4016
rect 916 3996 923 4133
rect 936 3987 943 4153
rect 956 3963 963 4173
rect 976 4167 983 4183
rect 996 4147 1003 4253
rect 1036 4167 1043 4233
rect 1076 4196 1083 4373
rect 1156 4227 1163 4463
rect 1196 4447 1203 4733
rect 1176 4327 1183 4353
rect 1196 4227 1203 4413
rect 1216 4347 1223 4713
rect 1236 4676 1243 4733
rect 1276 4676 1303 4683
rect 1256 4647 1263 4663
rect 1276 4496 1283 4676
rect 1336 4503 1343 4773
rect 1316 4496 1343 4503
rect 1316 4463 1323 4496
rect 1376 4476 1383 4873
rect 1436 4643 1443 4693
rect 1416 4636 1443 4643
rect 1456 4583 1463 4953
rect 1496 4827 1503 4953
rect 1496 4707 1503 4813
rect 1456 4576 1483 4583
rect 1436 4496 1443 4533
rect 1256 4387 1263 4463
rect 1296 4456 1323 4463
rect 1236 4347 1243 4373
rect 1056 4123 1063 4183
rect 1056 4116 1083 4123
rect 996 3996 1023 4003
rect 1056 3996 1063 4073
rect 956 3956 983 3963
rect 896 3727 903 3813
rect 916 3716 923 3753
rect 896 3667 903 3683
rect 936 3567 943 3873
rect 956 3587 963 3773
rect 976 3747 983 3956
rect 1016 3907 1023 3996
rect 1076 3987 1083 4116
rect 996 3716 1003 3753
rect 1016 3747 1023 3893
rect 1016 3647 1023 3703
rect 1056 3687 1063 3703
rect 1036 3647 1043 3673
rect 1076 3607 1083 3713
rect 1096 3667 1103 4213
rect 1216 4196 1223 4313
rect 1276 4283 1283 4433
rect 1296 4307 1303 4456
rect 1396 4443 1403 4463
rect 1456 4443 1463 4463
rect 1396 4436 1463 4443
rect 1476 4407 1483 4576
rect 1496 4403 1503 4673
rect 1536 4663 1543 4793
rect 1516 4647 1523 4663
rect 1536 4656 1563 4663
rect 1556 4507 1563 4656
rect 1576 4547 1583 4833
rect 1596 4527 1603 4943
rect 1676 4543 1683 4633
rect 1696 4567 1703 4653
rect 1736 4647 1743 4956
rect 1776 4676 1783 4933
rect 1936 4727 1943 4943
rect 1676 4536 1703 4543
rect 1536 4476 1543 4493
rect 1556 4447 1563 4463
rect 1536 4407 1543 4433
rect 1496 4396 1523 4403
rect 1316 4307 1323 4353
rect 1256 4276 1283 4283
rect 1256 4207 1263 4276
rect 1116 4167 1123 4183
rect 1176 4147 1183 4183
rect 1116 3827 1123 4113
rect 1176 3996 1183 4093
rect 1196 4047 1203 4193
rect 1236 4176 1263 4183
rect 1136 3867 1143 3893
rect 1116 3767 1123 3813
rect 1136 3716 1143 3773
rect 1156 3743 1163 3953
rect 1176 3927 1183 3953
rect 1176 3867 1183 3913
rect 1196 3807 1203 3983
rect 1236 3747 1243 4053
rect 1256 4047 1263 4176
rect 1276 4067 1283 4253
rect 1356 4207 1363 4253
rect 1296 4127 1303 4153
rect 1336 4147 1343 4183
rect 1376 4167 1383 4183
rect 1356 4127 1363 4153
rect 1396 4147 1403 4393
rect 1416 4147 1423 4233
rect 1296 4016 1303 4033
rect 1256 3987 1263 4013
rect 1316 3996 1323 4013
rect 1256 3787 1263 3953
rect 1296 3767 1303 3873
rect 1156 3736 1183 3743
rect 1176 3716 1183 3736
rect 1296 3727 1303 3753
rect 1156 3607 1163 3703
rect 1196 3667 1203 3703
rect 1316 3703 1323 3873
rect 1336 3767 1343 4113
rect 1436 4107 1443 4373
rect 1496 4196 1503 4373
rect 1516 4227 1523 4396
rect 1556 4387 1563 4433
rect 1536 4227 1543 4293
rect 1356 3887 1363 4053
rect 1396 4023 1403 4073
rect 1396 4016 1423 4023
rect 1416 4003 1423 4016
rect 1416 3996 1443 4003
rect 1376 3887 1383 3983
rect 1356 3767 1363 3853
rect 1376 3807 1383 3853
rect 1296 3696 1323 3703
rect 976 3527 983 3533
rect 996 3516 1003 3533
rect 856 3367 863 3393
rect 876 3287 883 3293
rect 716 3167 723 3223
rect 756 3216 783 3223
rect 676 3036 683 3073
rect 696 3003 703 3113
rect 676 2996 703 3003
rect 636 2856 663 2863
rect 556 2556 563 2573
rect 396 2276 403 2293
rect 416 2247 423 2263
rect 356 2236 383 2243
rect 356 2076 363 2113
rect 376 2107 383 2236
rect 396 2076 403 2173
rect 296 1927 303 2033
rect 136 1287 143 1303
rect 96 807 103 823
rect 96 636 103 653
rect 116 407 123 1113
rect 136 1107 143 1273
rect 136 767 143 813
rect 136 647 143 753
rect 156 687 163 1413
rect 176 1223 183 1553
rect 196 1487 203 1573
rect 236 1547 243 1583
rect 216 1307 223 1493
rect 176 1216 203 1223
rect 176 827 183 1093
rect 196 1067 203 1216
rect 236 1103 243 1173
rect 256 1127 263 1393
rect 276 1127 283 1893
rect 316 1787 323 2013
rect 336 1747 343 1783
rect 296 1567 303 1693
rect 356 1627 363 2013
rect 376 1967 383 2063
rect 376 1767 383 1783
rect 316 1207 323 1613
rect 336 1596 343 1613
rect 396 1587 403 1733
rect 416 1707 423 2213
rect 436 2087 443 2213
rect 456 2096 463 2263
rect 476 2107 483 2393
rect 496 2207 503 2393
rect 576 2363 583 2613
rect 596 2387 603 2713
rect 616 2587 623 2853
rect 636 2707 643 2743
rect 656 2647 663 2856
rect 676 2727 683 2996
rect 716 2947 723 3113
rect 796 3027 803 3233
rect 816 3187 823 3223
rect 876 3203 883 3273
rect 896 3227 903 3513
rect 976 3447 983 3513
rect 976 3367 983 3433
rect 916 3267 923 3293
rect 876 3196 903 3203
rect 816 3127 823 3173
rect 816 3016 823 3053
rect 836 3036 843 3073
rect 876 3036 883 3113
rect 756 2987 763 3013
rect 716 2736 743 2743
rect 736 2727 743 2736
rect 576 2356 603 2363
rect 556 2287 563 2313
rect 496 2187 503 2193
rect 456 2027 463 2053
rect 456 1827 463 1993
rect 476 1847 483 1893
rect 496 1807 503 2113
rect 516 2047 523 2273
rect 596 2267 603 2356
rect 576 2256 593 2263
rect 616 2247 623 2553
rect 656 2327 663 2573
rect 716 2567 723 2693
rect 516 1867 523 2033
rect 536 1967 543 2233
rect 576 2167 583 2233
rect 636 2227 643 2293
rect 696 2276 703 2493
rect 716 2303 723 2513
rect 736 2367 743 2633
rect 756 2447 763 2953
rect 776 2687 783 2933
rect 796 2787 803 2873
rect 836 2727 843 2913
rect 796 2667 803 2713
rect 796 2307 803 2563
rect 816 2447 823 2713
rect 856 2603 863 3013
rect 896 2967 903 3196
rect 916 3167 923 3223
rect 916 3036 923 3073
rect 956 3036 973 3043
rect 936 2947 943 3023
rect 996 2927 1003 3393
rect 1016 3147 1023 3593
rect 1036 3387 1043 3533
rect 1076 3467 1083 3523
rect 1036 3327 1043 3373
rect 1076 3303 1083 3453
rect 1056 3296 1083 3303
rect 1056 3283 1063 3296
rect 1036 3276 1063 3283
rect 1036 3256 1043 3276
rect 1076 3256 1083 3273
rect 1016 2967 1023 2973
rect 1056 2967 1063 3003
rect 1076 2863 1083 3213
rect 1096 3207 1103 3573
rect 1116 3527 1123 3553
rect 1136 3487 1143 3503
rect 1136 3467 1143 3473
rect 1196 3467 1203 3613
rect 1116 3067 1123 3233
rect 1136 3227 1143 3373
rect 1176 3227 1183 3453
rect 1216 3363 1223 3593
rect 1236 3587 1243 3693
rect 1256 3567 1263 3653
rect 1276 3587 1283 3673
rect 1296 3607 1303 3696
rect 1276 3536 1283 3553
rect 1236 3516 1263 3523
rect 1296 3516 1303 3593
rect 1236 3467 1243 3516
rect 1196 3356 1223 3363
rect 1196 3307 1203 3356
rect 1276 3347 1283 3493
rect 1216 3223 1223 3313
rect 1256 3247 1263 3313
rect 1196 3187 1203 3223
rect 1216 3216 1243 3223
rect 1136 3083 1143 3173
rect 1136 3076 1163 3083
rect 1096 2887 1103 3013
rect 1116 3007 1123 3033
rect 1136 2947 1143 3053
rect 1156 3036 1163 3076
rect 1196 3036 1203 3113
rect 1216 2987 1223 3193
rect 1256 3167 1263 3213
rect 1236 3067 1243 3093
rect 1276 3063 1283 3333
rect 1316 3067 1323 3153
rect 1256 3056 1283 3063
rect 1236 2967 1243 3033
rect 1256 3027 1263 3056
rect 1076 2856 1103 2863
rect 876 2723 883 2773
rect 916 2756 923 2853
rect 956 2756 963 2773
rect 1036 2756 1043 2773
rect 976 2727 983 2743
rect 876 2716 903 2723
rect 836 2596 863 2603
rect 716 2296 743 2303
rect 736 2287 743 2296
rect 776 2276 783 2293
rect 816 2287 823 2353
rect 836 2327 843 2596
rect 856 2547 863 2563
rect 896 2467 903 2716
rect 1016 2707 1023 2723
rect 1096 2707 1103 2856
rect 856 2287 863 2433
rect 876 2276 883 2333
rect 536 1887 543 1953
rect 456 1776 483 1783
rect 476 1727 483 1776
rect 356 1567 363 1583
rect 216 1096 243 1103
rect 256 1103 263 1113
rect 316 1107 323 1193
rect 356 1123 363 1553
rect 376 1287 383 1303
rect 396 1267 403 1453
rect 416 1227 423 1653
rect 436 1427 443 1613
rect 456 1567 463 1673
rect 496 1587 503 1773
rect 516 1747 523 1833
rect 556 1827 563 2093
rect 576 2076 583 2153
rect 596 2096 603 2133
rect 616 2107 623 2213
rect 636 2076 643 2193
rect 656 2127 663 2273
rect 676 2207 683 2263
rect 736 2256 763 2263
rect 736 2223 743 2256
rect 796 2247 803 2263
rect 716 2216 743 2223
rect 716 2207 723 2216
rect 676 2076 683 2153
rect 696 2087 703 2173
rect 736 2083 743 2193
rect 756 2187 763 2233
rect 716 2076 743 2083
rect 756 2076 763 2113
rect 776 2096 783 2213
rect 796 2107 803 2173
rect 796 2076 803 2093
rect 596 1907 603 2053
rect 656 1987 663 2063
rect 616 1796 623 1853
rect 676 1843 683 2033
rect 716 1987 723 2076
rect 696 1867 703 1953
rect 736 1927 743 2053
rect 676 1836 703 1843
rect 667 1816 683 1823
rect 676 1796 683 1816
rect 696 1807 703 1836
rect 536 1507 543 1633
rect 556 1596 563 1753
rect 596 1607 603 1783
rect 636 1767 643 1783
rect 656 1747 663 1793
rect 456 1296 463 1373
rect 336 1116 363 1123
rect 256 1096 283 1103
rect 216 816 223 1096
rect 236 827 243 1033
rect 216 567 223 643
rect 56 323 63 363
rect 96 356 103 373
rect 116 327 123 343
rect 56 316 83 323
rect 76 127 83 316
rect 96 156 103 313
rect 136 167 143 173
rect 176 167 183 343
rect 216 207 223 393
rect 256 383 263 873
rect 296 867 303 1083
rect 316 1047 323 1073
rect 336 1027 343 1116
rect 276 587 283 813
rect 296 807 303 823
rect 336 807 343 823
rect 356 787 363 1093
rect 376 887 383 1213
rect 476 1167 483 1313
rect 416 1136 423 1153
rect 396 1116 403 1133
rect 436 1116 463 1123
rect 376 867 383 873
rect 416 747 423 823
rect 436 707 443 933
rect 456 747 463 1116
rect 496 1116 503 1303
rect 536 1127 543 1253
rect 476 1107 483 1113
rect 556 1047 563 1193
rect 576 1107 583 1433
rect 596 1347 603 1373
rect 636 1343 643 1573
rect 636 1336 663 1343
rect 656 1207 663 1336
rect 616 1127 623 1133
rect 656 1116 663 1153
rect 676 1127 683 1693
rect 696 1687 703 1763
rect 696 1607 703 1673
rect 716 1667 723 1893
rect 776 1847 783 2013
rect 787 1836 793 1843
rect 816 1827 823 2233
rect 836 2187 843 2263
rect 856 2227 863 2243
rect 876 2207 883 2233
rect 836 2027 843 2113
rect 856 2076 863 2133
rect 896 2076 903 2193
rect 916 2047 923 2673
rect 936 2567 943 2613
rect 956 2487 963 2693
rect 996 2547 1003 2633
rect 956 2276 963 2453
rect 1056 2427 1063 2593
rect 1096 2556 1103 2653
rect 936 2227 943 2253
rect 976 2187 983 2333
rect 996 2307 1003 2413
rect 836 2007 843 2013
rect 736 1767 743 1783
rect 776 1767 783 1783
rect 736 1647 743 1753
rect 756 1647 763 1733
rect 696 1387 703 1563
rect 716 1316 723 1373
rect 756 1343 763 1633
rect 776 1527 783 1733
rect 796 1467 803 1813
rect 816 1603 823 1653
rect 836 1627 843 1753
rect 856 1707 863 2033
rect 936 2007 943 2113
rect 956 2067 963 2153
rect 996 2107 1003 2153
rect 976 2076 983 2093
rect 1016 2076 1023 2133
rect 1036 2107 1043 2313
rect 1076 2307 1083 2533
rect 1116 2407 1123 2913
rect 1136 2787 1143 2833
rect 1176 2807 1183 2853
rect 1156 2756 1163 2773
rect 1156 2556 1163 2673
rect 1176 2567 1183 2743
rect 1216 2707 1223 2733
rect 1236 2667 1243 2833
rect 1256 2787 1263 2913
rect 1296 2907 1303 3013
rect 1336 2783 1343 3733
rect 1356 3667 1363 3733
rect 1396 3716 1403 3833
rect 1416 3767 1423 3953
rect 1436 3927 1443 3953
rect 1476 3927 1483 4033
rect 1436 3716 1443 3833
rect 1476 3707 1483 3873
rect 1496 3807 1503 4133
rect 1516 4127 1523 4183
rect 1516 4107 1523 4113
rect 1536 4043 1543 4193
rect 1527 4036 1543 4043
rect 1516 3996 1523 4033
rect 1556 4027 1563 4273
rect 1596 4207 1603 4233
rect 1616 4227 1623 4533
rect 1636 4247 1643 4493
rect 1696 4476 1703 4536
rect 1656 4223 1663 4293
rect 1647 4216 1663 4223
rect 1676 4207 1683 4463
rect 1716 4443 1723 4453
rect 1716 4436 1743 4443
rect 1716 4243 1723 4413
rect 1736 4387 1743 4436
rect 1736 4267 1743 4373
rect 1716 4236 1743 4243
rect 1576 4047 1583 4153
rect 1616 4123 1623 4183
rect 1636 4143 1643 4193
rect 1656 4167 1663 4173
rect 1676 4147 1683 4163
rect 1636 4136 1663 4143
rect 1656 4123 1663 4136
rect 1616 4116 1643 4123
rect 1656 4116 1683 4123
rect 1496 3716 1503 3753
rect 1516 3747 1523 3913
rect 1536 3907 1543 4013
rect 1556 3996 1583 4003
rect 1576 3927 1583 3996
rect 1616 3947 1623 4013
rect 1636 3907 1643 4116
rect 1656 3996 1663 4053
rect 1676 4016 1683 4116
rect 1696 4067 1703 4173
rect 1716 4107 1723 4193
rect 1707 3996 1723 4003
rect 1716 3947 1723 3996
rect 1736 3907 1743 4236
rect 1756 4227 1763 4533
rect 1776 4247 1783 4633
rect 1816 4503 1823 4553
rect 1816 4496 1843 4503
rect 1856 4496 1863 4653
rect 1916 4623 1923 4713
rect 1896 4616 1923 4623
rect 1836 4447 1843 4496
rect 1856 4423 1863 4453
rect 1836 4416 1863 4423
rect 1816 4196 1823 4253
rect 1836 4227 1843 4416
rect 1856 4267 1863 4293
rect 1876 4243 1883 4453
rect 1867 4236 1883 4243
rect 1896 4227 1903 4616
rect 1916 4287 1923 4593
rect 1936 4227 1943 4663
rect 1956 4367 1963 4733
rect 1996 4667 2003 5013
rect 2036 4983 2043 5233
rect 2076 5136 2083 5233
rect 2196 5007 2203 5423
rect 2236 5183 2243 5513
rect 2316 5467 2323 5553
rect 2256 5436 2283 5443
rect 2256 5207 2263 5436
rect 2416 5427 2423 5713
rect 2616 5623 2623 5633
rect 2596 5607 2603 5623
rect 2616 5616 2643 5623
rect 2476 5487 2483 5573
rect 2476 5456 2483 5473
rect 2336 5407 2343 5423
rect 2396 5387 2403 5403
rect 2236 5176 2263 5183
rect 2256 5156 2263 5176
rect 2216 5143 2223 5153
rect 2216 5136 2243 5143
rect 2036 4976 2063 4983
rect 2116 4956 2123 4973
rect 2156 4956 2163 4993
rect 2176 4923 2183 4943
rect 2176 4916 2203 4923
rect 2016 4507 2023 4873
rect 2036 4507 2043 4693
rect 2076 4567 2083 4913
rect 2096 4696 2103 4813
rect 2116 4647 2123 4683
rect 2176 4676 2183 4713
rect 2196 4707 2203 4916
rect 2036 4476 2043 4493
rect 2076 4476 2083 4513
rect 2156 4507 2163 4663
rect 2196 4643 2203 4663
rect 2216 4647 2223 4683
rect 2176 4636 2203 4643
rect 2176 4547 2183 4636
rect 2236 4627 2243 4953
rect 2276 4727 2283 5143
rect 2336 5107 2343 5153
rect 2416 5127 2423 5413
rect 2436 5387 2443 5453
rect 2476 5167 2483 5413
rect 2496 5407 2503 5433
rect 2536 5416 2543 5453
rect 2576 5407 2583 5533
rect 2656 5436 2663 5653
rect 2696 5443 2703 5693
rect 2716 5607 2723 5916
rect 2816 5887 2823 5923
rect 2916 5887 2923 5913
rect 2936 5903 2943 5933
rect 2936 5896 2963 5903
rect 2996 5687 3003 5933
rect 3056 5916 3083 5923
rect 3076 5907 3083 5916
rect 3096 5847 3103 5993
rect 3116 5707 3123 5913
rect 3136 5887 3143 5903
rect 2816 5607 2823 5673
rect 2836 5587 2843 5653
rect 2896 5607 2903 5623
rect 2876 5587 2883 5603
rect 2696 5436 2723 5443
rect 2507 5396 2523 5403
rect 2676 5347 2683 5423
rect 2736 5347 2743 5423
rect 2776 5416 2783 5453
rect 2296 4956 2303 4993
rect 2316 4787 2323 4943
rect 2316 4707 2323 4773
rect 1996 4456 2003 4473
rect 2096 4456 2103 4473
rect 2016 4387 2023 4443
rect 2116 4387 2123 4493
rect 2136 4476 2163 4483
rect 2196 4476 2203 4613
rect 2256 4587 2263 4673
rect 2236 4476 2243 4513
rect 1976 4227 1983 4373
rect 1856 4183 1863 4213
rect 1996 4196 2003 4293
rect 2036 4247 2043 4353
rect 2056 4307 2063 4353
rect 1756 4167 1763 4183
rect 1796 4163 1803 4183
rect 1836 4176 1863 4183
rect 1796 4156 1813 4163
rect 1956 4163 1963 4183
rect 1956 4156 1983 4163
rect 1776 4027 1783 4153
rect 1756 3996 1763 4013
rect 1796 3996 1823 4003
rect 1376 3687 1383 3703
rect 1456 3696 1473 3703
rect 1356 3516 1363 3553
rect 1396 3516 1403 3553
rect 1436 3516 1443 3573
rect 1416 3487 1423 3503
rect 1356 3047 1363 3453
rect 1416 3347 1423 3473
rect 1456 3387 1463 3673
rect 1476 3527 1483 3673
rect 1516 3547 1523 3653
rect 1536 3647 1543 3893
rect 1776 3867 1783 3973
rect 1816 3967 1823 3996
rect 1836 3967 1843 4153
rect 1876 4067 1883 4153
rect 1896 3996 1903 4153
rect 1556 3667 1563 3813
rect 1596 3716 1603 3773
rect 1576 3643 1583 3703
rect 1556 3636 1583 3643
rect 1536 3516 1543 3553
rect 1476 3407 1483 3493
rect 1516 3407 1523 3473
rect 1456 3267 1463 3373
rect 1376 3107 1383 3253
rect 1416 3236 1423 3253
rect 1456 3236 1483 3243
rect 1396 3147 1403 3223
rect 1476 3147 1483 3236
rect 1496 3207 1503 3333
rect 1536 3327 1543 3473
rect 1556 3347 1563 3636
rect 1576 3516 1583 3533
rect 1596 3307 1603 3653
rect 1616 3587 1623 3753
rect 1656 3716 1663 3753
rect 1636 3687 1643 3703
rect 1676 3683 1683 3853
rect 1716 3716 1723 3813
rect 1756 3716 1763 3773
rect 1796 3727 1803 3773
rect 1836 3743 1843 3793
rect 1816 3736 1843 3743
rect 1776 3696 1803 3703
rect 1796 3687 1803 3696
rect 1676 3676 1703 3683
rect 1616 3367 1623 3553
rect 1676 3487 1683 3653
rect 1696 3627 1703 3676
rect 1756 3676 1773 3683
rect 1716 3536 1723 3673
rect 1756 3516 1763 3676
rect 1776 3527 1783 3553
rect 1796 3507 1803 3533
rect 1816 3527 1823 3736
rect 1856 3727 1863 3913
rect 1876 3903 1883 3983
rect 1916 3976 1923 4153
rect 1896 3927 1903 3953
rect 1936 3947 1943 4133
rect 1956 4047 1963 4113
rect 1976 4067 1983 4156
rect 1996 4087 2003 4133
rect 2016 4107 2023 4183
rect 2036 4147 2043 4173
rect 2056 4127 2063 4293
rect 2076 4107 2083 4273
rect 2096 4267 2103 4313
rect 2136 4307 2143 4476
rect 2176 4447 2183 4463
rect 2256 4443 2263 4473
rect 2236 4436 2263 4443
rect 2096 4216 2103 4233
rect 2136 4216 2143 4253
rect 2216 4227 2223 4373
rect 2236 4347 2243 4436
rect 2256 4287 2263 4413
rect 2256 4227 2263 4273
rect 2276 4267 2283 4693
rect 2336 4687 2343 4973
rect 2356 4956 2363 5093
rect 2416 4947 2423 5113
rect 2456 5107 2463 5123
rect 2476 4956 2483 5033
rect 2496 4887 2503 5143
rect 2516 4956 2523 5013
rect 2376 4627 2383 4733
rect 2396 4676 2403 4753
rect 2416 4547 2423 4633
rect 2376 4476 2383 4513
rect 2316 4447 2323 4463
rect 2356 4447 2363 4463
rect 2396 4447 2403 4533
rect 2416 4507 2423 4533
rect 2436 4456 2443 4593
rect 2456 4503 2463 4663
rect 2456 4496 2473 4503
rect 2496 4483 2503 4713
rect 2596 4707 2603 4963
rect 2616 4703 2623 5013
rect 2636 4987 2643 5333
rect 2676 5143 2683 5173
rect 2796 5167 2803 5433
rect 2816 5147 2823 5433
rect 2876 5156 2883 5193
rect 2916 5187 2923 5473
rect 2936 5436 2943 5473
rect 2936 5167 2943 5333
rect 2956 5187 2963 5453
rect 2976 5387 2983 5513
rect 3036 5407 3043 5633
rect 3056 5623 3063 5653
rect 3116 5647 3123 5693
rect 3136 5636 3143 5653
rect 3056 5616 3083 5623
rect 3076 5527 3083 5616
rect 3116 5567 3123 5603
rect 2656 5136 2683 5143
rect 2736 5136 2763 5143
rect 2756 5103 2763 5136
rect 2736 5096 2763 5103
rect 2736 4976 2743 5096
rect 2636 4956 2643 4973
rect 2616 4696 2643 4703
rect 2556 4656 2583 4663
rect 2476 4476 2503 4483
rect 2476 4467 2483 4476
rect 2556 4476 2563 4656
rect 2596 4487 2603 4673
rect 2636 4663 2643 4696
rect 2696 4667 2703 4793
rect 2616 4656 2643 4663
rect 2656 4496 2663 4653
rect 2716 4647 2723 4973
rect 2756 4687 2763 4943
rect 2776 4696 2783 4973
rect 2816 4956 2823 5113
rect 2896 4987 2903 5143
rect 2956 5107 2963 5123
rect 2976 5083 2983 5373
rect 3156 5347 3163 5693
rect 3176 5547 3183 5973
rect 3236 5927 3243 5953
rect 3216 5867 3223 5903
rect 3216 5587 3223 5643
rect 3276 5636 3283 5713
rect 3296 5707 3303 6153
rect 3416 6136 3443 6143
rect 3476 6136 3483 6153
rect 3356 6096 3383 6103
rect 3376 6027 3383 6096
rect 3336 5936 3343 6013
rect 3416 5947 3423 6136
rect 3456 6087 3463 6123
rect 3536 6116 3563 6123
rect 3596 6116 3603 6153
rect 3676 6136 3683 6153
rect 3716 6136 3723 6153
rect 3556 6083 3563 6116
rect 3556 6076 3583 6083
rect 3656 6007 3663 6093
rect 3756 6047 3763 6083
rect 3356 5907 3363 5933
rect 3416 5916 3443 5923
rect 3336 5643 3343 5853
rect 3316 5636 3343 5643
rect 3256 5607 3263 5623
rect 3316 5587 3323 5636
rect 3356 5623 3363 5653
rect 3436 5647 3443 5916
rect 3516 5916 3523 5993
rect 3816 5947 3823 6153
rect 3856 6096 3863 6153
rect 3936 6087 3943 6103
rect 3936 6067 3943 6073
rect 3576 5936 3623 5943
rect 3576 5867 3583 5936
rect 3616 5916 3623 5936
rect 3716 5936 3743 5943
rect 3596 5896 3603 5913
rect 3676 5907 3683 5933
rect 3736 5923 3743 5936
rect 3936 5927 3943 6053
rect 3736 5916 3763 5923
rect 3856 5916 3883 5923
rect 3696 5887 3703 5893
rect 3856 5867 3863 5916
rect 3596 5656 3623 5663
rect 3356 5616 3383 5623
rect 3016 5127 3023 5143
rect 3136 5143 3143 5173
rect 3136 5136 3163 5143
rect 2956 5076 2983 5083
rect 2956 4983 2963 5076
rect 2936 4976 2963 4983
rect 2896 4967 2903 4973
rect 2796 4703 2803 4953
rect 2896 4943 2903 4953
rect 2896 4936 2923 4943
rect 2956 4927 2963 4976
rect 3036 4956 3043 5123
rect 3156 4907 3163 4963
rect 2796 4696 2823 4703
rect 2736 4647 2743 4663
rect 2296 4327 2303 4373
rect 2296 4207 2303 4313
rect 2316 4227 2323 4433
rect 2016 4027 2023 4053
rect 1967 4016 2003 4023
rect 1916 3903 1923 3913
rect 1876 3896 1923 3903
rect 1916 3767 1923 3873
rect 1936 3827 1943 3893
rect 1956 3803 1963 3993
rect 1936 3796 1963 3803
rect 1896 3703 1903 3713
rect 1916 3707 1923 3753
rect 1936 3747 1943 3796
rect 1956 3727 1963 3753
rect 1976 3747 1983 3833
rect 1996 3763 2003 3973
rect 1996 3756 2023 3763
rect 1836 3647 1843 3703
rect 1876 3696 1903 3703
rect 1876 3643 1883 3696
rect 1936 3696 1963 3703
rect 1856 3636 1883 3643
rect 1856 3587 1863 3636
rect 1836 3536 1843 3553
rect 1856 3516 1863 3553
rect 1696 3407 1703 3503
rect 1736 3467 1743 3503
rect 1676 3327 1683 3393
rect 1576 3236 1583 3293
rect 1696 3247 1703 3333
rect 1716 3267 1723 3333
rect 1736 3267 1743 3353
rect 1596 3187 1603 3223
rect 1636 3207 1643 3223
rect 1656 3187 1663 3233
rect 1736 3223 1743 3253
rect 1716 3216 1743 3223
rect 1396 3087 1403 3113
rect 1396 3036 1403 3073
rect 1436 3036 1443 3053
rect 1476 3036 1483 3053
rect 1416 2947 1423 3033
rect 1316 2776 1343 2783
rect 1296 2727 1303 2773
rect 1256 2707 1263 2723
rect 1256 2647 1263 2693
rect 1136 2507 1143 2543
rect 1096 2327 1103 2393
rect 1056 2296 1073 2303
rect 1056 2276 1063 2296
rect 1116 2276 1123 2333
rect 1096 2127 1103 2273
rect 1136 2227 1143 2263
rect 1156 2207 1163 2353
rect 1196 2347 1203 2553
rect 1216 2467 1223 2543
rect 1116 2127 1123 2173
rect 1176 2163 1183 2293
rect 1196 2256 1203 2273
rect 1236 2227 1243 2513
rect 1256 2507 1263 2553
rect 1276 2507 1283 2543
rect 1256 2207 1263 2373
rect 1316 2303 1323 2776
rect 1336 2727 1343 2743
rect 1356 2627 1363 2693
rect 1376 2687 1383 2723
rect 1416 2707 1423 2893
rect 1416 2563 1423 2673
rect 1436 2607 1443 2973
rect 1456 2967 1463 3023
rect 1456 2787 1463 2813
rect 1476 2767 1483 2993
rect 1496 2987 1503 3023
rect 1536 3007 1543 3133
rect 1556 3007 1563 3033
rect 1516 2907 1523 2973
rect 1496 2727 1503 2833
rect 1596 2807 1603 3113
rect 1616 3036 1623 3053
rect 1656 3036 1683 3043
rect 1676 2987 1683 3036
rect 1696 2807 1703 3133
rect 1716 3127 1723 3216
rect 1756 3207 1763 3433
rect 1776 3287 1783 3493
rect 1836 3467 1843 3493
rect 1876 3467 1883 3613
rect 1896 3547 1903 3613
rect 1936 3563 1943 3673
rect 1956 3607 1963 3696
rect 1976 3607 1983 3693
rect 1956 3583 1963 3593
rect 1956 3576 1983 3583
rect 1936 3556 1963 3563
rect 1936 3516 1943 3533
rect 1796 3427 1803 3453
rect 1756 3027 1763 3113
rect 1776 2947 1783 3233
rect 1796 3227 1803 3373
rect 1816 3307 1823 3373
rect 1836 3247 1843 3453
rect 1956 3427 1963 3556
rect 1976 3447 1983 3576
rect 1996 3507 2003 3733
rect 2016 3561 2023 3756
rect 2036 3747 2043 4093
rect 2056 3996 2063 4073
rect 2076 4027 2083 4033
rect 2116 4027 2123 4193
rect 2136 4176 2163 4183
rect 2136 4107 2143 4176
rect 2236 4163 2243 4183
rect 2216 4156 2243 4163
rect 2136 4027 2143 4093
rect 2176 4047 2183 4153
rect 2196 4127 2203 4153
rect 2216 4127 2223 4156
rect 2256 4143 2263 4193
rect 2336 4187 2343 4333
rect 2287 4156 2303 4163
rect 2236 4136 2263 4143
rect 2096 3996 2123 4003
rect 2076 3847 2083 3973
rect 2116 3967 2123 3996
rect 2176 3996 2183 4033
rect 2216 4027 2223 4073
rect 2056 3716 2063 3793
rect 2116 3787 2123 3933
rect 2156 3907 2163 3983
rect 2076 3747 2083 3773
rect 2096 3716 2103 3773
rect 2196 3727 2203 3913
rect 2236 3887 2243 4136
rect 2316 4127 2323 4183
rect 2256 4067 2263 4073
rect 2256 4007 2263 4053
rect 2276 4027 2283 4053
rect 2316 4027 2323 4113
rect 2336 4067 2343 4173
rect 2356 4123 2363 4413
rect 2416 4127 2423 4183
rect 2436 4127 2443 4233
rect 2456 4216 2463 4433
rect 2476 4427 2483 4433
rect 2496 4407 2503 4453
rect 2536 4427 2543 4463
rect 2576 4443 2583 4463
rect 2636 4443 2643 4463
rect 2576 4436 2643 4443
rect 2656 4387 2663 4413
rect 2676 4387 2683 4473
rect 2496 4227 2503 4293
rect 2356 4116 2383 4123
rect 2276 4007 2283 4013
rect 2356 3996 2363 4093
rect 2216 3727 2223 3833
rect 2036 3587 2043 3703
rect 2076 3667 2083 3703
rect 2116 3696 2143 3703
rect 2176 3696 2203 3703
rect 2096 3516 2103 3553
rect 1876 3247 1883 3393
rect 1976 3367 1983 3413
rect 1796 2827 1803 3193
rect 1816 3187 1823 3223
rect 1876 3147 1883 3193
rect 1896 3147 1903 3353
rect 1996 3343 2003 3473
rect 2036 3467 2043 3503
rect 2056 3387 2063 3473
rect 1976 3336 2003 3343
rect 1936 3287 1943 3293
rect 1936 3236 1943 3273
rect 1976 3236 1983 3336
rect 1916 3207 1923 3233
rect 2016 3227 2023 3373
rect 1816 3067 1823 3093
rect 1836 3007 1843 3023
rect 1856 2927 1863 3073
rect 1716 2787 1723 2813
rect 1576 2776 1603 2783
rect 1516 2687 1523 2763
rect 1536 2727 1543 2773
rect 1556 2707 1563 2763
rect 1596 2747 1603 2776
rect 1616 2776 1643 2783
rect 1516 2567 1523 2613
rect 1356 2556 1383 2563
rect 1416 2556 1443 2563
rect 1356 2547 1363 2556
rect 1296 2296 1323 2303
rect 1276 2247 1283 2263
rect 1156 2156 1183 2163
rect 1156 2143 1163 2156
rect 1136 2136 1163 2143
rect 1036 2043 1043 2063
rect 1016 2036 1043 2043
rect 876 1796 883 1853
rect 896 1727 903 1773
rect 916 1747 923 1813
rect 936 1796 943 1993
rect 956 1767 963 1783
rect 876 1607 883 1613
rect 816 1596 843 1603
rect 916 1596 923 1693
rect 936 1643 943 1693
rect 956 1687 963 1753
rect 976 1667 983 2013
rect 996 1847 1003 2013
rect 1016 1927 1023 2036
rect 1036 1787 1043 1973
rect 1076 1823 1083 2093
rect 1136 1847 1143 2136
rect 1156 1967 1163 2113
rect 1136 1827 1143 1833
rect 1056 1816 1083 1823
rect 1056 1707 1063 1816
rect 1076 1663 1083 1733
rect 1096 1707 1103 1753
rect 1116 1727 1123 1783
rect 1176 1763 1183 1953
rect 1156 1756 1183 1763
rect 1056 1656 1083 1663
rect 936 1636 963 1643
rect 856 1547 863 1583
rect 736 1336 763 1343
rect 736 1167 743 1336
rect 816 1316 823 1533
rect 756 1287 763 1303
rect 756 1187 763 1273
rect 836 1267 843 1513
rect 856 1407 863 1453
rect 876 1363 883 1493
rect 896 1447 903 1573
rect 936 1367 943 1613
rect 956 1587 963 1636
rect 1016 1596 1023 1613
rect 1056 1596 1063 1656
rect 1076 1603 1083 1633
rect 1076 1596 1103 1603
rect 996 1567 1003 1583
rect 1036 1563 1043 1583
rect 1036 1556 1063 1563
rect 1056 1547 1063 1556
rect 876 1356 903 1363
rect 876 1316 883 1333
rect 896 1287 903 1356
rect 936 1316 943 1333
rect 976 1316 983 1353
rect 896 1187 903 1273
rect 916 1207 923 1303
rect 956 1247 963 1303
rect 296 547 303 673
rect 256 376 273 383
rect 236 343 243 373
rect 276 356 283 373
rect 236 336 263 343
rect 316 207 323 233
rect 216 147 223 163
rect 316 136 323 193
rect 336 167 343 573
rect 356 567 363 603
rect 356 307 363 473
rect 376 367 383 693
rect 416 636 423 653
rect 456 636 463 693
rect 476 687 483 953
rect 516 836 523 853
rect 536 843 543 933
rect 576 867 583 1093
rect 536 836 563 843
rect 476 636 483 673
rect 516 636 523 653
rect 536 547 543 773
rect 576 663 583 833
rect 596 807 603 1113
rect 616 847 623 1073
rect 656 1047 663 1073
rect 656 823 663 1033
rect 636 816 663 823
rect 556 656 583 663
rect 556 627 563 656
rect 616 636 623 693
rect 636 647 643 673
rect 656 627 663 816
rect 676 667 683 1113
rect 756 1087 763 1133
rect 856 1116 863 1133
rect 916 1116 923 1133
rect 736 927 743 1083
rect 776 887 783 1113
rect 836 1087 843 1103
rect 716 836 723 853
rect 696 787 703 823
rect 736 687 743 823
rect 596 587 603 623
rect 416 387 423 513
rect 416 356 423 373
rect 456 343 463 533
rect 396 307 403 323
rect 416 156 423 213
rect 436 207 443 343
rect 456 336 483 343
rect 476 267 483 336
rect 516 327 523 343
rect 536 327 543 533
rect 556 343 563 453
rect 616 447 623 593
rect 656 383 663 593
rect 676 467 683 653
rect 716 616 723 653
rect 756 647 763 713
rect 696 567 703 603
rect 756 487 763 633
rect 776 587 783 853
rect 796 647 803 893
rect 856 823 863 873
rect 896 867 903 1103
rect 936 1096 963 1103
rect 856 816 883 823
rect 916 767 923 823
rect 936 747 943 853
rect 956 847 963 1096
rect 976 987 983 1113
rect 996 1107 1003 1273
rect 1016 1116 1023 1333
rect 1036 1287 1043 1533
rect 1136 1527 1143 1693
rect 1156 1687 1163 1756
rect 1176 1603 1183 1733
rect 1196 1707 1203 2193
rect 1216 2076 1223 2133
rect 1216 1827 1223 2033
rect 1256 1927 1263 1993
rect 1256 1763 1263 1913
rect 1236 1756 1263 1763
rect 1156 1596 1183 1603
rect 1056 1327 1063 1353
rect 1076 1207 1083 1293
rect 1116 1287 1123 1303
rect 956 787 963 833
rect 996 816 1003 913
rect 1056 767 1063 1133
rect 1096 863 1103 1093
rect 1076 856 1103 863
rect 1076 836 1083 856
rect 1096 803 1103 823
rect 1076 796 1103 803
rect 836 636 843 673
rect 816 427 823 623
rect 856 616 863 653
rect 976 636 1003 643
rect 876 567 883 633
rect 956 607 963 623
rect 636 376 663 383
rect 636 347 643 376
rect 676 356 683 413
rect 556 336 583 343
rect 616 327 623 333
rect 336 127 343 153
rect 376 136 403 143
rect 376 107 383 136
rect 436 123 443 143
rect 476 123 483 193
rect 496 167 503 323
rect 536 136 543 233
rect 556 127 563 313
rect 596 307 603 323
rect 656 307 663 353
rect 856 347 863 453
rect 876 376 883 433
rect 696 307 703 323
rect 676 156 683 213
rect 696 167 703 293
rect 716 156 723 173
rect 756 167 763 343
rect 976 307 983 636
rect 1036 487 1043 673
rect 1056 627 1063 673
rect 1076 607 1083 796
rect 1116 667 1123 1113
rect 1136 1107 1143 1413
rect 1156 1247 1163 1596
rect 1176 1307 1183 1433
rect 1176 1123 1183 1153
rect 1196 1143 1203 1613
rect 1236 1367 1243 1756
rect 1276 1743 1283 2213
rect 1296 2147 1303 2296
rect 1336 2187 1343 2433
rect 1376 2267 1383 2333
rect 1396 2183 1403 2393
rect 1436 2287 1443 2303
rect 1496 2287 1503 2513
rect 1536 2383 1543 2693
rect 1556 2556 1563 2573
rect 1576 2487 1583 2733
rect 1616 2587 1623 2776
rect 1656 2747 1663 2763
rect 1696 2727 1703 2763
rect 1756 2747 1763 2783
rect 1796 2776 1803 2793
rect 1516 2376 1543 2383
rect 1376 2176 1403 2183
rect 1296 1767 1303 2113
rect 1316 1847 1323 1953
rect 1316 1796 1323 1833
rect 1336 1827 1343 2073
rect 1336 1747 1343 1773
rect 1276 1736 1303 1743
rect 1296 1727 1303 1736
rect 1236 1347 1243 1353
rect 1236 1303 1243 1333
rect 1216 1296 1243 1303
rect 1256 1247 1263 1303
rect 1276 1287 1283 1713
rect 1296 1467 1303 1693
rect 1316 1367 1323 1673
rect 1356 1627 1363 2133
rect 1376 1987 1383 2176
rect 1396 2087 1403 2153
rect 1416 2127 1423 2273
rect 1456 2267 1463 2283
rect 1456 2207 1463 2213
rect 1496 2207 1503 2273
rect 1516 2267 1523 2376
rect 1536 2296 1543 2333
rect 1576 2267 1583 2303
rect 1436 2076 1443 2113
rect 1376 1796 1383 1833
rect 1396 1823 1403 2033
rect 1416 1887 1423 2063
rect 1456 2056 1463 2193
rect 1596 2187 1603 2283
rect 1616 2247 1623 2553
rect 1636 2387 1643 2613
rect 1656 2507 1663 2633
rect 1676 2387 1683 2563
rect 1716 2427 1723 2573
rect 1736 2527 1743 2733
rect 1776 2507 1783 2753
rect 1816 2647 1823 2853
rect 1836 2807 1843 2913
rect 1876 2887 1883 3113
rect 1896 3036 1903 3133
rect 1956 3127 1963 3203
rect 1936 3036 1943 3073
rect 1996 3067 2003 3223
rect 2036 3223 2043 3373
rect 2076 3347 2083 3413
rect 2076 3236 2083 3333
rect 2096 3327 2103 3473
rect 2116 3327 2123 3673
rect 2136 3647 2143 3696
rect 2196 3687 2203 3696
rect 2156 3607 2163 3683
rect 2176 3667 2183 3673
rect 2236 3647 2243 3703
rect 2096 3287 2103 3313
rect 2136 3267 2143 3593
rect 2156 3516 2163 3553
rect 2176 3536 2183 3613
rect 2196 3547 2203 3573
rect 2196 3516 2203 3533
rect 2216 3527 2223 3593
rect 2236 3527 2243 3553
rect 2256 3547 2263 3973
rect 2296 3967 2303 3983
rect 2296 3887 2303 3953
rect 2336 3927 2343 3953
rect 2296 3747 2303 3773
rect 2336 3743 2343 3833
rect 2376 3747 2383 4116
rect 2416 4067 2423 4113
rect 2476 4087 2483 4173
rect 2496 4087 2503 4133
rect 2396 4007 2403 4013
rect 2476 3996 2483 4073
rect 2496 3987 2503 4013
rect 2396 3867 2403 3933
rect 2416 3907 2423 3983
rect 2416 3827 2423 3893
rect 2436 3843 2443 3893
rect 2456 3887 2463 3973
rect 2496 3927 2503 3953
rect 2476 3883 2483 3913
rect 2476 3876 2503 3883
rect 2436 3836 2463 3843
rect 2396 3787 2403 3813
rect 2316 3736 2343 3743
rect 2276 3716 2283 3733
rect 2236 3496 2243 3513
rect 2156 3263 2163 3313
rect 2176 3307 2183 3493
rect 2276 3483 2283 3653
rect 2296 3647 2303 3713
rect 2316 3587 2323 3736
rect 2396 3703 2403 3773
rect 2416 3727 2423 3733
rect 2376 3696 2403 3703
rect 2336 3643 2343 3673
rect 2356 3667 2363 3693
rect 2336 3636 2363 3643
rect 2356 3627 2363 3636
rect 2336 3543 2343 3613
rect 2336 3536 2363 3543
rect 2216 3463 2223 3483
rect 2216 3456 2243 3463
rect 2196 3307 2203 3453
rect 2236 3347 2243 3456
rect 2256 3447 2263 3483
rect 2276 3476 2303 3483
rect 2156 3256 2183 3263
rect 2176 3247 2183 3256
rect 2036 3216 2063 3223
rect 2056 3167 2063 3216
rect 1956 3036 1963 3053
rect 2016 3016 2043 3023
rect 2036 3007 2043 3016
rect 1836 2687 1843 2773
rect 1856 2747 1863 2793
rect 1876 2776 1883 2793
rect 1916 2787 1923 2933
rect 1796 2603 1803 2633
rect 1856 2607 1863 2733
rect 1896 2727 1903 2763
rect 1936 2707 1943 2773
rect 1956 2756 1963 2853
rect 2036 2827 2043 2833
rect 1796 2596 1823 2603
rect 1816 2587 1823 2596
rect 1796 2556 1803 2573
rect 1876 2563 1883 2673
rect 1896 2587 1903 2653
rect 1856 2556 1883 2563
rect 1676 2327 1683 2373
rect 1656 2207 1663 2303
rect 1576 2076 1583 2093
rect 1396 1816 1423 1823
rect 1396 1767 1403 1783
rect 1416 1707 1423 1816
rect 1436 1796 1443 1993
rect 1476 1947 1483 2073
rect 1496 1987 1503 2063
rect 1476 1783 1483 1853
rect 1496 1796 1503 1953
rect 1516 1827 1523 1873
rect 1456 1776 1483 1783
rect 1516 1767 1523 1783
rect 1336 1467 1343 1563
rect 1376 1547 1383 1563
rect 1336 1447 1343 1453
rect 1356 1447 1363 1533
rect 1376 1316 1383 1333
rect 1296 1287 1303 1303
rect 1396 1247 1403 1633
rect 1416 1607 1423 1613
rect 1476 1603 1483 1753
rect 1536 1627 1543 2033
rect 1596 1987 1603 2113
rect 1556 1827 1563 1933
rect 1576 1867 1583 1913
rect 1576 1827 1583 1853
rect 1596 1767 1603 1833
rect 1616 1827 1623 2133
rect 1636 2067 1643 2113
rect 1696 2096 1703 2153
rect 1716 2107 1723 2313
rect 1656 2023 1663 2093
rect 1696 2027 1703 2053
rect 1656 2016 1683 2023
rect 1476 1596 1503 1603
rect 1496 1467 1503 1596
rect 1596 1596 1603 1653
rect 1636 1583 1643 1753
rect 1656 1747 1663 1813
rect 1676 1787 1683 2016
rect 1696 1927 1703 2013
rect 1736 2007 1743 2453
rect 1756 2267 1763 2473
rect 1776 2296 1783 2433
rect 1796 2327 1803 2513
rect 1816 2323 1823 2553
rect 1856 2467 1863 2556
rect 1916 2547 1923 2673
rect 1936 2547 1943 2693
rect 1876 2536 1903 2543
rect 1816 2316 1843 2323
rect 1796 2187 1803 2283
rect 1756 2076 1763 2153
rect 1796 2076 1803 2153
rect 1816 2107 1823 2213
rect 1836 2147 1843 2316
rect 1856 2307 1863 2453
rect 1876 2387 1883 2536
rect 1876 2227 1883 2353
rect 1896 2347 1903 2493
rect 1916 2407 1923 2433
rect 1976 2387 1983 2713
rect 1996 2687 2003 2813
rect 2036 2727 2043 2813
rect 2056 2767 2063 3153
rect 2076 2863 2083 3133
rect 2096 3043 2103 3073
rect 2116 3063 2123 3133
rect 2136 3087 2143 3233
rect 2216 3223 2223 3333
rect 2156 3167 2163 3223
rect 2196 3216 2223 3223
rect 2196 3127 2203 3216
rect 2116 3056 2143 3063
rect 2096 3036 2123 3043
rect 2116 3027 2123 3036
rect 2136 2996 2143 3056
rect 2076 2856 2103 2863
rect 2076 2727 2083 2743
rect 2047 2716 2063 2723
rect 1996 2367 2003 2653
rect 2016 2367 2023 2533
rect 2036 2507 2043 2673
rect 2096 2567 2103 2856
rect 2116 2787 2123 2933
rect 2116 2756 2123 2773
rect 2136 2763 2143 2873
rect 2156 2807 2163 2833
rect 2176 2827 2183 3113
rect 2196 2987 2203 3073
rect 2196 2827 2203 2893
rect 2136 2756 2163 2763
rect 2156 2607 2163 2693
rect 2176 2687 2183 2783
rect 2216 2776 2223 2893
rect 2236 2867 2243 3293
rect 2276 3287 2283 3353
rect 2296 3327 2303 3476
rect 2316 3283 2323 3493
rect 2356 3387 2363 3536
rect 2376 3527 2383 3696
rect 2436 3687 2443 3813
rect 2456 3767 2463 3836
rect 2476 3747 2483 3853
rect 2496 3823 2503 3876
rect 2516 3867 2523 4313
rect 2696 4267 2703 4573
rect 2756 4527 2763 4653
rect 2736 4307 2743 4513
rect 2756 4327 2763 4453
rect 2776 4327 2783 4613
rect 2796 4587 2803 4663
rect 2796 4496 2803 4513
rect 2816 4507 2823 4696
rect 2836 4467 2843 4493
rect 2816 4407 2823 4463
rect 2536 3847 2543 4253
rect 2716 4227 2723 4253
rect 2616 4216 2643 4223
rect 2556 4167 2563 4193
rect 2616 4187 2623 4216
rect 2716 4207 2723 4213
rect 2696 4187 2703 4203
rect 2596 4147 2603 4163
rect 2556 3967 2563 4093
rect 2596 3976 2603 4053
rect 2556 3887 2563 3933
rect 2576 3863 2583 3963
rect 2556 3856 2583 3863
rect 2556 3823 2563 3856
rect 2496 3816 2523 3823
rect 2496 3767 2503 3793
rect 2516 3743 2523 3816
rect 2536 3816 2563 3823
rect 2536 3787 2543 3816
rect 2556 3747 2563 3773
rect 2496 3736 2523 3743
rect 2456 3716 2483 3723
rect 2396 3567 2403 3653
rect 2396 3496 2403 3533
rect 2416 3407 2423 3483
rect 2436 3427 2443 3613
rect 2456 3487 2463 3673
rect 2476 3667 2483 3716
rect 2476 3547 2483 3593
rect 2496 3547 2503 3736
rect 2516 3503 2523 3713
rect 2536 3527 2543 3653
rect 2556 3627 2563 3683
rect 2556 3547 2563 3553
rect 2496 3496 2523 3503
rect 2556 3487 2563 3513
rect 2336 3307 2343 3333
rect 2456 3323 2463 3473
rect 2476 3467 2483 3483
rect 2536 3447 2543 3453
rect 2436 3316 2463 3323
rect 2316 3276 2343 3283
rect 2256 3167 2263 3273
rect 2276 3256 2283 3273
rect 2256 3067 2263 3093
rect 2276 2927 2283 3213
rect 2336 3187 2343 3276
rect 2396 3236 2403 3293
rect 2356 3187 2363 3213
rect 2376 3207 2383 3223
rect 2336 3123 2343 3173
rect 2316 3116 2343 3123
rect 2296 3036 2303 3073
rect 2296 2807 2303 2993
rect 2316 2847 2323 3116
rect 2376 3027 2383 3033
rect 2196 2747 2203 2763
rect 2196 2607 2203 2733
rect 2216 2583 2223 2673
rect 2236 2627 2243 2793
rect 2316 2776 2323 2813
rect 2356 2787 2363 2893
rect 2396 2823 2403 3173
rect 2436 3107 2443 3316
rect 2456 3236 2463 3293
rect 2476 3267 2483 3373
rect 2556 3367 2563 3473
rect 2496 3227 2503 3273
rect 2516 3203 2523 3313
rect 2556 3236 2563 3293
rect 2576 3207 2583 3813
rect 2616 3807 2623 3933
rect 2596 3736 2603 3793
rect 2636 3787 2643 4013
rect 2656 3863 2663 4153
rect 2736 4063 2743 4253
rect 2816 4216 2823 4333
rect 2836 4307 2843 4353
rect 2756 4187 2763 4203
rect 2776 4187 2783 4213
rect 2756 4147 2763 4173
rect 2776 4067 2783 4133
rect 2716 4056 2743 4063
rect 2676 4027 2683 4053
rect 2716 4007 2723 4056
rect 2676 3947 2683 3963
rect 2716 3927 2723 3933
rect 2676 3896 2723 3903
rect 2676 3887 2683 3896
rect 2656 3856 2683 3863
rect 2656 3767 2663 3833
rect 2676 3787 2683 3856
rect 2696 3763 2703 3873
rect 2716 3767 2723 3896
rect 2736 3887 2743 4033
rect 2756 3987 2763 4033
rect 2816 4027 2823 4073
rect 2796 3976 2803 4013
rect 2756 3803 2763 3953
rect 2816 3947 2823 3963
rect 2776 3887 2783 3933
rect 2796 3907 2803 3933
rect 2836 3907 2843 4233
rect 2856 4227 2863 4513
rect 2876 4487 2883 4893
rect 2936 4696 2943 4713
rect 2996 4696 3023 4703
rect 2916 4507 2923 4683
rect 2956 4663 2963 4693
rect 2956 4656 2983 4663
rect 2956 4647 2963 4656
rect 2996 4647 3003 4696
rect 3076 4667 3083 4853
rect 3036 4527 3043 4663
rect 3096 4663 3103 4893
rect 3176 4807 3183 5173
rect 3196 5127 3203 5143
rect 3216 4847 3223 5133
rect 3236 5107 3243 5573
rect 3356 5567 3363 5616
rect 3436 5607 3443 5633
rect 3256 5436 3263 5473
rect 3296 5147 3303 5533
rect 3456 5487 3463 5623
rect 3596 5483 3603 5656
rect 3596 5476 3623 5483
rect 3336 5407 3343 5443
rect 3456 5436 3483 5443
rect 3496 5436 3503 5473
rect 3316 5207 3323 5273
rect 3396 5176 3403 5193
rect 3476 5147 3483 5436
rect 3516 5143 3523 5473
rect 3596 5443 3603 5453
rect 3576 5436 3603 5443
rect 3576 5167 3583 5413
rect 3616 5247 3623 5476
rect 3676 5467 3683 5833
rect 3696 5667 3703 5753
rect 3696 5607 3703 5653
rect 3756 5636 3763 5673
rect 3776 5607 3783 5623
rect 3936 5623 3943 5913
rect 3996 5847 4003 5883
rect 3916 5616 3943 5623
rect 3996 5616 4003 5633
rect 3776 5436 3783 5593
rect 3236 4956 3243 4973
rect 3276 4963 3283 5073
rect 3276 4956 3303 4963
rect 3296 4787 3303 4956
rect 3316 4727 3323 4963
rect 3176 4663 3183 4693
rect 3096 4656 3123 4663
rect 3156 4656 3183 4663
rect 3196 4647 3203 4713
rect 3216 4676 3223 4693
rect 3256 4627 3263 4663
rect 2916 4476 2963 4483
rect 2876 4207 2883 4353
rect 2856 4107 2863 4183
rect 2876 4067 2883 4163
rect 2896 4147 2903 4183
rect 2916 4167 2923 4433
rect 2956 4267 2963 4476
rect 2956 4247 2963 4253
rect 2976 4207 2983 4443
rect 3036 4363 3043 4493
rect 3076 4483 3083 4613
rect 3067 4476 3083 4483
rect 3116 4476 3123 4493
rect 3056 4447 3063 4473
rect 3016 4356 3043 4363
rect 2856 3947 2863 3963
rect 2916 3947 2923 4053
rect 2936 4043 2943 4193
rect 2996 4167 3003 4183
rect 2976 4047 2983 4153
rect 3016 4147 3023 4356
rect 3036 4087 3043 4333
rect 3076 4267 3083 4413
rect 3096 4407 3103 4463
rect 3156 4427 3163 4533
rect 3096 4216 3103 4233
rect 3076 4187 3083 4203
rect 3116 4147 3123 4353
rect 2936 4036 2963 4043
rect 2936 3887 2943 4013
rect 2756 3796 2783 3803
rect 2756 3767 2763 3773
rect 2676 3756 2703 3763
rect 2636 3667 2643 3713
rect 2656 3707 2663 3723
rect 2596 3287 2603 3653
rect 2636 3536 2643 3573
rect 2616 3467 2623 3493
rect 2616 3407 2623 3453
rect 2636 3427 2643 3473
rect 2656 3327 2663 3613
rect 2676 3507 2683 3756
rect 2776 3747 2783 3796
rect 2856 3747 2863 3853
rect 2736 3707 2743 3733
rect 2936 3727 2943 3833
rect 2676 3427 2683 3473
rect 2616 3247 2623 3313
rect 2476 3187 2483 3203
rect 2516 3196 2543 3203
rect 2476 3047 2483 3173
rect 2536 3087 2543 3196
rect 2596 3187 2603 3223
rect 2436 2827 2443 3043
rect 2516 3036 2523 3073
rect 2536 3007 2543 3073
rect 2556 3036 2563 3133
rect 2396 2816 2423 2823
rect 2416 2807 2423 2816
rect 2436 2776 2463 2783
rect 2256 2727 2263 2753
rect 2336 2723 2343 2773
rect 2456 2747 2463 2776
rect 2316 2716 2343 2723
rect 2216 2576 2243 2583
rect 2196 2527 2203 2553
rect 2036 2407 2043 2493
rect 2056 2427 2063 2523
rect 2136 2503 2143 2523
rect 2176 2507 2183 2523
rect 2236 2516 2243 2576
rect 2256 2547 2263 2593
rect 2316 2567 2323 2716
rect 2296 2523 2303 2553
rect 2276 2516 2303 2523
rect 2136 2496 2163 2503
rect 1896 2287 1903 2333
rect 2056 2287 2063 2373
rect 2156 2347 2163 2496
rect 2176 2467 2183 2493
rect 2136 2296 2143 2333
rect 1856 2147 1863 2193
rect 1756 1847 1763 2033
rect 1776 1987 1783 2063
rect 1656 1596 1663 1673
rect 1696 1647 1703 1833
rect 1796 1827 1803 2033
rect 1816 1987 1823 2063
rect 1736 1796 1763 1803
rect 1796 1796 1803 1813
rect 1716 1587 1723 1613
rect 1616 1576 1643 1583
rect 1616 1567 1623 1576
rect 1416 1307 1423 1313
rect 1236 1147 1243 1233
rect 1196 1136 1223 1143
rect 1176 1116 1203 1123
rect 1136 836 1143 1053
rect 1216 1007 1223 1136
rect 1236 1116 1243 1133
rect 1196 767 1203 823
rect 1156 643 1163 693
rect 1136 636 1163 643
rect 996 376 1003 433
rect 1036 376 1063 383
rect 816 163 823 293
rect 1056 287 1063 376
rect 1096 307 1103 323
rect 1116 247 1123 343
rect 796 156 823 163
rect 576 136 583 153
rect 436 116 483 123
rect 516 107 523 123
rect 856 107 863 233
rect 956 156 963 173
rect 1136 147 1143 636
rect 1196 623 1203 673
rect 1176 616 1203 623
rect 1216 467 1223 933
rect 1236 727 1243 823
rect 1256 767 1263 1233
rect 1456 1147 1463 1353
rect 1496 1147 1503 1303
rect 1516 1247 1523 1293
rect 1536 1247 1543 1303
rect 1336 1136 1363 1143
rect 1336 1123 1343 1136
rect 1316 1116 1343 1123
rect 1316 887 1323 1116
rect 1416 947 1423 1133
rect 1436 1116 1463 1123
rect 1436 1107 1443 1116
rect 1536 1116 1543 1173
rect 1436 1047 1443 1093
rect 1476 947 1483 1103
rect 1416 907 1423 933
rect 1396 887 1403 893
rect 1276 827 1283 873
rect 1236 687 1243 713
rect 1296 687 1303 823
rect 1336 727 1343 833
rect 1376 767 1383 793
rect 1356 707 1363 753
rect 1236 603 1243 633
rect 1276 616 1283 653
rect 1296 647 1303 673
rect 1316 656 1323 693
rect 1396 663 1403 873
rect 1416 856 1443 863
rect 1476 856 1483 873
rect 1416 687 1423 856
rect 1496 687 1503 1073
rect 1556 1067 1563 1253
rect 1576 1127 1583 1193
rect 1596 1147 1603 1473
rect 1616 1227 1623 1373
rect 1676 1367 1683 1573
rect 1736 1387 1743 1733
rect 1756 1667 1763 1796
rect 1816 1767 1823 1933
rect 1896 1887 1903 2253
rect 1936 2207 1943 2283
rect 1976 2276 2003 2283
rect 1996 2263 2003 2276
rect 1996 2256 2043 2263
rect 1916 1967 1923 2173
rect 1936 1887 1943 2093
rect 1956 1927 1963 1953
rect 1976 1903 1983 2233
rect 2036 2227 2043 2256
rect 2056 2183 2063 2253
rect 2076 2207 2083 2283
rect 2096 2207 2103 2253
rect 2136 2183 2143 2193
rect 2056 2176 2143 2183
rect 1996 2076 2003 2153
rect 2036 2076 2043 2093
rect 1996 1927 2003 1993
rect 1956 1896 1983 1903
rect 1776 1596 1783 1733
rect 1796 1667 1803 1713
rect 1836 1627 1843 1813
rect 1856 1796 1863 1853
rect 1876 1727 1883 1783
rect 1896 1727 1903 1853
rect 1936 1767 1943 1783
rect 1936 1643 1943 1753
rect 1916 1636 1943 1643
rect 1916 1616 1923 1636
rect 1856 1596 1883 1603
rect 1656 1316 1663 1333
rect 1676 1296 1693 1303
rect 1616 1116 1623 1153
rect 1656 1116 1663 1253
rect 1716 1187 1723 1333
rect 1756 1323 1763 1593
rect 1876 1583 1883 1596
rect 1836 1567 1843 1583
rect 1876 1576 1903 1583
rect 1816 1527 1823 1553
rect 1836 1507 1843 1553
rect 1936 1467 1943 1613
rect 1956 1487 1963 1896
rect 2016 1867 2023 2073
rect 2056 1987 2063 2133
rect 2076 1963 2083 2153
rect 2136 2027 2143 2133
rect 2116 1963 2123 1993
rect 2056 1956 2083 1963
rect 2096 1956 2123 1963
rect 2056 1867 2063 1956
rect 2036 1787 2043 1803
rect 1976 1707 1983 1783
rect 2016 1747 2023 1783
rect 1996 1647 2003 1673
rect 2036 1607 2043 1753
rect 2056 1747 2063 1813
rect 2076 1703 2083 1873
rect 2056 1696 2083 1703
rect 2056 1596 2063 1696
rect 1936 1427 1943 1453
rect 1976 1447 1983 1473
rect 1736 1316 1763 1323
rect 1736 1207 1743 1316
rect 1776 1307 1783 1333
rect 1816 1316 1823 1333
rect 1856 1327 1863 1393
rect 1756 1267 1763 1293
rect 1796 1283 1803 1303
rect 1796 1276 1823 1283
rect 1696 1163 1703 1173
rect 1696 1156 1743 1163
rect 1676 1116 1683 1153
rect 1707 1136 1723 1143
rect 1716 1116 1723 1136
rect 1736 1127 1743 1156
rect 1576 1096 1603 1103
rect 1516 747 1523 1053
rect 1576 947 1583 1096
rect 1536 836 1543 893
rect 1576 836 1583 893
rect 1616 847 1623 1073
rect 1636 1067 1643 1103
rect 1696 1047 1703 1103
rect 1756 1067 1763 1173
rect 1816 1136 1823 1276
rect 1836 1247 1843 1303
rect 1776 1123 1783 1133
rect 1776 1116 1803 1123
rect 1856 1087 1863 1273
rect 1896 1267 1903 1283
rect 1936 1143 1943 1373
rect 1956 1287 1963 1303
rect 1956 1167 1963 1253
rect 1976 1187 1983 1273
rect 1936 1136 1963 1143
rect 1876 1116 1903 1123
rect 1756 987 1763 1053
rect 1736 847 1743 973
rect 1776 907 1783 933
rect 1556 747 1563 803
rect 1656 803 1663 843
rect 1716 807 1723 823
rect 1656 796 1683 803
rect 1516 667 1523 733
rect 1376 656 1403 663
rect 1376 643 1383 656
rect 1356 636 1383 643
rect 1236 596 1263 603
rect 1236 387 1243 596
rect 1156 307 1163 333
rect 1176 227 1183 343
rect 1156 156 1163 193
rect 1196 156 1203 173
rect 1236 167 1243 373
rect 1256 347 1263 433
rect 1316 387 1323 613
rect 1356 607 1363 636
rect 1436 616 1443 653
rect 1556 636 1563 653
rect 1316 327 1323 343
rect 1296 307 1303 323
rect 1336 307 1343 413
rect 1356 187 1363 373
rect 1436 347 1443 533
rect 1456 507 1463 633
rect 1476 616 1503 623
rect 1476 387 1483 616
rect 1536 587 1543 623
rect 1496 407 1503 573
rect 1516 383 1523 573
rect 1576 547 1583 793
rect 1636 636 1653 643
rect 1616 567 1623 623
rect 1676 607 1683 796
rect 1696 627 1703 773
rect 1716 707 1723 773
rect 1736 747 1743 833
rect 1736 616 1743 653
rect 1756 627 1763 893
rect 1836 823 1843 933
rect 1816 816 1843 823
rect 1776 616 1783 733
rect 1796 587 1803 633
rect 1816 607 1823 816
rect 1856 707 1863 1073
rect 1876 967 1883 1116
rect 1936 867 1943 1033
rect 1956 947 1963 1136
rect 1976 1083 1983 1173
rect 1996 1147 2003 1233
rect 2016 1096 2023 1323
rect 2036 1267 2043 1453
rect 2076 1347 2083 1653
rect 2096 1307 2103 1956
rect 2156 1947 2163 2313
rect 2176 2287 2183 2353
rect 2256 2267 2263 2283
rect 2176 2147 2183 2253
rect 2207 2196 2223 2203
rect 2196 2076 2203 2153
rect 2176 2047 2183 2063
rect 2176 1927 2183 2033
rect 2116 1707 2123 1873
rect 2216 1867 2223 2196
rect 2236 2147 2243 2253
rect 2256 2167 2263 2253
rect 2256 2076 2263 2113
rect 2276 2087 2283 2453
rect 2316 2407 2323 2513
rect 2296 2307 2303 2393
rect 2336 2387 2343 2633
rect 2376 2576 2383 2633
rect 2396 2527 2403 2533
rect 2156 1796 2163 1853
rect 2136 1767 2143 1783
rect 2156 1343 2163 1693
rect 2176 1547 2183 1833
rect 2216 1796 2223 1813
rect 2196 1763 2203 1783
rect 2196 1756 2223 1763
rect 2196 1507 2203 1733
rect 2216 1727 2223 1756
rect 2236 1667 2243 1783
rect 2256 1723 2263 1773
rect 2276 1747 2283 1783
rect 2296 1767 2303 2153
rect 2316 1847 2323 2133
rect 2336 1987 2343 2353
rect 2356 2167 2363 2473
rect 2376 2307 2383 2493
rect 2436 2487 2443 2633
rect 2456 2587 2463 2693
rect 2476 2643 2483 2773
rect 2496 2667 2503 2993
rect 2516 2807 2523 2933
rect 2576 2807 2583 3153
rect 2616 3087 2623 3193
rect 2476 2636 2503 2643
rect 2476 2587 2483 2613
rect 2456 2487 2463 2553
rect 2376 2227 2383 2263
rect 2396 2247 2403 2413
rect 2456 2407 2463 2433
rect 2416 2307 2423 2393
rect 2436 2263 2443 2333
rect 2476 2327 2483 2573
rect 2496 2347 2503 2636
rect 2516 2607 2523 2713
rect 2556 2687 2563 2783
rect 2556 2607 2563 2673
rect 2596 2663 2603 2893
rect 2576 2656 2603 2663
rect 2576 2627 2583 2656
rect 2616 2643 2623 3053
rect 2636 3007 2643 3253
rect 2656 3207 2663 3223
rect 2656 3047 2663 3173
rect 2676 3087 2683 3273
rect 2696 3267 2703 3573
rect 2716 3567 2723 3653
rect 2736 3527 2743 3653
rect 2756 3627 2763 3723
rect 2756 3527 2763 3593
rect 2736 3496 2743 3513
rect 2776 3496 2783 3613
rect 2796 3607 2803 3693
rect 2716 3127 2723 3483
rect 2796 3407 2803 3533
rect 2816 3527 2823 3673
rect 2836 3647 2843 3723
rect 2916 3627 2923 3703
rect 2856 3516 2863 3533
rect 2896 3523 2903 3593
rect 2956 3587 2963 4036
rect 2996 4016 3003 4073
rect 3016 4007 3023 4033
rect 2976 3967 2983 3983
rect 3036 3976 3043 4013
rect 3056 4007 3063 4053
rect 3016 3947 3023 3953
rect 3056 3867 3063 3963
rect 2976 3787 2983 3853
rect 2976 3687 2983 3773
rect 2996 3736 3003 3773
rect 3036 3736 3043 3793
rect 3056 3607 3063 3833
rect 3076 3787 3083 4093
rect 3136 4027 3143 4273
rect 3156 4196 3163 4233
rect 3176 4107 3183 4293
rect 3196 4203 3203 4373
rect 3196 4196 3223 4203
rect 3216 4087 3223 4196
rect 3236 4067 3243 4553
rect 3256 4227 3263 4513
rect 3276 4496 3283 4633
rect 3316 4467 3323 4653
rect 3336 4647 3343 4833
rect 3356 4547 3363 5133
rect 3407 4956 3423 4963
rect 3436 4956 3443 4973
rect 3416 4887 3423 4956
rect 3456 4947 3463 5053
rect 3376 4696 3403 4703
rect 3376 4627 3383 4696
rect 3376 4483 3383 4613
rect 3356 4476 3383 4483
rect 3276 4407 3283 4453
rect 3296 4423 3303 4463
rect 3296 4416 3313 4423
rect 3276 4216 3283 4373
rect 3336 4247 3343 4473
rect 3356 4447 3363 4476
rect 3396 4443 3403 4463
rect 3436 4456 3443 4473
rect 3376 4436 3403 4443
rect 3376 4423 3383 4436
rect 3367 4416 3383 4423
rect 3356 4247 3363 4333
rect 3316 4167 3323 4223
rect 3336 4187 3343 4193
rect 3096 3767 3103 4013
rect 3156 4003 3163 4033
rect 3136 3996 3163 4003
rect 3136 3976 3143 3996
rect 3176 3967 3183 4013
rect 3156 3956 3173 3963
rect 3116 3743 3123 3853
rect 3096 3736 3123 3743
rect 3076 3607 3083 3713
rect 3096 3647 3103 3736
rect 3136 3627 3143 3913
rect 3196 3847 3203 4053
rect 3256 4027 3263 4053
rect 3236 3987 3243 3993
rect 3216 3947 3223 3963
rect 3156 3727 3163 3793
rect 2896 3516 2923 3523
rect 2936 3516 2943 3553
rect 2816 3367 2823 3493
rect 2876 3467 2883 3503
rect 2736 3036 2743 3233
rect 2756 3227 2763 3293
rect 2776 3267 2783 3353
rect 2836 3263 2843 3433
rect 2876 3287 2883 3373
rect 2816 3256 2843 3263
rect 2776 3236 2783 3253
rect 2636 2907 2643 2993
rect 2596 2636 2623 2643
rect 2516 2556 2523 2573
rect 2556 2556 2563 2573
rect 2596 2567 2603 2636
rect 2516 2427 2523 2513
rect 2416 2256 2443 2263
rect 2476 2247 2483 2273
rect 2376 2103 2383 2173
rect 2356 2096 2383 2103
rect 2356 2076 2363 2096
rect 2396 2076 2403 2213
rect 2416 2107 2423 2173
rect 2436 2107 2443 2233
rect 2496 2223 2503 2293
rect 2516 2287 2523 2413
rect 2536 2347 2543 2543
rect 2576 2447 2583 2543
rect 2596 2447 2603 2493
rect 2616 2467 2623 2613
rect 2656 2607 2663 2893
rect 2676 2867 2683 3023
rect 2716 3007 2723 3023
rect 2676 2787 2683 2853
rect 2696 2607 2703 2913
rect 2716 2707 2723 2743
rect 2736 2647 2743 2993
rect 2756 2967 2763 3073
rect 2756 2647 2763 2953
rect 2776 2863 2783 3193
rect 2796 3036 2803 3073
rect 2816 3067 2823 3256
rect 2836 3036 2843 3133
rect 2876 3067 2883 3253
rect 2896 2987 2903 3473
rect 2916 3387 2923 3516
rect 3016 3516 3023 3533
rect 2996 3487 3003 3503
rect 2996 3367 3003 3473
rect 2916 3236 2923 3273
rect 2936 3187 2943 3223
rect 2776 2856 2803 2863
rect 2796 2767 2803 2856
rect 2856 2847 2863 2853
rect 2916 2847 2923 3093
rect 2956 3087 2963 3253
rect 2976 3236 2983 3293
rect 3016 3227 3023 3273
rect 3036 3247 3043 3553
rect 3056 3267 3063 3573
rect 3056 3236 3083 3243
rect 2996 3207 3003 3223
rect 2976 3056 3003 3063
rect 3016 3056 3023 3173
rect 3076 3127 3083 3236
rect 2856 2756 2863 2833
rect 2796 2736 2803 2753
rect 2816 2736 2843 2743
rect 2636 2556 2643 2593
rect 2656 2576 2673 2583
rect 2696 2563 2703 2573
rect 2676 2556 2703 2563
rect 2716 2556 2723 2573
rect 2756 2556 2763 2593
rect 2596 2327 2603 2393
rect 2556 2276 2563 2293
rect 2536 2247 2543 2263
rect 2476 2216 2503 2223
rect 2436 2076 2443 2093
rect 2456 2067 2463 2153
rect 2476 2107 2483 2216
rect 2536 2207 2543 2233
rect 2556 2076 2563 2093
rect 2376 1927 2383 2063
rect 2416 2007 2423 2063
rect 2496 2043 2503 2063
rect 2476 2036 2503 2043
rect 2256 1716 2283 1723
rect 2216 1596 2223 1613
rect 2256 1596 2263 1653
rect 2276 1587 2283 1716
rect 2296 1607 2303 1713
rect 2236 1447 2243 1583
rect 2136 1336 2163 1343
rect 2076 1287 2083 1303
rect 1976 1076 2003 1083
rect 1976 887 1983 1076
rect 2007 1056 2023 1063
rect 1996 927 2003 953
rect 1876 836 1903 843
rect 1956 836 1963 853
rect 1876 727 1883 836
rect 1996 823 2003 913
rect 2016 867 2023 1056
rect 2056 927 2063 1153
rect 2076 887 2083 1193
rect 2076 836 2083 853
rect 2096 847 2103 1153
rect 2116 1116 2123 1193
rect 2136 1167 2143 1336
rect 2176 1316 2183 1353
rect 2156 1247 2163 1303
rect 2156 1127 2163 1193
rect 2196 1027 2203 1433
rect 2236 1316 2243 1373
rect 2256 1316 2263 1453
rect 2296 1423 2303 1573
rect 2316 1547 2323 1793
rect 2336 1587 2343 1733
rect 2376 1727 2383 1853
rect 2416 1796 2423 1853
rect 2396 1767 2403 1783
rect 2356 1596 2363 1613
rect 2396 1596 2403 1713
rect 2436 1687 2443 1993
rect 2456 1887 2463 2033
rect 2476 1927 2483 2036
rect 2476 1796 2483 1813
rect 2496 1787 2503 2013
rect 2516 1887 2523 2033
rect 2536 1987 2543 2063
rect 2456 1643 2463 1773
rect 2496 1707 2503 1753
rect 2516 1727 2523 1813
rect 2556 1807 2563 2033
rect 2576 1923 2583 2233
rect 2616 2123 2623 2393
rect 2636 2247 2643 2513
rect 2736 2487 2743 2543
rect 2716 2276 2723 2413
rect 2756 2307 2763 2473
rect 2656 2223 2663 2263
rect 2756 2263 2763 2273
rect 2736 2256 2763 2263
rect 2596 2116 2623 2123
rect 2636 2216 2663 2223
rect 2596 2076 2603 2116
rect 2636 2103 2643 2216
rect 2656 2167 2663 2193
rect 2676 2123 2683 2213
rect 2616 2096 2643 2103
rect 2656 2116 2683 2123
rect 2616 2007 2623 2053
rect 2656 1967 2663 2116
rect 2676 2067 2683 2093
rect 2696 2076 2703 2153
rect 2736 2076 2743 2093
rect 2776 2076 2783 2413
rect 2816 2387 2823 2736
rect 2896 2727 2903 2753
rect 2856 2563 2863 2633
rect 2876 2576 2883 2673
rect 2896 2567 2903 2573
rect 2836 2556 2863 2563
rect 2836 2407 2843 2556
rect 2576 1916 2603 1923
rect 2536 1767 2543 1783
rect 2556 1756 2573 1763
rect 2536 1647 2543 1673
rect 2436 1636 2463 1643
rect 2436 1596 2443 1636
rect 2476 1627 2483 1633
rect 2496 1616 2513 1623
rect 2316 1447 2323 1533
rect 2356 1527 2363 1553
rect 2336 1467 2343 1513
rect 2376 1467 2383 1583
rect 2416 1487 2423 1573
rect 2296 1416 2323 1423
rect 2316 1316 2323 1416
rect 2356 1307 2363 1413
rect 2216 1287 2223 1303
rect 2276 1227 2283 1303
rect 2216 1116 2223 1153
rect 2276 1107 2283 1173
rect 2236 987 2243 1103
rect 1916 807 1923 823
rect 1976 816 2003 823
rect 1916 747 1923 793
rect 1936 747 1943 773
rect 1676 447 1683 573
rect 1496 376 1523 383
rect 1496 356 1503 376
rect 1376 307 1383 333
rect 1396 183 1403 323
rect 1416 267 1423 343
rect 1476 327 1483 343
rect 1376 176 1403 183
rect 1356 167 1363 173
rect 1376 123 1383 176
rect 1396 156 1423 163
rect 1456 156 1463 193
rect 1536 167 1543 393
rect 1396 147 1403 156
rect 1556 147 1563 353
rect 1576 243 1583 393
rect 1616 356 1623 413
rect 1656 367 1663 373
rect 1696 367 1703 513
rect 1596 327 1603 343
rect 1576 236 1603 243
rect 1596 207 1603 236
rect 1636 227 1643 343
rect 1616 156 1623 213
rect 1656 156 1663 173
rect 1676 147 1683 343
rect 1696 247 1703 333
rect 1716 327 1723 573
rect 1816 527 1823 593
rect 1736 343 1743 513
rect 1816 356 1823 453
rect 1856 367 1863 613
rect 1896 407 1903 693
rect 1916 636 1923 673
rect 1936 547 1943 633
rect 1956 547 1963 653
rect 2016 643 2023 793
rect 1996 636 2023 643
rect 1736 336 1763 343
rect 1476 123 1483 143
rect 1756 127 1763 336
rect 1896 343 1903 353
rect 1876 336 1903 343
rect 1776 303 1783 323
rect 1776 296 1803 303
rect 1776 167 1783 273
rect 1796 267 1803 296
rect 1936 267 1943 343
rect 1976 227 1983 343
rect 1996 267 2003 363
rect 2016 347 2023 413
rect 2036 356 2043 713
rect 2096 667 2103 833
rect 2136 827 2143 873
rect 2296 823 2303 1133
rect 2316 1027 2323 1273
rect 2336 1267 2343 1303
rect 2356 1207 2363 1293
rect 2376 1187 2383 1393
rect 2416 1327 2423 1353
rect 2396 1223 2403 1273
rect 2416 1247 2423 1283
rect 2396 1216 2423 1223
rect 2396 1147 2403 1193
rect 2347 1136 2383 1143
rect 2376 1116 2383 1136
rect 2416 1127 2423 1216
rect 2436 1207 2443 1303
rect 2436 1167 2443 1173
rect 2456 1147 2463 1613
rect 2476 1596 2483 1613
rect 2536 1603 2543 1633
rect 2516 1596 2543 1603
rect 2556 1596 2563 1653
rect 2576 1627 2583 1733
rect 2596 1687 2603 1916
rect 2636 1796 2643 1813
rect 2676 1796 2683 1953
rect 2716 1947 2723 2063
rect 2756 2043 2763 2063
rect 2756 2036 2783 2043
rect 2776 2007 2783 2036
rect 2616 1767 2623 1783
rect 2656 1667 2663 1783
rect 2716 1727 2723 1793
rect 2736 1647 2743 1973
rect 2756 1796 2763 1953
rect 2776 1807 2783 1993
rect 2796 1927 2803 2333
rect 2836 2287 2843 2353
rect 2876 2347 2883 2433
rect 2856 2256 2883 2263
rect 2856 2243 2863 2256
rect 2836 2236 2863 2243
rect 2816 2127 2823 2153
rect 2836 2103 2843 2236
rect 2816 2096 2843 2103
rect 2856 2096 2863 2113
rect 2816 2027 2823 2096
rect 2876 2076 2883 2193
rect 2916 2167 2923 2773
rect 2936 2627 2943 3053
rect 2996 3047 3003 3056
rect 3036 3036 3043 3073
rect 3056 3027 3063 3113
rect 3096 3087 3103 3573
rect 3136 3516 3163 3523
rect 3136 3483 3143 3516
rect 3136 3476 3163 3483
rect 3116 3267 3123 3373
rect 3136 3236 3143 3273
rect 3116 3147 3123 3223
rect 3136 3167 3143 3193
rect 3156 3107 3163 3476
rect 3176 3387 3183 3753
rect 3216 3727 3223 3753
rect 3196 3587 3203 3633
rect 3236 3567 3243 3693
rect 3256 3647 3263 3733
rect 3276 3647 3283 4093
rect 3296 3996 3303 4033
rect 3316 4016 3323 4053
rect 3356 4047 3363 4213
rect 3376 4187 3383 4203
rect 3416 4196 3423 4233
rect 3456 4207 3463 4933
rect 3496 4627 3503 5143
rect 3516 5136 3543 5143
rect 3616 5136 3623 5173
rect 3516 5127 3523 5136
rect 3656 4987 3663 5423
rect 3856 5407 3863 5423
rect 3876 5407 3883 5453
rect 3916 5443 3923 5593
rect 3936 5487 3943 5616
rect 3896 5436 3923 5443
rect 3716 5276 3733 5283
rect 3716 5176 3723 5276
rect 3896 5167 3903 5436
rect 3936 5407 3943 5423
rect 3936 5167 3943 5393
rect 3956 5383 3963 5403
rect 3996 5387 4003 5403
rect 3956 5376 3983 5383
rect 3976 5367 3983 5376
rect 3616 4947 3623 4973
rect 3676 4956 3683 5133
rect 3536 4676 3543 4813
rect 3516 4507 3523 4673
rect 3576 4663 3583 4693
rect 3576 4656 3603 4663
rect 3576 4643 3583 4656
rect 3556 4636 3583 4643
rect 3496 4456 3503 4473
rect 3516 4407 3523 4443
rect 3396 4167 3403 4183
rect 3356 3983 3363 4033
rect 3356 3976 3383 3983
rect 3316 3963 3323 3973
rect 3316 3956 3343 3963
rect 3296 3907 3303 3913
rect 3296 3707 3303 3893
rect 3316 3716 3323 3813
rect 3336 3727 3343 3956
rect 3356 3787 3363 3976
rect 3396 3727 3403 4073
rect 3416 3927 3423 3983
rect 3196 3347 3203 3553
rect 3196 3236 3203 3313
rect 3236 3267 3243 3513
rect 3256 3447 3263 3593
rect 3276 3467 3283 3633
rect 3256 3267 3263 3413
rect 3296 3287 3303 3613
rect 3316 3607 3323 3673
rect 3336 3667 3343 3683
rect 3376 3567 3383 3703
rect 3396 3627 3403 3713
rect 3416 3563 3423 3813
rect 3396 3556 3423 3563
rect 3396 3543 3403 3556
rect 3376 3536 3403 3543
rect 3436 3543 3443 4173
rect 3476 4143 3483 4393
rect 3496 4196 3503 4333
rect 3516 4203 3523 4393
rect 3536 4227 3543 4453
rect 3556 4367 3563 4636
rect 3576 4456 3583 4493
rect 3596 4476 3603 4513
rect 3636 4487 3643 4633
rect 3656 4623 3663 4683
rect 3696 4623 3703 4943
rect 3656 4616 3703 4623
rect 3616 4447 3623 4463
rect 3676 4456 3683 4616
rect 3716 4467 3723 4813
rect 3736 4767 3743 4973
rect 3756 4827 3763 4943
rect 3796 4727 3803 4933
rect 3836 4867 3843 4953
rect 3856 4807 3863 5143
rect 3976 5067 3983 5353
rect 3996 5127 4003 5143
rect 4016 5043 4023 5793
rect 4036 5787 4043 5883
rect 4056 5807 4063 6133
rect 4516 6116 4523 6133
rect 4216 6103 4223 6113
rect 4156 6027 4163 6103
rect 4196 6096 4223 6103
rect 4196 6087 4203 6096
rect 4116 5916 4123 6013
rect 4256 5936 4263 6013
rect 4067 5776 4073 5783
rect 4036 5387 4043 5633
rect 4056 5407 4063 5653
rect 4116 5623 4123 5673
rect 4096 5616 4123 5623
rect 4096 5436 4123 5443
rect 4076 5147 4083 5153
rect 4096 5127 4103 5436
rect 4136 5327 4143 5893
rect 4196 5687 4203 5933
rect 4236 5916 4243 5933
rect 4276 5927 4283 5953
rect 4336 5936 4343 6073
rect 4296 5916 4323 5923
rect 4356 5916 4403 5923
rect 4216 5787 4223 5913
rect 4296 5887 4303 5916
rect 4156 5656 4183 5663
rect 4156 5623 4163 5656
rect 4276 5647 4283 5873
rect 4376 5867 4383 5916
rect 4476 5903 4483 6053
rect 4496 6027 4503 6113
rect 4576 6067 4583 6083
rect 4616 6067 4623 6103
rect 4636 6087 4643 6113
rect 4536 5916 4543 6033
rect 4576 6007 4583 6053
rect 4576 5916 4583 5953
rect 4616 5916 4623 6053
rect 4656 5916 4663 5933
rect 4416 5887 4423 5903
rect 4456 5896 4483 5903
rect 4516 5896 4523 5913
rect 4336 5636 4343 5673
rect 4156 5616 4183 5623
rect 4156 5436 4163 5473
rect 4176 5467 4183 5616
rect 4256 5443 4263 5493
rect 4356 5467 4363 5473
rect 4376 5467 4383 5853
rect 4416 5636 4423 5713
rect 4396 5607 4403 5623
rect 4436 5587 4443 5623
rect 4456 5547 4463 5643
rect 4476 5587 4483 5896
rect 4556 5687 4563 5903
rect 4676 5896 4683 5913
rect 4716 5907 4723 6073
rect 4736 6027 4743 6123
rect 4756 6007 4763 6143
rect 4796 6136 4803 6173
rect 4816 6027 4823 6113
rect 4856 6087 4863 6153
rect 4996 6136 5003 6153
rect 5036 6136 5063 6143
rect 5096 6136 5123 6143
rect 4896 6067 4903 6133
rect 4916 6067 4923 6103
rect 4816 5943 4823 6013
rect 4956 5967 4963 6053
rect 4796 5936 4823 5943
rect 4636 5767 4643 5893
rect 4756 5887 4763 5933
rect 4856 5927 4863 5933
rect 4916 5916 4943 5923
rect 4816 5883 4823 5913
rect 4816 5876 4843 5883
rect 4536 5587 4543 5623
rect 4576 5547 4583 5623
rect 4596 5587 4603 5753
rect 4616 5687 4623 5693
rect 4616 5623 4623 5673
rect 4776 5667 4783 5793
rect 4616 5616 4643 5623
rect 4676 5587 4683 5623
rect 4236 5436 4263 5443
rect 4236 5327 4243 5436
rect 4256 5347 4263 5413
rect 4276 5403 4283 5453
rect 4356 5403 4363 5453
rect 4396 5416 4403 5533
rect 4276 5396 4303 5403
rect 4336 5367 4343 5403
rect 4356 5396 4383 5403
rect 4416 5387 4423 5403
rect 4176 5276 4193 5283
rect 4127 5176 4143 5183
rect 4176 5176 4183 5276
rect 4116 5103 4123 5173
rect 4096 5096 4123 5103
rect 4016 5036 4043 5043
rect 3956 4956 3983 4963
rect 3896 4927 3903 4943
rect 3827 4796 3833 4803
rect 3816 4683 3823 4753
rect 3816 4676 3843 4683
rect 3876 4676 3883 4713
rect 3736 4607 3743 4663
rect 3776 4627 3783 4663
rect 3816 4647 3823 4676
rect 3916 4663 3923 4853
rect 3896 4656 3923 4663
rect 3936 4647 3943 4913
rect 3776 4476 3783 4593
rect 3856 4507 3863 4643
rect 3516 4196 3543 4203
rect 3556 4196 3563 4233
rect 3536 4163 3543 4196
rect 3516 4156 3543 4163
rect 3476 4136 3503 4143
rect 3456 3827 3463 4133
rect 3476 3667 3483 4113
rect 3496 3996 3503 4136
rect 3496 3667 3503 3703
rect 3436 3536 3463 3543
rect 3376 3523 3383 3536
rect 3356 3516 3383 3523
rect 3416 3516 3433 3523
rect 3356 3467 3363 3516
rect 3396 3407 3403 3473
rect 2976 2827 2983 3013
rect 3016 2987 3023 3013
rect 2956 2767 2963 2793
rect 2936 2527 2943 2573
rect 2936 2247 2943 2433
rect 2956 2247 2963 2263
rect 2956 2187 2963 2233
rect 2916 2076 2923 2093
rect 2956 2076 2963 2153
rect 2836 2047 2843 2063
rect 2856 2007 2863 2053
rect 2896 2047 2903 2063
rect 2827 1996 2833 2003
rect 2816 1796 2823 1833
rect 2776 1727 2783 1763
rect 2796 1707 2803 1783
rect 2836 1767 2843 1783
rect 2896 1727 2903 1813
rect 2596 1596 2603 1613
rect 2636 1596 2663 1603
rect 2536 1567 2543 1573
rect 2576 1567 2583 1583
rect 2616 1547 2623 1583
rect 2616 1527 2623 1533
rect 2656 1527 2663 1596
rect 2576 1487 2583 1493
rect 2516 1316 2523 1353
rect 2476 1287 2483 1313
rect 2576 1307 2583 1473
rect 2536 1296 2563 1303
rect 2556 1287 2563 1296
rect 2396 1083 2403 1103
rect 2387 1076 2403 1083
rect 2147 816 2163 823
rect 2196 807 2203 823
rect 2296 816 2323 823
rect 2056 636 2063 653
rect 2076 567 2083 623
rect 2076 323 2083 533
rect 2096 356 2103 593
rect 2156 347 2163 793
rect 2176 667 2183 803
rect 2216 636 2223 693
rect 2196 587 2203 623
rect 2236 547 2243 613
rect 2216 356 2223 393
rect 2236 387 2243 533
rect 2236 367 2243 373
rect 2056 316 2083 323
rect 1816 176 1823 193
rect 1916 156 1923 213
rect 1956 156 1963 173
rect 1996 167 2003 193
rect 2056 147 2063 316
rect 2116 287 2123 343
rect 2136 267 2143 333
rect 2156 307 2163 333
rect 2196 267 2203 323
rect 2256 287 2263 373
rect 1376 116 1483 123
rect 2056 107 2063 133
rect 2076 123 2083 253
rect 2136 143 2143 253
rect 2276 187 2283 673
rect 2336 667 2343 1033
rect 2376 907 2383 1073
rect 2416 967 2423 1073
rect 2396 827 2403 933
rect 2436 843 2443 1133
rect 2476 1096 2483 1213
rect 2536 1096 2543 1273
rect 2576 1087 2583 1293
rect 2456 1047 2463 1053
rect 2496 967 2503 993
rect 2516 927 2523 1053
rect 2436 836 2463 843
rect 2476 836 2483 913
rect 2356 687 2363 823
rect 2296 587 2303 653
rect 2436 636 2443 693
rect 2416 567 2423 613
rect 2356 343 2363 413
rect 2416 356 2423 553
rect 2336 336 2363 343
rect 2276 156 2283 173
rect 2296 163 2303 213
rect 2316 183 2323 323
rect 2316 176 2343 183
rect 2296 156 2323 163
rect 2156 143 2163 153
rect 2336 147 2343 176
rect 2136 136 2163 143
rect 2376 127 2383 353
rect 2456 343 2463 836
rect 2476 636 2483 673
rect 2496 607 2503 823
rect 2516 383 2523 873
rect 2536 836 2543 1053
rect 2556 1047 2563 1083
rect 2596 1067 2603 1433
rect 2656 1316 2663 1453
rect 2676 1387 2683 1633
rect 2716 1616 2743 1623
rect 2736 1607 2743 1616
rect 2696 1527 2703 1583
rect 2756 1527 2763 1673
rect 2796 1427 2803 1633
rect 2816 1596 2823 1613
rect 2756 1387 2763 1413
rect 2616 1207 2623 1293
rect 2636 1207 2643 1303
rect 2676 1187 2683 1303
rect 2616 1116 2623 1173
rect 2696 1167 2703 1333
rect 2716 1207 2723 1313
rect 2636 1027 2643 1103
rect 2656 1087 2663 1153
rect 2716 1127 2723 1153
rect 2556 867 2563 993
rect 2576 427 2583 893
rect 2596 827 2603 853
rect 2616 747 2623 823
rect 2676 787 2683 1053
rect 2696 1047 2703 1103
rect 2696 847 2703 1033
rect 2716 947 2723 1113
rect 2736 1027 2743 1373
rect 2816 1347 2823 1493
rect 2836 1447 2843 1613
rect 2856 1596 2863 1673
rect 2876 1587 2883 1713
rect 2916 1683 2923 1753
rect 2936 1727 2943 1793
rect 2896 1676 2923 1683
rect 2896 1607 2903 1676
rect 2816 1316 2823 1333
rect 2756 1247 2763 1303
rect 2796 1247 2803 1303
rect 2796 1187 2803 1193
rect 2756 1136 2763 1153
rect 2796 1067 2803 1173
rect 2816 1147 2823 1173
rect 2836 1167 2843 1303
rect 2856 1147 2863 1433
rect 2876 1327 2883 1573
rect 2916 1327 2923 1413
rect 2956 1347 2963 1693
rect 2976 1427 2983 2773
rect 3056 2756 3063 2793
rect 3076 2787 3083 3073
rect 3096 3036 3123 3043
rect 3156 3036 3163 3053
rect 3096 3007 3103 3036
rect 2996 2687 3003 2743
rect 3036 2727 3043 2743
rect 2996 2556 3003 2593
rect 3016 2587 3023 2613
rect 3036 2556 3043 2693
rect 3096 2667 3103 2723
rect 3016 2127 3023 2553
rect 3056 2407 3063 2573
rect 3076 2427 3083 2653
rect 3056 2267 3063 2373
rect 3116 2367 3123 2533
rect 3016 2087 3023 2113
rect 2996 2027 3003 2033
rect 2996 1827 3003 2013
rect 3016 1787 3023 2053
rect 2996 1667 3003 1783
rect 3036 1687 3043 1773
rect 3016 1596 3023 1633
rect 3056 1627 3063 2133
rect 3076 2127 3083 2353
rect 3136 2327 3143 2993
rect 3156 2576 3163 2673
rect 3176 2583 3183 3193
rect 3216 3167 3223 3223
rect 3256 3187 3263 3223
rect 3196 3036 3203 3113
rect 3296 3087 3303 3233
rect 3316 3087 3323 3353
rect 3356 3327 3363 3393
rect 3336 3236 3343 3313
rect 3356 3267 3363 3313
rect 3356 3167 3363 3223
rect 3236 3036 3243 3053
rect 3176 2576 3203 2583
rect 3116 2307 3123 2313
rect 3116 2276 3123 2293
rect 3076 2076 3083 2093
rect 3096 1903 3103 2253
rect 3116 2147 3123 2233
rect 3176 2227 3183 2413
rect 3196 2167 3203 2576
rect 3216 2327 3223 2753
rect 3236 2727 3243 2743
rect 3236 2556 3243 2613
rect 3256 2587 3263 2973
rect 3276 2727 3283 2743
rect 3276 2707 3283 2713
rect 3276 2587 3283 2673
rect 3296 2587 3303 3053
rect 3316 3027 3323 3053
rect 3336 3047 3343 3153
rect 3376 3067 3383 3273
rect 3416 3267 3423 3473
rect 3436 3427 3443 3433
rect 3436 3247 3443 3373
rect 3456 3223 3463 3536
rect 3476 3463 3483 3653
rect 3516 3567 3523 4156
rect 3536 3996 3543 4133
rect 3596 4127 3603 4413
rect 3656 4367 3663 4443
rect 3616 4167 3623 4213
rect 3656 4187 3663 4353
rect 3696 4247 3703 4433
rect 3756 4347 3763 4463
rect 3816 4447 3823 4473
rect 3716 4167 3723 4183
rect 3616 4087 3623 4153
rect 3556 3803 3563 3953
rect 3596 3823 3603 4013
rect 3636 3996 3663 4003
rect 3696 3996 3703 4153
rect 3736 4143 3743 4313
rect 3796 4176 3803 4353
rect 3716 4136 3743 4143
rect 3636 3963 3643 3996
rect 3636 3956 3663 3963
rect 3596 3816 3623 3823
rect 3556 3796 3583 3803
rect 3556 3703 3563 3773
rect 3536 3696 3563 3703
rect 3496 3487 3503 3553
rect 3536 3547 3543 3673
rect 3576 3563 3583 3796
rect 3616 3727 3623 3816
rect 3616 3696 3643 3703
rect 3556 3556 3583 3563
rect 3556 3527 3563 3556
rect 3516 3467 3523 3483
rect 3476 3456 3503 3463
rect 3396 3067 3403 3193
rect 3416 3087 3423 3223
rect 3436 3216 3463 3223
rect 3376 3036 3393 3043
rect 3316 2967 3323 3013
rect 3356 3007 3363 3023
rect 3396 2927 3403 2953
rect 3416 2887 3423 3033
rect 3276 2556 3293 2563
rect 3236 2287 3243 2453
rect 3256 2307 3263 2543
rect 3316 2487 3323 2853
rect 3356 2767 3363 2793
rect 3416 2787 3423 2873
rect 3436 2787 3443 3216
rect 3456 2807 3463 3193
rect 3476 3147 3483 3433
rect 3496 3367 3503 3456
rect 3516 3367 3523 3453
rect 3556 3447 3563 3483
rect 3496 3247 3503 3273
rect 3556 3263 3563 3313
rect 3576 3287 3583 3533
rect 3596 3267 3603 3593
rect 3636 3587 3643 3696
rect 3656 3687 3663 3956
rect 3716 3867 3723 4136
rect 3656 3536 3693 3543
rect 3616 3516 3623 3533
rect 3656 3516 3663 3536
rect 3636 3427 3643 3503
rect 3676 3347 3683 3503
rect 3556 3256 3583 3263
rect 3536 3236 3543 3253
rect 3576 3236 3583 3256
rect 3656 3227 3663 3293
rect 3476 3067 3483 3133
rect 3496 3056 3503 3213
rect 3516 3067 3523 3193
rect 3536 2987 3543 3193
rect 3556 3147 3563 3223
rect 3576 3056 3583 3113
rect 3616 3087 3623 3193
rect 3676 3127 3683 3273
rect 3696 3263 3703 3473
rect 3716 3287 3723 3553
rect 3696 3256 3723 3263
rect 3716 3236 3723 3256
rect 3556 3047 3563 3053
rect 3596 3036 3623 3043
rect 3636 3036 3643 3113
rect 3376 2743 3383 2773
rect 3376 2736 3403 2743
rect 3436 2707 3443 2743
rect 3336 2407 3343 2573
rect 3116 2083 3123 2133
rect 3116 2076 3143 2083
rect 3116 1927 3123 2033
rect 3076 1896 3103 1903
rect 3076 1603 3083 1896
rect 3116 1783 3123 1813
rect 3136 1807 3143 2076
rect 3116 1776 3143 1783
rect 3076 1596 3103 1603
rect 3116 1596 3123 1653
rect 3136 1643 3143 1776
rect 3156 1747 3163 2153
rect 3216 2083 3223 2263
rect 3256 2227 3263 2263
rect 3276 2127 3283 2333
rect 3296 2267 3303 2333
rect 3316 2327 3323 2393
rect 3356 2387 3363 2543
rect 3376 2327 3383 2513
rect 3396 2507 3403 2543
rect 3416 2467 3423 2513
rect 3436 2507 3443 2613
rect 3476 2587 3483 2953
rect 3576 2947 3583 3013
rect 3616 3007 3623 3036
rect 3496 2756 3503 2853
rect 3536 2767 3543 2873
rect 3496 2647 3503 2713
rect 3516 2667 3523 2733
rect 3576 2687 3583 2743
rect 3456 2556 3483 2563
rect 3416 2367 3423 2453
rect 3456 2447 3463 2556
rect 3556 2556 3563 2613
rect 3207 2076 3223 2083
rect 3236 2076 3243 2113
rect 3296 2103 3303 2233
rect 3316 2227 3323 2293
rect 3296 2096 3323 2103
rect 3276 2076 3283 2093
rect 3316 2087 3323 2096
rect 3156 1667 3163 1733
rect 3136 1636 3163 1643
rect 3156 1596 3163 1636
rect 3036 1567 3043 1583
rect 3076 1527 3083 1573
rect 2916 1187 2923 1293
rect 2876 1147 2883 1173
rect 2816 1116 2823 1133
rect 2696 827 2703 833
rect 2716 827 2723 913
rect 2736 907 2743 1013
rect 2836 987 2843 1093
rect 2736 807 2743 823
rect 2816 807 2823 953
rect 2916 947 2923 1173
rect 2936 1047 2943 1333
rect 2876 823 2883 933
rect 2896 836 2903 853
rect 2936 823 2943 853
rect 2856 816 2883 823
rect 2916 816 2943 823
rect 2676 636 2683 773
rect 2736 747 2743 793
rect 2716 627 2723 713
rect 2756 663 2763 803
rect 2736 656 2763 663
rect 2736 627 2743 656
rect 2796 636 2803 693
rect 2836 636 2863 643
rect 2596 616 2623 623
rect 2596 587 2603 616
rect 2856 623 2863 636
rect 2816 587 2823 623
rect 2856 616 2883 623
rect 2596 547 2603 573
rect 2516 376 2543 383
rect 2396 167 2403 343
rect 2436 336 2463 343
rect 2536 343 2543 376
rect 2576 356 2583 393
rect 2536 336 2563 343
rect 2436 327 2443 336
rect 2756 343 2763 413
rect 2796 347 2803 533
rect 2736 336 2763 343
rect 2596 176 2603 193
rect 2776 187 2783 343
rect 2816 207 2823 433
rect 2856 347 2863 553
rect 2916 447 2923 816
rect 2956 687 2963 1303
rect 2996 1296 3023 1303
rect 2976 1167 2983 1293
rect 3016 1116 3023 1296
rect 3056 1267 3063 1313
rect 3076 1207 3083 1513
rect 3056 1116 3063 1153
rect 3096 1147 3103 1596
rect 3116 1387 3123 1453
rect 3176 1387 3183 1913
rect 3236 1796 3243 1973
rect 3256 1847 3263 2063
rect 3296 1987 3303 2063
rect 3336 1927 3343 2313
rect 3416 2276 3423 2353
rect 3456 2287 3463 2413
rect 3476 2276 3483 2293
rect 3356 2247 3363 2263
rect 3376 2223 3383 2233
rect 3436 2227 3443 2263
rect 3356 2216 3383 2223
rect 3356 2027 3363 2216
rect 3376 2076 3383 2193
rect 3396 2096 3403 2173
rect 3436 2127 3443 2193
rect 3416 2076 3423 2093
rect 3216 1767 3223 1783
rect 3256 1767 3263 1813
rect 3296 1796 3313 1803
rect 3116 1116 3123 1373
rect 3156 1147 3163 1303
rect 3196 1243 3203 1733
rect 3316 1707 3323 1793
rect 3216 1507 3223 1653
rect 3236 1596 3243 1633
rect 3276 1596 3283 1633
rect 3336 1627 3343 1833
rect 3396 1787 3403 2053
rect 3436 1827 3443 2093
rect 3456 2087 3463 2233
rect 3456 2067 3463 2073
rect 3376 1643 3383 1783
rect 3376 1636 3403 1643
rect 3396 1607 3403 1636
rect 3436 1627 3443 1783
rect 3456 1607 3463 1993
rect 3476 1807 3483 2153
rect 3496 2107 3503 2413
rect 3536 2227 3543 2243
rect 3576 2187 3583 2453
rect 3596 2427 3603 2973
rect 3616 2827 3623 2993
rect 3656 2927 3663 3023
rect 3696 2967 3703 3023
rect 3636 2767 3643 2813
rect 3676 2743 3683 2833
rect 3656 2736 3683 2743
rect 3616 2587 3623 2713
rect 3696 2643 3703 2813
rect 3676 2636 3703 2643
rect 3636 2576 3643 2593
rect 3476 1727 3483 1773
rect 3496 1763 3503 2063
rect 3516 1887 3523 2013
rect 3536 1807 3543 2173
rect 3596 2127 3603 2393
rect 3616 2287 3623 2353
rect 3576 2076 3583 2113
rect 3596 2027 3603 2093
rect 3496 1756 3523 1763
rect 3496 1607 3503 1613
rect 3316 1596 3343 1603
rect 3336 1583 3343 1596
rect 3336 1576 3363 1583
rect 3296 1567 3303 1573
rect 3236 1316 3243 1333
rect 3216 1287 3223 1293
rect 3196 1236 3223 1243
rect 3176 1136 3183 1173
rect 3036 1087 3043 1103
rect 3016 856 3023 873
rect 2936 636 2963 643
rect 2936 567 2943 636
rect 2976 427 2983 623
rect 3036 407 3043 613
rect 3056 587 3063 933
rect 3096 847 3103 1073
rect 3176 1027 3183 1093
rect 3216 963 3223 1236
rect 3256 1183 3263 1373
rect 3336 1267 3343 1553
rect 3416 1487 3423 1583
rect 3476 1567 3483 1583
rect 3516 1487 3523 1756
rect 3536 1747 3543 1763
rect 3536 1567 3543 1713
rect 3556 1707 3563 1933
rect 3576 1787 3583 1853
rect 3596 1796 3603 2013
rect 3616 1987 3623 2193
rect 3656 2107 3663 2573
rect 3676 2487 3683 2636
rect 3636 2027 3643 2063
rect 3576 1683 3583 1753
rect 3556 1676 3583 1683
rect 3556 1667 3563 1676
rect 3596 1587 3603 1733
rect 3616 1727 3623 1783
rect 3636 1747 3643 1813
rect 3656 1796 3663 1973
rect 3676 1827 3683 2393
rect 3696 2147 3703 2263
rect 3716 2167 3723 2813
rect 3736 2807 3743 4073
rect 3816 3747 3823 4253
rect 3836 4207 3843 4453
rect 3856 4407 3863 4493
rect 3896 4456 3903 4633
rect 3916 4347 3923 4443
rect 3936 4203 3943 4453
rect 3916 4196 3943 4203
rect 3856 4027 3863 4183
rect 3876 3787 3883 4153
rect 3956 4043 3963 4773
rect 3976 4727 3983 4956
rect 4016 4696 4023 4713
rect 3976 4327 3983 4443
rect 4016 4427 4023 4443
rect 4036 4363 4043 5036
rect 4056 4587 4063 5053
rect 4096 4843 4103 5096
rect 4156 4956 4183 4963
rect 4176 4887 4183 4956
rect 4076 4836 4103 4843
rect 4076 4707 4083 4836
rect 4136 4696 4143 4713
rect 4116 4583 4123 4683
rect 4096 4576 4123 4583
rect 4076 4456 4083 4493
rect 4096 4487 4103 4576
rect 4156 4567 4163 4693
rect 4176 4607 4183 4873
rect 4116 4483 4123 4553
rect 4116 4476 4143 4483
rect 4056 4387 4063 4443
rect 4116 4427 4123 4476
rect 4036 4356 4063 4363
rect 4036 4147 4043 4183
rect 3956 4036 3983 4043
rect 3916 3867 3923 4013
rect 3976 4007 3983 4036
rect 3816 3727 3823 3733
rect 3796 3696 3823 3703
rect 3796 3683 3803 3696
rect 3776 3676 3803 3683
rect 3756 3516 3763 3533
rect 3796 3516 3803 3653
rect 3836 3516 3843 3613
rect 3776 3467 3783 3503
rect 3776 3236 3783 3253
rect 3796 3236 3803 3353
rect 3856 3263 3863 3733
rect 3876 3703 3883 3773
rect 3956 3707 3963 3973
rect 4056 3967 4063 4356
rect 4076 4167 4083 4183
rect 4076 3996 4083 4013
rect 4096 3947 4103 4193
rect 4116 4167 4123 4393
rect 4176 4367 4183 4573
rect 4196 4527 4203 5133
rect 4216 5107 4223 5313
rect 4296 5156 4303 5293
rect 4276 5127 4283 5143
rect 4336 5047 4343 5313
rect 4356 5147 4363 5273
rect 4376 5007 4383 5373
rect 4416 5156 4423 5213
rect 4396 5107 4403 5143
rect 4436 5067 4443 5453
rect 4456 5347 4463 5453
rect 4516 5447 4523 5513
rect 4536 5447 4543 5453
rect 4476 5327 4483 5423
rect 4496 5307 4503 5413
rect 4516 5407 4523 5433
rect 4656 5427 4663 5573
rect 4696 5527 4703 5653
rect 4776 5636 4783 5653
rect 4756 5607 4763 5613
rect 4736 5587 4743 5593
rect 4816 5587 4823 5643
rect 4836 5627 4843 5876
rect 4936 5767 4943 5916
rect 4956 5867 4963 5913
rect 4976 5687 4983 6093
rect 5016 6047 5023 6133
rect 5036 6127 5043 6136
rect 5016 5667 5023 5903
rect 5036 5727 5043 6093
rect 5076 5943 5083 6123
rect 5116 6103 5123 6136
rect 5196 6103 5203 6173
rect 5316 6136 5323 6173
rect 5096 6096 5123 6103
rect 5176 6096 5203 6103
rect 5096 6027 5103 6096
rect 5056 5936 5083 5943
rect 5096 5936 5103 5953
rect 5056 5787 5063 5936
rect 5116 5916 5123 6013
rect 5176 5936 5183 6033
rect 5156 5916 5163 5933
rect 5196 5916 5223 5923
rect 5036 5667 5043 5713
rect 4556 5407 4563 5423
rect 4596 5416 4623 5423
rect 4476 5187 4483 5233
rect 4556 5207 4563 5373
rect 4576 5347 4583 5393
rect 4616 5367 4623 5416
rect 4676 5416 4683 5433
rect 4716 5407 4723 5513
rect 4736 5436 4753 5443
rect 4496 5176 4513 5183
rect 4496 5163 4503 5176
rect 4556 5176 4563 5193
rect 4476 5156 4503 5163
rect 4456 4956 4463 5013
rect 4236 4927 4243 4953
rect 4476 4923 4483 5033
rect 4356 4823 4363 4923
rect 4456 4916 4483 4923
rect 4356 4816 4373 4823
rect 4387 4816 4403 4823
rect 4276 4796 4293 4803
rect 4276 4696 4283 4796
rect 4216 4483 4223 4593
rect 4296 4563 4303 4733
rect 4356 4676 4363 4753
rect 4396 4663 4403 4816
rect 4456 4687 4463 4916
rect 4376 4656 4403 4663
rect 4456 4567 4463 4673
rect 4496 4587 4503 5093
rect 4536 5067 4543 5163
rect 4596 4983 4603 5193
rect 4616 5187 4623 5253
rect 4656 5147 4663 5353
rect 4696 5307 4703 5403
rect 4676 5107 4683 5293
rect 4716 5156 4723 5193
rect 4736 5187 4743 5436
rect 4796 5436 4803 5513
rect 4776 5247 4783 5423
rect 4816 5416 4823 5513
rect 4836 5287 4843 5553
rect 4856 5547 4863 5623
rect 4856 5436 4863 5493
rect 4876 5403 4883 5473
rect 4896 5467 4903 5593
rect 4956 5587 4963 5653
rect 4916 5436 4923 5513
rect 4936 5403 4943 5573
rect 4996 5567 5003 5603
rect 5016 5587 5023 5623
rect 4956 5447 4963 5533
rect 4976 5407 4983 5513
rect 5036 5447 5043 5653
rect 5056 5647 5063 5753
rect 5216 5747 5223 5916
rect 5236 5896 5243 6103
rect 5296 5916 5303 5953
rect 5116 5667 5123 5693
rect 5096 5636 5103 5653
rect 5076 5587 5083 5623
rect 4876 5396 4903 5403
rect 4916 5396 4943 5403
rect 4856 5347 4863 5393
rect 4696 5047 4703 5143
rect 4756 5127 4763 5143
rect 4576 4976 4603 4983
rect 4516 4607 4523 4653
rect 4276 4556 4303 4563
rect 4196 4476 4223 4483
rect 4196 4407 4203 4476
rect 4236 4427 4243 4533
rect 4256 4476 4263 4493
rect 4187 4316 4193 4323
rect 4156 4176 4163 4253
rect 4196 4187 4203 4313
rect 4276 4223 4283 4556
rect 4316 4527 4323 4533
rect 4256 4216 4283 4223
rect 4216 4167 4223 4203
rect 4256 4196 4263 4216
rect 4116 4007 4123 4153
rect 4236 4147 4243 4183
rect 4216 4016 4243 4023
rect 4216 4003 4223 4016
rect 4196 3996 4223 4003
rect 3876 3696 3903 3703
rect 3916 3696 3943 3703
rect 3916 3536 3923 3696
rect 3956 3523 3963 3693
rect 3996 3603 4003 3753
rect 3976 3596 4003 3603
rect 3976 3547 3983 3596
rect 4016 3587 4023 3713
rect 4036 3643 4043 3873
rect 4176 3703 4183 3753
rect 4156 3696 4183 3703
rect 4036 3636 4063 3643
rect 3996 3547 4003 3573
rect 3876 3516 3903 3523
rect 3936 3516 3963 3523
rect 3876 3487 3883 3516
rect 3836 3256 3863 3263
rect 3756 2827 3763 3113
rect 3776 3056 3783 3153
rect 3796 3063 3803 3173
rect 3816 3167 3823 3223
rect 3836 3187 3843 3256
rect 3876 3207 3883 3213
rect 3896 3187 3903 3393
rect 3796 3056 3823 3063
rect 3776 2787 3783 2873
rect 3816 2827 3823 3056
rect 3836 3043 3843 3153
rect 3836 3036 3863 3043
rect 3836 2847 3843 3013
rect 3736 2583 3743 2773
rect 3816 2756 3823 2773
rect 3756 2707 3763 2743
rect 3796 2707 3803 2743
rect 3736 2576 3763 2583
rect 3716 2076 3723 2093
rect 3736 2007 3743 2093
rect 3196 956 3223 963
rect 3236 1176 3263 1183
rect 3116 643 3123 693
rect 3136 667 3143 853
rect 3156 687 3163 823
rect 3116 636 3143 643
rect 3176 636 3183 673
rect 3196 647 3203 956
rect 3236 863 3243 1176
rect 3256 1107 3263 1153
rect 3276 1096 3283 1213
rect 3296 1116 3303 1253
rect 3376 1187 3383 1303
rect 3416 1287 3423 1303
rect 3436 1267 3443 1323
rect 3456 1303 3463 1353
rect 3456 1296 3483 1303
rect 3336 1116 3343 1173
rect 3236 856 3263 863
rect 3236 816 3243 833
rect 3256 727 3263 856
rect 2896 207 2903 373
rect 2916 367 2923 393
rect 3116 376 3123 593
rect 3036 356 3043 373
rect 3156 367 3163 633
rect 3276 547 3283 1033
rect 3316 1007 3323 1103
rect 3356 1083 3363 1133
rect 3396 1096 3403 1253
rect 3436 1083 3443 1173
rect 3356 1076 3383 1083
rect 3416 1076 3443 1083
rect 3296 847 3303 893
rect 3356 867 3363 1076
rect 3416 887 3423 1076
rect 3456 1047 3463 1253
rect 3516 1187 3523 1303
rect 3536 1267 3543 1353
rect 3476 1116 3483 1173
rect 3516 1116 3523 1153
rect 3556 1107 3563 1333
rect 3576 1047 3583 1253
rect 3616 1167 3623 1693
rect 3636 1607 3643 1673
rect 3656 1563 3663 1753
rect 3676 1596 3683 1633
rect 3696 1627 3703 1813
rect 3716 1796 3723 1833
rect 3736 1807 3743 1953
rect 3756 1827 3763 2576
rect 3776 2563 3783 2633
rect 3796 2563 3803 2573
rect 3776 2556 3803 2563
rect 3796 2367 3803 2556
rect 3876 2527 3883 2913
rect 3896 2907 3903 3033
rect 3916 2927 3923 3473
rect 3936 3107 3943 3113
rect 3936 3036 3943 3093
rect 3956 3036 3983 3043
rect 3956 3007 3963 3036
rect 3916 2756 3923 2793
rect 3896 2367 3903 2723
rect 3936 2643 3943 2933
rect 3996 2907 4003 3313
rect 4016 3207 4023 3223
rect 4016 3127 4023 3193
rect 4036 3087 4043 3613
rect 4056 3267 4063 3636
rect 4076 3483 4083 3533
rect 4136 3523 4143 3683
rect 4216 3667 4223 3913
rect 4236 3747 4243 3833
rect 4256 3767 4263 3983
rect 4276 3927 4283 4153
rect 4236 3687 4243 3733
rect 4296 3716 4303 4293
rect 4316 4216 4323 4513
rect 4376 4247 4383 4453
rect 4396 4443 4403 4493
rect 4456 4483 4463 4553
rect 4536 4487 4543 4973
rect 4576 4783 4583 4976
rect 4596 4956 4623 4963
rect 4576 4776 4603 4783
rect 4456 4476 4483 4483
rect 4476 4456 4483 4476
rect 4396 4436 4423 4443
rect 4416 4287 4423 4436
rect 4496 4436 4503 4473
rect 4556 4447 4563 4713
rect 4596 4656 4603 4776
rect 4616 4667 4623 4956
rect 4676 4727 4683 4953
rect 4696 4767 4703 5033
rect 4756 4983 4763 5113
rect 4776 5023 4783 5153
rect 4816 5027 4823 5273
rect 4856 5156 4863 5333
rect 4776 5016 4803 5023
rect 4736 4976 4763 4983
rect 4736 4947 4743 4976
rect 4796 4967 4803 5016
rect 4736 4927 4743 4933
rect 4676 4607 4683 4663
rect 4736 4627 4743 4893
rect 4756 4687 4763 4933
rect 4816 4923 4823 4973
rect 4836 4967 4843 5143
rect 4876 5087 4883 5143
rect 4896 5067 4903 5163
rect 4916 5047 4923 5396
rect 4936 5247 4943 5373
rect 4936 4967 4943 5233
rect 4956 5127 4963 5173
rect 4976 5163 4983 5233
rect 4996 5187 5003 5403
rect 4976 5156 5003 5163
rect 4976 5067 4983 5156
rect 4956 4956 4963 5013
rect 4996 4967 5003 5093
rect 5036 5023 5043 5253
rect 5056 5187 5063 5553
rect 5076 5547 5083 5573
rect 5116 5447 5123 5623
rect 5136 5547 5143 5643
rect 5156 5567 5163 5653
rect 5176 5647 5183 5733
rect 5256 5663 5263 5673
rect 5196 5656 5223 5663
rect 5256 5656 5283 5663
rect 5196 5487 5203 5656
rect 5076 5416 5083 5433
rect 5136 5387 5143 5403
rect 5176 5403 5183 5473
rect 5216 5427 5223 5533
rect 5176 5396 5203 5403
rect 5116 5267 5123 5333
rect 5156 5327 5163 5393
rect 5256 5387 5263 5433
rect 5076 5176 5083 5253
rect 5116 5176 5143 5183
rect 5016 5016 5043 5023
rect 4816 4916 4843 4923
rect 4796 4676 4803 4853
rect 4576 4507 4583 4513
rect 4356 4216 4383 4223
rect 4336 4187 4343 4203
rect 4316 3687 4323 3703
rect 4136 3516 4163 3523
rect 4196 3516 4203 3533
rect 4236 3516 4243 3673
rect 4256 3527 4263 3593
rect 4076 3476 4103 3483
rect 4136 3383 4143 3483
rect 4156 3403 4163 3516
rect 4276 3503 4283 3653
rect 4336 3607 4343 3733
rect 4256 3496 4283 3503
rect 4156 3396 4183 3403
rect 4136 3376 4153 3383
rect 4056 3147 4063 3223
rect 3987 2876 3993 2883
rect 3916 2636 3943 2643
rect 3796 2267 3803 2333
rect 3816 2076 3823 2233
rect 3836 2147 3843 2353
rect 3876 2276 3883 2313
rect 3916 2307 3923 2636
rect 3956 2607 3963 2813
rect 3956 2567 3963 2593
rect 3856 2227 3863 2263
rect 3896 2227 3903 2263
rect 3856 2083 3863 2173
rect 3856 2076 3883 2083
rect 3916 2076 3923 2173
rect 3956 2107 3963 2353
rect 3976 2147 3983 2513
rect 3996 2327 4003 2613
rect 4036 2583 4043 2893
rect 4056 2627 4063 3073
rect 4116 3067 4123 3253
rect 4176 3227 4183 3396
rect 4256 3203 4263 3496
rect 4276 3207 4283 3223
rect 4236 3196 4263 3203
rect 4076 2747 4083 3053
rect 4176 3036 4183 3073
rect 4036 2576 4063 2583
rect 4016 2556 4023 2573
rect 3796 2047 3803 2063
rect 3836 1947 3843 2063
rect 3796 1783 3803 1853
rect 3816 1796 3823 1813
rect 3856 1807 3863 2013
rect 3896 1967 3903 2063
rect 3936 2047 3943 2063
rect 3956 1987 3963 2033
rect 3776 1776 3803 1783
rect 3796 1747 3803 1753
rect 3876 1747 3883 1783
rect 3896 1767 3903 1813
rect 3916 1796 3923 1893
rect 3976 1827 3983 2113
rect 3996 2107 4003 2233
rect 4036 2127 4043 2553
rect 4056 2407 4063 2576
rect 4096 2527 4103 2563
rect 4116 2447 4123 3023
rect 4236 3016 4243 3196
rect 4296 3083 4303 3233
rect 4316 3127 4323 3573
rect 4336 3516 4343 3533
rect 4356 3247 4363 4093
rect 4376 4087 4383 4216
rect 4456 4216 4463 4313
rect 4396 3567 4403 4203
rect 4436 4187 4443 4203
rect 4476 4163 4483 4413
rect 4536 4407 4543 4443
rect 4556 4387 4563 4433
rect 4596 4427 4603 4463
rect 4616 4387 4623 4473
rect 4636 4447 4643 4473
rect 4496 4187 4503 4333
rect 4556 4196 4563 4293
rect 4476 4156 4503 4163
rect 4436 3987 4443 4033
rect 4436 3703 4443 3973
rect 4456 3967 4463 3983
rect 4436 3696 4463 3703
rect 4376 3516 4403 3523
rect 4356 3216 4383 3223
rect 4276 3076 4303 3083
rect 4156 2727 4163 2743
rect 4016 2096 4023 2113
rect 4056 2076 4063 2273
rect 4076 2103 4083 2433
rect 4136 2307 4143 2673
rect 4176 2603 4183 2953
rect 4216 2887 4223 3003
rect 4256 2747 4263 3003
rect 4276 2787 4283 3076
rect 4336 3056 4343 3073
rect 4356 2967 4363 3173
rect 4376 2943 4383 3216
rect 4396 3207 4403 3516
rect 4416 3267 4423 3633
rect 4436 3183 4443 3353
rect 4476 3247 4483 3953
rect 4356 2936 4383 2943
rect 4416 3176 4443 3183
rect 4196 2707 4203 2743
rect 4176 2596 4203 2603
rect 4156 2276 4163 2543
rect 4196 2467 4203 2596
rect 4236 2536 4243 2653
rect 4256 2587 4263 2733
rect 4216 2287 4223 2513
rect 4256 2427 4263 2523
rect 4176 2223 4183 2263
rect 4196 2256 4223 2263
rect 4196 2247 4203 2256
rect 4176 2216 4203 2223
rect 4096 2127 4103 2133
rect 4076 2096 4103 2103
rect 3996 2056 4023 2063
rect 4016 2047 4023 2056
rect 3636 1556 3663 1563
rect 3636 1287 3643 1556
rect 3676 1327 3683 1413
rect 3696 1347 3703 1613
rect 3656 1287 3663 1303
rect 3436 856 3463 863
rect 3296 627 3303 653
rect 3316 636 3323 833
rect 3336 767 3343 823
rect 3376 807 3383 823
rect 3376 643 3383 793
rect 3456 787 3463 856
rect 3496 823 3503 993
rect 3476 816 3503 823
rect 3356 636 3383 643
rect 3396 627 3403 753
rect 3476 667 3483 816
rect 3496 667 3503 673
rect 3176 356 3203 363
rect 2996 347 3003 353
rect 3056 287 3063 323
rect 3196 207 3203 356
rect 3296 343 3303 393
rect 3336 376 3343 613
rect 3276 336 3303 343
rect 3316 327 3323 373
rect 3416 363 3423 453
rect 3356 356 3383 363
rect 3396 356 3423 363
rect 2827 196 2843 203
rect 2536 156 2563 163
rect 2556 143 2563 156
rect 2736 156 2743 173
rect 2836 163 2843 196
rect 2816 156 2843 163
rect 2516 127 2523 143
rect 2556 136 2583 143
rect 2076 116 2103 123
rect 2856 123 2863 153
rect 2936 123 2943 193
rect 3236 187 3243 273
rect 2996 156 3023 163
rect 3056 156 3063 173
rect 2996 147 3003 156
rect 3136 127 3143 163
rect 3236 136 3243 173
rect 3296 156 3303 193
rect 3376 187 3383 356
rect 3436 183 3443 653
rect 3456 636 3483 643
rect 3496 636 3503 653
rect 3476 627 3483 636
rect 3416 176 3443 183
rect 3376 156 3383 173
rect 3416 147 3423 176
rect 3476 163 3483 343
rect 3496 167 3503 593
rect 3516 487 3523 1033
rect 3596 1007 3603 1083
rect 3636 1076 3643 1133
rect 3656 1127 3663 1273
rect 3676 1147 3683 1313
rect 3696 1247 3703 1303
rect 3756 1267 3763 1733
rect 3776 1307 3783 1713
rect 3876 1596 3883 1693
rect 3896 1563 3903 1593
rect 3896 1556 3923 1563
rect 3796 1267 3803 1333
rect 3856 1316 3863 1333
rect 3916 1327 3923 1556
rect 3956 1367 3963 1753
rect 3536 827 3543 913
rect 3636 883 3643 893
rect 3656 883 3663 1053
rect 3636 876 3663 883
rect 3636 867 3643 876
rect 3676 863 3683 1093
rect 3696 927 3703 1103
rect 3716 1047 3723 1233
rect 3756 1107 3763 1213
rect 3796 1083 3803 1113
rect 3736 1067 3743 1083
rect 3776 1076 3803 1083
rect 3656 856 3683 863
rect 3536 807 3543 813
rect 3576 687 3583 833
rect 3536 343 3543 433
rect 3596 407 3603 853
rect 3616 647 3623 833
rect 3616 616 3623 633
rect 3636 607 3643 673
rect 3656 667 3663 856
rect 3736 827 3743 843
rect 3676 643 3683 813
rect 3716 787 3723 823
rect 3756 823 3763 1033
rect 3776 867 3783 1053
rect 3796 887 3803 1076
rect 3816 883 3823 1313
rect 3876 1247 3883 1303
rect 3896 1147 3903 1293
rect 3936 1267 3943 1303
rect 3956 1227 3963 1323
rect 3976 1207 3983 1313
rect 3996 1227 4003 2033
rect 4036 2027 4043 2053
rect 4016 1787 4023 1973
rect 4036 1727 4043 1993
rect 4056 1767 4063 2033
rect 4076 2007 4083 2073
rect 4076 1707 4083 1773
rect 4096 1747 4103 2096
rect 4116 2076 4123 2193
rect 4156 2076 4163 2113
rect 4196 2087 4203 2216
rect 4216 2096 4223 2213
rect 4136 1867 4143 2063
rect 4136 1816 4163 1823
rect 4036 1587 4043 1693
rect 4076 1583 4083 1673
rect 4056 1576 4083 1583
rect 4016 1307 4023 1573
rect 4076 1327 4083 1576
rect 4096 1447 4103 1693
rect 4116 1627 4123 1783
rect 4136 1667 4143 1816
rect 4156 1616 4163 1633
rect 4196 1583 4203 1653
rect 4176 1576 4203 1583
rect 4216 1567 4223 2033
rect 4236 1687 4243 1853
rect 4256 1816 4263 2293
rect 4276 2287 4283 2773
rect 4356 2527 4363 2936
rect 4416 2867 4423 3176
rect 4456 2827 4463 3233
rect 4476 3036 4483 3053
rect 4496 2927 4503 4156
rect 4536 4147 4543 4183
rect 4596 4183 4603 4373
rect 4636 4267 4643 4433
rect 4656 4243 4663 4453
rect 4676 4347 4683 4593
rect 4736 4427 4743 4443
rect 4696 4287 4703 4413
rect 4756 4307 4763 4673
rect 4776 4647 4783 4663
rect 4856 4627 4863 4663
rect 4876 4627 4883 4673
rect 4896 4667 4903 4913
rect 4916 4696 4923 4933
rect 4976 4903 4983 4933
rect 4956 4896 4983 4903
rect 4956 4747 4963 4896
rect 4936 4667 4943 4683
rect 4776 4367 4783 4413
rect 4836 4367 4843 4443
rect 4636 4236 4663 4243
rect 4596 4176 4623 4183
rect 4536 4016 4543 4073
rect 4556 3996 4563 4013
rect 4616 4003 4623 4176
rect 4636 4167 4643 4236
rect 4676 4227 4683 4273
rect 4656 4216 4673 4223
rect 4696 4083 4703 4273
rect 4716 4187 4723 4253
rect 4736 4196 4743 4213
rect 4676 4076 4703 4083
rect 4616 3996 4643 4003
rect 4516 3827 4523 3983
rect 4576 3967 4583 3983
rect 4536 3696 4543 3853
rect 4556 3807 4563 3953
rect 4636 3887 4643 3996
rect 4656 3847 4663 4013
rect 4676 3967 4683 4076
rect 4676 3907 4683 3953
rect 4596 3716 4603 3733
rect 4616 3567 4623 3683
rect 4516 3527 4523 3553
rect 4376 2587 4383 2733
rect 4396 2727 4403 2743
rect 4436 2687 4443 2743
rect 4396 2576 4403 2593
rect 4376 2556 4383 2573
rect 4436 2563 4443 2573
rect 4416 2556 4443 2563
rect 4276 2047 4283 2253
rect 4296 2247 4303 2263
rect 4296 2167 4303 2233
rect 4296 1847 4303 2133
rect 4316 2007 4323 2513
rect 4347 2416 4353 2423
rect 4356 2267 4363 2373
rect 4336 2207 4343 2263
rect 4336 2076 4343 2173
rect 4376 2076 4383 2173
rect 4416 2087 4423 2313
rect 4436 2147 4443 2556
rect 4356 1987 4363 2063
rect 4296 1816 4313 1823
rect 4036 1316 4063 1323
rect 4036 1287 4043 1316
rect 3916 1103 3923 1193
rect 3896 1096 3923 1103
rect 3936 1116 3963 1123
rect 4036 1116 4043 1133
rect 3816 876 3843 883
rect 3756 816 3783 823
rect 3656 636 3683 643
rect 3656 616 3663 636
rect 3516 336 3543 343
rect 3456 156 3483 163
rect 2856 116 2883 123
rect 2916 116 2943 123
rect 3456 -24 3463 156
rect 3507 156 3523 163
rect 3476 136 3503 143
rect 3476 127 3483 136
rect 3516 116 3523 156
rect 3536 136 3543 193
rect 3556 163 3563 343
rect 3596 307 3603 343
rect 3556 156 3583 163
rect 3576 -24 3583 156
rect 3616 127 3623 553
rect 3696 447 3703 633
rect 3756 587 3763 603
rect 3776 567 3783 816
rect 3796 607 3803 833
rect 3836 623 3843 876
rect 3856 827 3863 1073
rect 3816 616 3843 623
rect 3856 616 3863 753
rect 3896 627 3903 843
rect 3936 836 3943 1116
rect 3976 1047 3983 1103
rect 4016 1087 4023 1103
rect 4076 1047 4083 1083
rect 4136 927 4143 1553
rect 4236 1147 4243 1433
rect 4256 1407 4263 1713
rect 4276 1647 4283 1793
rect 4316 1783 4323 1813
rect 4316 1776 4343 1783
rect 4236 1123 4243 1133
rect 4236 1116 4263 1123
rect 4176 1096 4183 1113
rect 3916 636 3923 823
rect 3956 807 3963 823
rect 3936 636 3963 643
rect 3796 467 3803 593
rect 3876 587 3883 603
rect 3656 356 3683 363
rect 3676 187 3683 356
rect 3796 356 3803 413
rect 3836 347 3843 433
rect 3696 327 3703 343
rect 3736 323 3743 333
rect 3716 316 3743 323
rect 3776 307 3783 343
rect 3816 267 3823 343
rect 3876 327 3883 473
rect 3896 287 3903 613
rect 3916 376 3923 573
rect 3936 407 3943 636
rect 3976 507 3983 913
rect 4096 823 4103 873
rect 4036 807 4043 823
rect 4076 816 4103 823
rect 3636 156 3663 163
rect 3676 156 3703 163
rect 3816 156 3843 163
rect 3636 -24 3643 156
rect 3676 127 3683 156
rect 3836 -24 3843 156
rect 3916 -24 3923 173
rect 3936 136 3943 273
rect 3976 187 3983 393
rect 3996 387 4003 773
rect 4056 667 4063 803
rect 4116 787 4123 803
rect 4156 663 4163 1083
rect 4196 856 4203 1033
rect 4236 856 4243 1116
rect 4296 947 4303 1733
rect 4336 1587 4343 1776
rect 4356 1707 4363 1873
rect 4396 1783 4403 1993
rect 4376 1776 4403 1783
rect 4416 1747 4423 1833
rect 4436 1783 4443 2073
rect 4456 1867 4463 2813
rect 4516 2667 4523 3493
rect 4536 3387 4543 3533
rect 4616 3516 4623 3533
rect 4636 3507 4643 3813
rect 4656 3487 4663 3793
rect 4696 3736 4703 3773
rect 4756 3743 4763 4073
rect 4776 4047 4783 4353
rect 4856 4347 4863 4573
rect 4896 4483 4903 4653
rect 4976 4567 4983 4873
rect 4996 4607 5003 4913
rect 5016 4707 5023 5016
rect 5036 4936 5043 4993
rect 5056 4987 5063 5173
rect 5076 4936 5083 5013
rect 5116 4927 5123 4973
rect 4876 4476 4903 4483
rect 4876 4243 4883 4476
rect 4956 4443 4963 4493
rect 4896 4307 4903 4443
rect 4936 4436 4963 4443
rect 4896 4267 4903 4293
rect 4876 4236 4903 4243
rect 4856 4216 4883 4223
rect 4876 4207 4883 4216
rect 4796 4147 4803 4203
rect 4776 3996 4783 4013
rect 4736 3736 4763 3743
rect 4756 3547 4763 3736
rect 4776 3647 4783 3833
rect 4796 3787 4803 4013
rect 4816 3867 4823 4193
rect 4836 4167 4843 4203
rect 4856 4127 4863 4133
rect 4876 4003 4883 4173
rect 4856 3996 4883 4003
rect 4816 3736 4823 3773
rect 4836 3763 4843 3853
rect 4856 3787 4863 3996
rect 4896 3767 4903 4236
rect 4936 4183 4943 4253
rect 4956 4227 4963 4373
rect 4976 4267 4983 4553
rect 5016 4487 5023 4693
rect 5036 4627 5043 4663
rect 5016 4407 5023 4443
rect 5036 4347 5043 4413
rect 4996 4227 5003 4293
rect 4916 4176 4943 4183
rect 4936 4027 4943 4176
rect 4996 4067 5003 4213
rect 5016 4047 5023 4333
rect 5076 4287 5083 4893
rect 5096 4847 5103 4923
rect 5136 4807 5143 5176
rect 5156 5087 5163 5163
rect 5236 5147 5243 5353
rect 5256 5347 5263 5373
rect 5276 5227 5283 5656
rect 5316 5647 5323 6053
rect 5336 5907 5343 6033
rect 5376 5967 5383 6103
rect 5416 6047 5423 6103
rect 5476 6087 5483 6153
rect 5536 6136 5543 6153
rect 5416 5987 5423 6033
rect 5516 6007 5523 6123
rect 5616 6116 5623 6153
rect 5436 5936 5463 5943
rect 5416 5923 5423 5933
rect 5436 5923 5443 5936
rect 5416 5916 5443 5923
rect 5396 5883 5403 5913
rect 5436 5887 5443 5916
rect 5376 5876 5403 5883
rect 5376 5747 5383 5876
rect 5336 5607 5343 5623
rect 5316 5567 5323 5603
rect 5336 5587 5343 5593
rect 5376 5567 5383 5713
rect 5416 5636 5423 5693
rect 5456 5647 5463 5793
rect 5296 5407 5303 5493
rect 5336 5436 5343 5493
rect 5316 5416 5323 5433
rect 5356 5267 5363 5413
rect 5396 5367 5403 5573
rect 5436 5567 5443 5623
rect 5476 5607 5483 5623
rect 5416 5387 5423 5403
rect 5216 5127 5223 5143
rect 5176 4976 5183 4993
rect 5156 4783 5163 4953
rect 5196 4787 5203 4943
rect 5216 4907 5223 4993
rect 5236 4947 5243 5053
rect 5256 4827 5263 5213
rect 5316 5176 5323 5193
rect 5336 5187 5343 5253
rect 5396 5187 5403 5213
rect 5416 5187 5423 5373
rect 5456 5207 5463 5403
rect 5476 5247 5483 5433
rect 5296 5127 5303 5153
rect 5296 4936 5303 4953
rect 5276 4887 5283 4923
rect 5136 4776 5163 4783
rect 5096 4567 5103 4663
rect 5116 4483 5123 4593
rect 5136 4507 5143 4776
rect 5156 4696 5163 4753
rect 5236 4707 5243 4773
rect 5176 4667 5183 4683
rect 5196 4547 5203 4673
rect 5216 4667 5223 4683
rect 5256 4676 5263 4733
rect 5276 4707 5283 4793
rect 5236 4607 5243 4663
rect 5156 4483 5163 4493
rect 5096 4476 5123 4483
rect 5136 4476 5163 4483
rect 5036 4216 5043 4253
rect 5076 4247 5083 4253
rect 5056 4167 5063 4203
rect 5076 4167 5083 4173
rect 5056 4147 5063 4153
rect 5096 4107 5103 4476
rect 5136 4456 5143 4476
rect 5196 4467 5203 4533
rect 5216 4456 5223 4493
rect 5116 4427 5123 4443
rect 5116 4247 5123 4413
rect 5156 4307 5163 4443
rect 5196 4436 5203 4453
rect 5256 4447 5263 4553
rect 5276 4487 5283 4613
rect 5316 4527 5323 4773
rect 5336 4507 5343 5173
rect 5396 5156 5403 5173
rect 5456 5143 5463 5193
rect 5496 5187 5503 5913
rect 5536 5903 5543 5953
rect 5516 5896 5543 5903
rect 5576 5916 5603 5923
rect 5636 5916 5643 6033
rect 5676 6027 5683 6073
rect 5716 6067 5723 6103
rect 5736 6067 5743 6103
rect 5796 6047 5803 6123
rect 5916 6103 5923 6113
rect 6016 6107 6023 6133
rect 6116 6116 6123 6153
rect 6176 6136 6183 6153
rect 6216 6136 6243 6143
rect 5856 6047 5863 6103
rect 5896 6096 5923 6103
rect 5876 6047 5883 6083
rect 6036 6027 6043 6113
rect 6236 6107 6243 6136
rect 6276 6127 6283 6153
rect 6396 6127 6403 6153
rect 6056 6087 6063 6103
rect 6056 6067 6063 6073
rect 5656 5927 5663 5933
rect 5516 5587 5523 5873
rect 5576 5847 5583 5916
rect 5616 5887 5623 5903
rect 5656 5896 5663 5913
rect 5676 5887 5683 6013
rect 5696 5916 5703 5973
rect 5716 5887 5723 5893
rect 5616 5687 5623 5833
rect 5616 5656 5643 5663
rect 5536 5587 5543 5643
rect 5556 5607 5563 5623
rect 5556 5436 5563 5473
rect 5596 5427 5603 5593
rect 5436 5136 5463 5143
rect 5396 4956 5403 5013
rect 5416 5007 5423 5133
rect 5416 4936 5443 4943
rect 5396 4696 5403 4913
rect 5436 4767 5443 4936
rect 5456 4923 5463 5136
rect 5496 5127 5503 5143
rect 5516 5127 5523 5393
rect 5536 5227 5543 5423
rect 5616 5263 5623 5656
rect 5696 5647 5703 5873
rect 5776 5807 5783 5993
rect 5796 5916 5803 5973
rect 5816 5947 5823 6013
rect 5836 5916 5843 5973
rect 5816 5887 5823 5903
rect 5856 5896 5863 5933
rect 5716 5467 5723 5753
rect 5796 5656 5803 5673
rect 5736 5567 5743 5633
rect 5776 5587 5783 5643
rect 5636 5407 5643 5433
rect 5656 5367 5663 5453
rect 5736 5443 5743 5533
rect 5716 5436 5743 5443
rect 5616 5256 5643 5263
rect 5576 5156 5583 5213
rect 5556 5067 5563 5143
rect 5616 5127 5623 5163
rect 5536 4956 5563 4963
rect 5536 4923 5543 4956
rect 5456 4916 5483 4923
rect 5436 4696 5443 4713
rect 5456 4707 5463 4733
rect 5476 4727 5483 4916
rect 5516 4867 5523 4923
rect 5536 4916 5563 4923
rect 5556 4887 5563 4916
rect 5516 4696 5543 4703
rect 5416 4507 5423 4673
rect 5536 4667 5543 4696
rect 5556 4687 5563 4873
rect 5636 4747 5643 5256
rect 5696 5247 5703 5413
rect 5736 5387 5743 5436
rect 5716 5327 5723 5373
rect 5756 5263 5763 5573
rect 5816 5447 5823 5673
rect 5876 5667 5883 5993
rect 6036 5927 6043 5953
rect 6036 5896 6043 5913
rect 5836 5436 5843 5573
rect 5896 5563 5903 5623
rect 5956 5607 5963 5873
rect 6056 5847 6063 5883
rect 5916 5587 5923 5603
rect 5896 5556 5923 5563
rect 5876 5436 5883 5553
rect 5816 5387 5823 5403
rect 5756 5256 5783 5263
rect 5656 5047 5663 5143
rect 5696 5127 5703 5143
rect 5656 4947 5663 5033
rect 5716 5007 5723 5163
rect 5736 5067 5743 5233
rect 5756 5007 5763 5233
rect 5776 5207 5783 5256
rect 5816 5247 5823 5373
rect 5856 5367 5863 5423
rect 5836 5176 5843 5213
rect 5796 5147 5803 5173
rect 5816 5127 5823 5163
rect 5756 4967 5763 4993
rect 5676 4956 5703 4963
rect 5676 4867 5683 4956
rect 5796 4963 5803 5053
rect 5796 4956 5823 4963
rect 5856 4956 5863 4993
rect 5716 4907 5723 4953
rect 5796 4927 5803 4956
rect 5236 4243 5243 4443
rect 5276 4423 5283 4473
rect 5296 4456 5303 4493
rect 5356 4476 5383 4483
rect 5336 4447 5343 4463
rect 5316 4423 5323 4433
rect 5276 4416 5303 4423
rect 5316 4416 5343 4423
rect 5296 4407 5303 4416
rect 5256 4247 5263 4313
rect 5216 4236 5243 4243
rect 5216 4207 5223 4236
rect 5136 4187 5143 4203
rect 4956 4016 4963 4033
rect 4976 3996 4983 4013
rect 4936 3947 4943 3983
rect 4996 3967 5003 4033
rect 5076 4027 5083 4053
rect 5096 4003 5103 4093
rect 5156 4083 5163 4193
rect 5216 4167 5223 4193
rect 5236 4107 5243 4213
rect 5256 4196 5263 4233
rect 5296 4207 5303 4333
rect 5316 4167 5323 4183
rect 5156 4076 5183 4083
rect 5036 3996 5063 4003
rect 4936 3863 4943 3933
rect 4996 3867 5003 3953
rect 5016 3947 5023 3963
rect 5056 3927 5063 3996
rect 5076 3996 5103 4003
rect 4936 3856 4963 3863
rect 4836 3756 4863 3763
rect 4856 3736 4863 3756
rect 4956 3747 4963 3856
rect 4976 3767 4983 3793
rect 4996 3767 5003 3853
rect 4976 3743 4983 3753
rect 4976 3736 5003 3743
rect 4836 3627 4843 3723
rect 4876 3687 4883 3733
rect 4936 3716 4943 3733
rect 4996 3716 5003 3736
rect 4896 3667 4903 3713
rect 4756 3516 4783 3523
rect 4556 3236 4563 3273
rect 4596 3203 4603 3253
rect 4616 3247 4623 3473
rect 4676 3256 4703 3263
rect 4596 3196 4623 3203
rect 4576 3043 4583 3073
rect 4556 3036 4583 3043
rect 4496 2107 4503 2473
rect 4516 2187 4523 2263
rect 4516 2096 4523 2153
rect 4516 1807 4523 2033
rect 4436 1776 4463 1783
rect 4356 1607 4363 1633
rect 4316 1307 4323 1333
rect 4356 1303 4363 1593
rect 4396 1567 4403 1603
rect 4456 1576 4463 1653
rect 4536 1627 4543 2913
rect 4596 2663 4603 3173
rect 4576 2656 4603 2663
rect 4576 2536 4583 2656
rect 4556 2327 4563 2523
rect 4596 2423 4603 2523
rect 4616 2447 4623 3196
rect 4696 3087 4703 3256
rect 4716 3207 4723 3273
rect 4736 3267 4743 3353
rect 4776 3287 4783 3516
rect 4736 3227 4743 3253
rect 4716 3067 4723 3193
rect 4756 3187 4763 3243
rect 4796 3236 4803 3293
rect 4896 3227 4903 3653
rect 4916 3587 4923 3703
rect 4976 3687 4983 3703
rect 4916 3267 4923 3553
rect 4956 3496 4963 3633
rect 4776 3187 4783 3223
rect 4916 3187 4923 3223
rect 4656 2743 4663 3053
rect 4716 3036 4723 3053
rect 4636 2736 4663 2743
rect 4636 2727 4643 2736
rect 4636 2567 4643 2693
rect 4596 2416 4613 2423
rect 4556 2247 4563 2263
rect 4576 2167 4583 2313
rect 4556 1816 4563 2083
rect 4596 1847 4603 2273
rect 4636 2256 4643 2313
rect 4616 2043 4623 2093
rect 4636 2076 4643 2093
rect 4616 2036 4643 2043
rect 4596 1816 4623 1823
rect 4516 1567 4523 1593
rect 4536 1567 4543 1583
rect 4336 1296 4363 1303
rect 4316 1047 4323 1293
rect 4336 1127 4343 1296
rect 4376 1116 4383 1133
rect 4396 887 4403 1093
rect 4396 863 4403 873
rect 4396 856 4423 863
rect 4216 827 4223 843
rect 4296 683 4303 833
rect 4416 807 4423 856
rect 4296 676 4323 683
rect 4296 667 4303 676
rect 4136 656 4163 663
rect 4156 647 4163 656
rect 4316 656 4323 676
rect 4336 667 4343 793
rect 4436 747 4443 1393
rect 4516 1367 4523 1553
rect 4516 1336 4523 1353
rect 4456 867 4463 1313
rect 4556 1147 4563 1653
rect 4596 1407 4603 1773
rect 4616 1607 4623 1816
rect 4636 1727 4643 2036
rect 4656 1887 4663 2433
rect 4696 2327 4703 2833
rect 4736 2647 4743 3113
rect 4936 3063 4943 3483
rect 4976 3476 4983 3513
rect 4996 3503 5003 3593
rect 5016 3527 5023 3703
rect 5036 3647 5043 3713
rect 5056 3607 5063 3753
rect 5076 3607 5083 3996
rect 5116 3976 5123 4053
rect 5096 3947 5103 3963
rect 5136 3927 5143 3963
rect 5176 3947 5183 4076
rect 5216 4047 5223 4093
rect 5336 4087 5343 4416
rect 5356 4147 5363 4253
rect 5116 3716 5123 3833
rect 5136 3747 5143 3913
rect 5036 3516 5043 3553
rect 4996 3496 5023 3503
rect 5016 3347 5023 3496
rect 4956 3207 4963 3223
rect 5036 3216 5043 3273
rect 4956 3087 4963 3193
rect 4816 3056 4843 3063
rect 4916 3056 4943 3063
rect 4816 3043 4823 3056
rect 4796 3036 4823 3043
rect 4916 3016 4923 3056
rect 4956 2887 4963 3023
rect 5036 3016 5043 3173
rect 4847 2876 4853 2883
rect 4736 2556 4743 2593
rect 4756 2576 4763 2793
rect 4796 2756 4803 2873
rect 4856 2763 4863 2833
rect 4996 2783 5003 3013
rect 5056 2996 5063 3573
rect 5096 3516 5103 3573
rect 5116 3503 5123 3613
rect 5136 3523 5143 3703
rect 5156 3687 5163 3723
rect 5176 3567 5183 3753
rect 5196 3567 5203 4033
rect 5216 3947 5223 3963
rect 5216 3747 5223 3853
rect 5256 3736 5263 3753
rect 5256 3667 5263 3693
rect 5136 3516 5163 3523
rect 5156 3507 5163 3516
rect 5116 3496 5143 3503
rect 5176 3496 5183 3513
rect 5076 3467 5083 3483
rect 5196 3427 5203 3483
rect 5136 3267 5143 3333
rect 5116 3223 5123 3243
rect 5116 3216 5163 3223
rect 5196 3207 5203 3213
rect 5176 3063 5183 3203
rect 5216 3107 5223 3493
rect 5256 3447 5263 3573
rect 5276 3487 5283 3833
rect 5296 3827 5303 4013
rect 5316 3996 5323 4033
rect 5356 3996 5363 4033
rect 5376 4027 5383 4476
rect 5396 4447 5403 4493
rect 5436 4487 5443 4653
rect 5476 4476 5483 4513
rect 5516 4476 5523 4553
rect 5396 4247 5403 4413
rect 5416 4287 5423 4473
rect 5456 4447 5463 4463
rect 5456 4427 5463 4433
rect 5436 4207 5443 4373
rect 5476 4196 5483 4213
rect 5396 4176 5413 4183
rect 5336 3907 5343 3983
rect 5376 3976 5383 3993
rect 5396 3967 5403 4176
rect 5456 4047 5463 4183
rect 5496 4087 5503 4183
rect 5416 3976 5423 4033
rect 5436 3987 5443 4013
rect 5476 4003 5483 4053
rect 5536 4023 5543 4633
rect 5576 4627 5583 4683
rect 5556 4476 5563 4553
rect 5596 4483 5603 4693
rect 5656 4627 5663 4853
rect 5736 4747 5743 4923
rect 5716 4696 5723 4733
rect 5756 4647 5763 4913
rect 5816 4887 5823 4913
rect 5836 4867 5843 4933
rect 5796 4676 5803 4853
rect 5836 4667 5843 4683
rect 5776 4647 5783 4663
rect 5816 4627 5823 4663
rect 5576 4476 5603 4483
rect 5576 4447 5583 4476
rect 5656 4483 5663 4493
rect 5636 4476 5663 4483
rect 5696 4476 5703 4533
rect 5716 4487 5723 4513
rect 5587 4436 5603 4443
rect 5556 4227 5563 4433
rect 5556 4067 5563 4153
rect 5576 4127 5583 4183
rect 5596 4167 5603 4393
rect 5616 4327 5623 4433
rect 5636 4347 5643 4476
rect 5716 4456 5743 4463
rect 5736 4427 5743 4456
rect 5796 4463 5803 4493
rect 5816 4467 5823 4513
rect 5836 4487 5843 4653
rect 5856 4527 5863 4813
rect 5896 4787 5903 5313
rect 5916 5267 5923 5556
rect 5936 5416 5943 5473
rect 5976 5443 5983 5633
rect 5996 5607 6003 5713
rect 6076 5687 6083 5953
rect 6096 5947 6103 6103
rect 6136 5967 6143 6093
rect 6296 6027 6303 6073
rect 6356 6067 6363 6113
rect 6416 6067 6423 6123
rect 6436 6087 6443 6143
rect 6476 6136 6503 6143
rect 6496 6087 6503 6136
rect 6516 6047 6523 6113
rect 6536 6047 6543 6123
rect 6556 6067 6563 6103
rect 6096 5903 6103 5933
rect 6096 5896 6123 5903
rect 6156 5896 6163 5913
rect 6236 5907 6243 5933
rect 6416 5916 6423 5933
rect 6196 5896 6223 5903
rect 6196 5827 6203 5896
rect 6236 5876 6243 5893
rect 6016 5636 6023 5653
rect 6136 5623 6143 5733
rect 6196 5667 6203 5813
rect 6216 5656 6223 5673
rect 6236 5667 6243 5793
rect 6336 5747 6343 5913
rect 6256 5656 6283 5663
rect 6316 5656 6323 5713
rect 6376 5687 6383 5853
rect 6396 5827 6403 5903
rect 6476 5896 6503 5903
rect 6476 5727 6483 5896
rect 6516 5876 6523 5973
rect 6536 5927 6543 6033
rect 6676 6027 6683 6123
rect 6736 6087 6743 6123
rect 6756 6047 6763 6143
rect 6796 6136 6823 6143
rect 6816 6047 6823 6136
rect 6856 6087 6863 6123
rect 6876 6027 6883 6133
rect 7036 6116 7043 6153
rect 7096 6123 7103 6133
rect 7096 6116 7123 6123
rect 6616 5936 6623 5973
rect 6556 5867 6563 5883
rect 6116 5616 6143 5623
rect 6076 5487 6083 5603
rect 6176 5547 6183 5623
rect 6256 5527 6263 5656
rect 6376 5643 6383 5673
rect 6496 5656 6503 5833
rect 6556 5663 6563 5853
rect 6596 5847 6603 5893
rect 6536 5656 6563 5663
rect 6296 5587 6303 5643
rect 6376 5636 6403 5643
rect 6576 5623 6583 5773
rect 6636 5727 6643 5903
rect 6576 5616 6593 5623
rect 6656 5623 6663 5673
rect 6676 5663 6683 6013
rect 7136 5987 7143 6103
rect 7176 6007 7183 6103
rect 7236 6007 7243 6123
rect 7256 6047 7263 6143
rect 7296 6136 7323 6143
rect 7276 6087 7283 6113
rect 6756 5907 6763 5913
rect 6816 5903 6823 5913
rect 6776 5896 6803 5903
rect 6816 5896 6843 5903
rect 6696 5687 6703 5883
rect 6736 5807 6743 5883
rect 6776 5847 6783 5896
rect 7016 5896 7023 5973
rect 7036 5927 7043 5953
rect 7056 5896 7063 5973
rect 7076 5916 7083 5953
rect 7116 5916 7123 5933
rect 7156 5916 7163 5933
rect 6856 5683 6863 5883
rect 6856 5676 6883 5683
rect 6676 5656 6703 5663
rect 6716 5656 6723 5673
rect 6636 5616 6663 5623
rect 6056 5456 6063 5473
rect 5956 5436 5983 5443
rect 6096 5436 6123 5443
rect 6256 5436 6283 5443
rect 6316 5436 6343 5443
rect 5956 5407 5963 5436
rect 6076 5407 6083 5423
rect 5996 5207 6003 5403
rect 5916 5156 5923 5173
rect 5956 5167 5963 5193
rect 6116 5187 6123 5436
rect 6196 5307 6203 5403
rect 6236 5347 6243 5403
rect 6276 5307 6283 5436
rect 6296 5347 6303 5403
rect 6336 5227 6343 5436
rect 6396 5287 6403 5403
rect 6036 5127 6043 5163
rect 6196 5163 6203 5193
rect 6236 5167 6243 5183
rect 6296 5167 6303 5213
rect 6196 5156 6223 5163
rect 5916 4956 5923 4973
rect 5956 4956 5963 5113
rect 6036 5107 6043 5113
rect 6056 5047 6063 5143
rect 6156 5087 6163 5143
rect 5936 4907 5943 4943
rect 5916 4696 5923 4773
rect 5956 4696 5963 4813
rect 5996 4727 6003 4973
rect 6176 4956 6183 5153
rect 6296 5127 6303 5153
rect 6216 4956 6223 4993
rect 6316 4987 6323 5173
rect 6336 5156 6343 5193
rect 6416 5067 6423 5433
rect 6476 5403 6483 5453
rect 6576 5443 6583 5593
rect 6696 5567 6703 5656
rect 6576 5436 6603 5443
rect 6516 5416 6523 5433
rect 6596 5427 6603 5436
rect 6776 5436 6783 5613
rect 6796 5607 6803 5623
rect 6816 5463 6823 5603
rect 6856 5467 6863 5653
rect 6876 5487 6883 5676
rect 6956 5667 6963 5883
rect 7036 5847 7043 5893
rect 7016 5687 7023 5833
rect 7036 5656 7043 5673
rect 6916 5587 6923 5603
rect 6816 5456 6843 5463
rect 6836 5447 6843 5456
rect 6476 5396 6503 5403
rect 6436 5163 6443 5193
rect 6436 5156 6463 5163
rect 6476 5127 6483 5183
rect 6556 5183 6563 5413
rect 6596 5407 6603 5413
rect 6616 5407 6623 5423
rect 6636 5403 6643 5433
rect 6676 5416 6683 5433
rect 6636 5396 6663 5403
rect 6736 5187 6743 5213
rect 6536 5176 6563 5183
rect 6496 5107 6503 5153
rect 6536 5143 6543 5176
rect 6756 5183 6763 5433
rect 6856 5423 6863 5453
rect 6836 5416 6863 5423
rect 6896 5416 6903 5433
rect 6856 5227 6863 5416
rect 6876 5387 6883 5403
rect 6756 5176 6783 5183
rect 6676 5156 6703 5163
rect 6736 5156 6743 5173
rect 6536 5136 6563 5143
rect 6376 4976 6383 4993
rect 6316 4956 6343 4963
rect 6016 4923 6023 4953
rect 6016 4916 6043 4923
rect 6036 4907 6043 4916
rect 6076 4723 6083 4923
rect 6096 4723 6103 4953
rect 6156 4907 6163 4943
rect 6076 4716 6103 4723
rect 5996 4687 6003 4713
rect 6036 4647 6043 4693
rect 6056 4627 6063 4673
rect 6096 4607 6103 4716
rect 6176 4676 6183 4713
rect 6236 4667 6243 4683
rect 5896 4476 5923 4483
rect 5776 4456 5803 4463
rect 5616 4187 5623 4313
rect 5456 3996 5483 4003
rect 5516 4016 5543 4023
rect 5456 3976 5463 3996
rect 5356 3767 5363 3953
rect 5396 3927 5403 3933
rect 5476 3827 5483 3963
rect 5516 3943 5523 4016
rect 5536 3967 5543 3983
rect 5556 3976 5583 3983
rect 5496 3936 5523 3943
rect 5496 3847 5503 3936
rect 5556 3847 5563 3976
rect 5596 3967 5603 4153
rect 5636 4067 5643 4173
rect 5656 4147 5663 4203
rect 5696 4196 5703 4233
rect 5756 4207 5763 4453
rect 5816 4407 5823 4433
rect 5796 4196 5803 4273
rect 5676 4047 5683 4183
rect 5716 4007 5723 4183
rect 5736 4167 5743 4183
rect 5836 4183 5843 4413
rect 5896 4407 5903 4476
rect 5996 4476 6023 4483
rect 5936 4447 5943 4453
rect 6016 4447 6023 4476
rect 6016 4287 6023 4433
rect 6056 4423 6063 4593
rect 6196 4567 6203 4663
rect 6076 4467 6083 4493
rect 6196 4487 6203 4493
rect 6216 4476 6223 4513
rect 6256 4507 6263 4703
rect 6296 4696 6303 4733
rect 6316 4727 6323 4956
rect 6416 4936 6423 4993
rect 6456 4947 6463 4953
rect 6356 4927 6363 4933
rect 6316 4667 6323 4693
rect 6336 4687 6343 4713
rect 6396 4647 6403 4663
rect 6196 4456 6203 4473
rect 6276 4467 6283 4553
rect 6316 4487 6323 4633
rect 6376 4456 6383 4533
rect 6416 4447 6423 4733
rect 6436 4587 6443 4733
rect 6476 4727 6483 4923
rect 6496 4747 6503 5053
rect 6556 4967 6563 5136
rect 6616 5127 6623 5153
rect 6676 5087 6683 5156
rect 6596 4936 6603 4953
rect 6536 4847 6543 4923
rect 6576 4887 6583 4923
rect 6616 4916 6623 4973
rect 6636 4936 6643 5033
rect 6456 4667 6463 4713
rect 6576 4707 6583 4833
rect 6616 4767 6623 4873
rect 6536 4696 6563 4703
rect 6476 4547 6483 4673
rect 6516 4667 6523 4683
rect 6556 4627 6563 4696
rect 6616 4696 6623 4753
rect 6596 4647 6603 4673
rect 6636 4647 6643 4663
rect 6456 4467 6463 4473
rect 6476 4447 6483 4493
rect 6496 4487 6503 4553
rect 6496 4456 6503 4473
rect 6056 4416 6083 4423
rect 5816 4176 5843 4183
rect 5616 3976 5623 3993
rect 5296 3667 5303 3713
rect 5376 3707 5383 3723
rect 5356 3687 5363 3703
rect 5396 3703 5403 3813
rect 5436 3716 5443 3793
rect 5516 3747 5523 3833
rect 5576 3743 5583 3933
rect 5636 3907 5643 3963
rect 5656 3787 5663 3953
rect 5556 3736 5583 3743
rect 5636 3736 5643 3753
rect 5676 3747 5683 3933
rect 5756 3807 5763 3993
rect 5796 3976 5803 4013
rect 5856 4007 5863 4053
rect 5876 4003 5883 4193
rect 5896 4167 5903 4183
rect 5936 4107 5943 4183
rect 5916 4067 5923 4093
rect 5876 3996 5903 4003
rect 5936 3996 5943 4073
rect 5956 4027 5963 4203
rect 5996 4167 6003 4183
rect 6036 4087 6043 4183
rect 5776 3943 5783 3973
rect 5776 3936 5803 3943
rect 5776 3927 5783 3936
rect 5396 3696 5423 3703
rect 5296 3496 5303 3573
rect 5356 3523 5363 3573
rect 5416 3547 5423 3696
rect 5356 3516 5383 3523
rect 5436 3507 5443 3653
rect 5336 3487 5343 3493
rect 5276 3307 5283 3473
rect 5316 3256 5323 3273
rect 5396 3223 5403 3473
rect 5376 3216 5403 3223
rect 5436 3187 5443 3353
rect 5456 3267 5463 3673
rect 5496 3663 5503 3733
rect 5536 3707 5543 3723
rect 5476 3656 5503 3663
rect 5476 3467 5483 3656
rect 5496 3487 5503 3633
rect 5536 3496 5543 3513
rect 5516 3447 5523 3483
rect 5576 3287 5583 3736
rect 5776 3736 5783 3773
rect 5596 3536 5603 3613
rect 5656 3587 5663 3713
rect 5796 3707 5803 3936
rect 5836 3727 5843 3793
rect 5856 3767 5863 3963
rect 5876 3907 5883 3973
rect 5896 3967 5903 3996
rect 5996 3996 6023 4003
rect 5896 3723 5903 3813
rect 5956 3787 5963 3993
rect 6016 3967 6023 3996
rect 6056 3987 6063 4193
rect 6076 4127 6083 4416
rect 6136 4287 6143 4443
rect 6436 4427 6443 4443
rect 6136 4223 6143 4233
rect 6176 4227 6183 4353
rect 6116 4216 6143 4223
rect 6116 4187 6123 4216
rect 6296 4203 6303 4273
rect 6116 4147 6123 4173
rect 6156 4147 6163 4203
rect 6276 4196 6303 4203
rect 6256 4127 6263 4183
rect 6096 3976 6103 4013
rect 6136 3963 6143 4113
rect 6116 3956 6143 3963
rect 5876 3716 5903 3723
rect 5916 3703 5923 3733
rect 5956 3716 5963 3773
rect 5976 3727 5983 3793
rect 5996 3727 6003 3953
rect 6016 3727 6023 3813
rect 6116 3807 6123 3956
rect 6056 3716 6063 3733
rect 6116 3723 6123 3753
rect 6116 3716 6143 3723
rect 5616 3487 5623 3503
rect 5716 3496 5723 3513
rect 5756 3507 5763 3553
rect 5816 3547 5823 3693
rect 5856 3567 5863 3703
rect 5916 3696 5943 3703
rect 5776 3516 5783 3533
rect 5856 3307 5863 3513
rect 5996 3503 6003 3673
rect 6056 3507 6063 3533
rect 5976 3496 6003 3503
rect 5896 3467 5903 3473
rect 5936 3427 5943 3473
rect 6036 3447 6043 3483
rect 5816 3267 5823 3293
rect 6036 3283 6043 3433
rect 6027 3276 6043 3283
rect 5736 3256 5763 3263
rect 5456 3207 5463 3253
rect 5476 3187 5483 3233
rect 5496 3227 5503 3243
rect 5536 3236 5543 3253
rect 5636 3236 5643 3253
rect 5676 3227 5683 3243
rect 5516 3167 5523 3223
rect 5556 3187 5563 3223
rect 5596 3187 5603 3223
rect 5756 3127 5763 3256
rect 5856 3256 5863 3273
rect 5176 3056 5193 3063
rect 5336 3036 5343 3073
rect 5436 3056 5463 3063
rect 5436 3043 5443 3056
rect 5416 3036 5443 3043
rect 5516 3036 5543 3043
rect 5096 2847 5103 3003
rect 4976 2776 5003 2783
rect 4836 2756 4863 2763
rect 4896 2756 4903 2773
rect 4776 2707 4783 2743
rect 4776 2587 4783 2693
rect 4696 2256 4703 2293
rect 4736 1807 4743 2313
rect 4776 2107 4783 2263
rect 4676 1767 4683 1793
rect 4776 1787 4783 2093
rect 4716 1776 4743 1783
rect 4716 1707 4723 1776
rect 4636 1576 4643 1673
rect 4596 1316 4603 1373
rect 4616 1327 4623 1563
rect 4676 1563 4683 1593
rect 4756 1587 4763 1693
rect 4796 1623 4803 2633
rect 4816 2527 4823 2593
rect 4836 2587 4843 2713
rect 4936 2567 4943 2753
rect 4976 2747 4983 2776
rect 5196 2776 5223 2783
rect 5256 2776 5263 2793
rect 4856 2527 4863 2543
rect 4896 2536 4903 2553
rect 4827 2496 4843 2503
rect 4816 2247 4823 2263
rect 4836 2056 4843 2496
rect 4916 2327 4923 2553
rect 4936 2523 4943 2553
rect 5016 2523 5023 2763
rect 5056 2743 5063 2773
rect 5056 2736 5083 2743
rect 5196 2727 5203 2776
rect 5076 2556 5083 2593
rect 5096 2536 5103 2553
rect 4936 2516 4963 2523
rect 4996 2516 5023 2523
rect 4936 2243 4943 2283
rect 4976 2276 4983 2493
rect 4936 2236 4963 2243
rect 4816 1847 4823 2043
rect 4916 1827 4923 2083
rect 4936 1803 4943 1953
rect 4956 1807 4963 2236
rect 4996 2227 5003 2263
rect 4996 2076 5003 2093
rect 5016 1967 5023 2473
rect 5036 2076 5043 2253
rect 5116 2143 5123 2573
rect 5136 2347 5143 2553
rect 5176 2536 5183 2573
rect 5236 2567 5243 2763
rect 5416 2743 5423 3036
rect 5516 3027 5523 3036
rect 5616 3036 5643 3043
rect 5516 2783 5523 3013
rect 5556 2887 5563 3023
rect 5636 3007 5643 3036
rect 5656 2887 5663 3003
rect 5696 2987 5703 3003
rect 5547 2876 5553 2883
rect 5516 2776 5543 2783
rect 5356 2727 5363 2743
rect 5396 2736 5423 2743
rect 5536 2743 5543 2776
rect 5716 2747 5723 3073
rect 5736 3047 5743 3053
rect 5736 3016 5743 3033
rect 5756 2996 5763 3093
rect 5776 3027 5783 3253
rect 5876 3243 5883 3273
rect 5876 3236 5903 3243
rect 5916 3167 5923 3263
rect 5856 3056 5863 3093
rect 5816 3003 5823 3053
rect 5896 3036 5903 3073
rect 5996 3067 6003 3253
rect 6016 3243 6023 3273
rect 6076 3267 6083 3703
rect 6116 3687 6123 3716
rect 6216 3707 6223 3973
rect 6236 3967 6243 4053
rect 6256 3976 6263 4013
rect 6276 3983 6283 4196
rect 6376 4167 6383 4253
rect 6316 4067 6323 4163
rect 6416 4147 6423 4183
rect 6356 4027 6363 4073
rect 6276 3976 6293 3983
rect 6356 3976 6363 3993
rect 6376 3956 6383 4053
rect 6456 3976 6463 4133
rect 6476 3987 6483 4203
rect 6496 3976 6503 4013
rect 6516 4007 6523 4573
rect 6596 4476 6623 4483
rect 6536 4187 6543 4253
rect 6556 4147 6563 4203
rect 6596 4196 6603 4273
rect 6616 4227 6623 4476
rect 6636 4467 6643 4633
rect 6676 4547 6683 5053
rect 6716 4943 6723 5033
rect 6756 5007 6763 5143
rect 6776 5067 6783 5176
rect 6896 5176 6923 5183
rect 6836 5127 6843 5163
rect 6876 5087 6883 5163
rect 6796 4956 6803 4973
rect 6896 4967 6903 4993
rect 6916 4947 6923 5176
rect 6936 5147 6943 5593
rect 6976 5587 6983 5643
rect 6996 5507 7003 5653
rect 7056 5647 7063 5693
rect 7116 5683 7123 5713
rect 7136 5707 7143 5913
rect 7216 5903 7223 5973
rect 7316 5927 7323 6136
rect 7356 6047 7363 6083
rect 7396 5967 7403 6103
rect 7416 5927 7423 6173
rect 7656 6167 7663 6173
rect 7436 6083 7443 6113
rect 7516 6087 7523 6133
rect 7556 6116 7563 6153
rect 7616 6136 7663 6143
rect 7616 6127 7623 6136
rect 7656 6123 7663 6136
rect 7736 6136 7743 6173
rect 7656 6116 7683 6123
rect 7676 6107 7683 6116
rect 7436 6076 7463 6083
rect 7456 6007 7463 6076
rect 7536 5987 7543 6103
rect 7656 6087 7663 6093
rect 7696 6087 7703 6133
rect 7576 6067 7583 6083
rect 7716 6067 7723 6113
rect 7536 5936 7563 5943
rect 7216 5896 7243 5903
rect 7236 5867 7243 5896
rect 7256 5847 7263 5913
rect 7296 5876 7303 5913
rect 7376 5896 7383 5913
rect 7336 5707 7343 5883
rect 7356 5687 7363 5893
rect 7396 5876 7403 5893
rect 7116 5676 7143 5683
rect 7136 5656 7143 5676
rect 6956 5247 6963 5473
rect 7056 5447 7063 5633
rect 7076 5587 7083 5643
rect 6976 5407 6983 5423
rect 7016 5407 7023 5433
rect 7036 5403 7043 5413
rect 7036 5396 7063 5403
rect 6956 5207 6963 5213
rect 6956 5176 6963 5193
rect 6996 5187 7003 5233
rect 7076 5176 7083 5193
rect 6976 5147 6983 5163
rect 7056 5127 7063 5163
rect 7096 5007 7103 5393
rect 7116 5187 7123 5493
rect 7136 5423 7143 5613
rect 7156 5467 7163 5673
rect 7176 5627 7183 5643
rect 7256 5607 7263 5673
rect 7336 5656 7363 5663
rect 7276 5607 7283 5643
rect 7296 5547 7303 5633
rect 7316 5623 7323 5643
rect 7316 5616 7343 5623
rect 7336 5607 7343 5616
rect 7336 5587 7343 5593
rect 7356 5587 7363 5656
rect 7376 5647 7383 5653
rect 7416 5636 7423 5673
rect 7456 5647 7463 5913
rect 7556 5867 7563 5936
rect 7576 5887 7583 5973
rect 7676 5916 7683 5953
rect 7696 5916 7703 5953
rect 7836 5936 7843 5973
rect 7876 5947 7883 6103
rect 7876 5916 7903 5923
rect 7136 5416 7163 5423
rect 7176 5396 7183 5493
rect 7196 5416 7203 5433
rect 7116 5147 7123 5173
rect 7136 5107 7143 5373
rect 7216 5187 7223 5403
rect 7256 5227 7263 5493
rect 7276 5247 7283 5433
rect 7296 5427 7303 5533
rect 7476 5507 7483 5713
rect 7556 5687 7563 5853
rect 7496 5587 7503 5643
rect 7576 5623 7583 5653
rect 7316 5467 7323 5473
rect 7316 5436 7323 5453
rect 7376 5407 7383 5423
rect 7196 5176 7213 5183
rect 7296 5176 7323 5183
rect 7176 5127 7183 5163
rect 7236 5147 7243 5163
rect 6936 4967 6943 4993
rect 7116 4956 7123 4973
rect 7156 4956 7163 4973
rect 7216 4967 7223 5093
rect 7276 4976 7283 5013
rect 6716 4936 6743 4943
rect 6816 4936 6843 4943
rect 6696 4663 6703 4933
rect 6816 4867 6823 4936
rect 6927 4936 6943 4943
rect 7036 4936 7063 4943
rect 6896 4907 6903 4923
rect 6696 4656 6723 4663
rect 6696 4567 6703 4656
rect 6776 4627 6783 4683
rect 6816 4667 6823 4853
rect 6916 4747 6923 4913
rect 6996 4687 7003 4923
rect 7016 4887 7023 4933
rect 6876 4676 6903 4683
rect 6876 4647 6883 4676
rect 7016 4667 7023 4873
rect 7036 4867 7043 4936
rect 7136 4727 7143 4953
rect 7216 4936 7243 4943
rect 7236 4887 7243 4936
rect 7216 4707 7223 4713
rect 7036 4696 7063 4703
rect 6836 4627 6843 4643
rect 6716 4496 6723 4613
rect 6656 4476 6683 4483
rect 6656 4287 6663 4476
rect 6756 4463 6763 4513
rect 6736 4456 6763 4463
rect 6776 4456 6783 4613
rect 6916 4527 6923 4643
rect 7036 4587 7043 4696
rect 7096 4647 7103 4693
rect 7136 4683 7143 4693
rect 7116 4676 7143 4683
rect 7216 4676 7223 4693
rect 6816 4456 6823 4513
rect 6916 4463 6923 4473
rect 6936 4467 6943 4493
rect 6896 4456 6923 4463
rect 6796 4436 6803 4453
rect 6896 4447 6903 4456
rect 7056 4456 7063 4493
rect 7076 4467 7083 4473
rect 7096 4456 7103 4473
rect 6936 4436 6943 4453
rect 6656 4196 6663 4273
rect 6716 4203 6723 4253
rect 6696 4196 6723 4203
rect 6756 4196 6763 4233
rect 6796 4207 6803 4213
rect 6576 4127 6583 4183
rect 6836 4183 6843 4233
rect 6736 4167 6743 4183
rect 6536 3987 6543 4013
rect 6556 4003 6563 4113
rect 6556 3996 6583 4003
rect 6576 3987 6583 3996
rect 6596 3976 6603 4093
rect 6676 4016 6683 4093
rect 6716 3996 6723 4133
rect 6776 4067 6783 4183
rect 6816 4176 6843 4183
rect 6856 4147 6863 4413
rect 6976 4247 6983 4443
rect 6996 4427 7003 4453
rect 7076 4436 7083 4453
rect 6916 4196 6943 4203
rect 6436 3963 6443 3973
rect 6416 3956 6443 3963
rect 6236 3736 6243 3753
rect 6276 3736 6283 3813
rect 6356 3716 6363 3773
rect 6516 3763 6523 3963
rect 6576 3956 6583 3973
rect 6616 3767 6623 3963
rect 6496 3756 6523 3763
rect 6496 3743 6503 3756
rect 6536 3747 6543 3753
rect 6476 3736 6503 3743
rect 6476 3707 6483 3736
rect 6616 3736 6643 3743
rect 6096 3516 6103 3573
rect 6376 3563 6383 3703
rect 6516 3587 6523 3723
rect 6376 3556 6403 3563
rect 6236 3536 6263 3543
rect 6256 3527 6263 3536
rect 6016 3236 6043 3243
rect 6116 3223 6123 3253
rect 6156 3247 6163 3453
rect 6176 3267 6183 3513
rect 6216 3243 6223 3493
rect 6256 3447 6263 3513
rect 6336 3496 6343 3533
rect 6356 3496 6363 3513
rect 6276 3287 6283 3483
rect 6316 3476 6323 3493
rect 6376 3476 6383 3533
rect 6396 3507 6403 3556
rect 6556 3547 6563 3713
rect 6596 3707 6603 3713
rect 6416 3307 6423 3483
rect 6516 3467 6523 3503
rect 6536 3483 6543 3533
rect 6576 3496 6583 3513
rect 6616 3487 6623 3573
rect 6636 3547 6643 3736
rect 6716 3736 6743 3743
rect 6656 3707 6663 3723
rect 6536 3476 6563 3483
rect 6596 3476 6613 3483
rect 6656 3467 6663 3693
rect 6696 3687 6703 3713
rect 6736 3667 6743 3736
rect 6736 3467 6743 3483
rect 6476 3267 6483 3293
rect 6296 3256 6323 3263
rect 6196 3236 6223 3243
rect 6096 3216 6143 3223
rect 6176 3216 6193 3223
rect 5936 3036 5963 3043
rect 5936 3007 5943 3036
rect 6036 3023 6043 3113
rect 6056 3056 6083 3063
rect 6056 3047 6063 3056
rect 6016 3016 6043 3023
rect 6156 3007 6163 3073
rect 6196 3067 6203 3073
rect 6176 3027 6183 3033
rect 5796 2996 5823 3003
rect 6196 2996 6203 3053
rect 6216 3016 6223 3113
rect 6236 3067 6243 3233
rect 6256 3227 6263 3233
rect 6276 3227 6283 3243
rect 6316 3227 6323 3256
rect 6376 3256 6403 3263
rect 6376 3107 6383 3256
rect 6556 3256 6563 3273
rect 6676 3267 6683 3273
rect 6756 3267 6763 3313
rect 6776 3287 6783 3993
rect 6876 3976 6883 4033
rect 6896 3956 6903 4153
rect 6916 4047 6923 4196
rect 7036 4203 7043 4433
rect 7056 4207 7063 4413
rect 7016 4196 7043 4203
rect 7016 4167 7023 4196
rect 7076 4187 7083 4393
rect 7096 4187 7103 4233
rect 7116 4167 7123 4313
rect 7156 4267 7163 4453
rect 7196 4427 7203 4473
rect 7176 4187 7183 4203
rect 6956 4127 6963 4163
rect 6956 3987 6963 4113
rect 7016 4016 7023 4153
rect 7036 4047 7043 4163
rect 7036 4027 7043 4033
rect 7096 3996 7103 4053
rect 7156 3976 7183 3983
rect 6936 3747 6943 3963
rect 6796 3716 6803 3733
rect 6916 3667 6923 3723
rect 7076 3716 7103 3723
rect 6836 3547 6843 3573
rect 6796 3327 6803 3483
rect 6836 3476 6843 3533
rect 6856 3496 6863 3553
rect 6916 3496 6923 3513
rect 6936 3487 6943 3653
rect 6976 3547 6983 3703
rect 6996 3667 7003 3683
rect 6956 3496 6963 3533
rect 6996 3496 7003 3533
rect 6896 3307 6903 3483
rect 7016 3476 7023 3573
rect 7076 3567 7083 3716
rect 7176 3703 7183 3976
rect 7196 3767 7203 4173
rect 7216 4027 7223 4533
rect 7236 4527 7243 4663
rect 7256 4507 7263 4973
rect 7276 4847 7283 4913
rect 7276 4683 7283 4733
rect 7296 4727 7303 4943
rect 7316 4707 7323 5176
rect 7336 4687 7343 5393
rect 7356 4987 7363 5393
rect 7416 5387 7423 5403
rect 7476 5227 7483 5453
rect 7496 5416 7503 5473
rect 7516 5467 7523 5623
rect 7556 5616 7583 5623
rect 7536 5443 7543 5533
rect 7596 5487 7603 5913
rect 7796 5903 7803 5913
rect 7756 5896 7783 5903
rect 7796 5896 7823 5903
rect 7776 5867 7783 5896
rect 7856 5667 7863 5903
rect 7696 5643 7703 5653
rect 7676 5636 7703 5643
rect 7856 5636 7863 5653
rect 7516 5436 7543 5443
rect 7516 5396 7523 5436
rect 7376 5167 7383 5213
rect 7416 5167 7423 5213
rect 7556 5207 7563 5403
rect 7436 5107 7443 5143
rect 7376 4947 7383 4953
rect 7396 4927 7403 4973
rect 7416 4967 7423 5013
rect 7456 5007 7463 5193
rect 7576 5183 7583 5433
rect 7556 5176 7583 5183
rect 7496 5127 7503 5173
rect 7516 5147 7523 5163
rect 7416 4936 7423 4953
rect 7467 4936 7483 4943
rect 7356 4867 7363 4923
rect 7376 4687 7383 4873
rect 7276 4676 7303 4683
rect 7316 4547 7323 4663
rect 7356 4656 7373 4663
rect 7276 4476 7293 4483
rect 7316 4447 7323 4473
rect 7336 4456 7343 4473
rect 7356 4467 7363 4633
rect 7376 4456 7383 4573
rect 7416 4567 7423 4683
rect 7416 4527 7423 4533
rect 7256 4196 7263 4233
rect 7256 3767 7263 3993
rect 7276 3987 7283 4353
rect 7196 3707 7203 3723
rect 7156 3696 7183 3703
rect 7116 3496 7123 3553
rect 7156 3527 7163 3673
rect 7216 3536 7223 3553
rect 7276 3536 7283 3733
rect 7296 3543 7303 4213
rect 7336 4196 7343 4253
rect 7376 4227 7383 4373
rect 7316 3987 7323 4183
rect 7356 4147 7363 4163
rect 7336 3956 7343 4013
rect 7356 3736 7363 3753
rect 7296 3536 7323 3543
rect 7156 3496 7163 3513
rect 7256 3503 7263 3533
rect 7236 3496 7263 3503
rect 7056 3307 7063 3483
rect 6616 3256 6643 3263
rect 6316 3056 6363 3063
rect 6276 3036 6303 3043
rect 6276 3007 6283 3036
rect 6236 2987 6243 3003
rect 6247 2876 6263 2883
rect 5936 2807 5943 2873
rect 5896 2756 5903 2793
rect 6036 2767 6043 2773
rect 6116 2767 6123 2793
rect 6256 2776 6263 2876
rect 6356 2787 6363 3056
rect 6456 3027 6463 3243
rect 6616 3227 6623 3256
rect 6496 3056 6503 3073
rect 6536 3047 6543 3213
rect 6576 3167 6583 3223
rect 6616 3207 6623 3213
rect 6656 3187 6663 3243
rect 6756 3236 6763 3253
rect 6796 3243 6803 3293
rect 6796 3236 6823 3243
rect 6796 3223 6803 3236
rect 6776 3216 6803 3223
rect 6856 3167 6863 3243
rect 6576 3056 6583 3093
rect 6616 3036 6643 3043
rect 6536 3023 6543 3033
rect 6536 3016 6563 3023
rect 6636 3007 6643 3036
rect 6696 2996 6703 3093
rect 6756 3056 6783 3063
rect 6716 3016 6723 3033
rect 6756 3027 6763 3056
rect 6896 3043 6903 3273
rect 7096 3256 7123 3263
rect 6916 3236 6943 3243
rect 6916 3047 6923 3236
rect 7016 3207 7023 3253
rect 7036 3187 7043 3243
rect 7076 3067 7083 3193
rect 6876 3036 6903 3043
rect 6756 3003 6763 3013
rect 6736 2996 6763 3003
rect 5516 2736 5543 2743
rect 5636 2727 5643 2743
rect 5756 2736 5783 2743
rect 5776 2727 5783 2736
rect 5956 2727 5963 2743
rect 5276 2716 5293 2723
rect 5196 2507 5203 2523
rect 5216 2467 5223 2523
rect 5276 2487 5283 2716
rect 5296 2507 5303 2553
rect 5316 2467 5323 2633
rect 5376 2547 5383 2723
rect 5496 2627 5503 2723
rect 5336 2527 5343 2543
rect 5436 2536 5443 2573
rect 5496 2556 5503 2613
rect 5556 2576 5563 2633
rect 5576 2556 5583 2613
rect 5756 2576 5763 2613
rect 5676 2556 5723 2563
rect 5716 2347 5723 2556
rect 5916 2543 5923 2593
rect 5956 2567 5963 2613
rect 5976 2603 5983 2723
rect 5996 2703 6003 2743
rect 6236 2743 6243 2773
rect 6376 2756 6383 2813
rect 6216 2736 6243 2743
rect 6076 2707 6083 2723
rect 5996 2696 6013 2703
rect 5976 2596 6003 2603
rect 5996 2556 6003 2596
rect 5896 2536 5923 2543
rect 5916 2527 5923 2536
rect 5916 2416 5933 2423
rect 5236 2296 5243 2313
rect 5276 2296 5283 2333
rect 5756 2296 5783 2303
rect 5136 2227 5143 2293
rect 5176 2247 5183 2263
rect 5216 2227 5223 2263
rect 5096 2136 5123 2143
rect 5096 2067 5103 2136
rect 4916 1796 4943 1803
rect 4816 1647 4823 1773
rect 4856 1767 4863 1783
rect 4776 1616 4803 1623
rect 4756 1563 4763 1573
rect 4676 1556 4703 1563
rect 4736 1556 4763 1563
rect 4656 1363 4663 1553
rect 4776 1467 4783 1616
rect 4836 1603 4843 1613
rect 4796 1596 4823 1603
rect 4836 1596 4863 1603
rect 4816 1387 4823 1596
rect 4856 1467 4863 1596
rect 4916 1576 4923 1796
rect 5016 1576 5023 1733
rect 4656 1356 4683 1363
rect 4656 1267 4663 1333
rect 4676 1287 4683 1356
rect 4736 1336 4743 1353
rect 4816 1347 4823 1373
rect 4816 1316 4823 1333
rect 4616 1123 4623 1253
rect 4796 1207 4803 1303
rect 4876 1287 4883 1553
rect 4896 1327 4903 1563
rect 4976 1563 4983 1573
rect 5056 1563 5063 1813
rect 5116 1783 5123 2113
rect 5176 2076 5183 2113
rect 5216 2087 5223 2213
rect 5436 2107 5443 2263
rect 5516 2256 5543 2263
rect 5536 2223 5543 2256
rect 5516 2216 5543 2223
rect 5336 2076 5363 2083
rect 5396 2076 5423 2083
rect 5216 2047 5223 2073
rect 5116 1776 5143 1783
rect 4976 1556 5003 1563
rect 5036 1556 5063 1563
rect 5076 1547 5083 1573
rect 5156 1563 5163 1973
rect 5256 1787 5263 2043
rect 5216 1703 5223 1773
rect 5216 1696 5243 1703
rect 4936 1336 4943 1353
rect 5076 1347 5083 1473
rect 5096 1447 5103 1563
rect 5136 1556 5163 1563
rect 5136 1367 5143 1556
rect 5236 1563 5243 1696
rect 5276 1683 5283 2013
rect 5296 1827 5303 2033
rect 5336 2007 5343 2076
rect 5376 1827 5383 2053
rect 5416 2043 5423 2076
rect 5416 2036 5443 2043
rect 5436 2027 5443 2036
rect 5516 2043 5523 2216
rect 5556 2056 5563 2293
rect 5656 2276 5663 2293
rect 5576 2247 5583 2273
rect 5716 2267 5723 2283
rect 5756 2263 5763 2296
rect 5756 2256 5783 2263
rect 5516 2036 5543 2043
rect 5576 1987 5583 2043
rect 5256 1676 5283 1683
rect 5256 1567 5263 1676
rect 5276 1596 5283 1653
rect 5296 1647 5303 1813
rect 5396 1807 5403 1913
rect 5316 1747 5323 1803
rect 5336 1767 5343 1783
rect 5416 1627 5423 1813
rect 5516 1783 5523 1813
rect 5576 1783 5583 1793
rect 5496 1776 5523 1783
rect 5536 1767 5543 1783
rect 5576 1776 5603 1783
rect 5596 1727 5603 1776
rect 5216 1556 5243 1563
rect 5176 1387 5183 1553
rect 5296 1487 5303 1573
rect 5336 1567 5343 1583
rect 5336 1547 5343 1553
rect 5396 1547 5403 1613
rect 5476 1596 5503 1603
rect 5516 1596 5523 1633
rect 5456 1547 5463 1563
rect 4976 1336 5003 1343
rect 4996 1303 5003 1336
rect 5076 1316 5083 1333
rect 5116 1327 5123 1333
rect 4976 1296 5003 1303
rect 4516 1116 4543 1123
rect 4596 1116 4643 1123
rect 4516 1087 4523 1116
rect 4556 1076 4573 1083
rect 4496 663 4503 803
rect 4516 787 4523 823
rect 4556 787 4563 993
rect 4576 856 4583 1073
rect 4616 856 4623 1116
rect 4756 1116 4763 1193
rect 4956 1127 4963 1293
rect 4676 836 4683 1113
rect 4876 1107 4883 1123
rect 4976 1107 4983 1296
rect 5056 1127 5063 1303
rect 5136 1207 5143 1353
rect 5216 1336 5223 1373
rect 5236 1287 5243 1313
rect 5316 1296 5323 1333
rect 5116 1087 5123 1123
rect 5196 1116 5223 1123
rect 5116 1047 5123 1073
rect 4816 836 4823 853
rect 4876 836 4883 853
rect 5216 847 5223 1116
rect 5356 1087 5363 1193
rect 5376 1136 5383 1333
rect 5416 1103 5423 1313
rect 5456 1107 5463 1493
rect 5496 1287 5503 1596
rect 5596 1576 5603 1693
rect 5616 1607 5623 2233
rect 5636 2047 5643 2083
rect 5716 2076 5723 2093
rect 5776 2027 5783 2256
rect 5796 2247 5803 2273
rect 5876 2267 5883 2293
rect 5836 2096 5863 2103
rect 5836 2047 5843 2096
rect 5916 2076 5923 2416
rect 6016 2287 6023 2693
rect 6196 2627 6203 2723
rect 6356 2667 6363 2753
rect 6136 2576 6143 2593
rect 6096 2523 6103 2573
rect 6156 2556 6163 2573
rect 6356 2556 6363 2653
rect 6456 2563 6463 2573
rect 6436 2556 6463 2563
rect 6076 2516 6103 2523
rect 6096 2296 6103 2493
rect 6196 2307 6203 2543
rect 6496 2536 6503 2773
rect 6576 2747 6583 2873
rect 6596 2727 6603 2973
rect 6796 2807 6803 3023
rect 6656 2707 6663 2783
rect 6796 2776 6823 2783
rect 6676 2747 6683 2763
rect 6716 2756 6723 2773
rect 6816 2727 6823 2776
rect 6876 2767 6883 3036
rect 6956 3036 6983 3043
rect 6936 3007 6943 3023
rect 6916 2743 6923 2793
rect 6936 2747 6943 2993
rect 6976 2987 6983 3036
rect 7016 3036 7043 3043
rect 6996 2756 7003 2793
rect 7016 2787 7023 3036
rect 7116 3027 7123 3256
rect 7136 3243 7143 3353
rect 7176 3267 7183 3483
rect 7316 3247 7323 3536
rect 7336 3263 7343 3723
rect 7376 3567 7383 3963
rect 7396 3743 7403 4443
rect 7416 4227 7423 4493
rect 7436 4427 7443 4513
rect 7456 4487 7463 4853
rect 7476 4707 7483 4913
rect 7476 4667 7483 4693
rect 7476 4587 7483 4653
rect 7496 4503 7503 4913
rect 7516 4887 7523 5113
rect 7536 4987 7543 5013
rect 7556 4987 7563 5176
rect 7596 5167 7603 5233
rect 7596 5027 7603 5123
rect 7616 5107 7623 5143
rect 7636 5127 7643 5393
rect 7536 4923 7543 4953
rect 7536 4916 7563 4923
rect 7516 4527 7523 4833
rect 7536 4747 7543 4893
rect 7556 4867 7563 4916
rect 7596 4887 7603 4923
rect 7636 4916 7643 4973
rect 7656 4936 7663 5623
rect 7676 5007 7683 5613
rect 7696 5087 7703 5593
rect 7756 5587 7763 5603
rect 7716 5403 7723 5433
rect 7756 5427 7763 5473
rect 7776 5467 7783 5573
rect 7836 5527 7843 5603
rect 7776 5407 7783 5453
rect 7796 5447 7803 5513
rect 7796 5416 7803 5433
rect 7716 5396 7743 5403
rect 7716 5176 7723 5193
rect 7736 5147 7743 5163
rect 7776 5127 7783 5173
rect 7896 5167 7903 5916
rect 7696 4923 7703 4973
rect 7676 4916 7703 4923
rect 7536 4696 7543 4713
rect 7596 4687 7603 4713
rect 7636 4687 7643 4733
rect 7676 4727 7683 4916
rect 7736 4747 7743 5073
rect 7776 4956 7783 5093
rect 7796 4947 7803 5133
rect 7816 5107 7823 5163
rect 7916 5147 7923 5433
rect 7836 4987 7843 5143
rect 7816 4956 7823 4973
rect 7856 4956 7863 5073
rect 7876 4936 7883 5113
rect 7756 4887 7763 4923
rect 7676 4707 7683 4713
rect 7756 4696 7763 4753
rect 7556 4547 7563 4683
rect 7576 4547 7583 4653
rect 7556 4507 7563 4513
rect 7476 4496 7503 4503
rect 7476 4476 7483 4496
rect 7547 4476 7553 4483
rect 7436 4267 7443 4393
rect 7456 4207 7463 4453
rect 7476 4327 7483 4433
rect 7496 4427 7503 4463
rect 7536 4456 7563 4463
rect 7556 4407 7563 4456
rect 7476 4227 7483 4293
rect 7416 4127 7423 4193
rect 7476 4167 7483 4183
rect 7436 3976 7443 4153
rect 7456 4127 7463 4163
rect 7456 4007 7463 4113
rect 7496 4023 7503 4193
rect 7476 4016 7503 4023
rect 7416 3947 7423 3963
rect 7456 3927 7463 3953
rect 7476 3743 7483 4016
rect 7496 3967 7503 3993
rect 7516 3767 7523 4253
rect 7536 4227 7543 4393
rect 7556 4367 7563 4373
rect 7576 4227 7583 4513
rect 7596 4443 7603 4553
rect 7636 4503 7643 4573
rect 7656 4527 7663 4663
rect 7676 4647 7683 4693
rect 7696 4676 7723 4683
rect 7716 4667 7723 4676
rect 7696 4623 7703 4653
rect 7676 4616 7703 4623
rect 7636 4496 7663 4503
rect 7656 4456 7663 4496
rect 7676 4467 7683 4616
rect 7596 4436 7623 4443
rect 7596 4387 7603 4413
rect 7616 4307 7623 4436
rect 7636 4427 7643 4453
rect 7616 4203 7623 4233
rect 7636 4207 7643 4393
rect 7676 4247 7683 4273
rect 7596 4196 7623 4203
rect 7576 4007 7583 4183
rect 7596 4007 7603 4173
rect 7616 4103 7623 4173
rect 7616 4096 7643 4103
rect 7616 4007 7623 4013
rect 7547 3996 7553 4003
rect 7536 3947 7543 3973
rect 7556 3927 7563 3963
rect 7536 3787 7543 3913
rect 7567 3776 7573 3783
rect 7596 3767 7603 3833
rect 7616 3767 7623 3913
rect 7636 3747 7643 4096
rect 7656 3987 7663 4153
rect 7676 4027 7683 4213
rect 7696 4027 7703 4413
rect 7716 4267 7723 4443
rect 7716 4067 7723 4233
rect 7736 4147 7743 4493
rect 7756 4483 7763 4533
rect 7776 4507 7783 4733
rect 7796 4543 7803 4933
rect 7816 4707 7823 4913
rect 7856 4696 7863 4713
rect 7836 4543 7843 4683
rect 7796 4536 7823 4543
rect 7836 4536 7863 4543
rect 7816 4487 7823 4536
rect 7836 4496 7843 4513
rect 7856 4507 7863 4536
rect 7756 4476 7783 4483
rect 7756 4247 7763 4453
rect 7776 4227 7783 4433
rect 7816 4227 7823 4433
rect 7836 4227 7843 4453
rect 7856 4227 7863 4463
rect 7876 4407 7883 4513
rect 7896 4287 7903 4993
rect 7716 4016 7723 4033
rect 7736 4023 7743 4133
rect 7756 4047 7763 4173
rect 7736 4016 7763 4023
rect 7756 3987 7763 4016
rect 7776 4007 7783 4153
rect 7816 4147 7823 4183
rect 7816 4027 7823 4093
rect 7836 4047 7843 4173
rect 7856 4107 7863 4163
rect 7856 4027 7863 4053
rect 7656 3867 7663 3973
rect 7687 3956 7693 3963
rect 7396 3736 7423 3743
rect 7456 3736 7483 3743
rect 7396 3543 7403 3736
rect 7436 3567 7443 3723
rect 7476 3563 7483 3736
rect 7496 3736 7523 3743
rect 7496 3583 7503 3736
rect 7536 3716 7563 3723
rect 7556 3707 7563 3716
rect 7496 3576 7523 3583
rect 7476 3556 7503 3563
rect 7376 3536 7403 3543
rect 7336 3256 7363 3263
rect 7136 3236 7163 3243
rect 7096 3016 7113 3023
rect 7136 2996 7143 3053
rect 7176 3043 7183 3223
rect 7216 3207 7223 3223
rect 7236 3047 7243 3233
rect 7296 3207 7303 3223
rect 7356 3207 7363 3256
rect 7276 3187 7283 3203
rect 7176 3036 7203 3043
rect 7156 3016 7163 3033
rect 7056 2763 7063 2973
rect 7036 2756 7063 2763
rect 6896 2736 6923 2743
rect 6576 2587 6583 2633
rect 6296 2296 6323 2303
rect 6356 2296 6373 2303
rect 6296 2267 6303 2296
rect 5956 2107 5963 2263
rect 5996 2227 6003 2263
rect 6216 2247 6223 2263
rect 5556 1547 5563 1573
rect 5636 1563 5643 1873
rect 5676 1796 5683 1813
rect 5716 1767 5723 1783
rect 5736 1747 5743 1763
rect 5756 1687 5763 1833
rect 5776 1796 5803 1803
rect 5776 1747 5783 1796
rect 5896 1787 5903 1803
rect 5836 1767 5843 1783
rect 5816 1747 5823 1763
rect 5696 1616 5703 1653
rect 5876 1627 5883 1783
rect 5896 1747 5903 1773
rect 5576 1507 5583 1563
rect 5616 1556 5643 1563
rect 5636 1367 5643 1556
rect 5536 1303 5543 1333
rect 5536 1296 5563 1303
rect 5656 1303 5663 1553
rect 5676 1487 5683 1583
rect 5676 1347 5683 1473
rect 5696 1307 5703 1453
rect 5636 1296 5663 1303
rect 5656 1136 5683 1143
rect 5656 1127 5663 1136
rect 5396 1096 5423 1103
rect 5356 856 5363 1073
rect 5436 1047 5443 1083
rect 5476 1047 5483 1073
rect 5596 1067 5603 1103
rect 5656 1083 5663 1113
rect 5636 1076 5663 1083
rect 5596 987 5603 1053
rect 5136 807 5143 823
rect 5276 823 5283 853
rect 5256 816 5283 823
rect 4476 656 4503 663
rect 4076 636 4103 643
rect 4096 623 4103 636
rect 4356 636 4383 643
rect 4236 627 4243 633
rect 4096 616 4123 623
rect 4096 587 4103 616
rect 4236 603 4243 613
rect 4216 596 4243 603
rect 3996 363 4003 373
rect 3996 356 4023 363
rect 4056 356 4063 393
rect 4076 327 4083 343
rect 4096 307 4103 553
rect 4116 447 4123 573
rect 4376 567 4383 636
rect 4436 616 4443 653
rect 4056 136 4063 273
rect 4096 167 4103 293
rect 4116 247 4123 393
rect 4136 376 4143 433
rect 4176 376 4203 383
rect 4116 156 4123 233
rect 4156 187 4163 363
rect 4196 327 4203 376
rect 4216 356 4223 433
rect 4276 227 4283 343
rect 4296 207 4303 353
rect 4316 287 4323 373
rect 4356 356 4363 493
rect 4416 447 4423 603
rect 4456 596 4463 653
rect 4476 616 4483 656
rect 4516 643 4523 673
rect 4596 663 4603 773
rect 4576 656 4603 663
rect 4716 656 4723 693
rect 4496 636 4523 643
rect 4476 376 4483 453
rect 4496 407 4503 636
rect 4416 347 4423 363
rect 4336 267 4343 343
rect 4376 287 4383 323
rect 4176 136 4183 193
rect 4316 156 4323 193
rect 4436 187 4443 353
rect 4516 347 4523 593
rect 4576 487 4583 656
rect 4696 507 4703 623
rect 4776 547 4783 653
rect 4816 616 4823 633
rect 4376 156 4403 163
rect 4276 107 4283 143
rect 4396 -24 4403 156
rect 4456 156 4463 173
rect 4536 156 4543 253
rect 4576 247 4583 353
rect 4596 347 4603 383
rect 4636 363 4643 433
rect 4776 427 4783 513
rect 4616 356 4643 363
rect 4476 127 4483 143
rect 4556 123 4563 233
rect 4636 123 4643 293
rect 4676 187 4683 363
rect 4716 347 4723 373
rect 4736 356 4743 373
rect 4556 116 4583 123
rect 4616 116 4643 123
rect 4656 156 4683 163
rect 4656 -24 4663 156
rect 4696 147 4703 253
rect 4716 156 4723 253
rect 4756 127 4763 313
rect 4776 167 4783 413
rect 4796 407 4803 603
rect 4836 596 4843 693
rect 4976 636 4983 673
rect 4996 667 5003 713
rect 5076 656 5103 663
rect 4996 636 5003 653
rect 4856 616 4883 623
rect 4816 307 4823 573
rect 4876 527 4883 616
rect 4896 616 4923 623
rect 4896 587 4903 616
rect 4956 567 4963 623
rect 4836 376 4843 473
rect 4896 383 4903 533
rect 4876 376 4903 383
rect 4936 376 4943 413
rect 4896 327 4903 376
rect 4916 307 4923 343
rect 4956 267 4963 553
rect 4816 156 4823 253
rect 4856 156 4863 173
rect 4956 123 4963 213
rect 4976 187 4983 343
rect 4996 156 5003 453
rect 5016 227 5023 623
rect 5076 607 5083 656
rect 5076 447 5083 593
rect 5136 427 5143 653
rect 5176 507 5183 673
rect 5276 656 5283 816
rect 5196 636 5223 643
rect 5196 627 5203 636
rect 5356 636 5363 693
rect 5396 656 5403 713
rect 5436 647 5443 933
rect 5476 836 5483 973
rect 5516 847 5523 853
rect 5456 807 5463 823
rect 5176 403 5183 493
rect 5176 396 5203 403
rect 5056 227 5063 363
rect 5136 356 5143 393
rect 5156 287 5163 343
rect 5176 327 5183 373
rect 5136 167 5143 193
rect 5016 156 5043 163
rect 5076 156 5103 163
rect 4936 116 4963 123
rect 5016 -24 5023 156
rect 5076 127 5083 156
rect 5176 147 5183 253
rect 5196 163 5203 396
rect 5256 376 5263 533
rect 5296 527 5303 623
rect 5416 607 5423 623
rect 5456 607 5463 643
rect 5536 636 5543 813
rect 5556 627 5563 973
rect 5636 887 5643 1076
rect 5716 1067 5723 1303
rect 5736 1147 5743 1353
rect 5796 1327 5803 1593
rect 5836 1576 5843 1613
rect 5916 1567 5923 1973
rect 6016 1887 6023 2053
rect 6116 2043 6123 2173
rect 6216 2163 6223 2233
rect 6256 2227 6263 2263
rect 6376 2247 6383 2293
rect 6216 2156 6243 2163
rect 6216 2076 6223 2113
rect 6056 2027 6063 2043
rect 6096 2036 6123 2043
rect 6136 2056 6163 2063
rect 6136 1947 6143 2056
rect 6236 1987 6243 2156
rect 6396 2096 6403 2113
rect 6356 2076 6363 2093
rect 6416 2087 6423 2093
rect 6336 2047 6343 2073
rect 5996 1783 6003 1853
rect 6056 1847 6063 1853
rect 6016 1816 6023 1833
rect 6056 1816 6063 1833
rect 6036 1787 6043 1803
rect 6156 1796 6183 1803
rect 5936 1687 5943 1783
rect 5976 1776 6003 1783
rect 5936 1587 5943 1633
rect 5956 1596 5963 1633
rect 5976 1616 5983 1653
rect 6076 1647 6083 1793
rect 6136 1616 6143 1633
rect 6007 1596 6023 1603
rect 6016 1587 6023 1596
rect 6096 1596 6123 1603
rect 6156 1596 6163 1673
rect 6176 1627 6183 1796
rect 6196 1787 6203 1853
rect 6316 1843 6323 2033
rect 6316 1836 6343 1843
rect 6256 1783 6263 1813
rect 6256 1776 6283 1783
rect 6216 1667 6223 1763
rect 5876 1487 5883 1553
rect 5876 1303 5883 1473
rect 6096 1387 6103 1596
rect 6236 1576 6243 1613
rect 6276 1563 6283 1673
rect 6336 1667 6343 1836
rect 6376 1767 6383 1813
rect 6396 1607 6403 1993
rect 6436 1847 6443 2513
rect 6536 2427 6543 2543
rect 6487 2416 6493 2423
rect 6496 2296 6523 2303
rect 6516 2263 6523 2296
rect 6516 2256 6543 2263
rect 6516 2187 6523 2256
rect 6456 2076 6483 2083
rect 6536 2076 6543 2113
rect 6456 1807 6463 2076
rect 6476 1796 6483 1973
rect 6556 1816 6563 1833
rect 6416 1727 6423 1783
rect 6496 1767 6503 1793
rect 6576 1707 6583 2493
rect 6636 2263 6643 2653
rect 6656 2507 6663 2613
rect 6736 2576 6743 2613
rect 6616 2256 6643 2263
rect 6636 2147 6643 2256
rect 6636 2096 6643 2113
rect 6676 2063 6683 2333
rect 6756 2267 6763 2273
rect 6776 2267 6783 2573
rect 6796 2556 6803 2613
rect 6836 2556 6843 2633
rect 6896 2507 6903 2563
rect 6956 2547 6963 2753
rect 7016 2707 7023 2743
rect 7076 2736 7103 2743
rect 6976 2556 6983 2653
rect 7016 2556 7023 2613
rect 7076 2527 7083 2736
rect 7176 2667 7183 2743
rect 7196 2727 7203 3036
rect 7256 3016 7263 3073
rect 7216 3003 7223 3013
rect 7216 2996 7243 3003
rect 7276 2807 7283 2993
rect 6896 2296 6923 2303
rect 6956 2296 6963 2333
rect 7136 2307 7143 2573
rect 7176 2556 7183 2593
rect 7216 2556 7223 2613
rect 7296 2607 7303 3033
rect 7156 2487 7163 2553
rect 7236 2507 7243 2543
rect 7296 2536 7303 2573
rect 7316 2567 7323 2773
rect 7336 2527 7343 3093
rect 7376 3083 7383 3233
rect 7396 3223 7403 3513
rect 7416 3267 7423 3553
rect 7476 3516 7483 3533
rect 7496 3496 7503 3556
rect 7516 3307 7523 3576
rect 7556 3287 7563 3553
rect 7576 3527 7583 3693
rect 7596 3547 7603 3733
rect 7656 3716 7663 3833
rect 7676 3747 7683 3873
rect 7636 3547 7643 3683
rect 7596 3496 7603 3513
rect 7636 3483 7643 3533
rect 7616 3476 7643 3483
rect 7656 3483 7663 3533
rect 7676 3507 7683 3553
rect 7696 3527 7703 3933
rect 7716 3647 7723 3973
rect 7736 3947 7743 3983
rect 7716 3536 7723 3553
rect 7736 3547 7743 3853
rect 7756 3767 7763 3953
rect 7776 3887 7783 3993
rect 7796 3967 7803 4013
rect 7796 3827 7803 3933
rect 7836 3747 7843 3933
rect 7756 3547 7763 3733
rect 7816 3716 7823 3733
rect 7776 3527 7783 3693
rect 7796 3667 7803 3703
rect 7796 3527 7803 3633
rect 7736 3516 7763 3523
rect 7756 3507 7763 3516
rect 7836 3516 7843 3693
rect 7856 3567 7863 3953
rect 7876 3543 7883 4033
rect 7896 3707 7903 4213
rect 7916 3847 7923 4753
rect 7856 3536 7883 3543
rect 7656 3476 7683 3483
rect 7576 3263 7583 3473
rect 7396 3216 7423 3223
rect 7356 3076 7383 3083
rect 7356 3036 7363 3076
rect 7396 3036 7403 3073
rect 7416 3043 7423 3216
rect 7436 3067 7443 3203
rect 7456 3187 7463 3223
rect 7456 3067 7463 3173
rect 7476 3107 7483 3253
rect 7416 3036 7443 3043
rect 7476 3036 7493 3043
rect 7516 3023 7523 3263
rect 7556 3256 7583 3263
rect 7536 3087 7543 3243
rect 7596 3067 7603 3293
rect 7616 3067 7623 3253
rect 7636 3207 7643 3223
rect 7656 3087 7663 3453
rect 7676 3287 7683 3476
rect 7716 3267 7723 3493
rect 7676 3236 7683 3253
rect 7736 3236 7743 3453
rect 7496 3016 7523 3023
rect 7376 2756 7383 3013
rect 7516 2987 7523 3016
rect 7536 2927 7543 3013
rect 7447 2876 7463 2883
rect 7456 2776 7463 2876
rect 7496 2776 7503 2793
rect 7356 2727 7363 2743
rect 7416 2663 7423 2763
rect 7396 2656 7423 2663
rect 7396 2587 7403 2656
rect 7436 2607 7443 2613
rect 7316 2507 7323 2523
rect 6856 2276 6863 2293
rect 6827 2256 6843 2263
rect 6776 2123 6783 2253
rect 6876 2247 6883 2263
rect 6756 2116 6783 2123
rect 6756 2107 6763 2116
rect 6736 2067 6743 2093
rect 6756 2076 6763 2093
rect 6656 2056 6683 2063
rect 6656 1987 6663 2056
rect 6596 1807 6603 1973
rect 6696 1807 6703 2063
rect 6816 2043 6823 2233
rect 6856 2056 6863 2213
rect 6896 2127 6903 2296
rect 6976 2247 6983 2293
rect 7016 2247 7023 2283
rect 6916 2047 6923 2083
rect 6816 2036 6843 2043
rect 6616 1763 6623 1783
rect 6656 1767 6663 1773
rect 6616 1756 6643 1763
rect 6636 1667 6643 1756
rect 6476 1616 6483 1653
rect 6356 1596 6383 1603
rect 6216 1387 6223 1563
rect 6256 1556 6283 1563
rect 6376 1347 6383 1596
rect 6436 1596 6463 1603
rect 6496 1596 6503 1653
rect 6596 1616 6603 1633
rect 6636 1616 6643 1653
rect 6436 1587 6443 1596
rect 6556 1547 6563 1613
rect 6616 1596 6623 1613
rect 6656 1603 6663 1653
rect 6676 1647 6683 1803
rect 6716 1667 6723 2033
rect 6656 1596 6683 1603
rect 6676 1567 6683 1596
rect 6716 1576 6723 1633
rect 6736 1603 6743 1873
rect 6756 1796 6763 1813
rect 6796 1796 6803 1853
rect 6836 1783 6843 1813
rect 6876 1783 6883 1833
rect 6936 1783 6943 1853
rect 6976 1823 6983 2093
rect 6996 2076 7003 2133
rect 7036 2076 7043 2153
rect 7056 2087 7063 2293
rect 7136 2276 7143 2293
rect 7196 2243 7203 2493
rect 7236 2276 7243 2473
rect 7256 2243 7263 2333
rect 7316 2307 7323 2493
rect 7196 2236 7223 2243
rect 7256 2236 7283 2243
rect 6816 1776 6843 1783
rect 6856 1776 6883 1783
rect 6916 1776 6943 1783
rect 6956 1816 6983 1823
rect 7016 1823 7023 2033
rect 7016 1816 7043 1823
rect 6956 1627 6963 1816
rect 7036 1687 7043 1816
rect 7056 1807 7063 2053
rect 6736 1596 6763 1603
rect 6696 1547 6703 1563
rect 6296 1336 6323 1343
rect 6296 1323 6303 1336
rect 6276 1316 6303 1323
rect 5876 1296 5903 1303
rect 5936 1287 5943 1303
rect 5956 1296 5983 1303
rect 5776 1096 5783 1253
rect 5896 1116 5903 1153
rect 5756 1047 5763 1083
rect 5656 856 5663 953
rect 5796 947 5803 1073
rect 5876 1047 5883 1103
rect 5236 327 5243 363
rect 5196 156 5223 163
rect 5256 156 5263 233
rect 5316 187 5323 413
rect 5336 376 5343 573
rect 5556 407 5563 613
rect 5276 136 5283 173
rect 5456 167 5463 343
rect 5496 267 5503 343
rect 5516 327 5523 353
rect 5396 127 5403 163
rect 5476 156 5483 193
rect 5516 156 5523 273
rect 5576 247 5583 343
rect 5616 163 5623 373
rect 5636 207 5643 813
rect 5676 807 5683 833
rect 5756 816 5763 853
rect 5836 687 5843 813
rect 5856 603 5863 1033
rect 5936 887 5943 1273
rect 5956 1087 5963 1296
rect 6056 1247 6063 1303
rect 6076 1096 6083 1173
rect 6136 1136 6143 1173
rect 5836 596 5863 603
rect 5896 603 5903 853
rect 5936 616 5943 833
rect 5896 596 5923 603
rect 5856 487 5863 596
rect 5956 587 5963 603
rect 5976 547 5983 953
rect 5996 907 6003 1053
rect 6016 1023 6023 1083
rect 6036 1067 6043 1093
rect 6056 1023 6063 1083
rect 6096 1076 6103 1133
rect 6116 1096 6123 1133
rect 6156 1047 6163 1093
rect 6196 1067 6203 1313
rect 6296 1267 6303 1316
rect 6336 1267 6343 1323
rect 6436 1316 6463 1323
rect 6376 1287 6383 1313
rect 6416 1267 6423 1283
rect 6216 1116 6223 1153
rect 6296 1127 6303 1173
rect 6356 1136 6363 1173
rect 6376 1147 6383 1253
rect 6376 1116 6383 1133
rect 6396 1116 6403 1173
rect 6436 1116 6443 1213
rect 6456 1167 6463 1316
rect 6296 1047 6303 1113
rect 6016 1016 6063 1023
rect 6036 836 6043 893
rect 6156 823 6163 873
rect 6196 856 6223 863
rect 6136 816 6163 823
rect 6056 616 6063 793
rect 6016 603 6023 613
rect 6016 596 6043 603
rect 6096 587 6103 813
rect 6176 807 6183 823
rect 6196 807 6203 856
rect 6176 767 6183 793
rect 6236 727 6243 823
rect 6136 627 6143 653
rect 6196 636 6223 643
rect 6256 636 6263 1033
rect 6316 987 6323 1093
rect 6416 1087 6423 1103
rect 6456 1096 6483 1103
rect 6376 856 6403 863
rect 6376 827 6383 856
rect 6456 827 6463 953
rect 6476 847 6483 1096
rect 6496 967 6503 1333
rect 6616 1307 6623 1333
rect 6276 767 6283 823
rect 6316 807 6323 823
rect 6516 823 6523 873
rect 6536 867 6543 1293
rect 6696 1287 6703 1303
rect 6656 1096 6663 1253
rect 6696 1247 6703 1273
rect 6736 1227 6743 1303
rect 6556 1047 6563 1083
rect 6556 863 6563 1033
rect 6596 1007 6603 1083
rect 6636 1047 6643 1083
rect 6676 1047 6683 1083
rect 6556 856 6583 863
rect 6516 816 6533 823
rect 6296 707 6303 803
rect 5696 363 5703 473
rect 5856 387 5863 473
rect 5696 356 5723 363
rect 5756 356 5763 373
rect 5796 347 5803 353
rect 5676 307 5683 323
rect 5736 267 5743 343
rect 5776 336 5793 343
rect 5816 307 5823 373
rect 6036 356 6043 553
rect 6116 547 6123 603
rect 5836 247 5843 323
rect 5996 287 6003 343
rect 6076 227 6083 323
rect 5616 156 5643 163
rect 5716 156 5723 193
rect 5976 156 5983 193
rect 6136 187 6143 573
rect 6156 187 6163 603
rect 6196 567 6203 636
rect 6196 207 6203 323
rect 6236 307 6243 623
rect 6276 616 6283 633
rect 6316 627 6323 713
rect 6336 387 6343 593
rect 6416 463 6423 653
rect 6436 627 6443 653
rect 6456 636 6463 693
rect 6496 636 6503 713
rect 6396 456 6423 463
rect 6376 376 6383 413
rect 6316 323 6323 333
rect 6296 316 6323 323
rect 6356 176 6363 273
rect 6396 207 6403 456
rect 6556 447 6563 623
rect 6576 607 6583 856
rect 6596 816 6623 823
rect 6596 507 6603 816
rect 6676 787 6683 1033
rect 6716 1007 6723 1123
rect 6696 687 6703 823
rect 6736 743 6743 823
rect 6756 807 6763 1596
rect 6796 1596 6823 1603
rect 6836 1596 6863 1603
rect 6896 1596 6903 1613
rect 6796 1367 6803 1596
rect 6836 1263 6843 1596
rect 6836 1256 6863 1263
rect 6796 1116 6823 1123
rect 6716 736 6743 743
rect 6716 636 6723 736
rect 6456 376 6463 393
rect 6436 327 6443 363
rect 6476 327 6483 373
rect 6496 327 6503 393
rect 6556 356 6563 393
rect 6076 163 6083 173
rect 6056 156 6083 163
rect 6176 156 6183 173
rect 6256 156 6283 163
rect 6276 127 6283 156
rect 6296 147 6303 173
rect 6476 156 6483 273
rect 6576 263 6583 343
rect 6596 287 6603 433
rect 6616 403 6623 633
rect 6736 607 6743 623
rect 6776 607 6783 613
rect 6796 607 6803 1053
rect 6816 687 6823 1116
rect 6676 507 6683 603
rect 6616 396 6643 403
rect 6616 287 6623 373
rect 6636 347 6643 396
rect 6696 376 6703 573
rect 6736 407 6743 593
rect 6836 587 6843 1073
rect 6856 827 6863 1256
rect 6896 1047 6903 1293
rect 6916 1107 6923 1373
rect 6936 1287 6943 1303
rect 6956 1143 6963 1353
rect 7036 1287 7043 1633
rect 7056 1596 7063 1633
rect 6936 1136 6963 1143
rect 6936 1087 6943 1136
rect 7036 1127 7043 1273
rect 7056 1147 7063 1333
rect 7076 1327 7083 1753
rect 7136 1647 7143 2133
rect 7156 2047 7163 2083
rect 7196 1887 7203 2236
rect 7236 2076 7243 2133
rect 7156 1767 7163 1783
rect 7196 1747 7203 1783
rect 7156 1616 7183 1623
rect 7136 1547 7143 1603
rect 7156 1547 7163 1616
rect 7136 1336 7143 1373
rect 7216 1347 7223 1873
rect 7276 1767 7283 1783
rect 7236 1743 7243 1753
rect 7296 1747 7303 2113
rect 7336 1847 7343 2313
rect 7356 2267 7363 2553
rect 7376 2536 7383 2553
rect 7416 2536 7423 2593
rect 7456 2527 7463 2733
rect 7476 2607 7483 2763
rect 7516 2643 7523 2773
rect 7496 2636 7523 2643
rect 7496 2607 7503 2636
rect 7376 2127 7383 2493
rect 7436 2327 7443 2523
rect 7456 2303 7463 2493
rect 7476 2407 7483 2553
rect 7496 2547 7503 2563
rect 7436 2296 7463 2303
rect 7396 2227 7403 2283
rect 7436 2276 7443 2296
rect 7416 2167 7423 2263
rect 7476 2107 7483 2293
rect 7476 2076 7483 2093
rect 7496 2047 7503 2513
rect 7536 2347 7543 2893
rect 7556 2776 7563 2973
rect 7596 2776 7603 2913
rect 7556 2563 7563 2653
rect 7576 2583 7583 2763
rect 7616 2583 7623 3033
rect 7636 2787 7643 3053
rect 7676 2987 7683 3023
rect 7656 2756 7663 2873
rect 7696 2756 7703 3073
rect 7716 2783 7723 3093
rect 7756 3043 7763 3473
rect 7816 3467 7823 3493
rect 7827 3356 7843 3363
rect 7796 3067 7803 3273
rect 7816 3087 7823 3273
rect 7836 3256 7843 3356
rect 7856 3287 7863 3493
rect 7876 3487 7883 3503
rect 7856 3107 7863 3243
rect 7736 3036 7763 3043
rect 7736 2907 7743 3036
rect 7836 3036 7843 3053
rect 7856 3027 7863 3073
rect 7756 3016 7783 3023
rect 7756 2887 7763 3016
rect 7747 2876 7753 2883
rect 7796 2807 7803 2993
rect 7816 2787 7823 3013
rect 7716 2776 7743 2783
rect 7736 2743 7743 2776
rect 7576 2576 7603 2583
rect 7616 2576 7643 2583
rect 7556 2556 7583 2563
rect 7596 2327 7603 2576
rect 7636 2527 7643 2576
rect 7676 2567 7683 2743
rect 7716 2736 7743 2743
rect 7756 2567 7763 2773
rect 7836 2756 7843 2873
rect 7856 2727 7863 2743
rect 7776 2556 7783 2713
rect 7576 2296 7583 2313
rect 7616 2296 7623 2513
rect 7516 2096 7523 2113
rect 7576 2083 7583 2253
rect 7596 2127 7603 2283
rect 7576 2076 7603 2083
rect 7536 2047 7543 2063
rect 7316 1767 7323 1813
rect 7416 1796 7423 1853
rect 7336 1767 7343 1773
rect 7236 1736 7273 1743
rect 7327 1736 7333 1743
rect 7236 1596 7243 1613
rect 7316 1596 7343 1603
rect 7336 1567 7343 1596
rect 7356 1387 7363 1763
rect 7376 1747 7383 1783
rect 7396 1747 7403 1783
rect 7376 1587 7383 1613
rect 7336 1336 7343 1353
rect 7376 1336 7383 1533
rect 7396 1367 7403 1653
rect 7436 1627 7443 1783
rect 7476 1667 7483 1833
rect 7536 1827 7543 2033
rect 7576 1887 7583 2076
rect 7636 2067 7643 2313
rect 7456 1616 7463 1633
rect 7516 1603 7523 1633
rect 7576 1607 7583 1853
rect 7656 1827 7663 2333
rect 7736 2227 7743 2263
rect 7776 2147 7783 2263
rect 7676 2076 7683 2133
rect 7716 2076 7723 2113
rect 7516 1596 7543 1603
rect 7536 1587 7543 1596
rect 7556 1567 7563 1583
rect 7396 1336 7423 1343
rect 7456 1336 7483 1343
rect 6976 1067 6983 1103
rect 7056 1096 7063 1133
rect 7116 1067 7123 1273
rect 7136 1087 7143 1123
rect 7176 867 7183 1333
rect 7276 1316 7303 1323
rect 7196 1287 7203 1313
rect 7296 1267 7303 1316
rect 7356 1287 7363 1323
rect 7396 1287 7403 1336
rect 7196 1116 7223 1123
rect 7256 1116 7263 1133
rect 6996 856 7023 863
rect 7056 856 7083 863
rect 6876 616 6883 693
rect 6936 627 6943 653
rect 6916 587 6923 603
rect 6576 256 6603 263
rect 6556 207 6563 253
rect 6556 156 6563 193
rect 6576 176 6583 233
rect 6596 207 6603 256
rect 6596 156 6603 173
rect 6616 156 6623 213
rect 6636 203 6643 333
rect 6676 327 6683 363
rect 6676 227 6683 293
rect 6636 196 6663 203
rect 6656 156 6663 196
rect 6396 143 6403 153
rect 6676 147 6683 213
rect 6736 187 6743 373
rect 6756 287 6763 343
rect 6696 156 6703 173
rect 6776 167 6783 413
rect 6976 387 6983 853
rect 6996 827 7003 856
rect 7076 823 7083 856
rect 7076 816 7103 823
rect 6916 343 6923 373
rect 6856 287 6863 343
rect 6896 336 6923 343
rect 6936 327 6943 343
rect 6836 176 6843 253
rect 6996 167 7003 673
rect 7016 667 7023 813
rect 7016 603 7023 653
rect 7076 647 7083 816
rect 7116 607 7123 643
rect 7016 596 7043 603
rect 7156 407 7163 713
rect 7176 687 7183 823
rect 7196 687 7203 1116
rect 7196 636 7203 673
rect 7056 356 7063 373
rect 7096 343 7103 373
rect 7076 336 7103 343
rect 7116 343 7123 393
rect 7116 336 7143 343
rect 7216 327 7223 673
rect 7276 376 7303 383
rect 7296 367 7303 376
rect 7256 347 7263 363
rect 7316 327 7323 1113
rect 7356 827 7363 843
rect 7396 667 7403 1083
rect 7416 867 7423 1293
rect 7476 1267 7483 1336
rect 7496 1287 7503 1373
rect 7436 907 7443 1173
rect 7456 1087 7463 1193
rect 7476 1127 7483 1233
rect 7516 1227 7523 1353
rect 7556 1316 7563 1333
rect 7576 1307 7583 1573
rect 7596 1367 7603 1733
rect 7616 1367 7623 1813
rect 7636 1727 7643 1783
rect 7676 1747 7683 1783
rect 7776 1767 7783 2053
rect 7676 1596 7683 1713
rect 7736 1627 7743 1763
rect 7776 1623 7783 1733
rect 7796 1647 7803 2293
rect 7756 1616 7783 1623
rect 7716 1596 7723 1613
rect 7756 1567 7763 1616
rect 7596 1143 7603 1333
rect 7676 1303 7683 1333
rect 7696 1327 7703 1553
rect 7656 1296 7683 1303
rect 7616 1167 7623 1213
rect 7636 1163 7643 1283
rect 7636 1156 7653 1163
rect 7556 1136 7603 1143
rect 7496 1116 7503 1133
rect 7536 1116 7543 1133
rect 7556 1116 7563 1136
rect 7616 1123 7623 1133
rect 7596 1116 7623 1123
rect 7576 1087 7583 1103
rect 7336 427 7343 653
rect 7416 636 7423 653
rect 7376 376 7383 393
rect 7156 227 7163 323
rect 7396 207 7403 413
rect 7436 387 7443 873
rect 7456 867 7463 1073
rect 7476 847 7483 893
rect 7516 856 7523 873
rect 7556 856 7563 873
rect 7536 827 7543 843
rect 7476 727 7483 803
rect 7456 407 7463 653
rect 7496 643 7503 753
rect 7576 747 7583 853
rect 7476 636 7503 643
rect 7476 603 7483 636
rect 7576 623 7583 713
rect 7596 667 7603 1073
rect 7636 887 7643 1156
rect 7676 1136 7683 1173
rect 7716 1163 7723 1353
rect 7776 1303 7783 1573
rect 7816 1327 7823 2713
rect 7856 2287 7863 2543
rect 7876 2263 7883 2573
rect 7896 2307 7903 3673
rect 7916 3667 7923 3813
rect 7856 2256 7883 2263
rect 7856 2076 7863 2213
rect 7876 2107 7883 2256
rect 7896 2087 7903 2273
rect 7856 1807 7863 2033
rect 7876 1923 7883 2063
rect 7896 1947 7903 2033
rect 7876 1916 7893 1923
rect 7836 1747 7843 1783
rect 7856 1727 7863 1763
rect 7876 1627 7883 1753
rect 7896 1603 7903 1893
rect 7876 1596 7903 1603
rect 7736 1247 7743 1303
rect 7776 1296 7803 1303
rect 7796 1207 7803 1296
rect 7716 1156 7743 1163
rect 7656 1127 7663 1133
rect 7696 1116 7703 1133
rect 7716 863 7723 1133
rect 7736 867 7743 1156
rect 7796 1116 7803 1193
rect 7776 967 7783 1093
rect 7696 856 7723 863
rect 7636 767 7643 823
rect 7636 636 7643 653
rect 7656 647 7663 733
rect 7676 687 7683 813
rect 7696 667 7703 856
rect 7716 807 7723 823
rect 7756 807 7763 813
rect 7716 787 7723 793
rect 7736 727 7743 803
rect 7776 727 7783 933
rect 7796 827 7803 853
rect 7687 636 7703 643
rect 7556 616 7583 623
rect 7476 596 7503 603
rect 7556 467 7563 616
rect 7656 616 7683 623
rect 7656 607 7663 616
rect 7456 376 7483 383
rect 7416 343 7423 373
rect 7476 347 7483 376
rect 7416 336 7443 343
rect 7516 343 7523 453
rect 7496 336 7523 343
rect 7476 227 7483 333
rect 7596 307 7603 343
rect 7636 327 7643 343
rect 7656 327 7663 573
rect 7036 156 7043 193
rect 7136 163 7143 173
rect 7136 156 7163 163
rect 7456 156 7463 193
rect 7536 156 7563 163
rect 6376 136 6403 143
rect 6436 127 6443 143
rect 7556 107 7563 156
rect 7596 147 7603 193
rect 7676 187 7683 573
rect 7756 347 7763 653
rect 7776 647 7783 673
rect 7796 656 7803 793
rect 7816 687 7823 1313
rect 7836 1287 7843 1553
rect 7836 867 7843 1193
rect 7856 1187 7863 1573
rect 7896 1567 7903 1573
rect 7856 1136 7863 1153
rect 7876 1147 7883 1273
rect 7896 1207 7903 1283
rect 7856 947 7863 1093
rect 7876 1087 7883 1103
rect 7836 707 7843 823
rect 7856 787 7863 803
rect 7836 623 7843 673
rect 7856 656 7863 693
rect 7876 667 7883 813
rect 7836 616 7863 623
rect 7796 356 7803 493
rect 7856 347 7863 616
rect 7876 607 7883 613
rect 7896 507 7903 1173
rect 7896 367 7903 473
rect 7776 327 7783 343
rect 7916 307 7923 2733
rect 7687 176 7703 183
rect 7836 176 7843 213
rect 7716 156 7743 163
rect 7736 147 7743 156
rect 7736 127 7743 133
rect 7756 107 7763 143
<< m3contact >>
rect 13 6153 27 6167
rect 33 6133 47 6147
rect 213 6133 227 6147
rect 233 6133 247 6147
rect 313 6133 327 6147
rect 393 6133 407 6147
rect 413 6133 427 6147
rect 493 6133 507 6147
rect 553 6133 567 6147
rect 653 6133 667 6147
rect 1413 6133 1427 6147
rect 53 6093 67 6107
rect 93 6053 107 6067
rect 153 5973 167 5987
rect 13 5873 27 5887
rect 73 5913 87 5927
rect 113 5913 127 5927
rect 73 5873 87 5887
rect 53 5653 67 5667
rect 373 6113 387 6127
rect 313 5973 327 5987
rect 213 5953 227 5967
rect 253 5953 267 5967
rect 193 5673 207 5687
rect 253 5933 267 5947
rect 293 5933 307 5947
rect 273 5913 287 5927
rect 233 5893 247 5907
rect 113 5653 127 5667
rect 133 5653 147 5667
rect 53 5633 67 5647
rect 33 5473 47 5487
rect 173 5633 187 5647
rect 93 5473 107 5487
rect 133 5473 147 5487
rect 93 5453 107 5467
rect 353 5913 367 5927
rect 333 5893 347 5907
rect 373 5893 387 5907
rect 353 5673 367 5687
rect 493 5913 507 5927
rect 593 6113 607 6127
rect 693 6113 707 6127
rect 613 6093 627 6107
rect 633 6073 647 6087
rect 673 6073 687 6087
rect 733 6073 747 6087
rect 533 5933 547 5947
rect 613 5913 627 5927
rect 513 5893 527 5907
rect 573 5873 587 5887
rect 293 5653 307 5667
rect 333 5653 347 5667
rect 293 5633 307 5647
rect 313 5593 327 5607
rect 273 5473 287 5487
rect 173 5413 187 5427
rect 173 5373 187 5387
rect 313 5433 327 5447
rect 313 5253 327 5267
rect 253 5153 267 5167
rect 153 5133 167 5147
rect 273 5133 287 5147
rect 53 4953 67 4967
rect 153 4973 167 4987
rect 73 4933 87 4947
rect 253 4953 267 4967
rect 133 4933 147 4947
rect 233 4773 247 4787
rect 213 4653 227 4667
rect 133 4633 147 4647
rect 133 4613 147 4627
rect 113 4473 127 4487
rect 13 4333 27 4347
rect 53 4333 67 4347
rect 113 4293 127 4307
rect 93 4253 107 4267
rect 53 4233 67 4247
rect 33 4213 47 4227
rect 53 4193 67 4207
rect 93 4193 107 4207
rect 13 4153 27 4167
rect 93 4173 107 4187
rect 113 4173 127 4187
rect 53 4153 67 4167
rect 73 4153 87 4167
rect 53 4113 67 4127
rect 33 4093 47 4107
rect 13 4053 27 4067
rect 13 3453 27 3467
rect 13 3433 27 3447
rect 193 4573 207 4587
rect 213 4533 227 4547
rect 173 4453 187 4467
rect 153 4233 167 4247
rect 193 4213 207 4227
rect 253 4653 267 4667
rect 393 5633 407 5647
rect 413 5613 427 5627
rect 553 5613 567 5627
rect 553 5593 567 5607
rect 373 5533 387 5547
rect 433 5533 447 5547
rect 353 5433 367 5447
rect 513 5473 527 5487
rect 393 5433 407 5447
rect 433 5433 447 5447
rect 473 5433 487 5447
rect 413 5253 427 5267
rect 353 5133 367 5147
rect 373 5113 387 5127
rect 393 5113 407 5127
rect 373 4953 387 4967
rect 373 4913 387 4927
rect 273 4633 287 4647
rect 253 4573 267 4587
rect 373 4633 387 4647
rect 333 4593 347 4607
rect 373 4593 387 4607
rect 313 4533 327 4547
rect 273 4513 287 4527
rect 293 4493 307 4507
rect 393 4513 407 4527
rect 253 4453 267 4467
rect 233 4233 247 4247
rect 153 4193 167 4207
rect 93 3993 107 4007
rect 73 3773 87 3787
rect 93 3633 107 3647
rect 133 4013 147 4027
rect 133 3993 147 4007
rect 213 4173 227 4187
rect 173 4133 187 4147
rect 313 4333 327 4347
rect 353 4473 367 4487
rect 473 5153 487 5167
rect 473 4933 487 4947
rect 453 4653 467 4667
rect 593 5573 607 5587
rect 613 5533 627 5547
rect 593 5453 607 5467
rect 573 5433 587 5447
rect 613 5353 627 5367
rect 593 4933 607 4947
rect 613 4793 627 4807
rect 553 4773 567 4787
rect 493 4653 507 4667
rect 473 4613 487 4627
rect 453 4593 467 4607
rect 553 4613 567 4627
rect 413 4473 427 4487
rect 373 4453 387 4467
rect 413 4453 427 4467
rect 393 4433 407 4447
rect 313 4213 327 4227
rect 273 4193 287 4207
rect 313 4193 327 4207
rect 273 4173 287 4187
rect 233 4113 247 4127
rect 253 4113 267 4127
rect 333 4173 347 4187
rect 293 4133 307 4147
rect 293 4113 307 4127
rect 273 4073 287 4087
rect 233 4033 247 4047
rect 253 4033 267 4047
rect 173 4013 187 4027
rect 153 3973 167 3987
rect 153 3953 167 3967
rect 133 3693 147 3707
rect 153 3693 167 3707
rect 113 3593 127 3607
rect 93 3573 107 3587
rect 73 3553 87 3567
rect 33 3413 47 3427
rect 33 3393 47 3407
rect 153 3653 167 3667
rect 153 3533 167 3547
rect 113 3493 127 3507
rect 113 3433 127 3447
rect 113 3413 127 3427
rect 93 3193 107 3207
rect 73 3113 87 3127
rect 33 3033 47 3047
rect 93 3033 107 3047
rect 53 3013 67 3027
rect 33 2993 47 3007
rect 73 2993 87 3007
rect 73 2833 87 2847
rect 33 2773 47 2787
rect 33 2593 47 2607
rect 133 3373 147 3387
rect 153 3373 167 3387
rect 153 3313 167 3327
rect 133 3253 147 3267
rect 133 3213 147 3227
rect 153 3093 167 3107
rect 233 3973 247 3987
rect 273 3973 287 3987
rect 213 3773 227 3787
rect 213 3513 227 3527
rect 313 4073 327 4087
rect 373 4273 387 4287
rect 353 4153 367 4167
rect 333 4053 347 4067
rect 413 4233 427 4247
rect 393 4213 407 4227
rect 493 4553 507 4567
rect 533 4553 547 4567
rect 453 4513 467 4527
rect 493 4513 507 4527
rect 513 4493 527 4507
rect 473 4433 487 4447
rect 513 4433 527 4447
rect 533 4413 547 4427
rect 453 4293 467 4307
rect 453 4253 467 4267
rect 513 4253 527 4267
rect 433 4213 447 4227
rect 493 4233 507 4247
rect 433 4173 447 4187
rect 433 4153 447 4167
rect 453 4153 467 4167
rect 593 4633 607 4647
rect 653 6053 667 6067
rect 653 5953 667 5967
rect 713 5953 727 5967
rect 793 5933 807 5947
rect 873 6093 887 6107
rect 1053 6093 1067 6107
rect 1173 6093 1187 6107
rect 1273 6093 1287 6107
rect 1673 6153 1687 6167
rect 1793 6153 1807 6167
rect 2093 6153 2107 6167
rect 2173 6153 2187 6167
rect 1473 6133 1487 6147
rect 1393 6093 1407 6107
rect 1433 6093 1447 6107
rect 1493 6093 1507 6107
rect 1533 6093 1547 6107
rect 1613 6093 1627 6107
rect 833 6073 847 6087
rect 1093 6073 1107 6087
rect 1233 6033 1247 6047
rect 853 5973 867 5987
rect 913 5953 927 5967
rect 673 5853 687 5867
rect 673 5633 687 5647
rect 713 5633 727 5647
rect 673 5613 687 5627
rect 693 5613 707 5627
rect 733 5613 747 5627
rect 853 5613 867 5627
rect 793 5573 807 5587
rect 813 5573 827 5587
rect 793 5513 807 5527
rect 713 5493 727 5507
rect 693 5473 707 5487
rect 693 5453 707 5467
rect 673 5413 687 5427
rect 733 5453 747 5467
rect 753 5453 767 5467
rect 753 5153 767 5167
rect 733 5133 747 5147
rect 853 5553 867 5567
rect 893 5473 907 5487
rect 873 5453 887 5467
rect 893 5433 907 5447
rect 1013 5933 1027 5947
rect 1333 6073 1347 6087
rect 1453 6073 1467 6087
rect 1473 6073 1487 6087
rect 1513 6073 1527 6087
rect 1453 6053 1467 6067
rect 1513 5993 1527 6007
rect 1253 5953 1267 5967
rect 1353 5953 1367 5967
rect 1513 5953 1527 5967
rect 1313 5933 1327 5947
rect 1113 5893 1127 5907
rect 1153 5893 1167 5907
rect 1053 5873 1067 5887
rect 1093 5873 1107 5887
rect 1153 5713 1167 5727
rect 993 5653 1007 5667
rect 953 5593 967 5607
rect 953 5533 967 5547
rect 933 5433 947 5447
rect 1073 5633 1087 5647
rect 1253 5913 1267 5927
rect 1293 5913 1307 5927
rect 1273 5893 1287 5907
rect 1253 5873 1267 5887
rect 1333 5873 1347 5887
rect 1193 5653 1207 5667
rect 1213 5653 1227 5667
rect 1333 5673 1347 5687
rect 1053 5613 1067 5627
rect 1093 5613 1107 5627
rect 1193 5613 1207 5627
rect 1313 5653 1327 5667
rect 1053 5573 1067 5587
rect 1033 5533 1047 5547
rect 1013 5453 1027 5467
rect 1273 5553 1287 5567
rect 1413 5933 1427 5947
rect 1453 5933 1467 5947
rect 1473 5933 1487 5947
rect 1493 5933 1507 5947
rect 1453 5893 1467 5907
rect 1393 5673 1407 5687
rect 1373 5653 1387 5667
rect 1313 5553 1327 5567
rect 1293 5493 1307 5507
rect 1373 5633 1387 5647
rect 1353 5473 1367 5487
rect 1313 5433 1327 5447
rect 993 5413 1007 5427
rect 1193 5413 1207 5427
rect 1253 5413 1267 5427
rect 1293 5413 1307 5427
rect 1213 5393 1227 5407
rect 853 5153 867 5167
rect 913 5153 927 5167
rect 1293 5373 1307 5387
rect 913 5133 927 5147
rect 1033 5133 1047 5147
rect 1253 5133 1267 5147
rect 773 5113 787 5127
rect 813 5113 827 5127
rect 993 5113 1007 5127
rect 1153 5113 1167 5127
rect 973 5093 987 5107
rect 853 4953 867 4967
rect 953 4953 967 4967
rect 653 4833 667 4847
rect 633 4613 647 4627
rect 573 4593 587 4607
rect 573 4533 587 4547
rect 633 4493 647 4507
rect 693 4653 707 4667
rect 673 4573 687 4587
rect 653 4473 667 4487
rect 633 4453 647 4467
rect 593 4433 607 4447
rect 573 4393 587 4407
rect 653 4393 667 4407
rect 633 4373 647 4387
rect 593 4353 607 4367
rect 573 4313 587 4327
rect 553 4273 567 4287
rect 533 4193 547 4207
rect 513 4173 527 4187
rect 553 4173 567 4187
rect 393 4133 407 4147
rect 393 4073 407 4087
rect 353 4013 367 4027
rect 373 4013 387 4027
rect 313 3993 327 4007
rect 413 4013 427 4027
rect 433 4013 447 4027
rect 253 3833 267 3847
rect 253 3553 267 3567
rect 253 3533 267 3547
rect 233 3473 247 3487
rect 213 3233 227 3247
rect 213 3213 227 3227
rect 213 3093 227 3107
rect 173 3073 187 3087
rect 173 3053 187 3067
rect 193 3053 207 3067
rect 153 3033 167 3047
rect 133 3013 147 3027
rect 173 3013 187 3027
rect 153 2993 167 3007
rect 113 2813 127 2827
rect 93 2773 107 2787
rect 113 2773 127 2787
rect 93 2613 107 2627
rect 93 2573 107 2587
rect 73 2553 87 2567
rect 53 2533 67 2547
rect 33 2513 47 2527
rect 13 2493 27 2507
rect 33 2493 47 2507
rect 13 2453 27 2467
rect 73 2293 87 2307
rect 93 2233 107 2247
rect 133 2713 147 2727
rect 133 2593 147 2607
rect 313 3893 327 3907
rect 293 3853 307 3867
rect 373 3973 387 3987
rect 333 3873 347 3887
rect 393 3853 407 3867
rect 353 3813 367 3827
rect 373 3693 387 3707
rect 313 3673 327 3687
rect 353 3673 367 3687
rect 373 3673 387 3687
rect 293 3613 307 3627
rect 313 3553 327 3567
rect 293 3533 307 3547
rect 393 3653 407 3667
rect 433 3973 447 3987
rect 533 4133 547 4147
rect 473 4053 487 4067
rect 513 3993 527 4007
rect 613 4253 627 4267
rect 613 4153 627 4167
rect 593 4133 607 4147
rect 633 4133 647 4147
rect 613 4093 627 4107
rect 593 4073 607 4087
rect 573 4013 587 4027
rect 693 4493 707 4507
rect 813 4853 827 4867
rect 793 4673 807 4687
rect 753 4653 767 4667
rect 773 4613 787 4627
rect 933 4933 947 4947
rect 873 4673 887 4687
rect 833 4633 847 4647
rect 893 4653 907 4667
rect 873 4633 887 4647
rect 773 4553 787 4567
rect 813 4553 827 4567
rect 793 4513 807 4527
rect 833 4513 847 4527
rect 773 4473 787 4487
rect 753 4453 767 4467
rect 713 4353 727 4367
rect 713 4233 727 4247
rect 673 4153 687 4167
rect 693 4153 707 4167
rect 853 4493 867 4507
rect 833 4473 847 4487
rect 793 4453 807 4467
rect 833 4453 847 4467
rect 893 4573 907 4587
rect 893 4473 907 4487
rect 953 4753 967 4767
rect 1013 4953 1027 4967
rect 1053 4953 1067 4967
rect 1033 4773 1047 4787
rect 953 4673 967 4687
rect 973 4673 987 4687
rect 953 4633 967 4647
rect 973 4593 987 4607
rect 953 4553 967 4567
rect 933 4473 947 4487
rect 853 4433 867 4447
rect 893 4433 907 4447
rect 813 4373 827 4387
rect 833 4373 847 4387
rect 833 4333 847 4347
rect 893 4333 907 4347
rect 833 4293 847 4307
rect 773 4213 787 4227
rect 793 4213 807 4227
rect 773 4193 787 4207
rect 793 4193 807 4207
rect 733 4133 747 4147
rect 653 4073 667 4087
rect 713 4073 727 4087
rect 733 4073 747 4087
rect 613 4033 627 4047
rect 633 4013 647 4027
rect 653 4013 667 4027
rect 693 4013 707 4027
rect 613 3993 627 4007
rect 533 3973 547 3987
rect 593 3973 607 3987
rect 453 3953 467 3967
rect 493 3953 507 3967
rect 513 3953 527 3967
rect 433 3873 447 3887
rect 473 3873 487 3887
rect 453 3713 467 3727
rect 453 3693 467 3707
rect 553 3933 567 3947
rect 633 3953 647 3967
rect 593 3833 607 3847
rect 573 3793 587 3807
rect 553 3713 567 3727
rect 533 3693 547 3707
rect 493 3673 507 3687
rect 353 3533 367 3547
rect 373 3533 387 3547
rect 253 3433 267 3447
rect 293 3393 307 3407
rect 353 3493 367 3507
rect 373 3493 387 3507
rect 333 3353 347 3367
rect 333 3293 347 3307
rect 273 3273 287 3287
rect 293 3273 307 3287
rect 253 3253 267 3267
rect 313 3233 327 3247
rect 273 3213 287 3227
rect 313 3213 327 3227
rect 253 3053 267 3067
rect 293 3053 307 3067
rect 273 3013 287 3027
rect 333 3113 347 3127
rect 373 3433 387 3447
rect 473 3613 487 3627
rect 413 3593 427 3607
rect 393 3313 407 3327
rect 473 3573 487 3587
rect 553 3613 567 3627
rect 513 3593 527 3607
rect 493 3553 507 3567
rect 533 3573 547 3587
rect 513 3533 527 3547
rect 553 3553 567 3567
rect 433 3493 447 3507
rect 513 3493 527 3507
rect 473 3453 487 3467
rect 413 3253 427 3267
rect 513 3313 527 3327
rect 393 3233 407 3247
rect 433 3233 447 3247
rect 473 3233 487 3247
rect 513 3233 527 3247
rect 413 3193 427 3207
rect 433 3193 447 3207
rect 433 3153 447 3167
rect 533 3213 547 3227
rect 493 3173 507 3187
rect 513 3153 527 3167
rect 453 3133 467 3147
rect 253 2993 267 3007
rect 313 2993 327 3007
rect 233 2933 247 2947
rect 273 2893 287 2907
rect 233 2793 247 2807
rect 173 2753 187 2767
rect 213 2753 227 2767
rect 213 2733 227 2747
rect 173 2633 187 2647
rect 173 2613 187 2627
rect 153 2573 167 2587
rect 213 2573 227 2587
rect 153 2533 167 2547
rect 193 2533 207 2547
rect 153 2433 167 2447
rect 133 2293 147 2307
rect 133 2253 147 2267
rect 213 2413 227 2427
rect 173 2293 187 2307
rect 153 2213 167 2227
rect 113 2153 127 2167
rect 73 2133 87 2147
rect 153 2133 167 2147
rect 393 3113 407 3127
rect 413 3073 427 3087
rect 433 3073 447 3087
rect 533 3073 547 3087
rect 393 3033 407 3047
rect 373 2933 387 2947
rect 333 2833 347 2847
rect 353 2813 367 2827
rect 273 2773 287 2787
rect 333 2773 347 2787
rect 313 2753 327 2767
rect 253 2733 267 2747
rect 293 2733 307 2747
rect 293 2713 307 2727
rect 293 2693 307 2707
rect 273 2613 287 2627
rect 253 2533 267 2547
rect 273 2533 287 2547
rect 293 2533 307 2547
rect 253 2513 267 2527
rect 233 2293 247 2307
rect 213 2253 227 2267
rect 273 2273 287 2287
rect 293 2273 307 2287
rect 253 2253 267 2267
rect 293 2213 307 2227
rect 233 2193 247 2207
rect 273 2193 287 2207
rect 213 2173 227 2187
rect 73 2113 87 2127
rect 113 2113 127 2127
rect 33 2093 47 2107
rect 53 2093 67 2107
rect 173 2113 187 2127
rect 33 2053 47 2067
rect 53 2053 67 2067
rect 133 2053 147 2067
rect 73 2033 87 2047
rect 93 2033 107 2047
rect 73 1913 87 1927
rect 33 1813 47 1827
rect 233 2153 247 2167
rect 273 2153 287 2167
rect 253 2093 267 2107
rect 273 2093 287 2107
rect 233 2073 247 2087
rect 293 2073 307 2087
rect 233 2053 247 2067
rect 273 2053 287 2067
rect 253 2013 267 2027
rect 213 1933 227 1947
rect 213 1913 227 1927
rect 193 1893 207 1907
rect 93 1773 107 1787
rect 173 1773 187 1787
rect 133 1753 147 1767
rect 73 1673 87 1687
rect 73 1633 87 1647
rect 53 1613 67 1627
rect 93 1613 107 1627
rect 213 1733 227 1747
rect 153 1713 167 1727
rect 93 1533 107 1547
rect 73 1293 87 1307
rect 33 633 47 647
rect 173 1593 187 1607
rect 333 2733 347 2747
rect 333 2533 347 2547
rect 333 2473 347 2487
rect 353 2393 367 2407
rect 393 2813 407 2827
rect 453 3053 467 3067
rect 513 3033 527 3047
rect 513 2813 527 2827
rect 453 2793 467 2807
rect 493 2793 507 2807
rect 433 2773 447 2787
rect 473 2773 487 2787
rect 473 2753 487 2767
rect 493 2733 507 2747
rect 453 2713 467 2727
rect 413 2673 427 2687
rect 493 2633 507 2647
rect 453 2593 467 2607
rect 393 2533 407 2547
rect 393 2453 407 2467
rect 393 2373 407 2387
rect 473 2533 487 2547
rect 593 3773 607 3787
rect 613 3773 627 3787
rect 793 4153 807 4167
rect 813 4153 827 4167
rect 793 4073 807 4087
rect 853 4253 867 4267
rect 853 4153 867 4167
rect 873 4133 887 4147
rect 853 4053 867 4067
rect 753 4013 767 4027
rect 793 4013 807 4027
rect 833 4013 847 4027
rect 933 4393 947 4407
rect 933 4273 947 4287
rect 913 4193 927 4207
rect 933 4193 947 4207
rect 973 4493 987 4507
rect 1013 4633 1027 4647
rect 1213 5093 1227 5107
rect 1333 5113 1347 5127
rect 1293 5073 1307 5087
rect 1333 5033 1347 5047
rect 1413 5613 1427 5627
rect 1553 6013 1567 6027
rect 1533 5633 1547 5647
rect 1753 6133 1767 6147
rect 1833 6133 1847 6147
rect 1693 6033 1707 6047
rect 1833 6073 1847 6087
rect 1813 6033 1827 6047
rect 1733 6013 1747 6027
rect 1813 6013 1827 6027
rect 1633 5973 1647 5987
rect 1793 5973 1807 5987
rect 1653 5953 1667 5967
rect 1673 5953 1687 5967
rect 1573 5893 1587 5907
rect 1593 5633 1607 5647
rect 1613 5633 1627 5647
rect 1693 5933 1707 5947
rect 1713 5913 1727 5927
rect 1713 5873 1727 5887
rect 1713 5693 1727 5707
rect 1753 5673 1767 5687
rect 1513 5573 1527 5587
rect 1473 5553 1487 5567
rect 1453 5513 1467 5527
rect 1593 5593 1607 5607
rect 1733 5613 1747 5627
rect 1573 5553 1587 5567
rect 1673 5553 1687 5567
rect 1553 5513 1567 5527
rect 1473 5453 1487 5467
rect 1493 5433 1507 5447
rect 1553 5433 1567 5447
rect 1373 5413 1387 5427
rect 1453 5413 1467 5427
rect 1493 5133 1507 5147
rect 1553 5133 1567 5147
rect 1673 5473 1687 5487
rect 1713 5473 1727 5487
rect 1633 5433 1647 5447
rect 1693 5453 1707 5467
rect 1753 5473 1767 5487
rect 1613 5413 1627 5427
rect 1673 5393 1687 5407
rect 1653 5373 1667 5387
rect 1773 5413 1787 5427
rect 1793 5393 1807 5407
rect 1773 5373 1787 5387
rect 1893 6113 1907 6127
rect 1973 6113 1987 6127
rect 2013 6113 2027 6127
rect 1913 6073 1927 6087
rect 1853 5993 1867 6007
rect 1853 5933 1867 5947
rect 1833 5913 1847 5927
rect 2093 6113 2107 6127
rect 1993 6073 2007 6087
rect 2073 6073 2087 6087
rect 2033 6053 2047 6067
rect 2893 6133 2907 6147
rect 2153 6113 2167 6127
rect 2233 6113 2247 6127
rect 2113 6073 2127 6087
rect 2093 6033 2107 6047
rect 2153 6033 2167 6047
rect 2013 5953 2027 5967
rect 2053 5893 2067 5907
rect 1893 5873 1907 5887
rect 1973 5873 1987 5887
rect 2293 6093 2307 6107
rect 2273 6073 2287 6087
rect 2253 6053 2267 6067
rect 2233 5973 2247 5987
rect 2273 5913 2287 5927
rect 2093 5873 2107 5887
rect 2133 5873 2147 5887
rect 2173 5873 2187 5887
rect 2253 5873 2267 5887
rect 2273 5873 2287 5887
rect 2393 6113 2407 6127
rect 2433 6113 2447 6127
rect 2693 6113 2707 6127
rect 2373 6093 2387 6107
rect 2353 6073 2367 6087
rect 2393 6033 2407 6047
rect 2333 5973 2347 5987
rect 2313 5913 2327 5927
rect 2353 5913 2367 5927
rect 2293 5833 2307 5847
rect 2513 6093 2527 6107
rect 2553 6093 2567 6107
rect 2733 6093 2747 6107
rect 2553 5953 2567 5967
rect 2533 5933 2547 5947
rect 2593 5933 2607 5947
rect 2413 5913 2427 5927
rect 2573 5913 2587 5927
rect 2473 5893 2487 5907
rect 2513 5893 2527 5907
rect 2493 5873 2507 5887
rect 2453 5853 2467 5867
rect 2513 5853 2527 5867
rect 2693 5913 2707 5927
rect 2873 6013 2887 6027
rect 3033 6093 3047 6107
rect 4793 6173 4807 6187
rect 5193 6173 5207 6187
rect 5313 6173 5327 6187
rect 7413 6173 7427 6187
rect 7733 6173 7747 6187
rect 3293 6153 3307 6167
rect 3473 6153 3487 6167
rect 3593 6153 3607 6167
rect 3673 6153 3687 6167
rect 3713 6153 3727 6167
rect 3813 6153 3827 6167
rect 3853 6153 3867 6167
rect 2993 6073 3007 6087
rect 3233 6093 3247 6107
rect 3113 6073 3127 6087
rect 3273 6053 3287 6067
rect 3093 5993 3107 6007
rect 2973 5953 2987 5967
rect 2933 5933 2947 5947
rect 2993 5933 3007 5947
rect 3033 5933 3047 5947
rect 2593 5873 2607 5887
rect 2553 5833 2567 5847
rect 2153 5713 2167 5727
rect 2393 5713 2407 5727
rect 2413 5713 2427 5727
rect 2093 5693 2107 5707
rect 1853 5613 1867 5627
rect 2013 5653 2027 5667
rect 2053 5653 2067 5667
rect 1913 5613 1927 5627
rect 1973 5593 1987 5607
rect 1893 5573 1907 5587
rect 1913 5573 1927 5587
rect 1893 5553 1907 5567
rect 1853 5433 1867 5447
rect 1913 5533 1927 5547
rect 1833 5413 1847 5427
rect 1873 5413 1887 5427
rect 1953 5513 1967 5527
rect 2033 5633 2047 5647
rect 1993 5573 2007 5587
rect 2013 5553 2027 5567
rect 1973 5473 1987 5487
rect 1933 5413 1947 5427
rect 1993 5413 2007 5427
rect 1813 5353 1827 5367
rect 1833 5353 1847 5367
rect 1913 5353 1927 5367
rect 1373 5093 1387 5107
rect 1413 5033 1427 5047
rect 1373 4953 1387 4967
rect 1693 5053 1707 5067
rect 1853 5073 1867 5087
rect 1793 5033 1807 5047
rect 1793 5013 1807 5027
rect 2213 5673 2227 5687
rect 2373 5673 2387 5687
rect 2113 5613 2127 5627
rect 2153 5533 2167 5547
rect 2073 5473 2087 5487
rect 2113 5453 2127 5467
rect 2313 5633 2327 5647
rect 2273 5593 2287 5607
rect 2233 5573 2247 5587
rect 2393 5613 2407 5627
rect 2333 5593 2347 5607
rect 2393 5573 2407 5587
rect 2313 5553 2327 5567
rect 2193 5513 2207 5527
rect 2233 5513 2247 5527
rect 2173 5453 2187 5467
rect 2213 5453 2227 5467
rect 2093 5413 2107 5427
rect 2173 5413 2187 5427
rect 2133 5393 2147 5407
rect 2033 5333 2047 5347
rect 2033 5233 2047 5247
rect 2073 5233 2087 5247
rect 2013 5113 2027 5127
rect 1993 5013 2007 5027
rect 1953 4993 1967 5007
rect 1593 4973 1607 4987
rect 1793 4973 1807 4987
rect 1913 4973 1927 4987
rect 1453 4953 1467 4967
rect 1493 4953 1507 4967
rect 1573 4953 1587 4967
rect 1633 4953 1647 4967
rect 1353 4893 1367 4907
rect 1213 4873 1227 4887
rect 1373 4873 1387 4887
rect 1073 4833 1087 4847
rect 1333 4773 1347 4787
rect 1133 4733 1147 4747
rect 1193 4733 1207 4747
rect 1233 4733 1247 4747
rect 1053 4713 1067 4727
rect 1093 4693 1107 4707
rect 1113 4653 1127 4667
rect 1073 4613 1087 4627
rect 1093 4613 1107 4627
rect 1053 4533 1067 4547
rect 993 4473 1007 4487
rect 973 4453 987 4467
rect 993 4433 1007 4447
rect 993 4313 1007 4327
rect 973 4273 987 4287
rect 1033 4493 1047 4507
rect 1173 4613 1187 4627
rect 1153 4573 1167 4587
rect 1173 4533 1187 4547
rect 1113 4513 1127 4527
rect 1073 4473 1087 4487
rect 1093 4433 1107 4447
rect 1033 4413 1047 4427
rect 1133 4413 1147 4427
rect 1053 4373 1067 4387
rect 1073 4373 1087 4387
rect 1053 4313 1067 4327
rect 993 4253 1007 4267
rect 1013 4253 1027 4267
rect 953 4173 967 4187
rect 913 4153 927 4167
rect 933 4153 947 4167
rect 913 4133 927 4147
rect 733 3933 747 3947
rect 713 3793 727 3807
rect 713 3773 727 3787
rect 693 3753 707 3767
rect 673 3733 687 3747
rect 653 3713 667 3727
rect 613 3693 627 3707
rect 633 3693 647 3707
rect 653 3673 667 3687
rect 673 3673 687 3687
rect 713 3673 727 3687
rect 593 3653 607 3667
rect 573 3533 587 3547
rect 633 3613 647 3627
rect 613 3573 627 3587
rect 773 3973 787 3987
rect 773 3913 787 3927
rect 753 3833 767 3847
rect 753 3813 767 3827
rect 753 3733 767 3747
rect 773 3733 787 3747
rect 853 3953 867 3967
rect 813 3933 827 3947
rect 833 3933 847 3947
rect 833 3853 847 3867
rect 753 3713 767 3727
rect 793 3713 807 3727
rect 713 3593 727 3607
rect 733 3593 747 3607
rect 673 3573 687 3587
rect 633 3553 647 3567
rect 653 3553 667 3567
rect 613 3493 627 3507
rect 573 3313 587 3327
rect 613 3273 627 3287
rect 593 3233 607 3247
rect 573 3213 587 3227
rect 573 3193 587 3207
rect 613 3133 627 3147
rect 633 3053 647 3067
rect 633 3033 647 3047
rect 633 2993 647 3007
rect 553 2853 567 2867
rect 573 2813 587 2827
rect 533 2693 547 2707
rect 533 2673 547 2687
rect 513 2593 527 2607
rect 613 2853 627 2867
rect 673 3513 687 3527
rect 813 3693 827 3707
rect 793 3673 807 3687
rect 773 3653 787 3667
rect 793 3593 807 3607
rect 753 3573 767 3587
rect 753 3553 767 3567
rect 833 3653 847 3667
rect 853 3593 867 3607
rect 813 3533 827 3547
rect 833 3533 847 3547
rect 693 3493 707 3507
rect 673 3473 687 3487
rect 733 3473 747 3487
rect 813 3493 827 3507
rect 733 3413 747 3427
rect 773 3433 787 3447
rect 753 3253 767 3267
rect 733 3233 747 3247
rect 893 3973 907 3987
rect 933 3973 947 3987
rect 973 4153 987 4167
rect 1033 4233 1047 4247
rect 1013 4173 1027 4187
rect 1213 4713 1227 4727
rect 1193 4433 1207 4447
rect 1193 4413 1207 4427
rect 1173 4353 1187 4367
rect 1173 4313 1187 4327
rect 1253 4633 1267 4647
rect 1313 4653 1327 4667
rect 1233 4473 1247 4487
rect 1333 4473 1347 4487
rect 1433 4693 1447 4707
rect 1393 4673 1407 4687
rect 1573 4833 1587 4847
rect 1493 4813 1507 4827
rect 1533 4793 1547 4807
rect 1493 4693 1507 4707
rect 1493 4673 1507 4687
rect 1433 4533 1447 4547
rect 1413 4473 1427 4487
rect 1273 4433 1287 4447
rect 1233 4373 1247 4387
rect 1253 4373 1267 4387
rect 1213 4333 1227 4347
rect 1233 4333 1247 4347
rect 1213 4313 1227 4327
rect 1093 4213 1107 4227
rect 1153 4213 1167 4227
rect 1193 4213 1207 4227
rect 1033 4153 1047 4167
rect 993 4133 1007 4147
rect 1053 4073 1067 4087
rect 973 3973 987 3987
rect 933 3873 947 3887
rect 893 3813 907 3827
rect 913 3753 927 3767
rect 893 3713 907 3727
rect 893 3653 907 3667
rect 953 3773 967 3787
rect 1033 3973 1047 3987
rect 1073 3973 1087 3987
rect 1013 3893 1027 3907
rect 993 3753 1007 3767
rect 973 3733 987 3747
rect 1013 3733 1027 3747
rect 1033 3713 1047 3727
rect 1073 3713 1087 3727
rect 973 3693 987 3707
rect 1033 3673 1047 3687
rect 1053 3673 1067 3687
rect 1013 3633 1027 3647
rect 1033 3633 1047 3647
rect 1133 4193 1147 4207
rect 1153 4193 1167 4207
rect 1193 4193 1207 4207
rect 1353 4453 1367 4467
rect 1393 4393 1407 4407
rect 1473 4393 1487 4407
rect 1513 4633 1527 4647
rect 1573 4533 1587 4547
rect 1653 4933 1667 4947
rect 1713 4673 1727 4687
rect 1633 4653 1647 4667
rect 1693 4653 1707 4667
rect 1673 4633 1687 4647
rect 1613 4533 1627 4547
rect 1873 4953 1887 4967
rect 1773 4933 1787 4947
rect 1953 4733 1967 4747
rect 1913 4713 1927 4727
rect 1933 4713 1947 4727
rect 1753 4653 1767 4667
rect 1813 4653 1827 4667
rect 1853 4653 1867 4667
rect 1893 4653 1907 4667
rect 1733 4633 1747 4647
rect 1773 4633 1787 4647
rect 1693 4553 1707 4567
rect 1593 4513 1607 4527
rect 1533 4493 1547 4507
rect 1553 4493 1567 4507
rect 1573 4473 1587 4487
rect 1593 4453 1607 4467
rect 1533 4433 1547 4447
rect 1553 4433 1567 4447
rect 1313 4353 1327 4367
rect 1293 4293 1307 4307
rect 1313 4293 1327 4307
rect 1273 4253 1287 4267
rect 1353 4253 1367 4267
rect 1113 4153 1127 4167
rect 1173 4133 1187 4147
rect 1113 4113 1127 4127
rect 1173 4093 1187 4107
rect 1133 3993 1147 4007
rect 1233 4053 1247 4067
rect 1193 4033 1207 4047
rect 1213 3993 1227 4007
rect 1153 3973 1167 3987
rect 1153 3953 1167 3967
rect 1173 3953 1187 3967
rect 1133 3893 1147 3907
rect 1133 3853 1147 3867
rect 1113 3813 1127 3827
rect 1133 3773 1147 3787
rect 1113 3753 1127 3767
rect 1173 3913 1187 3927
rect 1173 3853 1187 3867
rect 1193 3793 1207 3807
rect 1313 4193 1327 4207
rect 1353 4193 1367 4207
rect 1293 4173 1307 4187
rect 1353 4153 1367 4167
rect 1373 4153 1387 4167
rect 1333 4133 1347 4147
rect 1433 4373 1447 4387
rect 1493 4373 1507 4387
rect 1413 4233 1427 4247
rect 1393 4133 1407 4147
rect 1413 4133 1427 4147
rect 1293 4113 1307 4127
rect 1333 4113 1347 4127
rect 1353 4113 1367 4127
rect 1273 4053 1287 4067
rect 1293 4033 1307 4047
rect 1253 4013 1267 4027
rect 1313 4013 1327 4027
rect 1273 3993 1287 4007
rect 1253 3973 1267 3987
rect 1293 3873 1307 3887
rect 1313 3873 1327 3887
rect 1253 3773 1267 3787
rect 1293 3753 1307 3767
rect 1233 3733 1247 3747
rect 1293 3713 1307 3727
rect 1113 3693 1127 3707
rect 1093 3653 1107 3667
rect 1233 3693 1247 3707
rect 1273 3693 1287 3707
rect 1453 4193 1467 4207
rect 1533 4393 1547 4407
rect 1553 4373 1567 4387
rect 1533 4293 1547 4307
rect 1553 4273 1567 4287
rect 1513 4213 1527 4227
rect 1533 4193 1547 4207
rect 1473 4173 1487 4187
rect 1493 4133 1507 4147
rect 1433 4093 1447 4107
rect 1393 4073 1407 4087
rect 1353 4053 1367 4067
rect 1473 4033 1487 4047
rect 1413 3953 1427 3967
rect 1433 3953 1447 3967
rect 1353 3873 1367 3887
rect 1373 3873 1387 3887
rect 1353 3853 1367 3867
rect 1373 3853 1387 3867
rect 1393 3833 1407 3847
rect 1373 3793 1387 3807
rect 1333 3753 1347 3767
rect 1333 3733 1347 3747
rect 1353 3733 1367 3747
rect 1193 3653 1207 3667
rect 1193 3613 1207 3627
rect 1013 3593 1027 3607
rect 1073 3593 1087 3607
rect 1153 3593 1167 3607
rect 953 3573 967 3587
rect 933 3553 947 3567
rect 973 3533 987 3547
rect 993 3533 1007 3547
rect 893 3513 907 3527
rect 953 3513 967 3527
rect 973 3513 987 3527
rect 873 3453 887 3467
rect 813 3393 827 3407
rect 853 3393 867 3407
rect 853 3353 867 3367
rect 873 3293 887 3307
rect 873 3273 887 3287
rect 793 3233 807 3247
rect 713 3153 727 3167
rect 693 3113 707 3127
rect 713 3113 727 3127
rect 673 3073 687 3087
rect 653 2913 667 2927
rect 593 2773 607 2787
rect 593 2733 607 2747
rect 593 2713 607 2727
rect 573 2613 587 2627
rect 553 2573 567 2587
rect 513 2553 527 2567
rect 473 2393 487 2407
rect 493 2393 507 2407
rect 453 2313 467 2327
rect 393 2293 407 2307
rect 433 2273 447 2287
rect 373 2253 387 2267
rect 333 2213 347 2227
rect 353 2113 367 2127
rect 413 2233 427 2247
rect 413 2213 427 2227
rect 433 2213 447 2227
rect 393 2173 407 2187
rect 373 2093 387 2107
rect 333 2053 347 2067
rect 293 2033 307 2047
rect 313 2033 327 2047
rect 273 1973 287 1987
rect 353 2013 367 2027
rect 293 1913 307 1927
rect 273 1893 287 1907
rect 253 1653 267 1667
rect 233 1613 247 1627
rect 253 1593 267 1607
rect 133 1573 147 1587
rect 193 1573 207 1587
rect 173 1553 187 1567
rect 153 1413 167 1427
rect 113 1273 127 1287
rect 133 1273 147 1287
rect 93 1233 107 1247
rect 113 1113 127 1127
rect 93 793 107 807
rect 93 653 107 667
rect 133 1093 147 1107
rect 133 813 147 827
rect 133 753 147 767
rect 233 1533 247 1547
rect 213 1493 227 1507
rect 193 1473 207 1487
rect 253 1393 267 1407
rect 213 1293 227 1307
rect 173 1093 187 1107
rect 233 1173 247 1187
rect 313 1773 327 1787
rect 333 1733 347 1747
rect 293 1693 307 1707
rect 373 1953 387 1967
rect 373 1753 387 1767
rect 393 1733 407 1747
rect 313 1613 327 1627
rect 333 1613 347 1627
rect 353 1613 367 1627
rect 293 1553 307 1567
rect 373 1593 387 1607
rect 633 2693 647 2707
rect 753 3033 767 3047
rect 853 3213 867 3227
rect 833 3193 847 3207
rect 973 3433 987 3447
rect 993 3393 1007 3407
rect 973 3353 987 3367
rect 913 3293 927 3307
rect 913 3253 927 3267
rect 933 3233 947 3247
rect 973 3233 987 3247
rect 893 3213 907 3227
rect 813 3173 827 3187
rect 813 3113 827 3127
rect 873 3113 887 3127
rect 833 3073 847 3087
rect 813 3053 827 3067
rect 753 3013 767 3027
rect 793 3013 807 3027
rect 853 3013 867 3027
rect 753 2973 767 2987
rect 753 2953 767 2967
rect 713 2933 727 2947
rect 673 2713 687 2727
rect 733 2713 747 2727
rect 713 2693 727 2707
rect 653 2633 667 2647
rect 613 2573 627 2587
rect 653 2573 667 2587
rect 613 2553 627 2567
rect 593 2373 607 2387
rect 553 2313 567 2327
rect 513 2273 527 2287
rect 553 2273 567 2287
rect 493 2193 507 2207
rect 493 2173 507 2187
rect 493 2113 507 2127
rect 433 2073 447 2087
rect 473 2073 487 2087
rect 453 2053 467 2067
rect 453 2013 467 2027
rect 453 1993 467 2007
rect 473 1893 487 1907
rect 473 1833 487 1847
rect 453 1813 467 1827
rect 533 2253 547 2267
rect 593 2253 607 2267
rect 733 2633 747 2647
rect 673 2553 687 2567
rect 713 2553 727 2567
rect 713 2513 727 2527
rect 693 2493 707 2507
rect 653 2313 667 2327
rect 633 2293 647 2307
rect 533 2233 547 2247
rect 573 2233 587 2247
rect 613 2233 627 2247
rect 513 2033 527 2047
rect 653 2273 667 2287
rect 773 2933 787 2947
rect 833 2913 847 2927
rect 793 2873 807 2887
rect 793 2773 807 2787
rect 813 2753 827 2767
rect 793 2713 807 2727
rect 813 2713 827 2727
rect 833 2713 847 2727
rect 773 2673 787 2687
rect 793 2653 807 2667
rect 753 2433 767 2447
rect 733 2353 747 2367
rect 953 3213 967 3227
rect 913 3153 927 3167
rect 913 3073 927 3087
rect 893 2953 907 2967
rect 973 3013 987 3027
rect 933 2933 947 2947
rect 1093 3573 1107 3587
rect 1033 3533 1047 3547
rect 1073 3453 1087 3467
rect 1033 3373 1047 3387
rect 1033 3313 1047 3327
rect 1073 3273 1087 3287
rect 1053 3233 1067 3247
rect 1073 3213 1087 3227
rect 1013 3133 1027 3147
rect 1033 3013 1047 3027
rect 1013 2993 1027 3007
rect 1013 2973 1027 2987
rect 1053 2953 1067 2967
rect 993 2913 1007 2927
rect 913 2853 927 2867
rect 1113 3553 1127 3567
rect 1113 3513 1127 3527
rect 1153 3513 1167 3527
rect 1173 3493 1187 3507
rect 1133 3473 1147 3487
rect 1213 3593 1227 3607
rect 1133 3453 1147 3467
rect 1173 3453 1187 3467
rect 1193 3453 1207 3467
rect 1133 3373 1147 3387
rect 1113 3233 1127 3247
rect 1093 3193 1107 3207
rect 1253 3673 1267 3687
rect 1273 3673 1287 3687
rect 1253 3653 1267 3667
rect 1233 3573 1247 3587
rect 1293 3593 1307 3607
rect 1273 3573 1287 3587
rect 1253 3553 1267 3567
rect 1273 3553 1287 3567
rect 1273 3493 1287 3507
rect 1233 3453 1247 3467
rect 1273 3333 1287 3347
rect 1213 3313 1227 3327
rect 1253 3313 1267 3327
rect 1193 3293 1207 3307
rect 1133 3213 1147 3227
rect 1173 3213 1187 3227
rect 1253 3233 1267 3247
rect 1253 3213 1267 3227
rect 1213 3193 1227 3207
rect 1133 3173 1147 3187
rect 1193 3173 1207 3187
rect 1193 3113 1207 3127
rect 1113 3053 1127 3067
rect 1133 3053 1147 3067
rect 1113 3033 1127 3047
rect 1093 3013 1107 3027
rect 1113 2993 1127 3007
rect 1173 3053 1187 3067
rect 1253 3153 1267 3167
rect 1233 3093 1247 3107
rect 1233 3053 1247 3067
rect 1313 3213 1327 3227
rect 1313 3153 1327 3167
rect 1233 3033 1247 3047
rect 1213 2973 1227 2987
rect 1313 3053 1327 3067
rect 1273 3033 1287 3047
rect 1313 3033 1327 3047
rect 1253 3013 1267 3027
rect 1293 3013 1307 3027
rect 1233 2953 1247 2967
rect 1133 2933 1147 2947
rect 1113 2913 1127 2927
rect 1253 2913 1267 2927
rect 1093 2873 1107 2887
rect 873 2773 887 2787
rect 953 2773 967 2787
rect 1033 2773 1047 2787
rect 993 2753 1007 2767
rect 893 2733 907 2747
rect 933 2733 947 2747
rect 1053 2733 1067 2747
rect 813 2433 827 2447
rect 813 2353 827 2367
rect 773 2293 787 2307
rect 793 2293 807 2307
rect 853 2533 867 2547
rect 973 2713 987 2727
rect 953 2693 967 2707
rect 1013 2693 1027 2707
rect 1093 2693 1107 2707
rect 913 2673 927 2687
rect 893 2453 907 2467
rect 853 2433 867 2447
rect 833 2313 847 2327
rect 873 2333 887 2347
rect 813 2273 827 2287
rect 853 2273 867 2287
rect 613 2213 627 2227
rect 633 2213 647 2227
rect 573 2153 587 2167
rect 533 1953 547 1967
rect 533 1873 547 1887
rect 513 1853 527 1867
rect 513 1833 527 1847
rect 493 1793 507 1807
rect 493 1773 507 1787
rect 473 1713 487 1727
rect 413 1693 427 1707
rect 453 1673 467 1687
rect 413 1653 427 1667
rect 393 1573 407 1587
rect 353 1553 367 1567
rect 333 1293 347 1307
rect 313 1193 327 1207
rect 253 1113 267 1127
rect 273 1113 287 1127
rect 393 1453 407 1467
rect 373 1273 387 1287
rect 393 1253 407 1267
rect 433 1613 447 1627
rect 593 2133 607 2147
rect 633 2193 647 2207
rect 613 2093 627 2107
rect 613 2073 627 2087
rect 713 2253 727 2267
rect 793 2233 807 2247
rect 813 2233 827 2247
rect 673 2193 687 2207
rect 713 2193 727 2207
rect 733 2193 747 2207
rect 693 2173 707 2187
rect 673 2153 687 2167
rect 653 2113 667 2127
rect 693 2073 707 2087
rect 773 2213 787 2227
rect 753 2173 767 2187
rect 753 2113 767 2127
rect 793 2173 807 2187
rect 793 2093 807 2107
rect 593 2053 607 2067
rect 693 2053 707 2067
rect 673 2033 687 2047
rect 653 1973 667 1987
rect 593 1893 607 1907
rect 613 1853 627 1867
rect 553 1813 567 1827
rect 573 1793 587 1807
rect 733 2053 747 2067
rect 713 1973 727 1987
rect 693 1953 707 1967
rect 773 2013 787 2027
rect 733 1913 747 1927
rect 713 1893 727 1907
rect 653 1793 667 1807
rect 693 1793 707 1807
rect 553 1773 567 1787
rect 553 1753 567 1767
rect 513 1733 527 1747
rect 533 1633 547 1647
rect 513 1593 527 1607
rect 493 1573 507 1587
rect 453 1553 467 1567
rect 653 1733 667 1747
rect 673 1693 687 1707
rect 593 1593 607 1607
rect 633 1593 647 1607
rect 633 1573 647 1587
rect 533 1493 547 1507
rect 573 1433 587 1447
rect 433 1413 447 1427
rect 453 1373 467 1387
rect 473 1313 487 1327
rect 513 1313 527 1327
rect 553 1313 567 1327
rect 373 1213 387 1227
rect 413 1213 427 1227
rect 193 1053 207 1067
rect 173 813 187 827
rect 253 1073 267 1087
rect 233 1033 247 1047
rect 253 873 267 887
rect 233 813 247 827
rect 153 673 167 687
rect 133 633 147 647
rect 213 553 227 567
rect 113 393 127 407
rect 213 393 227 407
rect 73 373 87 387
rect 93 373 107 387
rect 73 333 87 347
rect 133 333 147 347
rect 33 153 47 167
rect 93 313 107 327
rect 113 313 127 327
rect 153 313 167 327
rect 133 173 147 187
rect 233 373 247 387
rect 313 1073 327 1087
rect 313 1033 327 1047
rect 333 1013 347 1027
rect 293 853 307 867
rect 273 833 287 847
rect 313 833 327 847
rect 273 813 287 827
rect 293 793 307 807
rect 333 793 347 807
rect 413 1153 427 1167
rect 473 1153 487 1167
rect 393 1133 407 1147
rect 433 933 447 947
rect 373 873 387 887
rect 373 853 387 867
rect 373 813 387 827
rect 393 793 407 807
rect 353 773 367 787
rect 413 733 427 747
rect 473 1113 487 1127
rect 533 1293 547 1307
rect 533 1253 547 1267
rect 553 1193 567 1207
rect 533 1113 547 1127
rect 473 1093 487 1107
rect 513 1093 527 1107
rect 593 1373 607 1387
rect 593 1333 607 1347
rect 613 1313 627 1327
rect 653 1193 667 1207
rect 653 1153 667 1167
rect 613 1133 627 1147
rect 633 1133 647 1147
rect 593 1113 607 1127
rect 613 1113 627 1127
rect 693 1673 707 1687
rect 773 1833 787 1847
rect 873 2233 887 2247
rect 853 2213 867 2227
rect 873 2193 887 2207
rect 893 2193 907 2207
rect 833 2173 847 2187
rect 853 2133 867 2147
rect 833 2113 847 2127
rect 873 2093 887 2107
rect 933 2613 947 2627
rect 933 2553 947 2567
rect 1093 2653 1107 2667
rect 993 2633 1007 2647
rect 973 2553 987 2567
rect 1053 2593 1067 2607
rect 993 2533 1007 2547
rect 953 2473 967 2487
rect 953 2453 967 2467
rect 1073 2533 1087 2547
rect 993 2413 1007 2427
rect 1053 2413 1067 2427
rect 973 2333 987 2347
rect 933 2253 947 2267
rect 933 2213 947 2227
rect 1033 2313 1047 2327
rect 993 2293 1007 2307
rect 1013 2273 1027 2287
rect 993 2253 1007 2267
rect 973 2173 987 2187
rect 953 2153 967 2167
rect 993 2153 1007 2167
rect 933 2113 947 2127
rect 853 2033 867 2047
rect 913 2033 927 2047
rect 833 2013 847 2027
rect 833 1993 847 2007
rect 793 1813 807 1827
rect 813 1813 827 1827
rect 753 1753 767 1767
rect 713 1653 727 1667
rect 753 1733 767 1747
rect 773 1733 787 1747
rect 733 1633 747 1647
rect 753 1633 767 1647
rect 693 1593 707 1607
rect 713 1573 727 1587
rect 733 1553 747 1567
rect 693 1373 707 1387
rect 713 1373 727 1387
rect 773 1513 787 1527
rect 813 1793 827 1807
rect 833 1773 847 1787
rect 833 1753 847 1767
rect 813 1653 827 1667
rect 1013 2133 1027 2147
rect 973 2093 987 2107
rect 993 2093 1007 2107
rect 1173 2853 1187 2867
rect 1133 2833 1147 2847
rect 1233 2833 1247 2847
rect 1173 2793 1187 2807
rect 1133 2773 1147 2787
rect 1153 2773 1167 2787
rect 1193 2753 1207 2767
rect 1133 2733 1147 2747
rect 1153 2673 1167 2687
rect 1213 2733 1227 2747
rect 1213 2693 1227 2707
rect 1293 2893 1307 2907
rect 1293 2773 1307 2787
rect 1433 3913 1447 3927
rect 1473 3913 1487 3927
rect 1473 3873 1487 3887
rect 1433 3833 1447 3847
rect 1413 3753 1427 3767
rect 1513 4113 1527 4127
rect 1513 4093 1527 4107
rect 1513 4033 1527 4047
rect 1593 4233 1607 4247
rect 1633 4493 1647 4507
rect 1653 4473 1667 4487
rect 1753 4533 1767 4547
rect 1733 4473 1747 4487
rect 1653 4293 1667 4307
rect 1633 4233 1647 4247
rect 1613 4213 1627 4227
rect 1713 4453 1727 4467
rect 1713 4413 1727 4427
rect 1733 4373 1747 4387
rect 1733 4253 1747 4267
rect 1593 4193 1607 4207
rect 1633 4193 1647 4207
rect 1673 4193 1687 4207
rect 1713 4193 1727 4207
rect 1573 4173 1587 4187
rect 1593 4153 1607 4167
rect 1653 4173 1667 4187
rect 1693 4173 1707 4187
rect 1673 4133 1687 4147
rect 1573 4033 1587 4047
rect 1533 4013 1547 4027
rect 1553 4013 1567 4027
rect 1613 4013 1627 4027
rect 1513 3913 1527 3927
rect 1493 3793 1507 3807
rect 1493 3753 1507 3767
rect 1613 3933 1627 3947
rect 1573 3913 1587 3927
rect 1653 4053 1667 4067
rect 1713 4093 1727 4107
rect 1693 4053 1707 4067
rect 1693 3993 1707 4007
rect 1713 3933 1727 3947
rect 1813 4553 1827 4567
rect 1793 4453 1807 4467
rect 1853 4453 1867 4467
rect 1873 4453 1887 4467
rect 1833 4433 1847 4447
rect 1813 4253 1827 4267
rect 1773 4233 1787 4247
rect 1753 4213 1767 4227
rect 1773 4193 1787 4207
rect 1853 4293 1867 4307
rect 1853 4253 1867 4267
rect 1913 4593 1927 4607
rect 1913 4273 1927 4287
rect 2153 5153 2167 5167
rect 2133 5113 2147 5127
rect 2313 5453 2327 5467
rect 2693 5693 2707 5707
rect 2653 5653 2667 5667
rect 2433 5633 2447 5647
rect 2613 5633 2627 5647
rect 2513 5613 2527 5627
rect 2593 5593 2607 5607
rect 2473 5573 2487 5587
rect 2573 5533 2587 5547
rect 2473 5473 2487 5487
rect 2433 5453 2447 5467
rect 2533 5453 2547 5467
rect 2293 5413 2307 5427
rect 2373 5413 2387 5427
rect 2413 5413 2427 5427
rect 2333 5393 2347 5407
rect 2353 5393 2367 5407
rect 2253 5193 2267 5207
rect 2213 5153 2227 5167
rect 2293 5153 2307 5167
rect 2333 5153 2347 5167
rect 2373 5153 2387 5167
rect 2153 4993 2167 5007
rect 2193 4993 2207 5007
rect 2113 4973 2127 4987
rect 2193 4953 2207 4967
rect 2233 4953 2247 4967
rect 2033 4933 2047 4947
rect 2133 4933 2147 4947
rect 2073 4913 2087 4927
rect 2013 4873 2027 4887
rect 1993 4653 2007 4667
rect 2033 4693 2047 4707
rect 2093 4813 2107 4827
rect 2173 4713 2187 4727
rect 2133 4693 2147 4707
rect 2193 4693 2207 4707
rect 2113 4633 2127 4647
rect 2073 4553 2087 4567
rect 2073 4513 2087 4527
rect 2013 4493 2027 4507
rect 2033 4493 2047 4507
rect 1993 4473 2007 4487
rect 2213 4633 2227 4647
rect 2313 5133 2327 5147
rect 2493 5433 2507 5447
rect 2453 5413 2467 5427
rect 2473 5413 2487 5427
rect 2913 5913 2927 5927
rect 2873 5893 2887 5907
rect 2813 5873 2827 5887
rect 2853 5873 2867 5887
rect 2893 5873 2907 5887
rect 2913 5873 2927 5887
rect 3013 5913 3027 5927
rect 3073 5893 3087 5907
rect 3173 5973 3187 5987
rect 3153 5933 3167 5947
rect 3113 5913 3127 5927
rect 3093 5833 3107 5847
rect 3133 5873 3147 5887
rect 3113 5693 3127 5707
rect 3153 5693 3167 5707
rect 2813 5673 2827 5687
rect 2993 5673 3007 5687
rect 2753 5653 2767 5667
rect 2793 5653 2807 5667
rect 2773 5633 2787 5647
rect 2833 5653 2847 5667
rect 2913 5653 2927 5667
rect 2953 5653 2967 5667
rect 3053 5653 3067 5667
rect 2713 5593 2727 5607
rect 2813 5593 2827 5607
rect 2933 5633 2947 5647
rect 3013 5633 3027 5647
rect 3033 5633 3047 5647
rect 2853 5613 2867 5627
rect 2893 5593 2907 5607
rect 2993 5593 3007 5607
rect 2833 5573 2847 5587
rect 2873 5573 2887 5587
rect 2973 5513 2987 5527
rect 2913 5473 2927 5487
rect 2933 5473 2947 5487
rect 2773 5453 2787 5467
rect 2753 5433 2767 5447
rect 2633 5413 2647 5427
rect 2493 5393 2507 5407
rect 2553 5393 2567 5407
rect 2573 5393 2587 5407
rect 2793 5433 2807 5447
rect 2813 5433 2827 5447
rect 2893 5433 2907 5447
rect 2633 5333 2647 5347
rect 2673 5333 2687 5347
rect 2733 5333 2747 5347
rect 2433 5153 2447 5167
rect 2473 5153 2487 5167
rect 2353 5113 2367 5127
rect 2413 5113 2427 5127
rect 2333 5093 2347 5107
rect 2353 5093 2367 5107
rect 2293 4993 2307 5007
rect 2333 4973 2347 4987
rect 2313 4773 2327 4787
rect 2273 4713 2287 4727
rect 2273 4693 2287 4707
rect 2313 4693 2327 4707
rect 2253 4673 2267 4687
rect 2193 4613 2207 4627
rect 2233 4613 2247 4627
rect 2173 4533 2187 4547
rect 2113 4493 2127 4507
rect 2153 4493 2167 4507
rect 2093 4473 2107 4487
rect 2053 4453 2067 4467
rect 1973 4433 1987 4447
rect 2253 4573 2267 4587
rect 2233 4513 2247 4527
rect 1973 4373 1987 4387
rect 2013 4373 2027 4387
rect 2113 4373 2127 4387
rect 1953 4353 1967 4367
rect 2033 4353 2047 4367
rect 2053 4353 2067 4367
rect 1993 4293 2007 4307
rect 1833 4213 1847 4227
rect 1853 4213 1867 4227
rect 1893 4213 1907 4227
rect 1933 4213 1947 4227
rect 1973 4213 1987 4227
rect 1893 4193 1907 4207
rect 1933 4193 1947 4207
rect 2093 4313 2107 4327
rect 2053 4293 2067 4307
rect 2033 4233 2047 4247
rect 2033 4193 2047 4207
rect 1753 4153 1767 4167
rect 1773 4153 1787 4167
rect 1873 4173 1887 4187
rect 1913 4173 1927 4187
rect 1813 4153 1827 4167
rect 1833 4153 1847 4167
rect 1893 4153 1907 4167
rect 1913 4153 1927 4167
rect 1973 4173 1987 4187
rect 1753 4013 1767 4027
rect 1773 4013 1787 4027
rect 1773 3973 1787 3987
rect 1533 3893 1547 3907
rect 1633 3893 1647 3907
rect 1733 3893 1747 3907
rect 1413 3693 1427 3707
rect 1473 3693 1487 3707
rect 1453 3673 1467 3687
rect 1473 3673 1487 3687
rect 1513 3673 1527 3687
rect 1353 3653 1367 3667
rect 1433 3573 1447 3587
rect 1353 3553 1367 3567
rect 1393 3553 1407 3567
rect 1373 3493 1387 3507
rect 1413 3473 1427 3487
rect 1353 3453 1367 3467
rect 1873 4053 1887 4067
rect 1853 3993 1867 4007
rect 1813 3953 1827 3967
rect 1833 3953 1847 3967
rect 1853 3913 1867 3927
rect 1673 3853 1687 3867
rect 1773 3853 1787 3867
rect 1553 3813 1567 3827
rect 1593 3773 1607 3787
rect 1613 3753 1627 3767
rect 1653 3753 1667 3767
rect 1553 3653 1567 3667
rect 1533 3633 1547 3647
rect 1593 3653 1607 3667
rect 1533 3553 1547 3567
rect 1513 3533 1527 3547
rect 1473 3513 1487 3527
rect 1473 3493 1487 3507
rect 1513 3473 1527 3487
rect 1533 3473 1547 3487
rect 1473 3393 1487 3407
rect 1513 3393 1527 3407
rect 1453 3373 1467 3387
rect 1413 3333 1427 3347
rect 1493 3333 1507 3347
rect 1373 3253 1387 3267
rect 1433 3193 1447 3207
rect 1573 3533 1587 3547
rect 1553 3333 1567 3347
rect 1533 3313 1547 3327
rect 1633 3673 1647 3687
rect 1713 3813 1727 3827
rect 1833 3793 1847 3807
rect 1753 3773 1767 3787
rect 1793 3773 1807 3787
rect 1693 3693 1707 3707
rect 1733 3693 1747 3707
rect 1673 3653 1687 3667
rect 1613 3573 1627 3587
rect 1613 3553 1627 3567
rect 1653 3513 1667 3527
rect 1713 3673 1727 3687
rect 1693 3613 1707 3627
rect 1793 3673 1807 3687
rect 1773 3553 1787 3567
rect 1793 3533 1807 3547
rect 1933 4133 1947 4147
rect 1893 3953 1907 3967
rect 1953 4113 1967 4127
rect 1993 4133 2007 4147
rect 2033 4173 2047 4187
rect 2033 4133 2047 4147
rect 2073 4273 2087 4287
rect 2053 4113 2067 4127
rect 2253 4473 2267 4487
rect 2213 4453 2227 4467
rect 2173 4433 2187 4447
rect 2213 4373 2227 4387
rect 2133 4293 2147 4307
rect 2093 4253 2107 4267
rect 2133 4253 2147 4267
rect 2093 4233 2107 4247
rect 2253 4413 2267 4427
rect 2233 4333 2247 4347
rect 2253 4273 2267 4287
rect 2453 5093 2467 5107
rect 2473 5033 2487 5047
rect 2373 4933 2387 4947
rect 2413 4933 2427 4947
rect 2613 5133 2627 5147
rect 2513 5013 2527 5027
rect 2613 5013 2627 5027
rect 2493 4873 2507 4887
rect 2393 4753 2407 4767
rect 2373 4733 2387 4747
rect 2293 4673 2307 4687
rect 2333 4673 2347 4687
rect 2353 4653 2367 4667
rect 2313 4633 2327 4647
rect 2493 4713 2507 4727
rect 2433 4673 2447 4687
rect 2413 4633 2427 4647
rect 2373 4613 2387 4627
rect 2433 4593 2447 4607
rect 2393 4533 2407 4547
rect 2413 4533 2427 4547
rect 2373 4513 2387 4527
rect 2293 4473 2307 4487
rect 2333 4473 2347 4487
rect 2413 4493 2427 4507
rect 2593 4693 2607 4707
rect 2673 5173 2687 5187
rect 2793 5153 2807 5167
rect 2873 5193 2887 5207
rect 2833 5153 2847 5167
rect 2953 5453 2967 5467
rect 2933 5333 2947 5347
rect 2913 5173 2927 5187
rect 3013 5433 3027 5447
rect 3133 5653 3147 5667
rect 3093 5633 3107 5647
rect 3113 5633 3127 5647
rect 3113 5553 3127 5567
rect 3073 5513 3087 5527
rect 3073 5453 3087 5467
rect 3093 5413 3107 5427
rect 3033 5393 3047 5407
rect 2973 5373 2987 5387
rect 2953 5173 2967 5187
rect 2933 5153 2947 5167
rect 2813 5133 2827 5147
rect 2853 5133 2867 5147
rect 2813 5113 2827 5127
rect 2633 4973 2647 4987
rect 2713 4973 2727 4987
rect 2773 4973 2787 4987
rect 2693 4953 2707 4967
rect 2673 4913 2687 4927
rect 2693 4793 2707 4807
rect 2593 4673 2607 4687
rect 2513 4473 2527 4487
rect 2653 4653 2667 4667
rect 2693 4653 2707 4667
rect 2793 4953 2807 4967
rect 2953 5093 2967 5107
rect 3233 5953 3247 5967
rect 3193 5913 3207 5927
rect 3233 5913 3247 5927
rect 3253 5893 3267 5907
rect 3213 5853 3227 5867
rect 3273 5713 3287 5727
rect 3193 5653 3207 5667
rect 3233 5653 3247 5667
rect 3333 6013 3347 6027
rect 3373 6013 3387 6027
rect 3453 6073 3467 6087
rect 3513 6073 3527 6087
rect 3693 6113 3707 6127
rect 3733 6113 3747 6127
rect 3773 6113 3787 6127
rect 3653 6093 3667 6107
rect 3793 6093 3807 6107
rect 3753 6033 3767 6047
rect 3513 5993 3527 6007
rect 3653 5993 3667 6007
rect 3353 5933 3367 5947
rect 3413 5933 3427 5947
rect 3493 5933 3507 5947
rect 3313 5893 3327 5907
rect 3353 5893 3367 5907
rect 3393 5893 3407 5907
rect 3333 5853 3347 5867
rect 3293 5693 3307 5707
rect 3353 5653 3367 5667
rect 3293 5613 3307 5627
rect 3253 5593 3267 5607
rect 3473 5913 3487 5927
rect 4053 6133 4067 6147
rect 4513 6133 4527 6147
rect 3973 6093 3987 6107
rect 3933 6073 3947 6087
rect 3933 6053 3947 6067
rect 3593 5913 3607 5927
rect 3673 5933 3687 5947
rect 3653 5913 3667 5927
rect 3813 5933 3827 5947
rect 3833 5913 3847 5927
rect 3633 5893 3647 5907
rect 3673 5893 3687 5907
rect 3693 5893 3707 5907
rect 3693 5873 3707 5887
rect 3933 5913 3947 5927
rect 3573 5853 3587 5867
rect 3853 5853 3867 5867
rect 3673 5833 3687 5847
rect 3433 5633 3447 5647
rect 3213 5573 3227 5587
rect 3233 5573 3247 5587
rect 3313 5573 3327 5587
rect 3173 5533 3187 5547
rect 3213 5433 3227 5447
rect 3153 5333 3167 5347
rect 3133 5173 3147 5187
rect 3173 5173 3187 5187
rect 3053 5133 3067 5147
rect 3013 5113 3027 5127
rect 2833 4973 2847 4987
rect 2893 4973 2907 4987
rect 2853 4953 2867 4967
rect 2893 4953 2907 4967
rect 3073 4953 3087 4967
rect 2953 4913 2967 4927
rect 2873 4893 2887 4907
rect 3093 4893 3107 4907
rect 3153 4893 3167 4907
rect 2753 4673 2767 4687
rect 2753 4653 2767 4667
rect 2713 4633 2727 4647
rect 2733 4633 2747 4647
rect 2693 4573 2707 4587
rect 2593 4473 2607 4487
rect 2673 4473 2687 4487
rect 2473 4453 2487 4467
rect 2493 4453 2507 4467
rect 2313 4433 2327 4447
rect 2353 4433 2367 4447
rect 2393 4433 2407 4447
rect 2413 4433 2427 4447
rect 2453 4433 2467 4447
rect 2293 4373 2307 4387
rect 2293 4313 2307 4327
rect 2273 4253 2287 4267
rect 2213 4213 2227 4227
rect 2353 4413 2367 4427
rect 2333 4333 2347 4347
rect 2313 4213 2327 4227
rect 2113 4193 2127 4207
rect 2173 4193 2187 4207
rect 2213 4193 2227 4207
rect 2253 4193 2267 4207
rect 2293 4193 2307 4207
rect 2013 4093 2027 4107
rect 2033 4093 2047 4107
rect 2073 4093 2087 4107
rect 1993 4073 2007 4087
rect 1973 4053 1987 4067
rect 2013 4053 2027 4067
rect 1953 4013 1967 4027
rect 2013 4013 2027 4027
rect 1953 3993 1967 4007
rect 1973 3993 1987 4007
rect 2013 3993 2027 4007
rect 1933 3933 1947 3947
rect 1893 3913 1907 3927
rect 1933 3893 1947 3907
rect 1913 3873 1927 3887
rect 1933 3813 1947 3827
rect 1993 3973 2007 3987
rect 1973 3833 1987 3847
rect 1913 3753 1927 3767
rect 1853 3713 1867 3727
rect 1893 3713 1907 3727
rect 1953 3753 1967 3767
rect 1933 3733 1947 3747
rect 1973 3733 1987 3747
rect 1993 3733 2007 3747
rect 1953 3713 1967 3727
rect 1853 3673 1867 3687
rect 1833 3633 1847 3647
rect 1913 3693 1927 3707
rect 1933 3673 1947 3687
rect 1873 3613 1887 3627
rect 1893 3613 1907 3627
rect 1853 3573 1867 3587
rect 1833 3553 1847 3567
rect 1853 3553 1867 3567
rect 1813 3513 1827 3527
rect 1673 3473 1687 3487
rect 1773 3493 1787 3507
rect 1793 3493 1807 3507
rect 1833 3493 1847 3507
rect 1733 3453 1747 3467
rect 1753 3433 1767 3447
rect 1673 3393 1687 3407
rect 1693 3393 1707 3407
rect 1613 3353 1627 3367
rect 1733 3353 1747 3367
rect 1693 3333 1707 3347
rect 1713 3333 1727 3347
rect 1673 3313 1687 3327
rect 1573 3293 1587 3307
rect 1593 3293 1607 3307
rect 1513 3233 1527 3247
rect 1713 3253 1727 3267
rect 1733 3253 1747 3267
rect 1613 3233 1627 3247
rect 1653 3233 1667 3247
rect 1693 3233 1707 3247
rect 1553 3213 1567 3227
rect 1493 3193 1507 3207
rect 1533 3193 1547 3207
rect 1633 3193 1647 3207
rect 1673 3213 1687 3227
rect 1693 3193 1707 3207
rect 1593 3173 1607 3187
rect 1653 3173 1667 3187
rect 1393 3133 1407 3147
rect 1473 3133 1487 3147
rect 1533 3133 1547 3147
rect 1693 3133 1707 3147
rect 1393 3113 1407 3127
rect 1373 3093 1387 3107
rect 1393 3073 1407 3087
rect 1373 3053 1387 3067
rect 1353 3033 1367 3047
rect 1433 3053 1447 3067
rect 1473 3053 1487 3067
rect 1413 3033 1427 3047
rect 1513 3033 1527 3047
rect 1433 2973 1447 2987
rect 1413 2933 1427 2947
rect 1413 2893 1427 2907
rect 1273 2753 1287 2767
rect 1293 2713 1307 2727
rect 1233 2653 1247 2667
rect 1253 2633 1267 2647
rect 1173 2553 1187 2567
rect 1193 2553 1207 2567
rect 1233 2553 1247 2567
rect 1253 2553 1267 2567
rect 1293 2553 1307 2567
rect 1133 2493 1147 2507
rect 1093 2393 1107 2407
rect 1113 2393 1127 2407
rect 1153 2353 1167 2367
rect 1113 2333 1127 2347
rect 1093 2313 1107 2327
rect 1073 2293 1087 2307
rect 1093 2273 1107 2287
rect 1073 2253 1087 2267
rect 1133 2213 1147 2227
rect 1233 2513 1247 2527
rect 1213 2453 1227 2467
rect 1193 2333 1207 2347
rect 1173 2293 1187 2307
rect 1153 2193 1167 2207
rect 1113 2173 1127 2187
rect 1193 2273 1207 2287
rect 1253 2493 1267 2507
rect 1273 2493 1287 2507
rect 1253 2373 1267 2387
rect 1233 2213 1247 2227
rect 1353 2753 1367 2767
rect 1393 2753 1407 2767
rect 1333 2713 1347 2727
rect 1353 2693 1367 2707
rect 1413 2693 1427 2707
rect 1373 2673 1387 2687
rect 1413 2673 1427 2687
rect 1353 2613 1367 2627
rect 1333 2553 1347 2567
rect 1473 2993 1487 3007
rect 1453 2953 1467 2967
rect 1453 2813 1467 2827
rect 1453 2773 1467 2787
rect 1593 3113 1607 3127
rect 1553 3033 1567 3047
rect 1533 2993 1547 3007
rect 1553 2993 1567 3007
rect 1493 2973 1507 2987
rect 1513 2973 1527 2987
rect 1513 2893 1527 2907
rect 1493 2833 1507 2847
rect 1473 2753 1487 2767
rect 1613 3053 1627 3067
rect 1673 2973 1687 2987
rect 1973 3693 1987 3707
rect 1953 3593 1967 3607
rect 1973 3593 1987 3607
rect 1893 3533 1907 3547
rect 1913 3533 1927 3547
rect 1893 3513 1907 3527
rect 1833 3453 1847 3467
rect 1873 3453 1887 3467
rect 1793 3413 1807 3427
rect 1793 3373 1807 3387
rect 1813 3373 1827 3387
rect 1773 3273 1787 3287
rect 1773 3233 1787 3247
rect 1753 3193 1767 3207
rect 1713 3113 1727 3127
rect 1753 3113 1767 3127
rect 1733 3033 1747 3047
rect 1753 3013 1767 3027
rect 1813 3293 1827 3307
rect 2053 4073 2067 4087
rect 2073 4033 2087 4047
rect 2193 4173 2207 4187
rect 2173 4153 2187 4167
rect 2193 4153 2207 4167
rect 2133 4093 2147 4107
rect 2273 4173 2287 4187
rect 2193 4113 2207 4127
rect 2213 4113 2227 4127
rect 2213 4073 2227 4087
rect 2173 4033 2187 4047
rect 2073 4013 2087 4027
rect 2113 4013 2127 4027
rect 2073 3973 2087 3987
rect 2133 3993 2147 4007
rect 2213 3993 2227 4007
rect 2113 3953 2127 3967
rect 2073 3833 2087 3847
rect 2053 3793 2067 3807
rect 2033 3733 2047 3747
rect 2193 3973 2207 3987
rect 2193 3913 2207 3927
rect 2153 3893 2167 3907
rect 2073 3773 2087 3787
rect 2093 3773 2107 3787
rect 2113 3773 2127 3787
rect 2073 3733 2087 3747
rect 2333 4173 2347 4187
rect 2313 4113 2327 4127
rect 2253 4073 2267 4087
rect 2253 4053 2267 4067
rect 2273 4053 2287 4067
rect 2433 4233 2447 4247
rect 2373 4173 2387 4187
rect 2393 4153 2407 4167
rect 2473 4413 2487 4427
rect 2533 4413 2547 4427
rect 2653 4413 2667 4427
rect 2493 4393 2507 4407
rect 2653 4373 2667 4387
rect 2673 4373 2687 4387
rect 2513 4313 2527 4327
rect 2493 4293 2507 4307
rect 2493 4213 2507 4227
rect 2473 4193 2487 4207
rect 2473 4173 2487 4187
rect 2353 4093 2367 4107
rect 2333 4053 2347 4067
rect 2313 4013 2327 4027
rect 2253 3993 2267 4007
rect 2273 3993 2287 4007
rect 2313 3993 2327 4007
rect 2253 3973 2267 3987
rect 2233 3873 2247 3887
rect 2213 3833 2227 3847
rect 2213 3713 2227 3727
rect 2113 3673 2127 3687
rect 2073 3653 2087 3667
rect 2033 3573 2047 3587
rect 2013 3547 2027 3561
rect 2093 3553 2107 3567
rect 2013 3513 2027 3527
rect 2053 3513 2067 3527
rect 1993 3473 2007 3487
rect 1973 3433 1987 3447
rect 1953 3413 1967 3427
rect 1873 3393 1887 3407
rect 1893 3353 1907 3367
rect 1973 3353 1987 3367
rect 1833 3233 1847 3247
rect 1873 3233 1887 3247
rect 1793 3213 1807 3227
rect 1793 3193 1807 3207
rect 1773 2933 1787 2947
rect 1853 3193 1867 3207
rect 1873 3193 1887 3207
rect 1813 3173 1827 3187
rect 2073 3493 2087 3507
rect 2053 3473 2067 3487
rect 2093 3473 2107 3487
rect 2033 3453 2047 3467
rect 2073 3413 2087 3427
rect 2013 3373 2027 3387
rect 2033 3373 2047 3387
rect 2053 3373 2067 3387
rect 1933 3293 1947 3307
rect 1933 3273 1947 3287
rect 1913 3233 1927 3247
rect 1913 3193 1927 3207
rect 1873 3133 1887 3147
rect 1893 3133 1907 3147
rect 1873 3113 1887 3127
rect 1813 3093 1827 3107
rect 1853 3073 1867 3087
rect 1813 3053 1827 3067
rect 1833 2993 1847 3007
rect 1833 2913 1847 2927
rect 1853 2913 1867 2927
rect 1813 2853 1827 2867
rect 1713 2813 1727 2827
rect 1793 2813 1807 2827
rect 1593 2793 1607 2807
rect 1693 2793 1707 2807
rect 1793 2793 1807 2807
rect 1533 2773 1547 2787
rect 1453 2713 1467 2727
rect 1493 2713 1507 2727
rect 1533 2713 1547 2727
rect 1573 2733 1587 2747
rect 1593 2733 1607 2747
rect 1533 2693 1547 2707
rect 1553 2693 1567 2707
rect 1513 2673 1527 2687
rect 1513 2613 1527 2627
rect 1433 2593 1447 2607
rect 1513 2553 1527 2567
rect 1353 2533 1367 2547
rect 1493 2513 1507 2527
rect 1333 2433 1347 2447
rect 1273 2233 1287 2247
rect 1273 2213 1287 2227
rect 1193 2193 1207 2207
rect 1253 2193 1267 2207
rect 1093 2113 1107 2127
rect 1113 2113 1127 2127
rect 1033 2093 1047 2107
rect 1073 2093 1087 2107
rect 1113 2093 1127 2107
rect 1053 2073 1067 2087
rect 953 2053 967 2067
rect 993 2053 1007 2067
rect 973 2013 987 2027
rect 993 2013 1007 2027
rect 933 1993 947 2007
rect 873 1853 887 1867
rect 913 1813 927 1827
rect 893 1773 907 1787
rect 953 1753 967 1767
rect 913 1733 927 1747
rect 893 1713 907 1727
rect 853 1693 867 1707
rect 913 1693 927 1707
rect 933 1693 947 1707
rect 833 1613 847 1627
rect 873 1613 887 1627
rect 873 1593 887 1607
rect 953 1673 967 1687
rect 1033 1973 1047 1987
rect 1013 1913 1027 1927
rect 993 1833 1007 1847
rect 993 1793 1007 1807
rect 1093 2053 1107 2067
rect 1153 2113 1167 2127
rect 1153 1953 1167 1967
rect 1173 1953 1187 1967
rect 1133 1833 1147 1847
rect 1013 1773 1027 1787
rect 1033 1773 1047 1787
rect 1133 1813 1147 1827
rect 1093 1793 1107 1807
rect 1133 1793 1147 1807
rect 1073 1773 1087 1787
rect 1093 1753 1107 1767
rect 1073 1733 1087 1747
rect 1053 1693 1067 1707
rect 973 1653 987 1667
rect 1153 1773 1167 1787
rect 1113 1713 1127 1727
rect 1093 1693 1107 1707
rect 1133 1693 1147 1707
rect 933 1613 947 1627
rect 813 1573 827 1587
rect 893 1573 907 1587
rect 813 1533 827 1547
rect 853 1533 867 1547
rect 793 1453 807 1467
rect 693 1293 707 1307
rect 773 1313 787 1327
rect 833 1513 847 1527
rect 753 1273 767 1287
rect 793 1273 807 1287
rect 873 1493 887 1507
rect 853 1453 867 1467
rect 853 1393 867 1407
rect 893 1433 907 1447
rect 1013 1613 1027 1627
rect 973 1593 987 1607
rect 1073 1633 1087 1647
rect 953 1573 967 1587
rect 993 1553 1007 1567
rect 1033 1533 1047 1547
rect 1053 1533 1067 1547
rect 873 1333 887 1347
rect 933 1353 947 1367
rect 973 1353 987 1367
rect 933 1333 947 1347
rect 1013 1333 1027 1347
rect 853 1273 867 1287
rect 893 1273 907 1287
rect 833 1253 847 1267
rect 993 1293 1007 1307
rect 953 1233 967 1247
rect 913 1193 927 1207
rect 753 1173 767 1187
rect 893 1173 907 1187
rect 733 1153 747 1167
rect 753 1133 767 1147
rect 853 1133 867 1147
rect 913 1133 927 1147
rect 673 1113 687 1127
rect 573 1093 587 1107
rect 553 1033 567 1047
rect 473 953 487 967
rect 453 733 467 747
rect 373 693 387 707
rect 433 693 447 707
rect 453 693 467 707
rect 293 673 307 687
rect 273 573 287 587
rect 333 613 347 627
rect 313 593 327 607
rect 333 573 347 587
rect 293 533 307 547
rect 313 353 327 367
rect 293 313 307 327
rect 313 233 327 247
rect 213 193 227 207
rect 313 193 327 207
rect 133 153 147 167
rect 173 153 187 167
rect 213 133 227 147
rect 353 553 367 567
rect 353 473 367 487
rect 413 653 427 667
rect 533 933 547 947
rect 513 853 527 867
rect 573 853 587 867
rect 573 833 587 847
rect 493 813 507 827
rect 533 793 547 807
rect 533 773 547 787
rect 473 673 487 687
rect 493 653 507 667
rect 513 653 527 667
rect 393 613 407 627
rect 433 613 447 627
rect 613 1073 627 1087
rect 653 1073 667 1087
rect 653 1033 667 1047
rect 613 833 627 847
rect 593 793 607 807
rect 613 693 627 707
rect 573 633 587 647
rect 633 673 647 687
rect 713 1093 727 1107
rect 773 1113 787 1127
rect 813 1113 827 1127
rect 873 1113 887 1127
rect 973 1113 987 1127
rect 693 1073 707 1087
rect 753 1073 767 1087
rect 733 913 747 927
rect 793 1093 807 1107
rect 833 1073 847 1087
rect 793 893 807 907
rect 773 873 787 887
rect 713 853 727 867
rect 773 853 787 867
rect 753 833 767 847
rect 693 773 707 787
rect 753 713 767 727
rect 733 673 747 687
rect 673 653 687 667
rect 713 653 727 667
rect 553 613 567 627
rect 633 613 647 627
rect 653 613 667 627
rect 613 593 627 607
rect 593 573 607 587
rect 453 533 467 547
rect 533 533 547 547
rect 413 513 427 527
rect 373 353 387 367
rect 353 293 367 307
rect 393 293 407 307
rect 413 213 427 227
rect 333 153 347 167
rect 553 453 567 467
rect 613 433 627 447
rect 753 633 767 647
rect 733 593 747 607
rect 693 553 707 567
rect 853 873 867 887
rect 893 853 907 867
rect 933 853 947 867
rect 913 753 927 767
rect 1153 1673 1167 1687
rect 1213 2133 1227 2147
rect 1253 2073 1267 2087
rect 1213 2033 1227 2047
rect 1253 1993 1267 2007
rect 1253 1913 1267 1927
rect 1233 1793 1247 1807
rect 1213 1753 1227 1767
rect 1193 1693 1207 1707
rect 1193 1613 1207 1627
rect 1133 1513 1147 1527
rect 1133 1413 1147 1427
rect 1053 1353 1067 1367
rect 1053 1313 1067 1327
rect 1073 1293 1087 1307
rect 1093 1273 1107 1287
rect 1113 1273 1127 1287
rect 1073 1193 1087 1207
rect 1053 1133 1067 1147
rect 993 1093 1007 1107
rect 1033 1093 1047 1107
rect 973 973 987 987
rect 993 913 1007 927
rect 953 833 967 847
rect 953 773 967 787
rect 1073 1113 1087 1127
rect 1113 1113 1127 1127
rect 1093 1093 1107 1107
rect 1053 753 1067 767
rect 933 733 947 747
rect 833 673 847 687
rect 1033 673 1047 687
rect 1053 673 1067 687
rect 793 633 807 647
rect 853 653 867 667
rect 773 573 787 587
rect 753 473 767 487
rect 673 453 687 467
rect 873 633 887 647
rect 933 633 947 647
rect 953 593 967 607
rect 873 553 887 567
rect 853 453 867 467
rect 673 413 687 427
rect 813 413 827 427
rect 653 353 667 367
rect 733 353 747 367
rect 773 353 787 367
rect 613 333 627 347
rect 633 333 647 347
rect 473 253 487 267
rect 433 193 447 207
rect 473 193 487 207
rect 453 153 467 167
rect 353 133 367 147
rect 73 113 87 127
rect 293 113 307 127
rect 333 113 347 127
rect 533 313 547 327
rect 533 233 547 247
rect 493 153 507 167
rect 613 313 627 327
rect 873 433 887 447
rect 913 373 927 387
rect 893 353 907 367
rect 713 333 727 347
rect 593 293 607 307
rect 653 293 667 307
rect 693 293 707 307
rect 673 213 687 227
rect 573 153 587 167
rect 713 173 727 187
rect 693 153 707 167
rect 853 333 867 347
rect 1013 613 1027 627
rect 1053 613 1067 627
rect 1173 1433 1187 1447
rect 1173 1293 1187 1307
rect 1153 1233 1167 1247
rect 1173 1153 1187 1167
rect 1213 1593 1227 1607
rect 1313 2253 1327 2267
rect 1393 2393 1407 2407
rect 1373 2333 1387 2347
rect 1373 2253 1387 2267
rect 1333 2173 1347 2187
rect 1473 2293 1487 2307
rect 1553 2573 1567 2587
rect 1673 2773 1687 2787
rect 1713 2773 1727 2787
rect 1653 2733 1667 2747
rect 1733 2753 1747 2767
rect 1773 2753 1787 2767
rect 1733 2733 1747 2747
rect 1753 2733 1767 2747
rect 1693 2713 1707 2727
rect 1653 2633 1667 2647
rect 1633 2613 1647 2627
rect 1613 2573 1627 2587
rect 1613 2553 1627 2567
rect 1573 2473 1587 2487
rect 1413 2273 1427 2287
rect 1433 2273 1447 2287
rect 1293 2133 1307 2147
rect 1353 2133 1367 2147
rect 1293 2113 1307 2127
rect 1333 2073 1347 2087
rect 1313 1953 1327 1967
rect 1313 1833 1327 1847
rect 1333 1813 1347 1827
rect 1333 1773 1347 1787
rect 1293 1753 1307 1767
rect 1333 1733 1347 1747
rect 1273 1713 1287 1727
rect 1293 1713 1307 1727
rect 1233 1353 1247 1367
rect 1233 1333 1247 1347
rect 1293 1693 1307 1707
rect 1313 1673 1327 1687
rect 1293 1453 1307 1467
rect 1393 2153 1407 2167
rect 1493 2273 1507 2287
rect 1453 2253 1467 2267
rect 1453 2213 1467 2227
rect 1533 2333 1547 2347
rect 1553 2273 1567 2287
rect 1513 2253 1527 2267
rect 1573 2253 1587 2267
rect 1453 2193 1467 2207
rect 1493 2193 1507 2207
rect 1413 2113 1427 2127
rect 1433 2113 1447 2127
rect 1393 2073 1407 2087
rect 1393 2033 1407 2047
rect 1373 1973 1387 1987
rect 1373 1833 1387 1847
rect 1713 2573 1727 2587
rect 1653 2493 1667 2507
rect 1753 2553 1767 2567
rect 1733 2513 1747 2527
rect 1953 3113 1967 3127
rect 1933 3073 1947 3087
rect 1913 3053 1927 3067
rect 2013 3213 2027 3227
rect 2073 3333 2087 3347
rect 2133 3633 2147 3647
rect 2193 3673 2207 3687
rect 2213 3673 2227 3687
rect 2173 3653 2187 3667
rect 2233 3633 2247 3647
rect 2173 3613 2187 3627
rect 2133 3593 2147 3607
rect 2153 3593 2167 3607
rect 2093 3313 2107 3327
rect 2113 3313 2127 3327
rect 2093 3273 2107 3287
rect 2153 3553 2167 3567
rect 2213 3593 2227 3607
rect 2193 3573 2207 3587
rect 2193 3533 2207 3547
rect 2233 3553 2247 3567
rect 2333 3973 2347 3987
rect 2293 3953 2307 3967
rect 2333 3953 2347 3967
rect 2333 3913 2347 3927
rect 2293 3873 2307 3887
rect 2333 3833 2347 3847
rect 2293 3773 2307 3787
rect 2273 3733 2287 3747
rect 2413 4113 2427 4127
rect 2433 4113 2447 4127
rect 2493 4133 2507 4147
rect 2473 4073 2487 4087
rect 2493 4073 2507 4087
rect 2413 4053 2427 4067
rect 2393 4013 2407 4027
rect 2393 3993 2407 4007
rect 2433 3993 2447 4007
rect 2493 4013 2507 4027
rect 2393 3933 2407 3947
rect 2453 3973 2467 3987
rect 2413 3893 2427 3907
rect 2433 3893 2447 3907
rect 2393 3853 2407 3867
rect 2493 3953 2507 3967
rect 2473 3913 2487 3927
rect 2493 3913 2507 3927
rect 2453 3873 2467 3887
rect 2473 3853 2487 3867
rect 2393 3813 2407 3827
rect 2413 3813 2427 3827
rect 2433 3813 2447 3827
rect 2393 3773 2407 3787
rect 2293 3713 2307 3727
rect 2273 3653 2287 3667
rect 2253 3533 2267 3547
rect 2213 3513 2227 3527
rect 2233 3513 2247 3527
rect 2173 3493 2187 3507
rect 2153 3313 2167 3327
rect 2133 3253 2147 3267
rect 2293 3633 2307 3647
rect 2373 3733 2387 3747
rect 2353 3713 2367 3727
rect 2353 3693 2367 3707
rect 2413 3733 2427 3747
rect 2413 3713 2427 3727
rect 2353 3653 2367 3667
rect 2333 3613 2347 3627
rect 2353 3613 2367 3627
rect 2313 3573 2327 3587
rect 2313 3533 2327 3547
rect 2293 3513 2307 3527
rect 2333 3513 2347 3527
rect 2313 3493 2327 3507
rect 2193 3453 2207 3467
rect 2253 3433 2267 3447
rect 2273 3353 2287 3367
rect 2213 3333 2227 3347
rect 2233 3333 2247 3347
rect 2173 3293 2187 3307
rect 2193 3293 2207 3307
rect 2113 3233 2127 3247
rect 2133 3233 2147 3247
rect 2173 3233 2187 3247
rect 2093 3213 2107 3227
rect 2053 3153 2067 3167
rect 1953 3053 1967 3067
rect 1993 3053 2007 3067
rect 1993 3033 2007 3047
rect 1973 3013 1987 3027
rect 2033 2993 2047 3007
rect 1913 2933 1927 2947
rect 1873 2873 1887 2887
rect 1853 2793 1867 2807
rect 1833 2773 1847 2787
rect 1953 2853 1967 2867
rect 1913 2773 1927 2787
rect 1933 2773 1947 2787
rect 1853 2733 1867 2747
rect 1833 2673 1847 2687
rect 1793 2633 1807 2647
rect 1813 2633 1827 2647
rect 1893 2713 1907 2727
rect 2033 2833 2047 2847
rect 1993 2813 2007 2827
rect 2033 2813 2047 2827
rect 1973 2733 1987 2747
rect 1973 2713 1987 2727
rect 1933 2693 1947 2707
rect 1873 2673 1887 2687
rect 1913 2673 1927 2687
rect 1853 2593 1867 2607
rect 1793 2573 1807 2587
rect 1813 2573 1827 2587
rect 1813 2553 1827 2567
rect 1893 2653 1907 2667
rect 1893 2573 1907 2587
rect 1793 2513 1807 2527
rect 1773 2493 1787 2507
rect 1753 2473 1767 2487
rect 1733 2453 1747 2467
rect 1713 2413 1727 2427
rect 1633 2373 1647 2387
rect 1673 2373 1687 2387
rect 1673 2313 1687 2327
rect 1713 2313 1727 2327
rect 1633 2273 1647 2287
rect 1613 2233 1627 2247
rect 1693 2293 1707 2307
rect 1673 2273 1687 2287
rect 1653 2193 1667 2207
rect 1593 2173 1607 2187
rect 1693 2153 1707 2167
rect 1613 2133 1627 2147
rect 1593 2113 1607 2127
rect 1573 2093 1587 2107
rect 1473 2073 1487 2087
rect 1513 2073 1527 2087
rect 1433 1993 1447 2007
rect 1413 1873 1427 1887
rect 1393 1753 1407 1767
rect 1553 2053 1567 2067
rect 1533 2033 1547 2047
rect 1493 1973 1507 1987
rect 1493 1953 1507 1967
rect 1473 1933 1487 1947
rect 1473 1853 1487 1867
rect 1513 1873 1527 1887
rect 1513 1813 1527 1827
rect 1473 1753 1487 1767
rect 1513 1753 1527 1767
rect 1413 1693 1427 1707
rect 1393 1633 1407 1647
rect 1353 1613 1367 1627
rect 1353 1573 1367 1587
rect 1353 1533 1367 1547
rect 1333 1453 1347 1467
rect 1333 1433 1347 1447
rect 1353 1433 1367 1447
rect 1313 1353 1327 1367
rect 1373 1333 1387 1347
rect 1313 1313 1327 1327
rect 1353 1293 1367 1307
rect 1273 1273 1287 1287
rect 1293 1273 1307 1287
rect 1413 1613 1427 1627
rect 1433 1593 1447 1607
rect 1593 1973 1607 1987
rect 1553 1933 1567 1947
rect 1573 1913 1587 1927
rect 1573 1853 1587 1867
rect 1593 1833 1607 1847
rect 1553 1813 1567 1827
rect 1573 1813 1587 1827
rect 1553 1793 1567 1807
rect 1573 1773 1587 1787
rect 1633 2113 1647 2127
rect 1653 2093 1667 2107
rect 1713 2093 1727 2107
rect 1633 2053 1647 2067
rect 1673 2073 1687 2087
rect 1713 2073 1727 2087
rect 1693 2053 1707 2067
rect 1613 1813 1627 1827
rect 1653 1813 1667 1827
rect 1613 1793 1627 1807
rect 1633 1773 1647 1787
rect 1593 1753 1607 1767
rect 1633 1753 1647 1767
rect 1593 1653 1607 1667
rect 1533 1613 1547 1627
rect 1413 1573 1427 1587
rect 1453 1573 1467 1587
rect 1533 1593 1547 1607
rect 1553 1573 1567 1587
rect 1693 2013 1707 2027
rect 1773 2433 1787 2447
rect 1793 2313 1807 2327
rect 1853 2453 1867 2467
rect 1813 2293 1827 2307
rect 1753 2253 1767 2267
rect 1813 2213 1827 2227
rect 1793 2173 1807 2187
rect 1753 2153 1767 2167
rect 1793 2153 1807 2167
rect 1913 2533 1927 2547
rect 1933 2533 1947 2547
rect 1913 2513 1927 2527
rect 1953 2513 1967 2527
rect 1893 2493 1907 2507
rect 1873 2373 1887 2387
rect 1873 2353 1887 2367
rect 1853 2293 1867 2307
rect 1913 2433 1927 2447
rect 1913 2393 1927 2407
rect 2073 3133 2087 3147
rect 2113 3133 2127 3147
rect 2093 3073 2107 3087
rect 2233 3293 2247 3307
rect 2173 3193 2187 3207
rect 2153 3153 2167 3167
rect 2173 3113 2187 3127
rect 2193 3113 2207 3127
rect 2133 3073 2147 3087
rect 2113 3013 2127 3027
rect 2093 2993 2107 3007
rect 2153 3013 2167 3027
rect 2113 2933 2127 2947
rect 2053 2753 2067 2767
rect 2033 2713 2047 2727
rect 2073 2713 2087 2727
rect 1993 2673 2007 2687
rect 2033 2673 2047 2687
rect 1993 2653 2007 2667
rect 1973 2373 1987 2387
rect 2013 2533 2027 2547
rect 2133 2873 2147 2887
rect 2113 2773 2127 2787
rect 2153 2833 2167 2847
rect 2193 3073 2207 3087
rect 2193 2973 2207 2987
rect 2193 2893 2207 2907
rect 2213 2893 2227 2907
rect 2173 2813 2187 2827
rect 2193 2813 2207 2827
rect 2153 2793 2167 2807
rect 2153 2693 2167 2707
rect 2293 3313 2307 3327
rect 2253 3273 2267 3287
rect 2273 3273 2287 3287
rect 2453 3753 2467 3767
rect 2773 4613 2787 4627
rect 2733 4513 2747 4527
rect 2753 4513 2767 4527
rect 2713 4453 2727 4467
rect 2753 4453 2767 4467
rect 2793 4573 2807 4587
rect 2793 4513 2807 4527
rect 2853 4513 2867 4527
rect 2813 4493 2827 4507
rect 2833 4493 2847 4507
rect 2833 4453 2847 4467
rect 2813 4393 2827 4407
rect 2833 4353 2847 4367
rect 2813 4333 2827 4347
rect 2753 4313 2767 4327
rect 2773 4313 2787 4327
rect 2733 4293 2747 4307
rect 2533 4253 2547 4267
rect 2713 4253 2727 4267
rect 2513 3853 2527 3867
rect 2553 4193 2567 4207
rect 2573 4193 2587 4207
rect 2673 4213 2687 4227
rect 2713 4213 2727 4227
rect 2653 4193 2667 4207
rect 2713 4193 2727 4207
rect 2613 4173 2627 4187
rect 2553 4153 2567 4167
rect 2653 4153 2667 4167
rect 2593 4133 2607 4147
rect 2553 4093 2567 4107
rect 2593 4053 2607 4067
rect 2633 4013 2647 4027
rect 2553 3953 2567 3967
rect 2553 3873 2567 3887
rect 2613 3953 2627 3967
rect 2533 3833 2547 3847
rect 2493 3793 2507 3807
rect 2493 3753 2507 3767
rect 2473 3733 2487 3747
rect 2573 3813 2587 3827
rect 2533 3773 2547 3787
rect 2553 3773 2567 3787
rect 2433 3673 2447 3687
rect 2453 3673 2467 3687
rect 2393 3653 2407 3667
rect 2433 3613 2447 3627
rect 2393 3553 2407 3567
rect 2393 3533 2407 3547
rect 2373 3513 2387 3527
rect 2373 3473 2387 3487
rect 2473 3653 2487 3667
rect 2473 3593 2487 3607
rect 2513 3713 2527 3727
rect 2533 3713 2547 3727
rect 2473 3533 2487 3547
rect 2493 3533 2507 3547
rect 2533 3653 2547 3667
rect 2553 3613 2567 3627
rect 2553 3553 2567 3567
rect 2533 3513 2547 3527
rect 2553 3513 2567 3527
rect 2533 3493 2547 3507
rect 2453 3473 2467 3487
rect 2433 3413 2447 3427
rect 2413 3393 2427 3407
rect 2353 3373 2367 3387
rect 2333 3333 2347 3347
rect 2513 3473 2527 3487
rect 2553 3473 2567 3487
rect 2473 3453 2487 3467
rect 2533 3453 2547 3467
rect 2473 3373 2487 3387
rect 2393 3293 2407 3307
rect 2313 3253 2327 3267
rect 2293 3233 2307 3247
rect 2273 3213 2287 3227
rect 2253 3153 2267 3167
rect 2253 3093 2267 3107
rect 2253 3053 2267 3067
rect 2253 3033 2267 3047
rect 2353 3233 2367 3247
rect 2413 3213 2427 3227
rect 2373 3193 2387 3207
rect 2333 3173 2347 3187
rect 2353 3173 2367 3187
rect 2393 3173 2407 3187
rect 2293 3073 2307 3087
rect 2293 2993 2307 3007
rect 2273 2913 2287 2927
rect 2233 2853 2247 2867
rect 2373 3033 2387 3047
rect 2373 3013 2387 3027
rect 2353 2893 2367 2907
rect 2313 2833 2327 2847
rect 2313 2813 2327 2827
rect 2233 2793 2247 2807
rect 2293 2793 2307 2807
rect 2193 2733 2207 2747
rect 2173 2673 2187 2687
rect 2213 2673 2227 2687
rect 2153 2593 2167 2607
rect 2193 2593 2207 2607
rect 2273 2773 2287 2787
rect 2453 3293 2467 3307
rect 2553 3353 2567 3367
rect 2513 3313 2527 3327
rect 2493 3273 2507 3287
rect 2473 3253 2487 3267
rect 2493 3213 2507 3227
rect 2553 3293 2567 3307
rect 2533 3213 2547 3227
rect 2593 3793 2607 3807
rect 2613 3793 2627 3807
rect 2673 4053 2687 4067
rect 2773 4213 2787 4227
rect 2833 4293 2847 4307
rect 2833 4233 2847 4247
rect 2793 4193 2807 4207
rect 2753 4173 2767 4187
rect 2753 4133 2767 4147
rect 2773 4133 2787 4147
rect 2813 4073 2827 4087
rect 2773 4053 2787 4067
rect 2733 4033 2747 4047
rect 2753 4033 2767 4047
rect 2713 3993 2727 4007
rect 2693 3973 2707 3987
rect 2713 3953 2727 3967
rect 2713 3933 2727 3947
rect 2673 3873 2687 3887
rect 2693 3873 2707 3887
rect 2653 3833 2667 3847
rect 2633 3773 2647 3787
rect 2673 3773 2687 3787
rect 2653 3753 2667 3767
rect 2793 4013 2807 4027
rect 2813 4013 2827 4027
rect 2753 3953 2767 3967
rect 2773 3953 2787 3967
rect 2733 3873 2747 3887
rect 2773 3933 2787 3947
rect 2793 3933 2807 3947
rect 2813 3933 2827 3947
rect 3073 4853 3087 4867
rect 2933 4713 2947 4727
rect 2893 4693 2907 4707
rect 2953 4693 2967 4707
rect 2953 4633 2967 4647
rect 2993 4633 3007 4647
rect 3073 4653 3087 4667
rect 3213 5133 3227 5147
rect 3193 5113 3207 5127
rect 3433 5593 3447 5607
rect 3353 5553 3367 5567
rect 3293 5533 3307 5547
rect 3253 5473 3267 5487
rect 3493 5613 3507 5627
rect 3453 5473 3467 5487
rect 3493 5473 3507 5487
rect 3513 5473 3527 5487
rect 3653 5653 3667 5667
rect 3633 5633 3647 5647
rect 3333 5393 3347 5407
rect 3313 5193 3327 5207
rect 3393 5193 3407 5207
rect 3353 5173 3367 5187
rect 3373 5153 3387 5167
rect 3273 5133 3287 5147
rect 3293 5133 3307 5147
rect 3353 5133 3367 5147
rect 3473 5133 3487 5147
rect 3593 5453 3607 5467
rect 3573 5413 3587 5427
rect 3753 5673 3767 5687
rect 3693 5653 3707 5667
rect 3713 5633 3727 5647
rect 3733 5613 3747 5627
rect 3873 5613 3887 5627
rect 4013 5893 4027 5907
rect 3993 5833 4007 5847
rect 4013 5793 4027 5807
rect 3993 5633 4007 5647
rect 3693 5593 3707 5607
rect 3773 5593 3787 5607
rect 3913 5593 3927 5607
rect 3673 5453 3687 5467
rect 3733 5433 3747 5447
rect 3873 5453 3887 5467
rect 3833 5433 3847 5447
rect 3613 5233 3627 5247
rect 3613 5173 3627 5187
rect 3573 5153 3587 5167
rect 3233 5093 3247 5107
rect 3273 5073 3287 5087
rect 3233 4973 3247 4987
rect 3253 4973 3267 4987
rect 3213 4833 3227 4847
rect 3173 4793 3187 4807
rect 3293 4773 3307 4787
rect 3333 4833 3347 4847
rect 3193 4713 3207 4727
rect 3313 4713 3327 4727
rect 3173 4693 3187 4707
rect 3213 4693 3227 4707
rect 3273 4673 3287 4687
rect 3313 4673 3327 4687
rect 3133 4633 3147 4647
rect 3193 4633 3207 4647
rect 3233 4633 3247 4647
rect 3293 4653 3307 4667
rect 3313 4653 3327 4667
rect 3273 4633 3287 4647
rect 3073 4613 3087 4627
rect 3253 4613 3267 4627
rect 3033 4513 3047 4527
rect 2913 4493 2927 4507
rect 3033 4493 3047 4507
rect 2873 4473 2887 4487
rect 2893 4453 2907 4467
rect 2933 4453 2947 4467
rect 2913 4433 2927 4447
rect 2873 4353 2887 4367
rect 2853 4213 2867 4227
rect 2873 4193 2887 4207
rect 2853 4093 2867 4107
rect 2993 4453 3007 4467
rect 2953 4253 2967 4267
rect 2953 4233 2967 4247
rect 3013 4433 3027 4447
rect 3053 4473 3067 4487
rect 3233 4553 3247 4567
rect 3153 4533 3167 4547
rect 3113 4493 3127 4507
rect 3053 4433 3067 4447
rect 3073 4413 3087 4427
rect 2933 4193 2947 4207
rect 2973 4193 2987 4207
rect 2913 4153 2927 4167
rect 2893 4133 2907 4147
rect 2873 4053 2887 4067
rect 2913 4053 2927 4067
rect 2873 3973 2887 3987
rect 2893 3953 2907 3967
rect 2953 4173 2967 4187
rect 2973 4153 2987 4167
rect 2993 4153 3007 4167
rect 3033 4333 3047 4347
rect 3013 4133 3027 4147
rect 3133 4453 3147 4467
rect 3193 4453 3207 4467
rect 3173 4433 3187 4447
rect 3213 4433 3227 4447
rect 3153 4413 3167 4427
rect 3093 4393 3107 4407
rect 3193 4373 3207 4387
rect 3113 4353 3127 4367
rect 3073 4253 3087 4267
rect 3093 4233 3107 4247
rect 3053 4213 3067 4227
rect 3073 4173 3087 4187
rect 3173 4293 3187 4307
rect 3133 4273 3147 4287
rect 3113 4133 3127 4147
rect 3073 4093 3087 4107
rect 2993 4073 3007 4087
rect 3033 4073 3047 4087
rect 2933 4013 2947 4027
rect 2853 3933 2867 3947
rect 2913 3933 2927 3947
rect 2793 3893 2807 3907
rect 2833 3893 2847 3907
rect 2773 3873 2787 3887
rect 2933 3873 2947 3887
rect 2853 3853 2867 3867
rect 2633 3733 2647 3747
rect 2613 3713 2627 3727
rect 2633 3713 2647 3727
rect 2653 3693 2667 3707
rect 2633 3653 2647 3667
rect 2653 3613 2667 3627
rect 2633 3573 2647 3587
rect 2613 3493 2627 3507
rect 2613 3453 2627 3467
rect 2633 3413 2647 3427
rect 2613 3393 2627 3407
rect 2713 3753 2727 3767
rect 2753 3753 2767 3767
rect 2933 3833 2947 3847
rect 2693 3733 2707 3747
rect 2733 3733 2747 3747
rect 2773 3733 2787 3747
rect 2813 3733 2827 3747
rect 2853 3733 2867 3747
rect 2713 3713 2727 3727
rect 2733 3693 2747 3707
rect 2713 3653 2727 3667
rect 2733 3653 2747 3667
rect 2693 3573 2707 3587
rect 2673 3493 2687 3507
rect 2673 3473 2687 3487
rect 2673 3413 2687 3427
rect 2613 3313 2627 3327
rect 2653 3313 2667 3327
rect 2593 3273 2607 3287
rect 2673 3273 2687 3287
rect 2633 3253 2647 3267
rect 2613 3233 2627 3247
rect 2473 3173 2487 3187
rect 2433 3093 2447 3107
rect 2573 3193 2587 3207
rect 2613 3193 2627 3207
rect 2593 3173 2607 3187
rect 2573 3153 2587 3167
rect 2553 3133 2567 3147
rect 2513 3073 2527 3087
rect 2533 3073 2547 3087
rect 2473 3033 2487 3047
rect 2493 2993 2507 3007
rect 2533 2993 2547 3007
rect 2433 2813 2447 2827
rect 2413 2793 2427 2807
rect 2333 2773 2347 2787
rect 2353 2773 2367 2787
rect 2393 2773 2407 2787
rect 2253 2753 2267 2767
rect 2293 2753 2307 2767
rect 2253 2713 2267 2727
rect 2373 2753 2387 2767
rect 2413 2753 2427 2767
rect 2473 2773 2487 2787
rect 2453 2733 2467 2747
rect 2233 2613 2247 2627
rect 2253 2593 2267 2607
rect 2093 2553 2107 2567
rect 2193 2553 2207 2567
rect 2073 2533 2087 2547
rect 2113 2533 2127 2547
rect 2153 2533 2167 2547
rect 2213 2533 2227 2547
rect 2033 2493 2047 2507
rect 2093 2513 2107 2527
rect 2193 2513 2207 2527
rect 2453 2693 2467 2707
rect 2333 2633 2347 2647
rect 2373 2633 2387 2647
rect 2433 2633 2447 2647
rect 2293 2553 2307 2567
rect 2313 2553 2327 2567
rect 2253 2533 2267 2547
rect 2313 2513 2327 2527
rect 2053 2413 2067 2427
rect 2033 2393 2047 2407
rect 2053 2373 2067 2387
rect 1993 2353 2007 2367
rect 2013 2353 2027 2367
rect 1893 2333 1907 2347
rect 1913 2293 1927 2307
rect 1953 2293 1967 2307
rect 1993 2293 2007 2307
rect 2033 2293 2047 2307
rect 2173 2493 2187 2507
rect 2173 2453 2187 2467
rect 2273 2453 2287 2467
rect 2173 2353 2187 2367
rect 2133 2333 2147 2347
rect 2093 2293 2107 2307
rect 2153 2313 2167 2327
rect 1893 2273 1907 2287
rect 1893 2253 1907 2267
rect 1873 2213 1887 2227
rect 1853 2193 1867 2207
rect 1833 2133 1847 2147
rect 1853 2133 1867 2147
rect 1813 2093 1827 2107
rect 1853 2093 1867 2107
rect 1833 2073 1847 2087
rect 1753 2033 1767 2047
rect 1733 1993 1747 2007
rect 1693 1913 1707 1927
rect 1793 2033 1807 2047
rect 1773 1973 1787 1987
rect 1693 1833 1707 1847
rect 1753 1833 1767 1847
rect 1673 1773 1687 1787
rect 1653 1733 1667 1747
rect 1653 1673 1667 1687
rect 1873 2053 1887 2067
rect 1813 1973 1827 1987
rect 1813 1933 1827 1947
rect 1793 1813 1807 1827
rect 1713 1773 1727 1787
rect 1733 1733 1747 1747
rect 1693 1633 1707 1647
rect 1673 1613 1687 1627
rect 1713 1613 1727 1627
rect 1693 1593 1707 1607
rect 1673 1573 1687 1587
rect 1713 1573 1727 1587
rect 1613 1553 1627 1567
rect 1593 1473 1607 1487
rect 1493 1453 1507 1467
rect 1453 1353 1467 1367
rect 1413 1313 1427 1327
rect 1413 1293 1427 1307
rect 1233 1233 1247 1247
rect 1253 1233 1267 1247
rect 1393 1233 1407 1247
rect 1133 1093 1147 1107
rect 1133 1053 1147 1067
rect 1233 1133 1247 1147
rect 1213 993 1227 1007
rect 1213 933 1227 947
rect 1153 813 1167 827
rect 1193 753 1207 767
rect 1153 693 1167 707
rect 1113 653 1127 667
rect 1093 633 1107 647
rect 1193 673 1207 687
rect 1113 613 1127 627
rect 1073 593 1087 607
rect 1033 473 1047 487
rect 993 433 1007 447
rect 1013 353 1027 367
rect 813 293 827 307
rect 973 293 987 307
rect 753 153 767 167
rect 1073 333 1087 347
rect 1093 293 1107 307
rect 1053 273 1067 287
rect 853 233 867 247
rect 1113 233 1127 247
rect 553 113 567 127
rect 953 173 967 187
rect 913 153 927 167
rect 1033 153 1047 167
rect 1513 1293 1527 1307
rect 1553 1253 1567 1267
rect 1513 1233 1527 1247
rect 1533 1233 1547 1247
rect 1533 1173 1547 1187
rect 1413 1133 1427 1147
rect 1453 1133 1467 1147
rect 1493 1133 1507 1147
rect 1373 1093 1387 1107
rect 1493 1113 1507 1127
rect 1433 1093 1447 1107
rect 1433 1033 1447 1047
rect 1513 1093 1527 1107
rect 1493 1073 1507 1087
rect 1413 933 1427 947
rect 1473 933 1487 947
rect 1393 893 1407 907
rect 1413 893 1427 907
rect 1273 873 1287 887
rect 1313 873 1327 887
rect 1393 873 1407 887
rect 1473 873 1487 887
rect 1313 833 1327 847
rect 1333 833 1347 847
rect 1373 833 1387 847
rect 1273 813 1287 827
rect 1253 753 1267 767
rect 1233 713 1247 727
rect 1353 813 1367 827
rect 1373 793 1387 807
rect 1353 753 1367 767
rect 1373 753 1387 767
rect 1333 713 1347 727
rect 1313 693 1327 707
rect 1353 693 1367 707
rect 1233 673 1247 687
rect 1293 673 1307 687
rect 1273 653 1287 667
rect 1233 633 1247 647
rect 1453 833 1467 847
rect 1573 1193 1587 1207
rect 1613 1373 1627 1387
rect 1773 1773 1787 1787
rect 2013 2273 2027 2287
rect 2053 2273 2067 2287
rect 1973 2233 1987 2247
rect 1933 2193 1947 2207
rect 1913 2173 1927 2187
rect 1933 2093 1947 2107
rect 1913 1953 1927 1967
rect 1953 1953 1967 1967
rect 1953 1913 1967 1927
rect 2053 2253 2067 2267
rect 2113 2273 2127 2287
rect 2073 2193 2087 2207
rect 2093 2193 2107 2207
rect 1993 2153 2007 2167
rect 2073 2153 2087 2167
rect 2053 2133 2067 2147
rect 2033 2093 2047 2107
rect 2013 2073 2027 2087
rect 1993 1993 2007 2007
rect 1993 1913 2007 1927
rect 1893 1873 1907 1887
rect 1933 1873 1947 1887
rect 1853 1853 1867 1867
rect 1893 1853 1907 1867
rect 1833 1813 1847 1827
rect 1813 1753 1827 1767
rect 1773 1733 1787 1747
rect 1753 1653 1767 1667
rect 1753 1593 1767 1607
rect 1793 1713 1807 1727
rect 1793 1653 1807 1667
rect 1913 1793 1927 1807
rect 1933 1753 1947 1767
rect 1873 1713 1887 1727
rect 1893 1713 1907 1727
rect 1833 1613 1847 1627
rect 1933 1613 1947 1627
rect 1813 1593 1827 1607
rect 1733 1373 1747 1387
rect 1673 1353 1687 1367
rect 1653 1333 1667 1347
rect 1713 1333 1727 1347
rect 1693 1313 1707 1327
rect 1633 1293 1647 1307
rect 1653 1253 1667 1267
rect 1613 1213 1627 1227
rect 1613 1153 1627 1167
rect 1593 1133 1607 1147
rect 1573 1113 1587 1127
rect 1793 1573 1807 1587
rect 1813 1553 1827 1567
rect 1833 1553 1847 1567
rect 1813 1513 1827 1527
rect 1833 1493 1847 1507
rect 2053 1973 2067 1987
rect 2133 2133 2147 2147
rect 2113 2073 2127 2087
rect 2133 2013 2147 2027
rect 2113 1993 2127 2007
rect 2073 1873 2087 1887
rect 2013 1853 2027 1867
rect 2053 1853 2067 1867
rect 2053 1813 2067 1827
rect 1993 1793 2007 1807
rect 2033 1773 2047 1787
rect 2033 1753 2047 1767
rect 2013 1733 2027 1747
rect 1973 1693 1987 1707
rect 1993 1673 2007 1687
rect 1993 1633 2007 1647
rect 2053 1733 2067 1747
rect 2013 1593 2027 1607
rect 2033 1593 2047 1607
rect 2073 1653 2087 1667
rect 1953 1473 1967 1487
rect 1973 1473 1987 1487
rect 1933 1453 1947 1467
rect 2033 1453 2047 1467
rect 1973 1433 1987 1447
rect 1933 1413 1947 1427
rect 1853 1393 1867 1407
rect 1773 1333 1787 1347
rect 1813 1333 1827 1347
rect 1933 1373 1947 1387
rect 1853 1313 1867 1327
rect 1913 1313 1927 1327
rect 1753 1293 1767 1307
rect 1753 1253 1767 1267
rect 1733 1193 1747 1207
rect 1693 1173 1707 1187
rect 1713 1173 1727 1187
rect 1753 1173 1767 1187
rect 1673 1153 1687 1167
rect 1693 1133 1707 1147
rect 1733 1113 1747 1127
rect 1513 1053 1527 1067
rect 1553 1053 1567 1067
rect 1613 1073 1627 1087
rect 1573 933 1587 947
rect 1533 893 1547 907
rect 1573 893 1587 907
rect 1633 1053 1647 1067
rect 1733 1093 1747 1107
rect 1773 1133 1787 1147
rect 1873 1293 1887 1307
rect 1853 1273 1867 1287
rect 1833 1233 1847 1247
rect 1833 1113 1847 1127
rect 1893 1253 1907 1267
rect 1913 1133 1927 1147
rect 1973 1313 1987 1327
rect 1993 1293 2007 1307
rect 1953 1273 1967 1287
rect 1973 1273 1987 1287
rect 1953 1253 1967 1267
rect 1993 1233 2007 1247
rect 1973 1173 1987 1187
rect 1953 1153 1967 1167
rect 1853 1073 1867 1087
rect 1753 1053 1767 1067
rect 1693 1033 1707 1047
rect 1733 973 1747 987
rect 1753 973 1767 987
rect 1773 933 1787 947
rect 1833 933 1847 947
rect 1753 893 1767 907
rect 1773 893 1787 907
rect 1613 833 1627 847
rect 1593 813 1607 827
rect 1573 793 1587 807
rect 1693 833 1707 847
rect 1733 833 1747 847
rect 1673 813 1687 827
rect 1513 733 1527 747
rect 1553 733 1567 747
rect 1413 673 1427 687
rect 1493 673 1507 687
rect 1293 633 1307 647
rect 1433 653 1447 667
rect 1513 653 1527 667
rect 1553 653 1567 667
rect 1313 613 1327 627
rect 1333 613 1347 627
rect 1213 453 1227 467
rect 1293 593 1307 607
rect 1253 433 1267 447
rect 1233 373 1247 387
rect 1153 353 1167 367
rect 1193 353 1207 367
rect 1153 333 1167 347
rect 1153 293 1167 307
rect 1213 333 1227 347
rect 1173 213 1187 227
rect 1153 193 1167 207
rect 1193 173 1207 187
rect 1413 633 1427 647
rect 1393 613 1407 627
rect 1453 633 1467 647
rect 1513 633 1527 647
rect 1353 593 1367 607
rect 1433 533 1447 547
rect 1333 413 1347 427
rect 1313 373 1327 387
rect 1253 333 1267 347
rect 1273 333 1287 347
rect 1313 313 1327 327
rect 1353 373 1367 387
rect 1293 293 1307 307
rect 1333 293 1347 307
rect 1453 493 1467 507
rect 1493 573 1507 587
rect 1513 573 1527 587
rect 1533 573 1547 587
rect 1493 393 1507 407
rect 1473 373 1487 387
rect 1593 633 1607 647
rect 1653 613 1667 627
rect 1713 793 1727 807
rect 1693 773 1707 787
rect 1713 773 1727 787
rect 1733 733 1747 747
rect 1713 693 1727 707
rect 1733 653 1747 667
rect 1693 613 1707 627
rect 1773 813 1787 827
rect 1793 793 1807 807
rect 1773 733 1787 747
rect 1753 613 1767 627
rect 1793 633 1807 647
rect 1673 593 1687 607
rect 1713 593 1727 607
rect 1753 593 1767 607
rect 1933 1113 1947 1127
rect 1933 1033 1947 1047
rect 1873 953 1887 967
rect 2073 1333 2087 1347
rect 2193 2293 2207 2307
rect 2233 2293 2247 2307
rect 2173 2273 2187 2287
rect 2213 2273 2227 2287
rect 2233 2253 2247 2267
rect 2253 2253 2267 2267
rect 2193 2153 2207 2167
rect 2173 2133 2187 2147
rect 2173 2033 2187 2047
rect 2153 1933 2167 1947
rect 2173 1913 2187 1927
rect 2113 1873 2127 1887
rect 2253 2153 2267 2167
rect 2233 2133 2247 2147
rect 2253 2113 2267 2127
rect 2293 2393 2307 2407
rect 2313 2393 2327 2407
rect 2413 2553 2427 2567
rect 2353 2533 2367 2547
rect 2393 2533 2407 2547
rect 2393 2513 2407 2527
rect 2373 2493 2387 2507
rect 2353 2473 2367 2487
rect 2333 2373 2347 2387
rect 2333 2353 2347 2367
rect 2293 2293 2307 2307
rect 2293 2253 2307 2267
rect 2293 2153 2307 2167
rect 2273 2073 2287 2087
rect 2233 2053 2247 2067
rect 2153 1853 2167 1867
rect 2213 1853 2227 1867
rect 2173 1833 2187 1847
rect 2133 1753 2147 1767
rect 2113 1693 2127 1707
rect 2153 1693 2167 1707
rect 2133 1593 2147 1607
rect 2213 1813 2227 1827
rect 2193 1733 2207 1747
rect 2173 1533 2187 1547
rect 2213 1713 2227 1727
rect 2253 1773 2267 1787
rect 2313 2133 2327 2147
rect 2513 2933 2527 2947
rect 2613 3073 2627 3087
rect 2613 3053 2627 3067
rect 2593 2893 2607 2907
rect 2513 2793 2527 2807
rect 2573 2793 2587 2807
rect 2513 2773 2527 2787
rect 2533 2753 2547 2767
rect 2513 2713 2527 2727
rect 2493 2653 2507 2667
rect 2473 2613 2487 2627
rect 2473 2573 2487 2587
rect 2453 2553 2467 2567
rect 2433 2473 2447 2487
rect 2453 2473 2467 2487
rect 2453 2433 2467 2447
rect 2393 2413 2407 2427
rect 2373 2293 2387 2307
rect 2413 2393 2427 2407
rect 2453 2393 2467 2407
rect 2433 2333 2447 2347
rect 2413 2293 2427 2307
rect 2573 2753 2587 2767
rect 2553 2673 2567 2687
rect 2653 3193 2667 3207
rect 2653 3173 2667 3187
rect 2753 3613 2767 3627
rect 2773 3613 2787 3627
rect 2753 3593 2767 3607
rect 2733 3513 2747 3527
rect 2753 3513 2767 3527
rect 2813 3673 2827 3687
rect 2793 3593 2807 3607
rect 2793 3533 2807 3547
rect 2693 3253 2707 3267
rect 2693 3213 2707 3227
rect 2753 3473 2767 3487
rect 2933 3713 2947 3727
rect 2833 3633 2847 3647
rect 2913 3613 2927 3627
rect 2893 3593 2907 3607
rect 2853 3533 2867 3547
rect 2973 4033 2987 4047
rect 3053 4053 3067 4067
rect 3013 4033 3027 4047
rect 3033 4013 3047 4027
rect 3013 3993 3027 4007
rect 3053 3993 3067 4007
rect 2973 3953 2987 3967
rect 3013 3953 3027 3967
rect 3013 3933 3027 3947
rect 2973 3853 2987 3867
rect 3053 3853 3067 3867
rect 3053 3833 3067 3847
rect 3033 3793 3047 3807
rect 2973 3773 2987 3787
rect 2993 3773 3007 3787
rect 3013 3713 3027 3727
rect 2973 3673 2987 3687
rect 3153 4233 3167 4247
rect 3173 4093 3187 4107
rect 3213 4073 3227 4087
rect 3253 4513 3267 4527
rect 3333 4633 3347 4647
rect 3453 5053 3467 5067
rect 3433 4973 3447 4987
rect 3393 4953 3407 4967
rect 3453 4933 3467 4947
rect 3413 4873 3427 4887
rect 3433 4693 3447 4707
rect 3413 4673 3427 4687
rect 3373 4613 3387 4627
rect 3353 4533 3367 4547
rect 3333 4473 3347 4487
rect 3273 4453 3287 4467
rect 3313 4453 3327 4467
rect 3273 4393 3287 4407
rect 3273 4373 3287 4387
rect 3253 4213 3267 4227
rect 3413 4473 3427 4487
rect 3433 4473 3447 4487
rect 3353 4433 3367 4447
rect 3353 4333 3367 4347
rect 3333 4233 3347 4247
rect 3413 4233 3427 4247
rect 3293 4193 3307 4207
rect 3353 4213 3367 4227
rect 3333 4193 3347 4207
rect 3333 4173 3347 4187
rect 3313 4153 3327 4167
rect 3273 4093 3287 4107
rect 3193 4053 3207 4067
rect 3233 4053 3247 4067
rect 3253 4053 3267 4067
rect 3153 4033 3167 4047
rect 3093 4013 3107 4027
rect 3133 4013 3147 4027
rect 3073 3773 3087 3787
rect 3173 4013 3187 4027
rect 3113 3953 3127 3967
rect 3173 3953 3187 3967
rect 3133 3913 3147 3927
rect 3113 3853 3127 3867
rect 3093 3753 3107 3767
rect 3073 3713 3087 3727
rect 3113 3713 3127 3727
rect 3093 3633 3107 3647
rect 3253 4013 3267 4027
rect 3233 3993 3247 4007
rect 3233 3973 3247 3987
rect 3253 3953 3267 3967
rect 3213 3933 3227 3947
rect 3193 3833 3207 3847
rect 3153 3793 3167 3807
rect 3173 3753 3187 3767
rect 3213 3753 3227 3767
rect 3153 3713 3167 3727
rect 3133 3613 3147 3627
rect 3053 3593 3067 3607
rect 3073 3593 3087 3607
rect 2953 3573 2967 3587
rect 3053 3573 3067 3587
rect 3093 3573 3107 3587
rect 2933 3553 2947 3567
rect 3033 3553 3047 3567
rect 3013 3533 3027 3547
rect 2813 3493 2827 3507
rect 2833 3493 2847 3507
rect 2793 3393 2807 3407
rect 2893 3473 2907 3487
rect 2873 3453 2887 3467
rect 2773 3353 2787 3367
rect 2813 3353 2827 3367
rect 2753 3293 2767 3307
rect 2733 3233 2747 3247
rect 2713 3113 2727 3127
rect 2673 3073 2687 3087
rect 2653 3033 2667 3047
rect 2693 3033 2707 3047
rect 2773 3253 2787 3267
rect 2873 3373 2887 3387
rect 2873 3273 2887 3287
rect 2753 3213 2767 3227
rect 2793 3213 2807 3227
rect 2773 3193 2787 3207
rect 2753 3073 2767 3087
rect 2633 2993 2647 3007
rect 2633 2893 2647 2907
rect 2653 2893 2667 2907
rect 2573 2613 2587 2627
rect 2513 2593 2527 2607
rect 2553 2593 2567 2607
rect 2553 2573 2567 2587
rect 2613 2613 2627 2627
rect 2593 2553 2607 2567
rect 2513 2513 2527 2527
rect 2513 2413 2527 2427
rect 2493 2333 2507 2347
rect 2473 2313 2487 2327
rect 2493 2293 2507 2307
rect 2473 2273 2487 2287
rect 2393 2233 2407 2247
rect 2433 2233 2447 2247
rect 2473 2233 2487 2247
rect 2373 2213 2387 2227
rect 2393 2213 2407 2227
rect 2373 2173 2387 2187
rect 2353 2153 2367 2167
rect 2413 2173 2427 2187
rect 2593 2493 2607 2507
rect 2713 2993 2727 3007
rect 2733 2993 2747 3007
rect 2693 2913 2707 2927
rect 2673 2853 2687 2867
rect 2673 2773 2687 2787
rect 2673 2733 2687 2747
rect 2713 2693 2727 2707
rect 2753 2953 2767 2967
rect 2793 3073 2807 3087
rect 2873 3253 2887 3267
rect 2833 3233 2847 3247
rect 2853 3213 2867 3227
rect 2833 3133 2847 3147
rect 2813 3053 2827 3067
rect 2873 3033 2887 3047
rect 2813 3013 2827 3027
rect 2853 3013 2867 3027
rect 2973 3513 2987 3527
rect 2953 3493 2967 3507
rect 2993 3473 3007 3487
rect 2913 3373 2927 3387
rect 2993 3353 3007 3367
rect 2973 3293 2987 3307
rect 2913 3273 2927 3287
rect 2953 3253 2967 3267
rect 2933 3173 2947 3187
rect 2913 3093 2927 3107
rect 2893 2973 2907 2987
rect 2853 2853 2867 2867
rect 3013 3273 3027 3287
rect 3053 3253 3067 3267
rect 3033 3233 3047 3247
rect 3013 3213 3027 3227
rect 2993 3193 3007 3207
rect 3033 3193 3047 3207
rect 3013 3173 3027 3187
rect 2953 3073 2967 3087
rect 3053 3113 3067 3127
rect 3073 3113 3087 3127
rect 2853 2833 2867 2847
rect 2913 2833 2927 2847
rect 2793 2753 2807 2767
rect 2913 2773 2927 2787
rect 2893 2753 2907 2767
rect 2733 2633 2747 2647
rect 2753 2633 2767 2647
rect 2633 2593 2647 2607
rect 2653 2593 2667 2607
rect 2693 2593 2707 2607
rect 2753 2593 2767 2607
rect 2693 2573 2707 2587
rect 2793 2553 2807 2567
rect 2633 2513 2647 2527
rect 2613 2453 2627 2467
rect 2573 2433 2587 2447
rect 2593 2433 2607 2447
rect 2593 2393 2607 2407
rect 2613 2393 2627 2407
rect 2533 2333 2547 2347
rect 2593 2313 2607 2327
rect 2553 2293 2567 2307
rect 2513 2273 2527 2287
rect 2593 2273 2607 2287
rect 2573 2253 2587 2267
rect 2533 2233 2547 2247
rect 2573 2233 2587 2247
rect 2453 2153 2467 2167
rect 2413 2093 2427 2107
rect 2433 2093 2447 2107
rect 2533 2193 2547 2207
rect 2553 2093 2567 2107
rect 2473 2073 2487 2087
rect 2513 2073 2527 2087
rect 2333 1973 2347 1987
rect 2453 2053 2467 2067
rect 2413 1993 2427 2007
rect 2433 1993 2447 2007
rect 2373 1913 2387 1927
rect 2373 1853 2387 1867
rect 2413 1853 2427 1867
rect 2313 1833 2327 1847
rect 2313 1793 2327 1807
rect 2333 1793 2347 1807
rect 2293 1753 2307 1767
rect 2273 1733 2287 1747
rect 2233 1653 2247 1667
rect 2253 1653 2267 1667
rect 2213 1613 2227 1627
rect 2293 1713 2307 1727
rect 2293 1593 2307 1607
rect 2193 1493 2207 1507
rect 2273 1573 2287 1587
rect 2253 1453 2267 1467
rect 2193 1433 2207 1447
rect 2233 1433 2247 1447
rect 2173 1353 2187 1367
rect 2093 1293 2107 1307
rect 2113 1293 2127 1307
rect 2073 1273 2087 1287
rect 2033 1253 2047 1267
rect 2073 1193 2087 1207
rect 2113 1193 2127 1207
rect 2053 1153 2067 1167
rect 1953 933 1967 947
rect 2033 1073 2047 1087
rect 1993 953 2007 967
rect 1993 913 2007 927
rect 1973 873 1987 887
rect 1933 853 1947 867
rect 1953 853 1967 867
rect 2053 913 2067 927
rect 2093 1153 2107 1167
rect 2073 873 2087 887
rect 2013 853 2027 867
rect 2073 853 2087 867
rect 2153 1233 2167 1247
rect 2153 1193 2167 1207
rect 2133 1153 2147 1167
rect 2133 1133 2147 1147
rect 2153 1113 2167 1127
rect 2233 1373 2247 1387
rect 2353 1753 2367 1767
rect 2333 1733 2347 1747
rect 2393 1753 2407 1767
rect 2373 1713 2387 1727
rect 2393 1713 2407 1727
rect 2513 2033 2527 2047
rect 2493 2013 2507 2027
rect 2473 1913 2487 1927
rect 2453 1873 2467 1887
rect 2473 1813 2487 1827
rect 2553 2033 2567 2047
rect 2533 1973 2547 1987
rect 2513 1873 2527 1887
rect 2513 1813 2527 1827
rect 2453 1773 2467 1787
rect 2493 1773 2507 1787
rect 2433 1673 2447 1687
rect 2493 1753 2507 1767
rect 2773 2533 2787 2547
rect 2733 2473 2747 2487
rect 2753 2473 2767 2487
rect 2713 2413 2727 2427
rect 2673 2273 2687 2287
rect 2773 2413 2787 2427
rect 2753 2293 2767 2307
rect 2753 2273 2767 2287
rect 2633 2233 2647 2247
rect 2693 2253 2707 2267
rect 2673 2213 2687 2227
rect 2653 2193 2667 2207
rect 2653 2153 2667 2167
rect 2693 2153 2707 2167
rect 2633 2073 2647 2087
rect 2613 2053 2627 2067
rect 2613 1993 2627 2007
rect 2673 2093 2687 2107
rect 2733 2093 2747 2107
rect 2873 2733 2887 2747
rect 2893 2713 2907 2727
rect 2873 2673 2887 2687
rect 2853 2633 2867 2647
rect 2893 2573 2907 2587
rect 2893 2553 2907 2567
rect 2873 2433 2887 2447
rect 2833 2393 2847 2407
rect 2813 2373 2827 2387
rect 2833 2353 2847 2367
rect 2793 2333 2807 2347
rect 2673 2053 2687 2067
rect 2653 1953 2667 1967
rect 2673 1953 2687 1967
rect 2553 1793 2567 1807
rect 2573 1773 2587 1787
rect 2533 1753 2547 1767
rect 2573 1733 2587 1747
rect 2513 1713 2527 1727
rect 2493 1693 2507 1707
rect 2533 1673 2547 1687
rect 2553 1653 2567 1667
rect 2473 1633 2487 1647
rect 2533 1633 2547 1647
rect 2453 1613 2467 1627
rect 2473 1613 2487 1627
rect 2333 1573 2347 1587
rect 2353 1553 2367 1567
rect 2313 1533 2327 1547
rect 2333 1513 2347 1527
rect 2353 1513 2367 1527
rect 2413 1573 2427 1587
rect 2413 1473 2427 1487
rect 2333 1453 2347 1467
rect 2373 1453 2387 1467
rect 2313 1433 2327 1447
rect 2353 1413 2367 1427
rect 2373 1393 2387 1407
rect 2213 1273 2227 1287
rect 2313 1273 2327 1287
rect 2273 1213 2287 1227
rect 2273 1173 2287 1187
rect 2213 1153 2227 1167
rect 2253 1113 2267 1127
rect 2193 1013 2207 1027
rect 2273 1093 2287 1107
rect 2233 973 2247 987
rect 2133 873 2147 887
rect 2093 833 2107 847
rect 1913 793 1927 807
rect 2013 793 2027 807
rect 2053 793 2067 807
rect 1933 773 1947 787
rect 1913 733 1927 747
rect 1933 733 1947 747
rect 1873 713 1887 727
rect 1853 693 1867 707
rect 1893 693 1907 707
rect 1873 633 1887 647
rect 1853 613 1867 627
rect 1813 593 1827 607
rect 1713 573 1727 587
rect 1793 573 1807 587
rect 1613 553 1627 567
rect 1573 533 1587 547
rect 1693 513 1707 527
rect 1673 433 1687 447
rect 1613 413 1627 427
rect 1533 393 1547 407
rect 1573 393 1587 407
rect 1453 353 1467 367
rect 1373 333 1387 347
rect 1373 293 1387 307
rect 1313 173 1327 187
rect 1353 173 1367 187
rect 1433 333 1447 347
rect 1513 333 1527 347
rect 1473 313 1487 327
rect 1413 253 1427 267
rect 1453 193 1467 207
rect 1233 153 1247 167
rect 1273 153 1287 167
rect 1353 153 1367 167
rect 1133 133 1147 147
rect 1333 133 1347 147
rect 1553 353 1567 367
rect 1493 153 1507 167
rect 1533 153 1547 167
rect 1653 373 1667 387
rect 1653 353 1667 367
rect 1693 353 1707 367
rect 1593 313 1607 327
rect 1613 213 1627 227
rect 1633 213 1647 227
rect 1593 193 1607 207
rect 1653 173 1667 187
rect 1693 333 1707 347
rect 1733 513 1747 527
rect 1813 513 1827 527
rect 1813 453 1827 467
rect 1913 673 1927 687
rect 1953 653 1967 667
rect 1933 633 1947 647
rect 2033 713 2047 727
rect 1933 533 1947 547
rect 1953 533 1967 547
rect 2013 413 2027 427
rect 1893 393 1907 407
rect 1853 353 1867 367
rect 1893 353 1907 367
rect 1953 353 1967 367
rect 1713 313 1727 327
rect 1693 233 1707 247
rect 1733 153 1747 167
rect 1393 133 1407 147
rect 1433 133 1447 147
rect 1553 133 1567 147
rect 1673 133 1687 147
rect 1793 333 1807 347
rect 1833 313 1847 327
rect 1773 273 1787 287
rect 1793 253 1807 267
rect 1933 253 1947 267
rect 2133 813 2147 827
rect 2353 1293 2367 1307
rect 2333 1253 2347 1267
rect 2353 1193 2367 1207
rect 2413 1353 2427 1367
rect 2413 1313 2427 1327
rect 2393 1293 2407 1307
rect 2393 1273 2407 1287
rect 2413 1233 2427 1247
rect 2393 1193 2407 1207
rect 2373 1173 2387 1187
rect 2333 1113 2347 1127
rect 2393 1133 2407 1147
rect 2433 1193 2447 1207
rect 2433 1173 2447 1187
rect 2633 1813 2647 1827
rect 2773 1993 2787 2007
rect 2733 1973 2747 1987
rect 2713 1933 2727 1947
rect 2713 1793 2727 1807
rect 2593 1673 2607 1687
rect 2693 1773 2707 1787
rect 2713 1713 2727 1727
rect 2653 1653 2667 1667
rect 2753 1953 2767 1967
rect 2873 2333 2887 2347
rect 2813 2273 2827 2287
rect 2833 2273 2847 2287
rect 2813 2153 2827 2167
rect 2873 2193 2887 2207
rect 2853 2113 2867 2127
rect 2993 3033 3007 3047
rect 3113 3513 3127 3527
rect 3113 3373 3127 3387
rect 3133 3273 3147 3287
rect 3113 3253 3127 3267
rect 3133 3193 3147 3207
rect 3133 3153 3147 3167
rect 3113 3133 3127 3147
rect 3253 3733 3267 3747
rect 3213 3713 3227 3727
rect 3193 3693 3207 3707
rect 3233 3693 3247 3707
rect 3213 3673 3227 3687
rect 3193 3633 3207 3647
rect 3193 3573 3207 3587
rect 3313 4053 3327 4067
rect 3293 4033 3307 4047
rect 3513 5113 3527 5127
rect 3713 5413 3727 5427
rect 3753 5413 3767 5427
rect 3933 5473 3947 5487
rect 3853 5393 3867 5407
rect 3873 5393 3887 5407
rect 3673 5173 3687 5187
rect 3973 5413 3987 5427
rect 3933 5393 3947 5407
rect 3993 5373 4007 5387
rect 3973 5353 3987 5367
rect 3693 5153 3707 5167
rect 3793 5153 3807 5167
rect 3833 5153 3847 5167
rect 3893 5153 3907 5167
rect 3933 5153 3947 5167
rect 3673 5133 3687 5147
rect 3813 5133 3827 5147
rect 3613 4973 3627 4987
rect 3653 4973 3667 4987
rect 3553 4953 3567 4967
rect 3633 4953 3647 4967
rect 3733 4973 3747 4987
rect 3773 4973 3787 4987
rect 3713 4953 3727 4967
rect 3533 4933 3547 4947
rect 3613 4933 3627 4947
rect 3653 4933 3667 4947
rect 3533 4813 3547 4827
rect 3513 4673 3527 4687
rect 3573 4693 3587 4707
rect 3493 4613 3507 4627
rect 3613 4673 3627 4687
rect 3633 4653 3647 4667
rect 3513 4493 3527 4507
rect 3493 4473 3507 4487
rect 3533 4453 3547 4467
rect 3473 4433 3487 4447
rect 3473 4393 3487 4407
rect 3513 4393 3527 4407
rect 3453 4193 3467 4207
rect 3433 4173 3447 4187
rect 3393 4153 3407 4167
rect 3393 4073 3407 4087
rect 3353 4033 3367 4047
rect 3333 3993 3347 4007
rect 3313 3973 3327 3987
rect 3293 3913 3307 3927
rect 3293 3893 3307 3907
rect 3313 3813 3327 3827
rect 3353 3773 3367 3787
rect 3413 3913 3427 3927
rect 3413 3813 3427 3827
rect 3333 3713 3347 3727
rect 3353 3713 3367 3727
rect 3393 3713 3407 3727
rect 3293 3693 3307 3707
rect 3313 3673 3327 3687
rect 3253 3633 3267 3647
rect 3273 3633 3287 3647
rect 3253 3593 3267 3607
rect 3193 3553 3207 3567
rect 3233 3553 3247 3567
rect 3173 3373 3187 3387
rect 3233 3513 3247 3527
rect 3193 3333 3207 3347
rect 3193 3313 3207 3327
rect 3293 3613 3307 3627
rect 3273 3453 3287 3467
rect 3253 3433 3267 3447
rect 3253 3413 3267 3427
rect 3333 3653 3347 3667
rect 3313 3593 3327 3607
rect 3393 3613 3407 3627
rect 3373 3553 3387 3567
rect 3313 3533 3327 3547
rect 3453 4133 3467 4147
rect 3493 4333 3507 4347
rect 3633 4633 3647 4647
rect 3593 4513 3607 4527
rect 3573 4493 3587 4507
rect 3713 4813 3727 4827
rect 3633 4473 3647 4487
rect 3813 4953 3827 4967
rect 3833 4953 3847 4967
rect 3793 4933 3807 4947
rect 3753 4813 3767 4827
rect 3733 4753 3747 4767
rect 3833 4853 3847 4867
rect 3953 5133 3967 5147
rect 3993 5113 4007 5127
rect 3973 5053 3987 5067
rect 4213 6113 4227 6127
rect 4373 6113 4387 6127
rect 4493 6113 4507 6127
rect 4553 6113 4567 6127
rect 4593 6113 4607 6127
rect 4633 6113 4647 6127
rect 4693 6113 4707 6127
rect 4273 6093 4287 6107
rect 4193 6073 4207 6087
rect 4333 6073 4347 6087
rect 4113 6013 4127 6027
rect 4153 6013 4167 6027
rect 4253 6013 4267 6027
rect 4273 5953 4287 5967
rect 4153 5913 4167 5927
rect 4093 5893 4107 5907
rect 4133 5893 4147 5907
rect 4053 5793 4067 5807
rect 4033 5773 4047 5787
rect 4053 5773 4067 5787
rect 4113 5673 4127 5687
rect 4053 5653 4067 5667
rect 4033 5633 4047 5647
rect 4073 5633 4087 5647
rect 4053 5393 4067 5407
rect 4033 5373 4047 5387
rect 4073 5153 4087 5167
rect 4073 5133 4087 5147
rect 4213 5913 4227 5927
rect 4473 6053 4487 6067
rect 4273 5913 4287 5927
rect 4273 5873 4287 5887
rect 4293 5873 4307 5887
rect 4193 5673 4207 5687
rect 4213 5653 4227 5667
rect 4433 5913 4447 5927
rect 4633 6073 4647 6087
rect 4673 6073 4687 6087
rect 4713 6073 4727 6087
rect 4573 6053 4587 6067
rect 4613 6053 4627 6067
rect 4533 6033 4547 6047
rect 4493 6013 4507 6027
rect 4513 5913 4527 5927
rect 4573 5993 4587 6007
rect 4573 5953 4587 5967
rect 4653 5933 4667 5947
rect 4673 5913 4687 5927
rect 4413 5873 4427 5887
rect 4373 5853 4387 5867
rect 4333 5673 4347 5687
rect 4193 5633 4207 5647
rect 4273 5633 4287 5647
rect 4293 5633 4307 5647
rect 4153 5473 4167 5487
rect 4313 5613 4327 5627
rect 4353 5613 4367 5627
rect 4253 5493 4267 5507
rect 4173 5453 4187 5467
rect 4353 5473 4367 5487
rect 4413 5713 4427 5727
rect 4393 5593 4407 5607
rect 4433 5573 4447 5587
rect 4633 5893 4647 5907
rect 4733 6013 4747 6027
rect 4853 6153 4867 6167
rect 4993 6153 5007 6167
rect 4773 6113 4787 6127
rect 4813 6113 4827 6127
rect 4893 6133 4907 6147
rect 4953 6133 4967 6147
rect 5013 6133 5027 6147
rect 4873 6113 4887 6127
rect 4853 6073 4867 6087
rect 4973 6113 4987 6127
rect 4973 6093 4987 6107
rect 4933 6073 4947 6087
rect 4893 6053 4907 6067
rect 4913 6053 4927 6067
rect 4953 6053 4967 6067
rect 4813 6013 4827 6027
rect 4753 5993 4767 6007
rect 4753 5933 4767 5947
rect 4953 5953 4967 5967
rect 4853 5933 4867 5947
rect 4713 5893 4727 5907
rect 4733 5893 4747 5907
rect 4773 5913 4787 5927
rect 4813 5913 4827 5927
rect 4853 5913 4867 5927
rect 4753 5873 4767 5887
rect 4773 5793 4787 5807
rect 4593 5753 4607 5767
rect 4633 5753 4647 5767
rect 4553 5673 4567 5687
rect 4513 5633 4527 5647
rect 4553 5633 4567 5647
rect 4473 5573 4487 5587
rect 4533 5573 4547 5587
rect 4613 5693 4627 5707
rect 4613 5673 4627 5687
rect 4693 5653 4707 5667
rect 4773 5653 4787 5667
rect 4653 5593 4667 5607
rect 4593 5573 4607 5587
rect 4653 5573 4667 5587
rect 4673 5573 4687 5587
rect 4393 5533 4407 5547
rect 4453 5533 4467 5547
rect 4573 5533 4587 5547
rect 4273 5453 4287 5467
rect 4353 5453 4367 5467
rect 4373 5453 4387 5467
rect 4253 5413 4267 5427
rect 4313 5413 4327 5427
rect 4513 5513 4527 5527
rect 4433 5453 4447 5467
rect 4453 5453 4467 5467
rect 4493 5453 4507 5467
rect 4373 5373 4387 5387
rect 4413 5373 4427 5387
rect 4333 5353 4347 5367
rect 4253 5333 4267 5347
rect 4133 5313 4147 5327
rect 4213 5313 4227 5327
rect 4233 5313 4247 5327
rect 4333 5313 4347 5327
rect 4113 5173 4127 5187
rect 4093 5113 4107 5127
rect 4153 5153 4167 5167
rect 4193 5133 4207 5147
rect 4053 5053 4067 5067
rect 4013 4973 4027 4987
rect 3873 4953 3887 4967
rect 3913 4953 3927 4967
rect 3933 4933 3947 4947
rect 3893 4913 3907 4927
rect 3933 4913 3947 4927
rect 3913 4853 3927 4867
rect 3833 4793 3847 4807
rect 3853 4793 3867 4807
rect 3813 4753 3827 4767
rect 3793 4713 3807 4727
rect 3753 4673 3767 4687
rect 3793 4673 3807 4687
rect 3873 4713 3887 4727
rect 3953 4773 3967 4787
rect 3813 4633 3827 4647
rect 3773 4613 3787 4627
rect 3733 4593 3747 4607
rect 3773 4593 3787 4607
rect 3733 4473 3747 4487
rect 3893 4633 3907 4647
rect 3933 4633 3947 4647
rect 3853 4493 3867 4507
rect 3813 4473 3827 4487
rect 3713 4453 3727 4467
rect 3613 4433 3627 4447
rect 3593 4413 3607 4427
rect 3553 4353 3567 4367
rect 3553 4233 3567 4247
rect 3533 4213 3547 4227
rect 3473 4113 3487 4127
rect 3453 3813 3467 3827
rect 3473 3653 3487 3667
rect 3493 3653 3507 3667
rect 3333 3493 3347 3507
rect 3393 3493 3407 3507
rect 3433 3493 3447 3507
rect 3393 3473 3407 3487
rect 3413 3473 3427 3487
rect 3353 3453 3367 3467
rect 3353 3393 3367 3407
rect 3393 3393 3407 3407
rect 3313 3353 3327 3367
rect 3293 3273 3307 3287
rect 3233 3253 3247 3267
rect 3253 3253 3267 3267
rect 3233 3233 3247 3247
rect 3273 3233 3287 3247
rect 3293 3233 3307 3247
rect 3173 3213 3187 3227
rect 3173 3193 3187 3207
rect 3153 3093 3167 3107
rect 3073 3073 3087 3087
rect 2953 3013 2967 3027
rect 2973 3013 2987 3027
rect 3013 3013 3027 3027
rect 3053 3013 3067 3027
rect 3013 2973 3027 2987
rect 2973 2813 2987 2827
rect 2953 2793 2967 2807
rect 3053 2793 3067 2807
rect 2973 2773 2987 2787
rect 2953 2753 2967 2767
rect 2933 2613 2947 2627
rect 2933 2573 2947 2587
rect 2933 2513 2947 2527
rect 2933 2433 2947 2447
rect 2933 2233 2947 2247
rect 2953 2233 2967 2247
rect 2953 2173 2967 2187
rect 2913 2153 2927 2167
rect 2953 2153 2967 2167
rect 2913 2093 2927 2107
rect 2853 2053 2867 2067
rect 2833 2033 2847 2047
rect 2813 2013 2827 2027
rect 2933 2053 2947 2067
rect 2893 2033 2907 2047
rect 2833 1993 2847 2007
rect 2853 1993 2867 2007
rect 2793 1913 2807 1927
rect 2813 1833 2827 1847
rect 2773 1793 2787 1807
rect 2893 1813 2907 1827
rect 2853 1793 2867 1807
rect 2773 1713 2787 1727
rect 2873 1773 2887 1787
rect 2833 1753 2847 1767
rect 2933 1793 2947 1807
rect 2913 1753 2927 1767
rect 2873 1713 2887 1727
rect 2893 1713 2907 1727
rect 2793 1693 2807 1707
rect 2753 1673 2767 1687
rect 2853 1673 2867 1687
rect 2673 1633 2687 1647
rect 2733 1633 2747 1647
rect 2573 1613 2587 1627
rect 2593 1613 2607 1627
rect 2533 1553 2547 1567
rect 2573 1553 2587 1567
rect 2613 1533 2627 1547
rect 2613 1513 2627 1527
rect 2653 1513 2667 1527
rect 2573 1493 2587 1507
rect 2573 1473 2587 1487
rect 2513 1353 2527 1367
rect 2473 1313 2487 1327
rect 2553 1313 2567 1327
rect 2653 1453 2667 1467
rect 2593 1433 2607 1447
rect 2493 1293 2507 1307
rect 2573 1293 2587 1307
rect 2473 1273 2487 1287
rect 2533 1273 2547 1287
rect 2553 1273 2567 1287
rect 2473 1213 2487 1227
rect 2433 1133 2447 1147
rect 2453 1133 2467 1147
rect 2413 1113 2427 1127
rect 2353 1093 2367 1107
rect 2373 1073 2387 1087
rect 2413 1073 2427 1087
rect 2333 1033 2347 1047
rect 2313 1013 2327 1027
rect 2153 793 2167 807
rect 2053 653 2067 667
rect 2093 653 2107 667
rect 2093 633 2107 647
rect 2113 613 2127 627
rect 2093 593 2107 607
rect 2073 553 2087 567
rect 2073 533 2087 547
rect 2013 333 2027 347
rect 2053 333 2067 347
rect 2193 793 2207 807
rect 2213 693 2227 707
rect 2173 653 2187 667
rect 2173 633 2187 647
rect 2273 673 2287 687
rect 2253 633 2267 647
rect 2233 613 2247 627
rect 2193 573 2207 587
rect 2233 533 2247 547
rect 2213 393 2227 407
rect 2233 373 2247 387
rect 2253 373 2267 387
rect 2233 353 2247 367
rect 1993 253 2007 267
rect 1913 213 1927 227
rect 1973 213 1987 227
rect 1813 193 1827 207
rect 1773 153 1787 167
rect 1993 193 2007 207
rect 1953 173 1967 187
rect 1993 153 2007 167
rect 2033 153 2047 167
rect 2133 333 2147 347
rect 2153 333 2167 347
rect 2113 273 2127 287
rect 2153 293 2167 307
rect 2253 273 2267 287
rect 2073 253 2087 267
rect 2133 253 2147 267
rect 2193 253 2207 267
rect 1793 133 1807 147
rect 2053 133 2067 147
rect 1753 113 1767 127
rect 2113 133 2127 147
rect 2413 953 2427 967
rect 2393 933 2407 947
rect 2373 893 2387 907
rect 2453 1073 2467 1087
rect 2493 1073 2507 1087
rect 2513 1073 2527 1087
rect 2513 1053 2527 1067
rect 2533 1053 2547 1067
rect 2453 1033 2467 1047
rect 2493 993 2507 1007
rect 2493 953 2507 967
rect 2473 913 2487 927
rect 2513 913 2527 927
rect 2513 873 2527 887
rect 2393 813 2407 827
rect 2433 813 2447 827
rect 2433 693 2447 707
rect 2353 673 2367 687
rect 2293 653 2307 667
rect 2333 653 2347 667
rect 2313 613 2327 627
rect 2413 613 2427 627
rect 2293 573 2307 587
rect 2413 553 2427 567
rect 2353 413 2367 427
rect 2293 333 2307 347
rect 2373 353 2387 367
rect 2293 213 2307 227
rect 2273 173 2287 187
rect 2153 153 2167 167
rect 2193 153 2207 167
rect 2333 133 2347 147
rect 2473 673 2487 687
rect 2493 593 2507 607
rect 2473 373 2487 387
rect 2573 1073 2587 1087
rect 2613 1313 2627 1327
rect 2733 1593 2747 1607
rect 2793 1633 2807 1647
rect 2693 1513 2707 1527
rect 2753 1513 2767 1527
rect 2813 1613 2827 1627
rect 2833 1613 2847 1627
rect 2813 1493 2827 1507
rect 2753 1413 2767 1427
rect 2793 1413 2807 1427
rect 2673 1373 2687 1387
rect 2733 1373 2747 1387
rect 2753 1373 2767 1387
rect 2693 1333 2707 1347
rect 2613 1293 2627 1307
rect 2613 1193 2627 1207
rect 2633 1193 2647 1207
rect 2613 1173 2627 1187
rect 2673 1173 2687 1187
rect 2713 1313 2727 1327
rect 2713 1193 2727 1207
rect 2653 1153 2667 1167
rect 2693 1153 2707 1167
rect 2593 1053 2607 1067
rect 2553 1033 2567 1047
rect 2673 1113 2687 1127
rect 2713 1113 2727 1127
rect 2653 1073 2667 1087
rect 2673 1053 2687 1067
rect 2633 1013 2647 1027
rect 2553 993 2567 1007
rect 2573 893 2587 907
rect 2553 853 2567 867
rect 2553 813 2567 827
rect 2553 633 2567 647
rect 2593 853 2607 867
rect 2593 813 2607 827
rect 2653 813 2667 827
rect 2693 1033 2707 1047
rect 2933 1713 2947 1727
rect 2953 1693 2967 1707
rect 2893 1593 2907 1607
rect 2933 1593 2947 1607
rect 2873 1573 2887 1587
rect 2833 1433 2847 1447
rect 2853 1433 2867 1447
rect 2813 1333 2827 1347
rect 2773 1313 2787 1327
rect 2753 1233 2767 1247
rect 2793 1233 2807 1247
rect 2793 1193 2807 1207
rect 2793 1173 2807 1187
rect 2813 1173 2827 1187
rect 2773 1093 2787 1107
rect 2833 1153 2847 1167
rect 2913 1413 2927 1427
rect 3013 2753 3027 2767
rect 3133 3053 3147 3067
rect 3153 3053 3167 3067
rect 3093 2993 3107 3007
rect 3133 2993 3147 3007
rect 3073 2773 3087 2787
rect 3113 2753 3127 2767
rect 3073 2733 3087 2747
rect 3033 2713 3047 2727
rect 3033 2693 3047 2707
rect 2993 2673 3007 2687
rect 3013 2613 3027 2627
rect 2993 2593 3007 2607
rect 3013 2573 3027 2587
rect 3013 2553 3027 2567
rect 3073 2653 3087 2667
rect 3093 2653 3107 2667
rect 3053 2573 3067 2587
rect 2993 2253 3007 2267
rect 3113 2553 3127 2567
rect 3113 2533 3127 2547
rect 3073 2413 3087 2427
rect 3053 2393 3067 2407
rect 3053 2373 3067 2387
rect 3073 2353 3087 2367
rect 3113 2353 3127 2367
rect 3053 2253 3067 2267
rect 3053 2133 3067 2147
rect 3013 2113 3027 2127
rect 3013 2073 3027 2087
rect 3013 2053 3027 2067
rect 2993 2033 3007 2047
rect 2993 2013 3007 2027
rect 2993 1813 3007 1827
rect 3013 1773 3027 1787
rect 3033 1773 3047 1787
rect 3033 1673 3047 1687
rect 2993 1653 3007 1667
rect 3013 1633 3027 1647
rect 3153 2673 3167 2687
rect 3253 3173 3267 3187
rect 3213 3153 3227 3167
rect 3193 3113 3207 3127
rect 3333 3313 3347 3327
rect 3353 3313 3367 3327
rect 3373 3273 3387 3287
rect 3353 3253 3367 3267
rect 3333 3153 3347 3167
rect 3353 3153 3367 3167
rect 3293 3073 3307 3087
rect 3233 3053 3247 3067
rect 3313 3053 3327 3067
rect 3273 3033 3287 3047
rect 3213 3013 3227 3027
rect 3253 3013 3267 3027
rect 3253 2973 3267 2987
rect 3213 2753 3227 2767
rect 3173 2533 3187 2547
rect 3173 2413 3187 2427
rect 3113 2313 3127 2327
rect 3133 2313 3147 2327
rect 3113 2293 3127 2307
rect 3153 2273 3167 2287
rect 3093 2253 3107 2267
rect 3133 2253 3147 2267
rect 3073 2113 3087 2127
rect 3073 2093 3087 2107
rect 3113 2233 3127 2247
rect 3173 2213 3187 2227
rect 3233 2713 3247 2727
rect 3233 2613 3247 2627
rect 3273 2713 3287 2727
rect 3273 2693 3287 2707
rect 3273 2673 3287 2687
rect 3433 3413 3447 3427
rect 3433 3373 3447 3387
rect 3413 3253 3427 3267
rect 3393 3233 3407 3247
rect 3433 3233 3447 3247
rect 3573 4153 3587 4167
rect 3533 4133 3547 4147
rect 3693 4433 3707 4447
rect 3653 4353 3667 4367
rect 3613 4213 3627 4227
rect 3793 4453 3807 4467
rect 3833 4453 3847 4467
rect 3813 4433 3827 4447
rect 3793 4353 3807 4367
rect 3753 4333 3767 4347
rect 3733 4313 3747 4327
rect 3693 4233 3707 4247
rect 3653 4173 3667 4187
rect 3673 4173 3687 4187
rect 3613 4153 3627 4167
rect 3693 4153 3707 4167
rect 3713 4153 3727 4167
rect 3593 4113 3607 4127
rect 3613 4073 3627 4087
rect 3593 4013 3607 4027
rect 3553 3953 3567 3967
rect 3813 4253 3827 4267
rect 3553 3773 3567 3787
rect 3533 3673 3547 3687
rect 3493 3553 3507 3567
rect 3513 3553 3527 3567
rect 3613 3713 3627 3727
rect 3593 3593 3607 3607
rect 3533 3533 3547 3547
rect 3573 3533 3587 3547
rect 3553 3513 3567 3527
rect 3533 3493 3547 3507
rect 3493 3473 3507 3487
rect 3473 3433 3487 3447
rect 3393 3193 3407 3207
rect 3413 3073 3427 3087
rect 3373 3053 3387 3067
rect 3393 3053 3407 3067
rect 3333 3033 3347 3047
rect 3413 3033 3427 3047
rect 3313 3013 3327 3027
rect 3393 3013 3407 3027
rect 3353 2993 3367 3007
rect 3313 2953 3327 2967
rect 3393 2913 3407 2927
rect 3413 2873 3427 2887
rect 3313 2853 3327 2867
rect 3253 2573 3267 2587
rect 3273 2573 3287 2587
rect 3293 2573 3307 2587
rect 3233 2453 3247 2467
rect 3213 2313 3227 2327
rect 3293 2533 3307 2547
rect 3353 2793 3367 2807
rect 3453 3193 3467 3207
rect 3513 3453 3527 3467
rect 3553 3433 3567 3447
rect 3493 3353 3507 3367
rect 3513 3353 3527 3367
rect 3553 3313 3567 3327
rect 3493 3273 3507 3287
rect 3533 3253 3547 3267
rect 3573 3273 3587 3287
rect 3733 4073 3747 4087
rect 3713 3853 3727 3867
rect 3673 3693 3687 3707
rect 3713 3693 3727 3707
rect 3653 3673 3667 3687
rect 3693 3673 3707 3687
rect 3633 3573 3647 3587
rect 3713 3553 3727 3567
rect 3613 3533 3627 3547
rect 3693 3513 3707 3527
rect 3633 3413 3647 3427
rect 3693 3473 3707 3487
rect 3673 3333 3687 3347
rect 3653 3293 3667 3307
rect 3593 3253 3607 3267
rect 3633 3233 3647 3247
rect 3673 3273 3687 3287
rect 3493 3213 3507 3227
rect 3513 3213 3527 3227
rect 3473 3133 3487 3147
rect 3473 3053 3487 3067
rect 3533 3193 3547 3207
rect 3473 3033 3487 3047
rect 3513 3033 3527 3047
rect 3593 3213 3607 3227
rect 3653 3213 3667 3227
rect 3613 3193 3627 3207
rect 3553 3133 3567 3147
rect 3573 3113 3587 3127
rect 3713 3273 3727 3287
rect 3693 3213 3707 3227
rect 3633 3113 3647 3127
rect 3673 3113 3687 3127
rect 3613 3073 3627 3087
rect 3553 3033 3567 3047
rect 3573 3013 3587 3027
rect 3533 2973 3547 2987
rect 3473 2953 3487 2967
rect 3453 2793 3467 2807
rect 3373 2773 3387 2787
rect 3413 2773 3427 2787
rect 3433 2773 3447 2787
rect 3353 2753 3367 2767
rect 3353 2733 3367 2747
rect 3413 2753 3427 2767
rect 3453 2753 3467 2767
rect 3433 2693 3447 2707
rect 3433 2613 3447 2627
rect 3333 2573 3347 2587
rect 3373 2573 3387 2587
rect 3313 2473 3327 2487
rect 3413 2553 3427 2567
rect 3313 2393 3327 2407
rect 3333 2393 3347 2407
rect 3273 2333 3287 2347
rect 3293 2333 3307 2347
rect 3253 2293 3267 2307
rect 3233 2273 3247 2287
rect 3153 2153 3167 2167
rect 3193 2153 3207 2167
rect 3113 2133 3127 2147
rect 3113 2033 3127 2047
rect 3113 1913 3127 1927
rect 3053 1613 3067 1627
rect 3053 1593 3067 1607
rect 3113 1813 3127 1827
rect 3133 1793 3147 1807
rect 3113 1653 3127 1667
rect 3193 2073 3207 2087
rect 3233 2233 3247 2247
rect 3253 2213 3267 2227
rect 3353 2373 3367 2387
rect 3413 2513 3427 2527
rect 3393 2493 3407 2507
rect 3673 3033 3687 3047
rect 3713 3033 3727 3047
rect 3613 2993 3627 3007
rect 3593 2973 3607 2987
rect 3573 2933 3587 2947
rect 3533 2873 3547 2887
rect 3493 2853 3507 2867
rect 3533 2753 3547 2767
rect 3553 2753 3567 2767
rect 3513 2733 3527 2747
rect 3493 2713 3507 2727
rect 3573 2673 3587 2687
rect 3513 2653 3527 2667
rect 3493 2633 3507 2647
rect 3553 2613 3567 2627
rect 3473 2573 3487 2587
rect 3433 2493 3447 2507
rect 3413 2453 3427 2467
rect 3513 2553 3527 2567
rect 3493 2533 3507 2547
rect 3533 2533 3547 2547
rect 3573 2453 3587 2467
rect 3453 2433 3467 2447
rect 3453 2413 3467 2427
rect 3493 2413 3507 2427
rect 3413 2353 3427 2367
rect 3333 2313 3347 2327
rect 3373 2313 3387 2327
rect 3313 2293 3327 2307
rect 3293 2253 3307 2267
rect 3233 2113 3247 2127
rect 3273 2113 3287 2127
rect 3273 2093 3287 2107
rect 3313 2213 3327 2227
rect 3313 2073 3327 2087
rect 3233 1973 3247 1987
rect 3173 1913 3187 1927
rect 3153 1733 3167 1747
rect 3153 1653 3167 1667
rect 3133 1613 3147 1627
rect 2993 1573 3007 1587
rect 3073 1573 3087 1587
rect 3033 1553 3047 1567
rect 3073 1513 3087 1527
rect 2973 1413 2987 1427
rect 2933 1333 2947 1347
rect 2953 1333 2967 1347
rect 2873 1313 2887 1327
rect 2913 1313 2927 1327
rect 2873 1293 2887 1307
rect 2913 1293 2927 1307
rect 2873 1173 2887 1187
rect 2913 1173 2927 1187
rect 2813 1133 2827 1147
rect 2853 1133 2867 1147
rect 2873 1133 2887 1147
rect 2853 1113 2867 1127
rect 2833 1093 2847 1107
rect 2873 1093 2887 1107
rect 2793 1053 2807 1067
rect 2733 1013 2747 1027
rect 2713 933 2727 947
rect 2713 913 2727 927
rect 2693 833 2707 847
rect 2833 973 2847 987
rect 2813 953 2827 967
rect 2733 893 2747 907
rect 2693 813 2707 827
rect 2713 813 2727 827
rect 2773 813 2787 827
rect 3053 1313 3067 1327
rect 2933 1033 2947 1047
rect 2873 933 2887 947
rect 2913 933 2927 947
rect 2833 833 2847 847
rect 2893 853 2907 867
rect 2933 853 2947 867
rect 2733 793 2747 807
rect 2673 773 2687 787
rect 2613 733 2627 747
rect 2633 633 2647 647
rect 2733 733 2747 747
rect 2713 713 2727 727
rect 2813 793 2827 807
rect 2793 693 2807 707
rect 2753 633 2767 647
rect 2893 653 2907 667
rect 2653 613 2667 627
rect 2713 613 2727 627
rect 2733 613 2747 627
rect 2773 613 2787 627
rect 2593 573 2607 587
rect 2813 573 2827 587
rect 2853 553 2867 567
rect 2593 533 2607 547
rect 2793 533 2807 547
rect 2573 413 2587 427
rect 2753 413 2767 427
rect 2573 393 2587 407
rect 2493 353 2507 367
rect 2613 353 2627 367
rect 2593 333 2607 347
rect 2813 433 2827 447
rect 2433 313 2447 327
rect 2593 193 2607 207
rect 2793 333 2807 347
rect 2973 1293 2987 1307
rect 2973 1153 2987 1167
rect 2973 1113 2987 1127
rect 3053 1253 3067 1267
rect 3073 1193 3087 1207
rect 3053 1153 3067 1167
rect 3113 1453 3127 1467
rect 3293 1973 3307 1987
rect 3373 2273 3387 2287
rect 3473 2293 3487 2307
rect 3453 2273 3467 2287
rect 3393 2253 3407 2267
rect 3353 2233 3367 2247
rect 3373 2233 3387 2247
rect 3453 2233 3467 2247
rect 3433 2213 3447 2227
rect 3373 2193 3387 2207
rect 3433 2193 3447 2207
rect 3393 2173 3407 2187
rect 3433 2113 3447 2127
rect 3413 2093 3427 2107
rect 3433 2093 3447 2107
rect 3393 2053 3407 2067
rect 3353 2013 3367 2027
rect 3333 1913 3347 1927
rect 3253 1833 3267 1847
rect 3333 1833 3347 1847
rect 3253 1813 3267 1827
rect 3313 1793 3327 1807
rect 3273 1773 3287 1787
rect 3213 1753 3227 1767
rect 3253 1753 3267 1767
rect 3193 1733 3207 1747
rect 3113 1373 3127 1387
rect 3173 1373 3187 1387
rect 3093 1133 3107 1147
rect 3173 1313 3187 1327
rect 3313 1693 3327 1707
rect 3213 1653 3227 1667
rect 3233 1633 3247 1647
rect 3273 1633 3287 1647
rect 3353 1793 3367 1807
rect 3473 2153 3487 2167
rect 3453 2073 3467 2087
rect 3453 2053 3467 2067
rect 3453 1993 3467 2007
rect 3433 1813 3447 1827
rect 3413 1793 3427 1807
rect 3393 1773 3407 1787
rect 3373 1613 3387 1627
rect 3433 1613 3447 1627
rect 3513 2253 3527 2267
rect 3553 2253 3567 2267
rect 3533 2213 3547 2227
rect 3693 2953 3707 2967
rect 3653 2913 3667 2927
rect 3673 2833 3687 2847
rect 3613 2813 3627 2827
rect 3633 2813 3647 2827
rect 3633 2753 3647 2767
rect 3613 2733 3627 2747
rect 3693 2813 3707 2827
rect 3713 2813 3727 2827
rect 3613 2713 3627 2727
rect 3633 2713 3647 2727
rect 3633 2593 3647 2607
rect 3613 2573 3627 2587
rect 3653 2573 3667 2587
rect 3613 2533 3627 2547
rect 3593 2413 3607 2427
rect 3593 2393 3607 2407
rect 3533 2173 3547 2187
rect 3573 2173 3587 2187
rect 3493 2093 3507 2107
rect 3513 2073 3527 2087
rect 3473 1793 3487 1807
rect 3473 1773 3487 1787
rect 3513 2013 3527 2027
rect 3513 1873 3527 1887
rect 3613 2353 3627 2367
rect 3613 2273 3627 2287
rect 3613 2253 3627 2267
rect 3613 2193 3627 2207
rect 3573 2113 3587 2127
rect 3593 2113 3607 2127
rect 3593 2093 3607 2107
rect 3553 2053 3567 2067
rect 3593 2013 3607 2027
rect 3553 1933 3567 1947
rect 3513 1793 3527 1807
rect 3533 1793 3547 1807
rect 3473 1713 3487 1727
rect 3493 1613 3507 1627
rect 3253 1573 3267 1587
rect 3293 1573 3307 1587
rect 3393 1593 3407 1607
rect 3433 1593 3447 1607
rect 3453 1593 3467 1607
rect 3493 1593 3507 1607
rect 3293 1553 3307 1567
rect 3213 1493 3227 1507
rect 3253 1373 3267 1387
rect 3233 1333 3247 1347
rect 3213 1293 3227 1307
rect 3213 1273 3227 1287
rect 3173 1173 3187 1187
rect 3133 1133 3147 1147
rect 3153 1133 3167 1147
rect 3153 1113 3167 1127
rect 2993 1093 3007 1107
rect 3173 1093 3187 1107
rect 3193 1093 3207 1107
rect 3033 1073 3047 1087
rect 3093 1073 3107 1087
rect 3053 933 3067 947
rect 3013 873 3027 887
rect 2973 853 2987 867
rect 2993 833 3007 847
rect 2953 673 2967 687
rect 3013 633 3027 647
rect 2933 553 2947 567
rect 2913 433 2927 447
rect 3033 613 3047 627
rect 2973 413 2987 427
rect 3173 1013 3187 1027
rect 3313 1313 3327 1327
rect 3293 1273 3307 1287
rect 3473 1553 3487 1567
rect 3533 1733 3547 1747
rect 3533 1713 3547 1727
rect 3573 1853 3587 1867
rect 3673 2473 3687 2487
rect 3673 2393 3687 2407
rect 3653 2093 3667 2107
rect 3653 2073 3667 2087
rect 3633 2013 3647 2027
rect 3613 1973 3627 1987
rect 3653 1973 3667 1987
rect 3633 1813 3647 1827
rect 3573 1773 3587 1787
rect 3573 1753 3587 1767
rect 3553 1693 3567 1707
rect 3593 1733 3607 1747
rect 3553 1653 3567 1667
rect 3553 1593 3567 1607
rect 3773 3993 3787 4007
rect 3933 4453 3947 4467
rect 3873 4433 3887 4447
rect 3853 4393 3867 4407
rect 3913 4333 3927 4347
rect 3833 4193 3847 4207
rect 3873 4193 3887 4207
rect 3893 4173 3907 4187
rect 3873 4153 3887 4167
rect 3833 4013 3847 4027
rect 3853 4013 3867 4027
rect 3853 3973 3867 3987
rect 3993 4933 4007 4947
rect 3973 4713 3987 4727
rect 4013 4713 4027 4727
rect 3973 4693 3987 4707
rect 3993 4673 4007 4687
rect 3993 4453 4007 4467
rect 4013 4413 4027 4427
rect 4113 4953 4127 4967
rect 4173 4873 4187 4887
rect 4133 4713 4147 4727
rect 4073 4693 4087 4707
rect 4093 4693 4107 4707
rect 4153 4693 4167 4707
rect 4053 4573 4067 4587
rect 4073 4493 4087 4507
rect 4173 4593 4187 4607
rect 4173 4573 4187 4587
rect 4113 4553 4127 4567
rect 4153 4553 4167 4567
rect 4093 4473 4107 4487
rect 4093 4433 4107 4447
rect 4113 4413 4127 4427
rect 4113 4393 4127 4407
rect 4053 4373 4067 4387
rect 3973 4313 3987 4327
rect 4033 4133 4047 4147
rect 3913 4013 3927 4027
rect 3953 4013 3967 4027
rect 3933 3993 3947 4007
rect 3973 3993 3987 4007
rect 3953 3973 3967 3987
rect 3873 3773 3887 3787
rect 3813 3733 3827 3747
rect 3853 3733 3867 3747
rect 3753 3713 3767 3727
rect 3813 3713 3827 3727
rect 3793 3653 3807 3667
rect 3833 3613 3847 3627
rect 3813 3493 3827 3507
rect 3773 3453 3787 3467
rect 3793 3353 3807 3367
rect 3773 3253 3787 3267
rect 4093 4193 4107 4207
rect 4073 4153 4087 4167
rect 4073 4013 4087 4027
rect 4053 3953 4067 3967
rect 4293 5293 4307 5307
rect 4253 5153 4267 5167
rect 4313 5133 4327 5147
rect 4273 5113 4287 5127
rect 4213 5093 4227 5107
rect 4353 5133 4367 5147
rect 4333 5033 4347 5047
rect 4413 5213 4427 5227
rect 4393 5093 4407 5107
rect 4533 5453 4547 5467
rect 4513 5433 4527 5447
rect 4533 5433 4547 5447
rect 4573 5433 4587 5447
rect 4453 5333 4467 5347
rect 4493 5413 4507 5427
rect 4473 5313 4487 5327
rect 4713 5633 4727 5647
rect 4753 5613 4767 5627
rect 4793 5613 4807 5627
rect 4733 5593 4747 5607
rect 4753 5593 4767 5607
rect 4893 5873 4907 5887
rect 4953 5913 4967 5927
rect 4953 5853 4967 5867
rect 4933 5753 4947 5767
rect 5033 6113 5047 6127
rect 5033 6093 5047 6107
rect 5013 6033 5027 6047
rect 4993 5933 5007 5947
rect 4973 5673 4987 5687
rect 5213 6133 5227 6147
rect 5273 6133 5287 6147
rect 5473 6153 5487 6167
rect 5533 6153 5547 6167
rect 5613 6153 5627 6167
rect 6113 6153 6127 6167
rect 6173 6153 6187 6167
rect 6273 6153 6287 6167
rect 6393 6153 6407 6167
rect 7033 6153 7047 6167
rect 5293 6113 5307 6127
rect 5173 6033 5187 6047
rect 5093 6013 5107 6027
rect 5113 6013 5127 6027
rect 5093 5953 5107 5967
rect 5073 5913 5087 5927
rect 5153 5933 5167 5947
rect 5053 5773 5067 5787
rect 5033 5713 5047 5727
rect 4953 5653 4967 5667
rect 5013 5653 5027 5667
rect 5033 5653 5047 5667
rect 4873 5633 4887 5647
rect 4913 5633 4927 5647
rect 4833 5613 4847 5627
rect 4733 5573 4747 5587
rect 4813 5573 4827 5587
rect 4833 5553 4847 5567
rect 4693 5513 4707 5527
rect 4713 5513 4727 5527
rect 4793 5513 4807 5527
rect 4813 5513 4827 5527
rect 4673 5433 4687 5447
rect 4513 5393 4527 5407
rect 4553 5393 4567 5407
rect 4573 5393 4587 5407
rect 4553 5373 4567 5387
rect 4493 5293 4507 5307
rect 4473 5233 4487 5247
rect 4633 5413 4647 5427
rect 4653 5413 4667 5427
rect 4653 5393 4667 5407
rect 4613 5353 4627 5367
rect 4653 5353 4667 5367
rect 4573 5333 4587 5347
rect 4613 5253 4627 5267
rect 4553 5193 4567 5207
rect 4593 5193 4607 5207
rect 4473 5173 4487 5187
rect 4513 5173 4527 5187
rect 4453 5133 4467 5147
rect 4493 5093 4507 5107
rect 4433 5053 4447 5067
rect 4473 5033 4487 5047
rect 4453 5013 4467 5027
rect 4373 4993 4387 5007
rect 4233 4953 4247 4967
rect 4413 4953 4427 4967
rect 4333 4933 4347 4947
rect 4393 4933 4407 4947
rect 4433 4933 4447 4947
rect 4233 4913 4247 4927
rect 4313 4913 4327 4927
rect 4233 4693 4247 4707
rect 4353 4753 4367 4767
rect 4293 4733 4307 4747
rect 4253 4673 4267 4687
rect 4213 4593 4227 4607
rect 4193 4513 4207 4527
rect 4313 4673 4327 4687
rect 4333 4653 4347 4667
rect 4453 4673 4467 4687
rect 4473 4653 4487 4667
rect 4573 5133 4587 5147
rect 4533 5053 4547 5067
rect 4533 4973 4547 4987
rect 4613 5173 4627 5187
rect 4713 5393 4727 5407
rect 4673 5293 4687 5307
rect 4693 5293 4707 5307
rect 4633 5133 4647 5147
rect 4653 5133 4667 5147
rect 4713 5193 4727 5207
rect 4753 5433 4767 5447
rect 4893 5613 4907 5627
rect 4893 5593 4907 5607
rect 4853 5533 4867 5547
rect 4853 5493 4867 5507
rect 4873 5473 4887 5487
rect 4853 5393 4867 5407
rect 4973 5613 4987 5627
rect 4933 5573 4947 5587
rect 4953 5573 4967 5587
rect 4913 5513 4927 5527
rect 4893 5453 4907 5467
rect 5013 5573 5027 5587
rect 4993 5553 5007 5567
rect 4953 5533 4967 5547
rect 4973 5513 4987 5527
rect 4953 5433 4967 5447
rect 5313 6053 5327 6067
rect 5293 5953 5307 5967
rect 5253 5913 5267 5927
rect 5273 5893 5287 5907
rect 5173 5733 5187 5747
rect 5213 5733 5227 5747
rect 5113 5693 5127 5707
rect 5093 5653 5107 5667
rect 5113 5653 5127 5667
rect 5153 5653 5167 5667
rect 5053 5633 5067 5647
rect 5073 5573 5087 5587
rect 5053 5553 5067 5567
rect 5033 5433 5047 5447
rect 5013 5413 5027 5427
rect 4853 5333 4867 5347
rect 4833 5273 4847 5287
rect 4773 5233 4787 5247
rect 4733 5173 4747 5187
rect 4733 5153 4747 5167
rect 4773 5153 4787 5167
rect 4673 5093 4687 5107
rect 4753 5113 4767 5127
rect 4693 5033 4707 5047
rect 4513 4653 4527 4667
rect 4513 4593 4527 4607
rect 4493 4573 4507 4587
rect 4233 4533 4247 4547
rect 4253 4493 4267 4507
rect 4233 4413 4247 4427
rect 4193 4393 4207 4407
rect 4173 4353 4187 4367
rect 4173 4313 4187 4327
rect 4153 4253 4167 4267
rect 4453 4553 4467 4567
rect 4313 4533 4327 4547
rect 4313 4513 4327 4527
rect 4293 4293 4307 4307
rect 4193 4173 4207 4187
rect 4113 4153 4127 4167
rect 4213 4153 4227 4167
rect 4273 4173 4287 4187
rect 4273 4153 4287 4167
rect 4233 4133 4247 4147
rect 4113 3993 4127 4007
rect 4093 3933 4107 3947
rect 4213 3913 4227 3927
rect 4033 3873 4047 3887
rect 3993 3753 4007 3767
rect 3953 3693 3967 3707
rect 4013 3713 4027 3727
rect 4173 3753 4187 3767
rect 4053 3733 4067 3747
rect 4093 3733 4107 3747
rect 4073 3713 4087 3727
rect 4113 3693 4127 3707
rect 4033 3613 4047 3627
rect 3993 3573 4007 3587
rect 4013 3573 4027 3587
rect 3973 3533 3987 3547
rect 3993 3533 4007 3547
rect 4013 3493 4027 3507
rect 3873 3473 3887 3487
rect 3913 3473 3927 3487
rect 3893 3393 3907 3407
rect 3753 3213 3767 3227
rect 3793 3173 3807 3187
rect 3773 3153 3787 3167
rect 3753 3113 3767 3127
rect 3853 3233 3867 3247
rect 3873 3213 3887 3227
rect 3873 3193 3887 3207
rect 3833 3173 3847 3187
rect 3893 3173 3907 3187
rect 3813 3153 3827 3167
rect 3833 3153 3847 3167
rect 3793 3013 3807 3027
rect 3773 2873 3787 2887
rect 3753 2813 3767 2827
rect 3733 2793 3747 2807
rect 3893 3033 3907 3047
rect 3833 3013 3847 3027
rect 3873 2913 3887 2927
rect 3833 2833 3847 2847
rect 3813 2813 3827 2827
rect 3733 2773 3747 2787
rect 3773 2773 3787 2787
rect 3813 2773 3827 2787
rect 3773 2753 3787 2767
rect 3833 2733 3847 2747
rect 3753 2693 3767 2707
rect 3793 2693 3807 2707
rect 3773 2633 3787 2647
rect 3733 2553 3747 2567
rect 3733 2253 3747 2267
rect 3713 2153 3727 2167
rect 3693 2133 3707 2147
rect 3713 2093 3727 2107
rect 3733 2093 3747 2107
rect 3693 2053 3707 2067
rect 3733 1993 3747 2007
rect 3733 1953 3747 1967
rect 3713 1833 3727 1847
rect 3673 1813 3687 1827
rect 3693 1813 3707 1827
rect 3673 1773 3687 1787
rect 3653 1753 3667 1767
rect 3633 1733 3647 1747
rect 3613 1713 3627 1727
rect 3613 1693 3627 1707
rect 3593 1573 3607 1587
rect 3533 1553 3547 1567
rect 3413 1473 3427 1487
rect 3513 1473 3527 1487
rect 3453 1353 3467 1367
rect 3533 1353 3547 1367
rect 3393 1313 3407 1327
rect 3293 1253 3307 1267
rect 3333 1253 3347 1267
rect 3273 1213 3287 1227
rect 3133 853 3147 867
rect 3093 833 3107 847
rect 3113 813 3127 827
rect 3113 693 3127 707
rect 3153 673 3167 687
rect 3173 673 3187 687
rect 3133 653 3147 667
rect 3153 633 3167 647
rect 3253 1153 3267 1167
rect 3253 1093 3267 1107
rect 3413 1273 3427 1287
rect 3393 1253 3407 1267
rect 3433 1253 3447 1267
rect 3453 1253 3467 1267
rect 3333 1173 3347 1187
rect 3373 1173 3387 1187
rect 3353 1133 3367 1147
rect 3273 1033 3287 1047
rect 3233 833 3247 847
rect 3253 713 3267 727
rect 3193 633 3207 647
rect 3253 633 3267 647
rect 3113 593 3127 607
rect 3053 573 3067 587
rect 2913 393 2927 407
rect 3033 393 3047 407
rect 2893 373 2907 387
rect 2853 333 2867 347
rect 2933 373 2947 387
rect 2973 373 2987 387
rect 3033 373 3047 387
rect 3073 373 3087 387
rect 2913 353 2927 367
rect 2953 353 2967 367
rect 2993 353 3007 367
rect 3433 1173 3447 1187
rect 3313 993 3327 1007
rect 3293 893 3307 907
rect 3553 1333 3567 1347
rect 3533 1253 3547 1267
rect 3473 1173 3487 1187
rect 3513 1173 3527 1187
rect 3513 1153 3527 1167
rect 3573 1293 3587 1307
rect 3573 1253 3587 1267
rect 3493 1093 3507 1107
rect 3533 1093 3547 1107
rect 3553 1093 3567 1107
rect 3633 1673 3647 1687
rect 3633 1593 3647 1607
rect 3673 1633 3687 1647
rect 3793 2573 3807 2587
rect 3853 2553 3867 2567
rect 3993 3313 4007 3327
rect 3933 3213 3947 3227
rect 3933 3113 3947 3127
rect 3933 3093 3947 3107
rect 3953 2993 3967 3007
rect 3933 2933 3947 2947
rect 3913 2913 3927 2927
rect 3893 2893 3907 2907
rect 3913 2793 3927 2807
rect 3873 2513 3887 2527
rect 4013 3193 4027 3207
rect 4013 3113 4027 3127
rect 4073 3533 4087 3547
rect 4273 3913 4287 3927
rect 4253 3753 4267 3767
rect 4233 3733 4247 3747
rect 4253 3713 4267 3727
rect 4393 4493 4407 4507
rect 4373 4453 4387 4467
rect 4553 4953 4567 4967
rect 4553 4713 4567 4727
rect 4433 4453 4447 4467
rect 4493 4473 4507 4487
rect 4533 4473 4547 4487
rect 4453 4433 4467 4447
rect 4513 4453 4527 4467
rect 4673 4953 4687 4967
rect 4773 4973 4787 4987
rect 4813 5013 4827 5027
rect 4813 4973 4827 4987
rect 4793 4953 4807 4967
rect 4733 4933 4747 4947
rect 4753 4933 4767 4947
rect 4733 4913 4747 4927
rect 4733 4893 4747 4907
rect 4693 4753 4707 4767
rect 4673 4713 4687 4727
rect 4693 4673 4707 4687
rect 4613 4653 4627 4667
rect 4873 5073 4887 5087
rect 4893 5053 4907 5067
rect 4973 5393 4987 5407
rect 4933 5373 4947 5387
rect 4933 5233 4947 5247
rect 4973 5233 4987 5247
rect 4913 5033 4927 5047
rect 4953 5173 4967 5187
rect 5033 5393 5047 5407
rect 5033 5253 5047 5267
rect 4993 5173 5007 5187
rect 4953 5113 4967 5127
rect 5013 5113 5027 5127
rect 4993 5093 5007 5107
rect 4973 5053 4987 5067
rect 4953 5013 4967 5027
rect 4833 4953 4847 4967
rect 4853 4953 4867 4967
rect 4933 4953 4947 4967
rect 5073 5533 5087 5547
rect 5253 5673 5267 5687
rect 5173 5633 5187 5647
rect 5153 5553 5167 5567
rect 5133 5533 5147 5547
rect 5233 5633 5247 5647
rect 5213 5533 5227 5547
rect 5173 5473 5187 5487
rect 5193 5473 5207 5487
rect 5073 5433 5087 5447
rect 5113 5433 5127 5447
rect 5113 5413 5127 5427
rect 5093 5393 5107 5407
rect 5153 5393 5167 5407
rect 5253 5433 5267 5447
rect 5213 5413 5227 5427
rect 5233 5393 5247 5407
rect 5133 5373 5147 5387
rect 5113 5333 5127 5347
rect 5253 5373 5267 5387
rect 5233 5353 5247 5367
rect 5153 5313 5167 5327
rect 5073 5253 5087 5267
rect 5113 5253 5127 5267
rect 5053 5173 5067 5187
rect 4993 4953 5007 4967
rect 4913 4933 4927 4947
rect 4933 4933 4947 4947
rect 4973 4933 4987 4947
rect 4893 4913 4907 4927
rect 4793 4853 4807 4867
rect 4753 4673 4767 4687
rect 4833 4673 4847 4687
rect 4873 4673 4887 4687
rect 4733 4613 4747 4627
rect 4673 4593 4687 4607
rect 4573 4513 4587 4527
rect 4573 4493 4587 4507
rect 4613 4473 4627 4487
rect 4633 4473 4647 4487
rect 4473 4413 4487 4427
rect 4453 4313 4467 4327
rect 4413 4273 4427 4287
rect 4373 4233 4387 4247
rect 4333 4173 4347 4187
rect 4353 4093 4367 4107
rect 4313 3973 4327 3987
rect 4333 3733 4347 3747
rect 4273 3693 4287 3707
rect 4233 3673 4247 3687
rect 4313 3673 4327 3687
rect 4213 3653 4227 3667
rect 4193 3533 4207 3547
rect 4273 3653 4287 3667
rect 4253 3593 4267 3607
rect 4113 3493 4127 3507
rect 4253 3513 4267 3527
rect 4173 3493 4187 3507
rect 4213 3493 4227 3507
rect 4333 3593 4347 3607
rect 4313 3573 4327 3587
rect 4053 3253 4067 3267
rect 4113 3253 4127 3267
rect 4053 3133 4067 3147
rect 4033 3073 4047 3087
rect 4053 3073 4067 3087
rect 3993 2893 4007 2907
rect 4033 2893 4047 2907
rect 3993 2873 4007 2887
rect 3953 2813 3967 2827
rect 3793 2353 3807 2367
rect 3833 2353 3847 2367
rect 3893 2353 3907 2367
rect 3793 2333 3807 2347
rect 3793 2253 3807 2267
rect 3813 2233 3827 2247
rect 3773 2073 3787 2087
rect 3873 2313 3887 2327
rect 4013 2753 4027 2767
rect 3993 2713 4007 2727
rect 3993 2613 4007 2627
rect 3953 2593 3967 2607
rect 3953 2553 3967 2567
rect 3973 2553 3987 2567
rect 3973 2513 3987 2527
rect 3953 2353 3967 2367
rect 3913 2293 3927 2307
rect 3913 2273 3927 2287
rect 3933 2253 3947 2267
rect 3853 2213 3867 2227
rect 3893 2213 3907 2227
rect 3853 2173 3867 2187
rect 3913 2173 3927 2187
rect 3833 2133 3847 2147
rect 4013 2573 4027 2587
rect 4173 3213 4187 3227
rect 4233 3213 4247 3227
rect 4293 3233 4307 3247
rect 4173 3073 4187 3087
rect 4073 3053 4087 3067
rect 4113 3053 4127 3067
rect 4093 3033 4107 3047
rect 4133 3033 4147 3047
rect 4073 2733 4087 2747
rect 4053 2613 4067 2627
rect 4033 2553 4047 2567
rect 3993 2313 4007 2327
rect 4013 2273 4027 2287
rect 3993 2233 4007 2247
rect 3973 2133 3987 2147
rect 3973 2113 3987 2127
rect 3953 2073 3967 2087
rect 3793 2033 3807 2047
rect 3853 2013 3867 2027
rect 3833 1933 3847 1947
rect 3793 1853 3807 1867
rect 3753 1813 3767 1827
rect 3733 1793 3747 1807
rect 3753 1793 3767 1807
rect 3933 2033 3947 2047
rect 3953 2033 3967 2047
rect 3953 1973 3967 1987
rect 3893 1953 3907 1967
rect 3913 1893 3927 1907
rect 3893 1813 3907 1827
rect 3853 1793 3867 1807
rect 3733 1753 3747 1767
rect 3833 1753 3847 1767
rect 4093 2513 4107 2527
rect 4153 3013 4167 3027
rect 4273 3193 4287 3207
rect 4333 3533 4347 3547
rect 4413 4213 4427 4227
rect 4373 4073 4387 4087
rect 4433 4173 4447 4187
rect 4553 4433 4567 4447
rect 4533 4393 4547 4407
rect 4593 4413 4607 4427
rect 4653 4453 4667 4467
rect 4633 4433 4647 4447
rect 4553 4373 4567 4387
rect 4593 4373 4607 4387
rect 4613 4373 4627 4387
rect 4493 4333 4507 4347
rect 4553 4293 4567 4307
rect 4513 4193 4527 4207
rect 4493 4173 4507 4187
rect 4433 4033 4447 4047
rect 4433 3973 4447 3987
rect 4413 3693 4427 3707
rect 4453 3953 4467 3967
rect 4473 3953 4487 3967
rect 4413 3633 4427 3647
rect 4393 3553 4407 3567
rect 4353 3233 4367 3247
rect 4353 3173 4367 3187
rect 4313 3113 4327 3127
rect 4173 2953 4187 2967
rect 4153 2713 4167 2727
rect 4133 2673 4147 2687
rect 4073 2433 4087 2447
rect 4113 2433 4127 2447
rect 4053 2393 4067 2407
rect 4053 2273 4067 2287
rect 4013 2113 4027 2127
rect 4033 2113 4047 2127
rect 3993 2093 4007 2107
rect 4213 2873 4227 2887
rect 4333 3073 4347 3087
rect 4313 3013 4327 3027
rect 4353 2953 4367 2967
rect 4453 3513 4467 3527
rect 4433 3353 4447 3367
rect 4413 3253 4427 3267
rect 4413 3233 4427 3247
rect 4393 3193 4407 3207
rect 4453 3233 4467 3247
rect 4473 3233 4487 3247
rect 4273 2773 4287 2787
rect 4253 2733 4267 2747
rect 4193 2693 4207 2707
rect 4233 2653 4247 2667
rect 4173 2573 4187 2587
rect 4133 2293 4147 2307
rect 4113 2273 4127 2287
rect 4253 2573 4267 2587
rect 4213 2513 4227 2527
rect 4193 2453 4207 2467
rect 4253 2413 4267 2427
rect 4253 2293 4267 2307
rect 4213 2273 4227 2287
rect 4093 2253 4107 2267
rect 4133 2253 4147 2267
rect 4193 2233 4207 2247
rect 4113 2193 4127 2207
rect 4093 2133 4107 2147
rect 4033 2053 4047 2067
rect 4013 2033 4027 2047
rect 3973 1813 3987 1827
rect 3953 1793 3967 1807
rect 3973 1773 3987 1787
rect 3893 1753 3907 1767
rect 3933 1753 3947 1767
rect 3953 1753 3967 1767
rect 3753 1733 3767 1747
rect 3793 1733 3807 1747
rect 3873 1733 3887 1747
rect 3693 1613 3707 1627
rect 3673 1413 3687 1427
rect 3693 1333 3707 1347
rect 3673 1313 3687 1327
rect 3633 1273 3647 1287
rect 3653 1273 3667 1287
rect 3613 1153 3627 1167
rect 3633 1133 3647 1147
rect 3613 1093 3627 1107
rect 3453 1033 3467 1047
rect 3513 1033 3527 1047
rect 3573 1033 3587 1047
rect 3493 993 3507 1007
rect 3413 873 3427 887
rect 3353 853 3367 867
rect 3293 833 3307 847
rect 3313 833 3327 847
rect 3293 653 3307 667
rect 3413 813 3427 827
rect 3353 793 3367 807
rect 3373 793 3387 807
rect 3333 753 3347 767
rect 3333 653 3347 667
rect 3453 773 3467 787
rect 3393 753 3407 767
rect 3493 673 3507 687
rect 3433 653 3447 667
rect 3473 653 3487 667
rect 3493 653 3507 667
rect 3293 613 3307 627
rect 3333 613 3347 627
rect 3393 613 3407 627
rect 3273 533 3287 547
rect 3293 393 3307 407
rect 3093 353 3107 367
rect 3153 353 3167 367
rect 2993 333 3007 347
rect 3153 313 3167 327
rect 3053 273 3067 287
rect 3233 333 3247 347
rect 3313 373 3327 387
rect 3413 453 3427 467
rect 3373 373 3387 387
rect 3253 313 3267 327
rect 3313 313 3327 327
rect 3233 273 3247 287
rect 2813 193 2827 207
rect 2733 173 2747 187
rect 2773 173 2787 187
rect 2393 153 2407 167
rect 2453 153 2467 167
rect 2493 153 2507 167
rect 2473 133 2487 147
rect 2693 153 2707 167
rect 2893 193 2907 207
rect 2933 193 2947 207
rect 3193 193 3207 207
rect 2853 153 2867 167
rect 2133 113 2147 127
rect 2373 113 2387 127
rect 2513 113 2527 127
rect 2893 133 2907 147
rect 3293 193 3307 207
rect 3053 173 3067 187
rect 3233 173 3247 187
rect 2993 133 3007 147
rect 3253 153 3267 167
rect 3373 173 3387 187
rect 3473 613 3487 627
rect 3493 593 3507 607
rect 3433 153 3447 167
rect 3773 1713 3787 1727
rect 3873 1693 3887 1707
rect 3853 1613 3867 1627
rect 3833 1593 3847 1607
rect 3893 1593 3907 1607
rect 3913 1573 3927 1587
rect 3793 1333 3807 1347
rect 3853 1333 3867 1347
rect 3773 1293 3787 1307
rect 3813 1313 3827 1327
rect 3953 1353 3967 1367
rect 3913 1313 3927 1327
rect 3753 1253 3767 1267
rect 3793 1253 3807 1267
rect 3693 1233 3707 1247
rect 3713 1233 3727 1247
rect 3673 1133 3687 1147
rect 3653 1113 3667 1127
rect 3653 1093 3667 1107
rect 3673 1093 3687 1107
rect 3653 1053 3667 1067
rect 3593 993 3607 1007
rect 3533 913 3547 927
rect 3633 893 3647 907
rect 3553 853 3567 867
rect 3593 853 3607 867
rect 3633 853 3647 867
rect 3753 1213 3767 1227
rect 3793 1113 3807 1127
rect 3753 1093 3767 1107
rect 3733 1053 3747 1067
rect 3773 1053 3787 1067
rect 3713 1033 3727 1047
rect 3753 1033 3767 1047
rect 3693 913 3707 927
rect 3573 833 3587 847
rect 3533 813 3547 827
rect 3533 793 3547 807
rect 3573 673 3587 687
rect 3573 633 3587 647
rect 3513 473 3527 487
rect 3533 433 3547 447
rect 3613 833 3627 847
rect 3633 673 3647 687
rect 3613 633 3627 647
rect 3693 833 3707 847
rect 3673 813 3687 827
rect 3653 653 3667 667
rect 3733 813 3747 827
rect 3793 873 3807 887
rect 3833 1293 3847 1307
rect 3893 1293 3907 1307
rect 3873 1233 3887 1247
rect 3933 1253 3947 1267
rect 3973 1313 3987 1327
rect 3953 1213 3967 1227
rect 4053 2033 4067 2047
rect 4033 2013 4047 2027
rect 4033 1993 4047 2007
rect 4013 1973 4027 1987
rect 4013 1773 4027 1787
rect 4073 1993 4087 2007
rect 4073 1773 4087 1787
rect 4053 1753 4067 1767
rect 4033 1713 4047 1727
rect 4153 2113 4167 2127
rect 4213 2213 4227 2227
rect 4193 2073 4207 2087
rect 4173 2053 4187 2067
rect 4233 2053 4247 2067
rect 4213 2033 4227 2047
rect 4133 1853 4147 1867
rect 4093 1733 4107 1747
rect 4033 1693 4047 1707
rect 4073 1693 4087 1707
rect 4093 1693 4107 1707
rect 4073 1673 4087 1687
rect 4013 1573 4027 1587
rect 4033 1573 4047 1587
rect 4193 1813 4207 1827
rect 4173 1793 4187 1807
rect 4133 1653 4147 1667
rect 4193 1653 4207 1667
rect 4153 1633 4167 1647
rect 4113 1613 4127 1627
rect 4113 1593 4127 1607
rect 4133 1573 4147 1587
rect 4233 1853 4247 1867
rect 4313 2733 4327 2747
rect 4333 2573 4347 2587
rect 4313 2533 4327 2547
rect 4433 3033 4447 3047
rect 4413 2853 4427 2867
rect 4473 3053 4487 3067
rect 4573 4173 4587 4187
rect 4633 4253 4647 4267
rect 4713 4453 4727 4467
rect 4693 4433 4707 4447
rect 4693 4413 4707 4427
rect 4733 4413 4747 4427
rect 4673 4333 4687 4347
rect 4813 4653 4827 4667
rect 4773 4633 4787 4647
rect 4993 4913 5007 4927
rect 4973 4873 4987 4887
rect 4953 4733 4967 4747
rect 4953 4693 4967 4707
rect 4893 4653 4907 4667
rect 4933 4653 4947 4667
rect 4853 4613 4867 4627
rect 4873 4613 4887 4627
rect 4853 4573 4867 4587
rect 4773 4453 4787 4467
rect 4813 4453 4827 4467
rect 4793 4433 4807 4447
rect 4773 4413 4787 4427
rect 4773 4353 4787 4367
rect 4833 4353 4847 4367
rect 4753 4293 4767 4307
rect 4673 4273 4687 4287
rect 4693 4273 4707 4287
rect 4533 4133 4547 4147
rect 4533 4073 4547 4087
rect 4553 4013 4567 4027
rect 4593 3993 4607 4007
rect 4673 4213 4687 4227
rect 4673 4173 4687 4187
rect 4633 4153 4647 4167
rect 4713 4253 4727 4267
rect 4733 4213 4747 4227
rect 4713 4173 4727 4187
rect 4753 4153 4767 4167
rect 4653 4013 4667 4027
rect 4613 3973 4627 3987
rect 4553 3953 4567 3967
rect 4573 3953 4587 3967
rect 4533 3853 4547 3867
rect 4513 3813 4527 3827
rect 4633 3873 4647 3887
rect 4753 4073 4767 4087
rect 4733 3993 4747 4007
rect 4673 3953 4687 3967
rect 4673 3893 4687 3907
rect 4633 3813 4647 3827
rect 4553 3793 4567 3807
rect 4593 3733 4607 3747
rect 4513 3553 4527 3567
rect 4613 3553 4627 3567
rect 4533 3533 4547 3547
rect 4613 3533 4627 3547
rect 4513 3513 4527 3527
rect 4513 3493 4527 3507
rect 4493 2913 4507 2927
rect 4453 2813 4467 2827
rect 4373 2733 4387 2747
rect 4393 2713 4407 2727
rect 4433 2673 4447 2687
rect 4393 2593 4407 2607
rect 4373 2573 4387 2587
rect 4433 2573 4447 2587
rect 4313 2513 4327 2527
rect 4353 2513 4367 2527
rect 4273 2273 4287 2287
rect 4273 2253 4287 2267
rect 4293 2233 4307 2247
rect 4293 2153 4307 2167
rect 4293 2133 4307 2147
rect 4273 2033 4287 2047
rect 4333 2413 4347 2427
rect 4353 2373 4367 2387
rect 4413 2313 4427 2327
rect 4353 2253 4367 2267
rect 4333 2193 4347 2207
rect 4333 2173 4347 2187
rect 4373 2173 4387 2187
rect 4433 2133 4447 2147
rect 4413 2073 4427 2087
rect 4433 2073 4447 2087
rect 4313 1993 4327 2007
rect 4393 2053 4407 2067
rect 4393 1993 4407 2007
rect 4353 1973 4367 1987
rect 4353 1873 4367 1887
rect 4293 1833 4307 1847
rect 4313 1813 4327 1827
rect 4273 1793 4287 1807
rect 4253 1713 4267 1727
rect 4233 1673 4247 1687
rect 4133 1553 4147 1567
rect 4213 1553 4227 1567
rect 4093 1433 4107 1447
rect 4013 1293 4027 1307
rect 4073 1313 4087 1327
rect 4033 1273 4047 1287
rect 3993 1213 4007 1227
rect 3913 1193 3927 1207
rect 3973 1193 3987 1207
rect 3873 1133 3887 1147
rect 3893 1133 3907 1147
rect 3833 1113 3847 1127
rect 3853 1093 3867 1107
rect 3993 1133 4007 1147
rect 4033 1133 4047 1147
rect 3853 1073 3867 1087
rect 3773 853 3787 867
rect 3813 853 3827 867
rect 3793 833 3807 847
rect 3713 773 3727 787
rect 3693 633 3707 647
rect 3633 593 3647 607
rect 3673 593 3687 607
rect 3613 553 3627 567
rect 3593 393 3607 407
rect 3533 193 3547 207
rect 3273 133 3287 147
rect 3413 133 3427 147
rect 3133 113 3147 127
rect 3393 113 3407 127
rect 373 93 387 107
rect 513 93 527 107
rect 853 93 867 107
rect 2053 93 2067 107
rect 3493 153 3507 167
rect 3473 113 3487 127
rect 3593 293 3607 307
rect 3553 113 3567 127
rect 3733 613 3747 627
rect 3713 593 3727 607
rect 3753 573 3767 587
rect 3853 813 3867 827
rect 3853 753 3867 767
rect 4093 1113 4107 1127
rect 4013 1073 4027 1087
rect 3973 1033 3987 1047
rect 4073 1033 4087 1047
rect 4233 1433 4247 1447
rect 4193 1313 4207 1327
rect 4293 1733 4307 1747
rect 4273 1633 4287 1647
rect 4273 1593 4287 1607
rect 4253 1393 4267 1407
rect 4253 1293 4267 1307
rect 4233 1133 4247 1147
rect 4173 1113 4187 1127
rect 4213 1093 4227 1107
rect 3973 913 3987 927
rect 4133 913 4147 927
rect 3953 793 3967 807
rect 3893 613 3907 627
rect 3793 593 3807 607
rect 3833 593 3847 607
rect 3773 553 3787 567
rect 3873 573 3887 587
rect 3873 473 3887 487
rect 3793 453 3807 467
rect 3693 433 3707 447
rect 3833 433 3847 447
rect 3793 413 3807 427
rect 3753 353 3767 367
rect 3733 333 3747 347
rect 3693 313 3707 327
rect 3773 293 3787 307
rect 3833 333 3847 347
rect 3873 313 3887 327
rect 3913 573 3927 587
rect 4093 873 4107 887
rect 4133 833 4147 847
rect 4033 793 4047 807
rect 3993 773 4007 787
rect 3973 493 3987 507
rect 3933 393 3947 407
rect 3973 393 3987 407
rect 3953 373 3967 387
rect 3933 353 3947 367
rect 3893 273 3907 287
rect 3933 273 3947 287
rect 3813 253 3827 267
rect 3673 173 3687 187
rect 3713 173 3727 187
rect 3913 173 3927 187
rect 3613 113 3627 127
rect 3733 133 3747 147
rect 3673 113 3687 127
rect 3853 153 3867 167
rect 4113 773 4127 787
rect 4053 653 4067 667
rect 4193 1073 4207 1087
rect 4193 1033 4207 1047
rect 4313 1593 4327 1607
rect 4413 1833 4427 1847
rect 4573 3513 4587 3527
rect 4653 3793 4667 3807
rect 4553 3493 4567 3507
rect 4593 3493 4607 3507
rect 4633 3493 4647 3507
rect 4693 3773 4707 3787
rect 5033 4993 5047 5007
rect 5093 5153 5107 5167
rect 5073 5013 5087 5027
rect 5053 4973 5067 4987
rect 5113 4973 5127 4987
rect 5053 4913 5067 4927
rect 5073 4893 5087 4907
rect 5013 4693 5027 4707
rect 5053 4693 5067 4707
rect 4993 4593 5007 4607
rect 4973 4553 4987 4567
rect 4953 4493 4967 4507
rect 4853 4333 4867 4347
rect 4913 4453 4927 4467
rect 4953 4373 4967 4387
rect 4893 4293 4907 4307
rect 4893 4253 4907 4267
rect 4933 4253 4947 4267
rect 4813 4213 4827 4227
rect 4813 4193 4827 4207
rect 4793 4133 4807 4147
rect 4773 4033 4787 4047
rect 4773 4013 4787 4027
rect 4793 4013 4807 4027
rect 4713 3713 4727 3727
rect 4873 4173 4887 4187
rect 4833 4153 4847 4167
rect 4853 4113 4867 4127
rect 4813 3853 4827 3867
rect 4833 3853 4847 3867
rect 4793 3773 4807 3787
rect 4813 3773 4827 3787
rect 4853 3773 4867 3787
rect 5033 4613 5047 4627
rect 5013 4473 5027 4487
rect 5033 4453 5047 4467
rect 5053 4433 5067 4447
rect 5033 4413 5047 4427
rect 5013 4393 5027 4407
rect 5013 4333 5027 4347
rect 5033 4333 5047 4347
rect 4993 4293 5007 4307
rect 4973 4253 4987 4267
rect 4953 4213 4967 4227
rect 4993 4213 5007 4227
rect 4973 4173 4987 4187
rect 4993 4053 5007 4067
rect 5113 4913 5127 4927
rect 5093 4833 5107 4847
rect 5193 5153 5207 5167
rect 5253 5333 5267 5347
rect 5333 6033 5347 6047
rect 5393 6073 5407 6087
rect 5493 6133 5507 6147
rect 5473 6073 5487 6087
rect 5413 6033 5427 6047
rect 6013 6133 6027 6147
rect 5753 6113 5767 6127
rect 5673 6093 5687 6107
rect 5633 6073 5647 6087
rect 5673 6073 5687 6087
rect 5693 6073 5707 6087
rect 5633 6033 5647 6047
rect 5513 5993 5527 6007
rect 5413 5973 5427 5987
rect 5373 5953 5387 5967
rect 5533 5953 5547 5967
rect 5413 5933 5427 5947
rect 5353 5913 5367 5927
rect 5393 5913 5407 5927
rect 5333 5893 5347 5907
rect 5473 5913 5487 5927
rect 5493 5913 5507 5927
rect 5433 5873 5447 5887
rect 5453 5793 5467 5807
rect 5373 5733 5387 5747
rect 5373 5713 5387 5727
rect 5313 5633 5327 5647
rect 5293 5613 5307 5627
rect 5333 5593 5347 5607
rect 5333 5573 5347 5587
rect 5413 5693 5427 5707
rect 5453 5633 5467 5647
rect 5393 5613 5407 5627
rect 5393 5573 5407 5587
rect 5313 5553 5327 5567
rect 5373 5553 5387 5567
rect 5293 5493 5307 5507
rect 5333 5493 5347 5507
rect 5313 5433 5327 5447
rect 5373 5433 5387 5447
rect 5353 5413 5367 5427
rect 5293 5393 5307 5407
rect 5473 5593 5487 5607
rect 5433 5553 5447 5567
rect 5473 5433 5487 5447
rect 5433 5413 5447 5427
rect 5413 5373 5427 5387
rect 5393 5353 5407 5367
rect 5333 5253 5347 5267
rect 5353 5253 5367 5267
rect 5253 5213 5267 5227
rect 5273 5213 5287 5227
rect 5173 5133 5187 5147
rect 5233 5133 5247 5147
rect 5213 5113 5227 5127
rect 5153 5073 5167 5087
rect 5233 5053 5247 5067
rect 5173 4993 5187 5007
rect 5213 4993 5227 5007
rect 5153 4953 5167 4967
rect 5133 4793 5147 4807
rect 5233 4933 5247 4947
rect 5213 4893 5227 4907
rect 5313 5193 5327 5207
rect 5273 5173 5287 5187
rect 5393 5213 5407 5227
rect 5473 5233 5487 5247
rect 5453 5193 5467 5207
rect 5333 5173 5347 5187
rect 5393 5173 5407 5187
rect 5413 5173 5427 5187
rect 5293 5153 5307 5167
rect 5293 5113 5307 5127
rect 5293 4953 5307 4967
rect 5313 4913 5327 4927
rect 5273 4873 5287 4887
rect 5253 4813 5267 4827
rect 5273 4793 5287 4807
rect 5113 4593 5127 4607
rect 5093 4553 5107 4567
rect 5193 4773 5207 4787
rect 5233 4773 5247 4787
rect 5153 4753 5167 4767
rect 5253 4733 5267 4747
rect 5193 4693 5207 4707
rect 5233 4693 5247 4707
rect 5193 4673 5207 4687
rect 5173 4653 5187 4667
rect 5313 4773 5327 4787
rect 5273 4693 5287 4707
rect 5293 4673 5307 4687
rect 5213 4653 5227 4667
rect 5273 4653 5287 4667
rect 5273 4613 5287 4627
rect 5233 4593 5247 4607
rect 5253 4553 5267 4567
rect 5193 4533 5207 4547
rect 5133 4493 5147 4507
rect 5153 4493 5167 4507
rect 5073 4273 5087 4287
rect 5033 4253 5047 4267
rect 5073 4253 5087 4267
rect 5073 4213 5087 4227
rect 5073 4173 5087 4187
rect 5053 4153 5067 4167
rect 5053 4133 5067 4147
rect 5213 4493 5227 4507
rect 5173 4453 5187 4467
rect 5193 4453 5207 4467
rect 5113 4413 5127 4427
rect 5313 4513 5327 4527
rect 5353 5153 5367 5167
rect 5373 5133 5387 5147
rect 5413 5133 5427 5147
rect 5773 6093 5787 6107
rect 5713 6053 5727 6067
rect 5733 6053 5747 6067
rect 5913 6113 5927 6127
rect 5973 6113 5987 6127
rect 6033 6113 6047 6127
rect 6073 6113 6087 6127
rect 6193 6113 6207 6127
rect 6013 6093 6027 6107
rect 5953 6073 5967 6087
rect 5793 6033 5807 6047
rect 5853 6033 5867 6047
rect 5873 6033 5887 6047
rect 6273 6113 6287 6127
rect 6313 6113 6327 6127
rect 6353 6113 6367 6127
rect 6393 6113 6407 6127
rect 6053 6073 6067 6087
rect 6053 6053 6067 6067
rect 5673 6013 5687 6027
rect 5813 6013 5827 6027
rect 6033 6013 6047 6027
rect 5653 5933 5667 5947
rect 5513 5873 5527 5887
rect 5653 5913 5667 5927
rect 5773 5993 5787 6007
rect 5693 5973 5707 5987
rect 5733 5913 5747 5927
rect 5713 5893 5727 5907
rect 5753 5893 5767 5907
rect 5613 5873 5627 5887
rect 5673 5873 5687 5887
rect 5693 5873 5707 5887
rect 5713 5873 5727 5887
rect 5573 5833 5587 5847
rect 5613 5833 5627 5847
rect 5573 5633 5587 5647
rect 5593 5613 5607 5627
rect 5553 5593 5567 5607
rect 5513 5573 5527 5587
rect 5533 5573 5547 5587
rect 5553 5473 5567 5487
rect 5513 5433 5527 5447
rect 5513 5393 5527 5407
rect 5473 5173 5487 5187
rect 5493 5173 5507 5187
rect 5393 5013 5407 5027
rect 5353 4953 5367 4967
rect 5413 4993 5427 5007
rect 5373 4933 5387 4947
rect 5393 4913 5407 4927
rect 5573 5413 5587 5427
rect 5593 5413 5607 5427
rect 5673 5653 5687 5667
rect 5793 5973 5807 5987
rect 5873 5993 5887 6007
rect 5833 5973 5847 5987
rect 5813 5933 5827 5947
rect 5853 5933 5867 5947
rect 5813 5873 5827 5887
rect 5773 5793 5787 5807
rect 5713 5753 5727 5767
rect 5653 5633 5667 5647
rect 5693 5633 5707 5647
rect 5793 5673 5807 5687
rect 5813 5673 5827 5687
rect 5753 5653 5767 5667
rect 5733 5633 5747 5647
rect 5753 5573 5767 5587
rect 5773 5573 5787 5587
rect 5733 5553 5747 5567
rect 5733 5533 5747 5547
rect 5653 5453 5667 5467
rect 5693 5453 5707 5467
rect 5713 5453 5727 5467
rect 5633 5433 5647 5447
rect 5633 5393 5647 5407
rect 5673 5433 5687 5447
rect 5693 5413 5707 5427
rect 5653 5353 5667 5367
rect 5533 5213 5547 5227
rect 5573 5213 5587 5227
rect 5493 5113 5507 5127
rect 5513 5113 5527 5127
rect 5593 5133 5607 5147
rect 5613 5113 5627 5127
rect 5553 5053 5567 5067
rect 5493 4933 5507 4947
rect 5613 4953 5627 4967
rect 5433 4753 5447 4767
rect 5453 4733 5467 4747
rect 5433 4713 5447 4727
rect 5593 4913 5607 4927
rect 5553 4873 5567 4887
rect 5513 4853 5527 4867
rect 5473 4713 5487 4727
rect 5453 4693 5467 4707
rect 5473 4693 5487 4707
rect 5413 4673 5427 4687
rect 5493 4673 5507 4687
rect 5713 5373 5727 5387
rect 5733 5373 5747 5387
rect 5713 5313 5727 5327
rect 6033 5953 6047 5967
rect 6073 5953 6087 5967
rect 5933 5933 5947 5947
rect 6033 5913 6047 5927
rect 5913 5893 5927 5907
rect 5993 5893 6007 5907
rect 5953 5873 5967 5887
rect 6013 5873 6027 5887
rect 5873 5653 5887 5667
rect 5833 5633 5847 5647
rect 5873 5633 5887 5647
rect 5933 5633 5947 5647
rect 5853 5613 5867 5627
rect 5833 5573 5847 5587
rect 5813 5433 5827 5447
rect 5873 5553 5887 5567
rect 6053 5833 6067 5847
rect 5993 5713 6007 5727
rect 5973 5633 5987 5647
rect 5953 5593 5967 5607
rect 5913 5573 5927 5587
rect 5793 5413 5807 5427
rect 5773 5393 5787 5407
rect 5813 5373 5827 5387
rect 5693 5233 5707 5247
rect 5733 5233 5747 5247
rect 5753 5233 5767 5247
rect 5673 5153 5687 5167
rect 5693 5113 5707 5127
rect 5653 5033 5667 5047
rect 5733 5053 5747 5067
rect 5893 5413 5907 5427
rect 5853 5353 5867 5367
rect 5893 5313 5907 5327
rect 5813 5233 5827 5247
rect 5833 5213 5847 5227
rect 5773 5193 5787 5207
rect 5793 5173 5807 5187
rect 5773 5153 5787 5167
rect 5793 5133 5807 5147
rect 5813 5113 5827 5127
rect 5793 5053 5807 5067
rect 5713 4993 5727 5007
rect 5753 4993 5767 5007
rect 5653 4933 5667 4947
rect 5713 4953 5727 4967
rect 5753 4953 5767 4967
rect 5853 4993 5867 5007
rect 5833 4933 5847 4947
rect 5873 4933 5887 4947
rect 5713 4893 5727 4907
rect 5653 4853 5667 4867
rect 5673 4853 5687 4867
rect 5633 4733 5647 4747
rect 5593 4693 5607 4707
rect 5633 4693 5647 4707
rect 5553 4673 5567 4687
rect 5433 4653 5447 4667
rect 5533 4653 5547 4667
rect 5293 4493 5307 4507
rect 5333 4493 5347 4507
rect 5393 4493 5407 4507
rect 5273 4473 5287 4487
rect 5153 4293 5167 4307
rect 5113 4233 5127 4247
rect 5253 4433 5267 4447
rect 5313 4473 5327 4487
rect 5313 4433 5327 4447
rect 5333 4433 5347 4447
rect 5293 4393 5307 4407
rect 5293 4333 5307 4347
rect 5253 4313 5267 4327
rect 5153 4213 5167 4227
rect 5193 4213 5207 4227
rect 5253 4233 5267 4247
rect 5233 4213 5247 4227
rect 5153 4193 5167 4207
rect 5173 4193 5187 4207
rect 5213 4193 5227 4207
rect 5133 4173 5147 4187
rect 5093 4093 5107 4107
rect 5073 4053 5087 4067
rect 4953 4033 4967 4047
rect 4993 4033 5007 4047
rect 5013 4033 5027 4047
rect 4933 4013 4947 4027
rect 4973 4013 4987 4027
rect 5213 4153 5227 4167
rect 5293 4193 5307 4207
rect 5273 4153 5287 4167
rect 5313 4153 5327 4167
rect 5213 4093 5227 4107
rect 5233 4093 5247 4107
rect 5113 4053 5127 4067
rect 4993 3953 5007 3967
rect 4933 3933 4947 3947
rect 5013 3933 5027 3947
rect 5053 3913 5067 3927
rect 4893 3753 4907 3767
rect 4993 3853 5007 3867
rect 4973 3793 4987 3807
rect 4973 3753 4987 3767
rect 4993 3753 5007 3767
rect 5053 3753 5067 3767
rect 4873 3733 4887 3747
rect 4933 3733 4947 3747
rect 4953 3733 4967 3747
rect 4773 3633 4787 3647
rect 4893 3713 4907 3727
rect 5033 3713 5047 3727
rect 4873 3673 4887 3687
rect 4893 3653 4907 3667
rect 4833 3613 4847 3627
rect 4753 3533 4767 3547
rect 4713 3513 4727 3527
rect 4613 3473 4627 3487
rect 4653 3473 4667 3487
rect 4553 3273 4567 3287
rect 4593 3253 4607 3267
rect 4713 3273 4727 3287
rect 4633 3253 4647 3267
rect 4613 3233 4627 3247
rect 4653 3233 4667 3247
rect 4593 3173 4607 3187
rect 4573 3073 4587 3087
rect 4533 2913 4547 2927
rect 4513 2653 4527 2667
rect 4473 2573 4487 2587
rect 4493 2533 4507 2547
rect 4493 2473 4507 2487
rect 4513 2173 4527 2187
rect 4513 2153 4527 2167
rect 4493 2093 4507 2107
rect 4493 2053 4507 2067
rect 4513 2033 4527 2047
rect 4453 1853 4467 1867
rect 4473 1793 4487 1807
rect 4513 1793 4527 1807
rect 4493 1753 4507 1767
rect 4413 1733 4427 1747
rect 4353 1693 4367 1707
rect 4453 1653 4467 1667
rect 4353 1633 4367 1647
rect 4353 1593 4367 1607
rect 4333 1573 4347 1587
rect 4313 1333 4327 1347
rect 4313 1293 4327 1307
rect 4553 2733 4567 2747
rect 4833 3513 4847 3527
rect 4793 3293 4807 3307
rect 4773 3273 4787 3287
rect 4733 3253 4747 3267
rect 4733 3213 4747 3227
rect 4713 3193 4727 3207
rect 4693 3073 4707 3087
rect 4953 3693 4967 3707
rect 4973 3673 4987 3687
rect 4953 3633 4967 3647
rect 4913 3573 4927 3587
rect 4913 3553 4927 3567
rect 4993 3593 5007 3607
rect 4973 3513 4987 3527
rect 4913 3253 4927 3267
rect 4813 3213 4827 3227
rect 4893 3213 4907 3227
rect 4753 3173 4767 3187
rect 4773 3173 4787 3187
rect 4913 3173 4927 3187
rect 4733 3113 4747 3127
rect 4653 3053 4667 3067
rect 4713 3053 4727 3067
rect 4673 3033 4687 3047
rect 4693 2833 4707 2847
rect 4673 2733 4687 2747
rect 4633 2713 4647 2727
rect 4633 2693 4647 2707
rect 4653 2573 4667 2587
rect 4633 2553 4647 2567
rect 4673 2553 4687 2567
rect 4613 2433 4627 2447
rect 4653 2433 4667 2447
rect 4553 2313 4567 2327
rect 4573 2313 4587 2327
rect 4633 2313 4647 2327
rect 4553 2233 4567 2247
rect 4593 2273 4607 2287
rect 4573 2153 4587 2167
rect 4613 2093 4627 2107
rect 4633 2093 4647 2107
rect 4593 1833 4607 1847
rect 4573 1793 4587 1807
rect 4593 1773 4607 1787
rect 4553 1653 4567 1667
rect 4533 1613 4547 1627
rect 4513 1593 4527 1607
rect 4393 1553 4407 1567
rect 4433 1553 4447 1567
rect 4473 1553 4487 1567
rect 4513 1553 4527 1567
rect 4533 1553 4547 1567
rect 4433 1393 4447 1407
rect 4373 1293 4387 1307
rect 4373 1133 4387 1147
rect 4333 1113 4347 1127
rect 4393 1093 4407 1107
rect 4313 1033 4327 1047
rect 4293 933 4307 947
rect 4393 873 4407 887
rect 4293 833 4307 847
rect 4393 833 4407 847
rect 4213 813 4227 827
rect 4313 813 4327 827
rect 4353 813 4367 827
rect 4333 793 4347 807
rect 4373 793 4387 807
rect 4413 793 4427 807
rect 4293 653 4307 667
rect 4513 1353 4527 1367
rect 4473 1333 4487 1347
rect 4453 1313 4467 1327
rect 4493 1313 4507 1327
rect 4573 1573 4587 1587
rect 5033 3633 5047 3647
rect 5353 4253 5367 4267
rect 5353 4133 5367 4147
rect 5333 4073 5347 4087
rect 5193 4033 5207 4047
rect 5213 4033 5227 4047
rect 5313 4033 5327 4047
rect 5353 4033 5367 4047
rect 5133 3913 5147 3927
rect 5113 3833 5127 3847
rect 5173 3753 5187 3767
rect 5133 3733 5147 3747
rect 5093 3693 5107 3707
rect 5113 3613 5127 3627
rect 5053 3593 5067 3607
rect 5073 3593 5087 3607
rect 5053 3573 5067 3587
rect 5093 3573 5107 3587
rect 5033 3553 5047 3567
rect 5013 3513 5027 3527
rect 5013 3333 5027 3347
rect 5033 3273 5047 3287
rect 4953 3193 4967 3207
rect 5033 3173 5047 3187
rect 4953 3073 4967 3087
rect 4853 3013 4867 3027
rect 4933 3033 4947 3047
rect 4973 3033 4987 3047
rect 4993 3013 5007 3027
rect 4793 2873 4807 2887
rect 4833 2873 4847 2887
rect 4753 2793 4767 2807
rect 4733 2633 4747 2647
rect 4733 2593 4747 2607
rect 4853 2833 4867 2847
rect 4893 2773 4907 2787
rect 5153 3673 5167 3687
rect 5293 4013 5307 4027
rect 5233 3973 5247 3987
rect 5253 3953 5267 3967
rect 5213 3853 5227 3867
rect 5273 3833 5287 3847
rect 5253 3753 5267 3767
rect 5213 3733 5227 3747
rect 5233 3713 5247 3727
rect 5253 3693 5267 3707
rect 5253 3653 5267 3667
rect 5253 3573 5267 3587
rect 5173 3553 5187 3567
rect 5193 3553 5207 3567
rect 5173 3513 5187 3527
rect 5153 3493 5167 3507
rect 5213 3493 5227 3507
rect 5153 3473 5167 3487
rect 5073 3453 5087 3467
rect 5193 3413 5207 3427
rect 5133 3333 5147 3347
rect 5093 3253 5107 3267
rect 5133 3253 5147 3267
rect 5193 3213 5207 3227
rect 5193 3193 5207 3207
rect 5533 4633 5547 4647
rect 5513 4553 5527 4567
rect 5473 4513 5487 4527
rect 5413 4473 5427 4487
rect 5433 4473 5447 4487
rect 5393 4433 5407 4447
rect 5493 4453 5507 4467
rect 5453 4433 5467 4447
rect 5453 4413 5467 4427
rect 5433 4373 5447 4387
rect 5413 4273 5427 4287
rect 5393 4233 5407 4247
rect 5473 4213 5487 4227
rect 5433 4193 5447 4207
rect 5373 4013 5387 4027
rect 5413 4173 5427 4187
rect 5513 4173 5527 4187
rect 5493 4073 5507 4087
rect 5473 4053 5487 4067
rect 5413 4033 5427 4047
rect 5453 4033 5467 4047
rect 5433 4013 5447 4027
rect 5573 4613 5587 4627
rect 5553 4553 5567 4567
rect 5613 4673 5627 4687
rect 5753 4913 5767 4927
rect 5793 4913 5807 4927
rect 5813 4913 5827 4927
rect 5713 4733 5727 4747
rect 5733 4733 5747 4747
rect 5673 4653 5687 4667
rect 5733 4653 5747 4667
rect 5813 4873 5827 4887
rect 5793 4853 5807 4867
rect 5833 4853 5847 4867
rect 5853 4813 5867 4827
rect 5753 4633 5767 4647
rect 5773 4633 5787 4647
rect 5833 4653 5847 4667
rect 5653 4613 5667 4627
rect 5813 4613 5827 4627
rect 5693 4533 5707 4547
rect 5653 4493 5667 4507
rect 5613 4473 5627 4487
rect 5713 4513 5727 4527
rect 5813 4513 5827 4527
rect 5753 4493 5767 4507
rect 5793 4493 5807 4507
rect 5553 4433 5567 4447
rect 5573 4433 5587 4447
rect 5613 4433 5627 4447
rect 5593 4393 5607 4407
rect 5553 4213 5567 4227
rect 5553 4153 5567 4167
rect 5713 4473 5727 4487
rect 5673 4453 5687 4467
rect 5753 4453 5767 4467
rect 5933 5473 5947 5487
rect 6133 6093 6147 6107
rect 6233 6093 6247 6107
rect 6333 6093 6347 6107
rect 6293 6073 6307 6087
rect 6453 6113 6467 6127
rect 6513 6113 6527 6127
rect 6433 6073 6447 6087
rect 6493 6073 6507 6087
rect 6353 6053 6367 6067
rect 6413 6053 6427 6067
rect 6573 6113 6587 6127
rect 6633 6113 6647 6127
rect 6593 6093 6607 6107
rect 6613 6093 6627 6107
rect 6653 6093 6667 6107
rect 6553 6053 6567 6067
rect 6513 6033 6527 6047
rect 6533 6033 6547 6047
rect 6293 6013 6307 6027
rect 6513 5973 6527 5987
rect 6133 5953 6147 5967
rect 6093 5933 6107 5947
rect 6233 5933 6247 5947
rect 6373 5933 6387 5947
rect 6413 5933 6427 5947
rect 6153 5913 6167 5927
rect 6333 5913 6347 5927
rect 6133 5873 6147 5887
rect 6173 5873 6187 5887
rect 6233 5893 6247 5907
rect 6253 5893 6267 5907
rect 6273 5873 6287 5887
rect 6193 5813 6207 5827
rect 6133 5733 6147 5747
rect 6073 5673 6087 5687
rect 6013 5653 6027 5667
rect 6053 5633 6067 5647
rect 6093 5633 6107 5647
rect 6233 5793 6247 5807
rect 6213 5673 6227 5687
rect 6193 5653 6207 5667
rect 6353 5893 6367 5907
rect 6373 5853 6387 5867
rect 6333 5733 6347 5747
rect 6313 5713 6327 5727
rect 6233 5653 6247 5667
rect 6393 5813 6407 5827
rect 6733 6073 6747 6087
rect 6773 6113 6787 6127
rect 6873 6133 6887 6147
rect 6913 6133 6927 6147
rect 6853 6073 6867 6087
rect 6753 6033 6767 6047
rect 6813 6033 6827 6047
rect 6893 6113 6907 6127
rect 6993 6113 7007 6127
rect 7093 6133 7107 6147
rect 7153 6113 7167 6127
rect 7053 6093 7067 6107
rect 7013 6073 7027 6087
rect 6673 6013 6687 6027
rect 6873 6013 6887 6027
rect 6613 5973 6627 5987
rect 6533 5913 6547 5927
rect 6653 5913 6667 5927
rect 6533 5893 6547 5907
rect 6593 5893 6607 5907
rect 6553 5853 6567 5867
rect 6493 5833 6507 5847
rect 6473 5713 6487 5727
rect 6373 5673 6387 5687
rect 5993 5593 6007 5607
rect 6033 5593 6047 5607
rect 6233 5613 6247 5627
rect 6173 5533 6187 5547
rect 6413 5653 6427 5667
rect 6453 5653 6467 5667
rect 6593 5833 6607 5847
rect 6573 5773 6587 5787
rect 6433 5633 6447 5647
rect 6513 5633 6527 5647
rect 6633 5713 6647 5727
rect 6653 5673 6667 5687
rect 6593 5613 6607 5627
rect 7273 6113 7287 6127
rect 7273 6073 7287 6087
rect 7253 6033 7267 6047
rect 7173 5993 7187 6007
rect 7233 5993 7247 6007
rect 7013 5973 7027 5987
rect 7053 5973 7067 5987
rect 7133 5973 7147 5987
rect 7213 5973 7227 5987
rect 6713 5893 6727 5907
rect 6753 5893 6767 5907
rect 6973 5893 6987 5907
rect 7033 5953 7047 5967
rect 7033 5893 7047 5907
rect 7073 5953 7087 5967
rect 7113 5933 7127 5947
rect 7153 5933 7167 5947
rect 7133 5913 7147 5927
rect 7193 5913 7207 5927
rect 7093 5893 7107 5907
rect 6813 5873 6827 5887
rect 6773 5833 6787 5847
rect 6733 5793 6747 5807
rect 6693 5673 6707 5687
rect 6713 5673 6727 5687
rect 6673 5613 6687 5627
rect 6573 5593 6587 5607
rect 6613 5593 6627 5607
rect 6293 5573 6307 5587
rect 6253 5513 6267 5527
rect 6053 5473 6067 5487
rect 6073 5473 6087 5487
rect 6473 5453 6487 5467
rect 6553 5453 6567 5467
rect 5973 5413 5987 5427
rect 6033 5413 6047 5427
rect 5953 5393 5967 5407
rect 5913 5253 5927 5267
rect 6073 5393 6087 5407
rect 5953 5193 5967 5207
rect 5993 5193 6007 5207
rect 5913 5173 5927 5187
rect 6213 5413 6227 5427
rect 6233 5333 6247 5347
rect 6293 5333 6307 5347
rect 6193 5293 6207 5307
rect 6273 5293 6287 5307
rect 6373 5433 6387 5447
rect 6413 5433 6427 5447
rect 6433 5433 6447 5447
rect 6393 5273 6407 5287
rect 6293 5213 6307 5227
rect 6333 5213 6347 5227
rect 6193 5193 6207 5207
rect 6113 5173 6127 5187
rect 5953 5153 5967 5167
rect 5973 5133 5987 5147
rect 6073 5153 6087 5167
rect 6133 5153 6147 5167
rect 6173 5153 6187 5167
rect 6273 5173 6287 5187
rect 6333 5193 6347 5207
rect 6313 5173 6327 5187
rect 6233 5153 6247 5167
rect 6253 5153 6267 5167
rect 6293 5153 6307 5167
rect 5933 5113 5947 5127
rect 5953 5113 5967 5127
rect 6033 5113 6047 5127
rect 5913 4973 5927 4987
rect 6033 5093 6047 5107
rect 6093 5133 6107 5147
rect 6113 5133 6127 5147
rect 6153 5073 6167 5087
rect 6053 5033 6067 5047
rect 5993 4973 6007 4987
rect 5973 4933 5987 4947
rect 5933 4893 5947 4907
rect 5953 4813 5967 4827
rect 5893 4773 5907 4787
rect 5913 4773 5927 4787
rect 6013 4953 6027 4967
rect 6093 4953 6107 4967
rect 6133 4953 6147 4967
rect 6293 5113 6307 5127
rect 6213 4993 6227 5007
rect 6373 5153 6387 5167
rect 6393 5133 6407 5147
rect 6353 5113 6367 5127
rect 6513 5433 6527 5447
rect 6853 5653 6867 5667
rect 6733 5613 6747 5627
rect 6773 5613 6787 5627
rect 6693 5553 6707 5567
rect 6633 5433 6647 5447
rect 6673 5433 6687 5447
rect 6753 5433 6767 5447
rect 6833 5613 6847 5627
rect 6793 5593 6807 5607
rect 6993 5873 7007 5887
rect 7033 5833 7047 5847
rect 7113 5713 7127 5727
rect 7053 5693 7067 5707
rect 7013 5673 7027 5687
rect 7033 5673 7047 5687
rect 6953 5653 6967 5667
rect 6993 5653 7007 5667
rect 6933 5633 6947 5647
rect 6933 5593 6947 5607
rect 6913 5573 6927 5587
rect 6873 5473 6887 5487
rect 6853 5453 6867 5467
rect 6813 5433 6827 5447
rect 6553 5413 6567 5427
rect 6593 5413 6607 5427
rect 6533 5393 6547 5407
rect 6433 5193 6447 5207
rect 6513 5173 6527 5187
rect 6593 5393 6607 5407
rect 6613 5393 6627 5407
rect 6693 5393 6707 5407
rect 6733 5213 6747 5227
rect 6493 5153 6507 5167
rect 6473 5113 6487 5127
rect 6733 5173 6747 5187
rect 6793 5413 6807 5427
rect 6893 5433 6907 5447
rect 6913 5393 6927 5407
rect 6853 5213 6867 5227
rect 6573 5153 6587 5167
rect 6613 5153 6627 5167
rect 6493 5093 6507 5107
rect 6413 5053 6427 5067
rect 6493 5053 6507 5067
rect 6373 4993 6387 5007
rect 6413 4993 6427 5007
rect 6253 4973 6267 4987
rect 6313 4973 6327 4987
rect 6053 4933 6067 4947
rect 6033 4893 6047 4907
rect 5993 4713 6007 4727
rect 6193 4933 6207 4947
rect 6273 4933 6287 4947
rect 6153 4893 6167 4907
rect 6293 4733 6307 4747
rect 6033 4693 6047 4707
rect 6073 4693 6087 4707
rect 5933 4673 5947 4687
rect 5993 4673 6007 4687
rect 6013 4673 6027 4687
rect 6053 4673 6067 4687
rect 6033 4633 6047 4647
rect 6053 4613 6067 4627
rect 6173 4713 6187 4727
rect 6133 4673 6147 4687
rect 6153 4633 6167 4647
rect 6053 4593 6067 4607
rect 6093 4593 6107 4607
rect 5853 4513 5867 4527
rect 5833 4473 5847 4487
rect 5813 4453 5827 4467
rect 5853 4453 5867 4467
rect 5733 4413 5747 4427
rect 5633 4333 5647 4347
rect 5613 4313 5627 4327
rect 5693 4233 5707 4247
rect 5613 4173 5627 4187
rect 5633 4173 5647 4187
rect 5593 4153 5607 4167
rect 5573 4113 5587 4127
rect 5553 4053 5567 4067
rect 5433 3973 5447 3987
rect 5353 3953 5367 3967
rect 5393 3953 5407 3967
rect 5433 3953 5447 3967
rect 5333 3893 5347 3907
rect 5293 3813 5307 3827
rect 5393 3913 5407 3927
rect 5553 4013 5567 4027
rect 5533 3953 5547 3967
rect 5813 4433 5827 4447
rect 5833 4433 5847 4447
rect 5873 4433 5887 4447
rect 5833 4413 5847 4427
rect 5813 4393 5827 4407
rect 5793 4273 5807 4287
rect 5753 4193 5767 4207
rect 5653 4133 5667 4147
rect 5633 4053 5647 4067
rect 5673 4033 5687 4047
rect 5773 4173 5787 4187
rect 5953 4473 5967 4487
rect 5933 4453 5947 4467
rect 5973 4453 5987 4467
rect 5933 4433 5947 4447
rect 6013 4433 6027 4447
rect 5893 4393 5907 4407
rect 6233 4653 6247 4667
rect 6193 4553 6207 4567
rect 6213 4513 6227 4527
rect 6073 4493 6087 4507
rect 6193 4493 6207 4507
rect 6193 4473 6207 4487
rect 6353 4933 6367 4947
rect 6393 4933 6407 4947
rect 6453 4953 6467 4967
rect 6453 4933 6467 4947
rect 6353 4913 6367 4927
rect 6433 4913 6447 4927
rect 6413 4733 6427 4747
rect 6433 4733 6447 4747
rect 6333 4713 6347 4727
rect 6313 4693 6327 4707
rect 6273 4673 6287 4687
rect 6333 4673 6347 4687
rect 6373 4673 6387 4687
rect 6313 4653 6327 4667
rect 6353 4633 6367 4647
rect 6393 4633 6407 4647
rect 6273 4553 6287 4567
rect 6253 4493 6267 4507
rect 6253 4473 6267 4487
rect 6073 4453 6087 4467
rect 6113 4453 6127 4467
rect 6373 4533 6387 4547
rect 6313 4473 6327 4487
rect 6353 4473 6367 4487
rect 6233 4453 6247 4467
rect 6273 4453 6287 4467
rect 6333 4453 6347 4467
rect 6593 5133 6607 5147
rect 6613 5113 6627 5127
rect 6713 5113 6727 5127
rect 6673 5073 6687 5087
rect 6673 5053 6687 5067
rect 6633 5033 6647 5047
rect 6613 4973 6627 4987
rect 6553 4953 6567 4967
rect 6593 4953 6607 4967
rect 6553 4933 6567 4947
rect 6653 4913 6667 4927
rect 6573 4873 6587 4887
rect 6613 4873 6627 4887
rect 6533 4833 6547 4847
rect 6573 4833 6587 4847
rect 6493 4733 6507 4747
rect 6453 4713 6467 4727
rect 6473 4713 6487 4727
rect 6613 4753 6627 4767
rect 6493 4693 6507 4707
rect 6473 4673 6487 4687
rect 6453 4653 6467 4667
rect 6433 4573 6447 4587
rect 6513 4653 6527 4667
rect 6573 4693 6587 4707
rect 6593 4673 6607 4687
rect 6573 4653 6587 4667
rect 6593 4633 6607 4647
rect 6633 4633 6647 4647
rect 6553 4613 6567 4627
rect 6513 4573 6527 4587
rect 6493 4553 6507 4567
rect 6473 4533 6487 4547
rect 6473 4493 6487 4507
rect 6453 4473 6467 4487
rect 6453 4453 6467 4467
rect 6493 4473 6507 4487
rect 6093 4433 6107 4447
rect 6013 4273 6027 4287
rect 5873 4193 5887 4207
rect 5913 4193 5927 4207
rect 5733 4153 5747 4167
rect 5853 4053 5867 4067
rect 5793 4013 5807 4027
rect 5613 3993 5627 4007
rect 5713 3993 5727 4007
rect 5753 3993 5767 4007
rect 5673 3973 5687 3987
rect 5713 3973 5727 3987
rect 5593 3953 5607 3967
rect 5573 3933 5587 3947
rect 5493 3833 5507 3847
rect 5513 3833 5527 3847
rect 5553 3833 5567 3847
rect 5393 3813 5407 3827
rect 5473 3813 5487 3827
rect 5353 3753 5367 3767
rect 5293 3713 5307 3727
rect 5333 3713 5347 3727
rect 5313 3693 5327 3707
rect 5373 3693 5387 3707
rect 5433 3793 5447 3807
rect 5493 3733 5507 3747
rect 5513 3733 5527 3747
rect 5653 3953 5667 3967
rect 5693 3953 5707 3967
rect 5733 3953 5747 3967
rect 5633 3893 5647 3907
rect 5673 3933 5687 3947
rect 5653 3773 5667 3787
rect 5633 3753 5647 3767
rect 5773 3973 5787 3987
rect 5853 3993 5867 4007
rect 5893 4153 5907 4167
rect 5913 4093 5927 4107
rect 5933 4093 5947 4107
rect 5933 4073 5947 4087
rect 5913 4053 5927 4067
rect 6013 4193 6027 4207
rect 6053 4193 6067 4207
rect 5993 4153 6007 4167
rect 6033 4073 6047 4087
rect 5953 4013 5967 4027
rect 5833 3973 5847 3987
rect 5873 3973 5887 3987
rect 5813 3953 5827 3967
rect 5773 3913 5787 3927
rect 5753 3793 5767 3807
rect 5773 3773 5787 3787
rect 5473 3713 5487 3727
rect 5353 3673 5367 3687
rect 5293 3653 5307 3667
rect 5293 3573 5307 3587
rect 5353 3573 5367 3587
rect 5313 3513 5327 3527
rect 5453 3693 5467 3707
rect 5453 3673 5467 3687
rect 5433 3653 5447 3667
rect 5413 3533 5427 3547
rect 5413 3513 5427 3527
rect 5333 3493 5347 3507
rect 5393 3493 5407 3507
rect 5433 3493 5447 3507
rect 5273 3473 5287 3487
rect 5333 3473 5347 3487
rect 5393 3473 5407 3487
rect 5253 3433 5267 3447
rect 5273 3293 5287 3307
rect 5313 3273 5327 3287
rect 5273 3253 5287 3267
rect 5293 3233 5307 3247
rect 5413 3233 5427 3247
rect 5353 3193 5367 3207
rect 5533 3693 5547 3707
rect 5493 3633 5507 3647
rect 5533 3513 5547 3527
rect 5493 3473 5507 3487
rect 5473 3453 5487 3467
rect 5553 3473 5567 3487
rect 5513 3433 5527 3447
rect 5673 3733 5687 3747
rect 5733 3733 5747 3747
rect 5653 3713 5667 3727
rect 5753 3713 5767 3727
rect 5593 3613 5607 3627
rect 5833 3793 5847 3807
rect 5953 3993 5967 4007
rect 5893 3953 5907 3967
rect 5873 3893 5887 3907
rect 5893 3813 5907 3827
rect 5853 3753 5867 3767
rect 5833 3713 5847 3727
rect 6413 4433 6427 4447
rect 6473 4433 6487 4447
rect 6433 4413 6447 4427
rect 6173 4353 6187 4367
rect 6133 4273 6147 4287
rect 6133 4233 6147 4247
rect 6293 4273 6307 4287
rect 6173 4213 6187 4227
rect 6233 4213 6247 4227
rect 6373 4253 6387 4267
rect 6113 4173 6127 4187
rect 6193 4173 6207 4187
rect 6113 4133 6127 4147
rect 6153 4133 6167 4147
rect 6073 4113 6087 4127
rect 6133 4113 6147 4127
rect 6253 4113 6267 4127
rect 6093 4013 6107 4027
rect 6053 3973 6067 3987
rect 5973 3953 5987 3967
rect 5993 3953 6007 3967
rect 6013 3953 6027 3967
rect 6073 3953 6087 3967
rect 6233 4053 6247 4067
rect 6153 4013 6167 4027
rect 6173 3973 6187 3987
rect 6213 3973 6227 3987
rect 5973 3793 5987 3807
rect 5953 3773 5967 3787
rect 5913 3733 5927 3747
rect 5793 3693 5807 3707
rect 5813 3693 5827 3707
rect 6013 3813 6027 3827
rect 6113 3793 6127 3807
rect 6113 3753 6127 3767
rect 6053 3733 6067 3747
rect 5973 3713 5987 3727
rect 5993 3713 6007 3727
rect 6013 3713 6027 3727
rect 6153 3733 6167 3747
rect 6193 3733 6207 3747
rect 5653 3573 5667 3587
rect 5753 3553 5767 3567
rect 5713 3513 5727 3527
rect 5673 3493 5687 3507
rect 5973 3673 5987 3687
rect 5993 3673 6007 3687
rect 6033 3673 6047 3687
rect 5853 3553 5867 3567
rect 5773 3533 5787 3547
rect 5813 3533 5827 3547
rect 5813 3513 5827 3527
rect 5853 3513 5867 3527
rect 5753 3493 5767 3507
rect 5793 3493 5807 3507
rect 5833 3493 5847 3507
rect 5613 3473 5627 3487
rect 5693 3473 5707 3487
rect 5733 3473 5747 3487
rect 5913 3493 5927 3507
rect 6053 3533 6067 3547
rect 6013 3493 6027 3507
rect 6053 3493 6067 3507
rect 5893 3473 5907 3487
rect 5933 3473 5947 3487
rect 5993 3473 6007 3487
rect 5893 3453 5907 3467
rect 6033 3433 6047 3447
rect 5933 3413 5947 3427
rect 5813 3293 5827 3307
rect 5853 3293 5867 3307
rect 5573 3273 5587 3287
rect 5853 3273 5867 3287
rect 5873 3273 5887 3287
rect 6013 3273 6027 3287
rect 5453 3253 5467 3267
rect 5533 3253 5547 3267
rect 5633 3253 5647 3267
rect 5693 3253 5707 3267
rect 5473 3233 5487 3247
rect 5453 3193 5467 3207
rect 5713 3233 5727 3247
rect 5493 3213 5507 3227
rect 5433 3173 5447 3187
rect 5473 3173 5487 3187
rect 5573 3193 5587 3207
rect 5673 3213 5687 3227
rect 5553 3173 5567 3187
rect 5593 3173 5607 3187
rect 5513 3153 5527 3167
rect 5773 3253 5787 3267
rect 5813 3253 5827 3267
rect 5753 3113 5767 3127
rect 5213 3093 5227 3107
rect 5753 3093 5767 3107
rect 5333 3073 5347 3087
rect 5713 3073 5727 3087
rect 5193 3053 5207 3067
rect 5293 3033 5307 3047
rect 5073 3013 5087 3027
rect 5173 3013 5187 3027
rect 5093 2833 5107 2847
rect 5253 2793 5267 2807
rect 4933 2753 4947 2767
rect 4813 2733 4827 2747
rect 4833 2713 4847 2727
rect 4873 2713 4887 2727
rect 4773 2693 4787 2707
rect 4793 2633 4807 2647
rect 4773 2573 4787 2587
rect 4773 2553 4787 2567
rect 4693 2313 4707 2327
rect 4733 2313 4747 2327
rect 4693 2293 4707 2307
rect 4673 2073 4687 2087
rect 4653 1873 4667 1887
rect 4653 1813 4667 1827
rect 4693 1813 4707 1827
rect 4773 2093 4787 2107
rect 4673 1793 4687 1807
rect 4733 1793 4747 1807
rect 4673 1753 4687 1767
rect 4633 1713 4647 1727
rect 4773 1773 4787 1787
rect 4713 1693 4727 1707
rect 4753 1693 4767 1707
rect 4633 1673 4647 1687
rect 4613 1593 4627 1607
rect 4673 1593 4687 1607
rect 4593 1393 4607 1407
rect 4593 1373 4607 1387
rect 4653 1553 4667 1567
rect 4813 2593 4827 2607
rect 5033 2773 5047 2787
rect 5053 2773 5067 2787
rect 4973 2733 4987 2747
rect 4833 2553 4847 2567
rect 4873 2553 4887 2567
rect 4913 2553 4927 2567
rect 4813 2513 4827 2527
rect 4853 2513 4867 2527
rect 4813 2233 4827 2247
rect 4973 2533 4987 2547
rect 5173 2753 5187 2767
rect 5113 2733 5127 2747
rect 5093 2713 5107 2727
rect 5153 2713 5167 2727
rect 5193 2713 5207 2727
rect 5073 2593 5087 2607
rect 5033 2553 5047 2567
rect 5113 2573 5127 2587
rect 5173 2573 5187 2587
rect 5093 2553 5107 2567
rect 5053 2533 5067 2547
rect 4973 2493 4987 2507
rect 4913 2313 4927 2327
rect 5013 2473 5027 2487
rect 4953 2253 4967 2267
rect 4853 2033 4867 2047
rect 4813 1833 4827 1847
rect 4933 1953 4947 1967
rect 4913 1813 4927 1827
rect 4993 2213 5007 2227
rect 4993 2093 5007 2107
rect 5053 2293 5067 2307
rect 5093 2293 5107 2307
rect 5073 2273 5087 2287
rect 5033 2253 5047 2267
rect 5133 2553 5147 2567
rect 5313 2753 5327 2767
rect 5573 3033 5587 3047
rect 5473 3013 5487 3027
rect 5513 3013 5527 3027
rect 5593 3013 5607 3027
rect 5673 3013 5687 3027
rect 5633 2993 5647 3007
rect 5693 2973 5707 2987
rect 5553 2873 5567 2887
rect 5653 2873 5667 2887
rect 5473 2733 5487 2747
rect 5733 3053 5747 3067
rect 5733 3033 5747 3047
rect 5833 3233 5847 3247
rect 5953 3253 5967 3267
rect 5993 3253 6007 3267
rect 5933 3233 5947 3247
rect 5913 3153 5927 3167
rect 5853 3093 5867 3107
rect 5813 3053 5827 3067
rect 5893 3073 5907 3087
rect 5773 3013 5787 3027
rect 6173 3713 6187 3727
rect 6253 4013 6267 4027
rect 6333 4193 6347 4207
rect 6353 4173 6367 4187
rect 6433 4193 6447 4207
rect 6373 4153 6387 4167
rect 6453 4173 6467 4187
rect 6413 4133 6427 4147
rect 6453 4133 6467 4147
rect 6353 4073 6367 4087
rect 6313 4053 6327 4067
rect 6373 4053 6387 4067
rect 6353 4013 6367 4027
rect 6353 3993 6367 4007
rect 6293 3973 6307 3987
rect 6233 3953 6247 3967
rect 6273 3953 6287 3967
rect 6313 3953 6327 3967
rect 6393 3973 6407 3987
rect 6433 3973 6447 3987
rect 6493 4013 6507 4027
rect 6473 3973 6487 3987
rect 6553 4493 6567 4507
rect 6533 4453 6547 4467
rect 6573 4453 6587 4467
rect 6593 4273 6607 4287
rect 6533 4253 6547 4267
rect 6533 4173 6547 4187
rect 6713 5033 6727 5047
rect 6693 4933 6707 4947
rect 6853 5173 6867 5187
rect 6833 5113 6847 5127
rect 6873 5073 6887 5087
rect 6773 5053 6787 5067
rect 6753 4993 6767 5007
rect 6893 4993 6907 5007
rect 6753 4973 6767 4987
rect 6793 4973 6807 4987
rect 6893 4953 6907 4967
rect 6973 5573 6987 5587
rect 7173 5893 7187 5907
rect 7333 6113 7347 6127
rect 7373 6113 7387 6127
rect 7353 6033 7367 6047
rect 7393 5953 7407 5967
rect 7553 6153 7567 6167
rect 7653 6153 7667 6167
rect 7513 6133 7527 6147
rect 7433 6113 7447 6127
rect 7473 6113 7487 6127
rect 7593 6113 7607 6127
rect 7613 6113 7627 6127
rect 7633 6113 7647 6127
rect 7693 6133 7707 6147
rect 7513 6073 7527 6087
rect 7453 5993 7467 6007
rect 7673 6093 7687 6107
rect 7713 6113 7727 6127
rect 7813 6113 7827 6127
rect 7853 6113 7867 6127
rect 7613 6073 7627 6087
rect 7653 6073 7667 6087
rect 7693 6073 7707 6087
rect 7833 6073 7847 6087
rect 7573 6053 7587 6067
rect 7713 6053 7727 6067
rect 7533 5973 7547 5987
rect 7573 5973 7587 5987
rect 7833 5973 7847 5987
rect 7253 5913 7267 5927
rect 7293 5913 7307 5927
rect 7313 5913 7327 5927
rect 7373 5913 7387 5927
rect 7413 5913 7427 5927
rect 7453 5913 7467 5927
rect 7233 5853 7247 5867
rect 7273 5893 7287 5907
rect 7313 5893 7327 5907
rect 7353 5893 7367 5907
rect 7393 5893 7407 5907
rect 7413 5893 7427 5907
rect 7253 5833 7267 5847
rect 7133 5693 7147 5707
rect 7333 5693 7347 5707
rect 7433 5873 7447 5887
rect 7093 5653 7107 5667
rect 7153 5673 7167 5687
rect 7253 5673 7267 5687
rect 7413 5673 7427 5687
rect 7013 5633 7027 5647
rect 7053 5633 7067 5647
rect 6993 5493 7007 5507
rect 6953 5473 6967 5487
rect 6993 5453 7007 5467
rect 7113 5633 7127 5647
rect 7133 5613 7147 5627
rect 7073 5573 7087 5587
rect 7113 5493 7127 5507
rect 7013 5433 7027 5447
rect 7053 5433 7067 5447
rect 7033 5413 7047 5427
rect 7073 5413 7087 5427
rect 6973 5393 6987 5407
rect 7013 5393 7027 5407
rect 7093 5393 7107 5407
rect 6953 5233 6967 5247
rect 6993 5233 7007 5247
rect 6953 5213 6967 5227
rect 6953 5193 6967 5207
rect 7073 5193 7087 5207
rect 6993 5173 7007 5187
rect 7033 5173 7047 5187
rect 7013 5153 7027 5167
rect 6933 5133 6947 5147
rect 6973 5133 6987 5147
rect 7053 5113 7067 5127
rect 7193 5653 7207 5667
rect 7233 5653 7247 5667
rect 7213 5633 7227 5647
rect 7173 5613 7187 5627
rect 7293 5653 7307 5667
rect 7293 5633 7307 5647
rect 7253 5593 7267 5607
rect 7273 5593 7287 5607
rect 7333 5593 7347 5607
rect 7373 5653 7387 5667
rect 7373 5633 7387 5647
rect 7513 5893 7527 5907
rect 7673 5953 7687 5967
rect 7693 5953 7707 5967
rect 7593 5913 7607 5927
rect 7633 5913 7647 5927
rect 7873 5933 7887 5947
rect 7733 5913 7747 5927
rect 7793 5913 7807 5927
rect 7573 5873 7587 5887
rect 7553 5853 7567 5867
rect 7473 5713 7487 5727
rect 7453 5633 7467 5647
rect 7433 5613 7447 5627
rect 7393 5593 7407 5607
rect 7353 5573 7367 5587
rect 7293 5533 7307 5547
rect 7173 5493 7187 5507
rect 7253 5493 7267 5507
rect 7153 5453 7167 5467
rect 7193 5433 7207 5447
rect 7133 5373 7147 5387
rect 7113 5173 7127 5187
rect 7113 5133 7127 5147
rect 7273 5433 7287 5447
rect 7553 5673 7567 5687
rect 7573 5653 7587 5667
rect 7533 5633 7547 5647
rect 7493 5573 7507 5587
rect 7473 5493 7487 5507
rect 7313 5473 7327 5487
rect 7493 5473 7507 5487
rect 7313 5453 7327 5467
rect 7473 5453 7487 5467
rect 7353 5433 7367 5447
rect 7393 5433 7407 5447
rect 7293 5413 7307 5427
rect 7333 5413 7347 5427
rect 7433 5413 7447 5427
rect 7333 5393 7347 5407
rect 7353 5393 7367 5407
rect 7373 5393 7387 5407
rect 7273 5233 7287 5247
rect 7253 5213 7267 5227
rect 7153 5173 7167 5187
rect 7213 5173 7227 5187
rect 7253 5173 7267 5187
rect 7273 5153 7287 5167
rect 7233 5133 7247 5147
rect 7173 5113 7187 5127
rect 7133 5093 7147 5107
rect 7213 5093 7227 5107
rect 6933 4993 6947 5007
rect 7093 4993 7107 5007
rect 7113 4973 7127 4987
rect 7153 4973 7167 4987
rect 7073 4953 7087 4967
rect 7133 4953 7147 4967
rect 7273 5013 7287 5027
rect 7253 4973 7267 4987
rect 7193 4953 7207 4967
rect 6773 4933 6787 4947
rect 6873 4933 6887 4947
rect 6913 4933 6927 4947
rect 6973 4933 6987 4947
rect 7013 4933 7027 4947
rect 6853 4913 6867 4927
rect 6953 4913 6967 4927
rect 6893 4893 6907 4907
rect 6813 4853 6827 4867
rect 6733 4673 6747 4687
rect 6753 4653 6767 4667
rect 6913 4733 6927 4747
rect 7013 4873 7027 4887
rect 6853 4673 6867 4687
rect 6813 4653 6827 4667
rect 6933 4673 6947 4687
rect 6993 4673 7007 4687
rect 7093 4933 7107 4947
rect 7033 4853 7047 4867
rect 7173 4933 7187 4947
rect 7233 4873 7247 4887
rect 7133 4713 7147 4727
rect 7213 4713 7227 4727
rect 6953 4653 6967 4667
rect 7013 4653 7027 4667
rect 6873 4633 6887 4647
rect 6713 4613 6727 4627
rect 6773 4613 6787 4627
rect 6833 4613 6847 4627
rect 6693 4553 6707 4567
rect 6673 4533 6687 4547
rect 6753 4513 6767 4527
rect 6633 4453 6647 4467
rect 6693 4453 6707 4467
rect 7093 4693 7107 4707
rect 7073 4673 7087 4687
rect 7173 4673 7187 4687
rect 7093 4633 7107 4647
rect 7193 4633 7207 4647
rect 7033 4573 7047 4587
rect 7213 4533 7227 4547
rect 6813 4513 6827 4527
rect 6913 4513 6927 4527
rect 6793 4453 6807 4467
rect 6933 4493 6947 4507
rect 7053 4493 7067 4507
rect 7133 4493 7147 4507
rect 6913 4473 6927 4487
rect 6933 4453 6947 4467
rect 6953 4453 6967 4467
rect 6993 4453 7007 4467
rect 7073 4473 7087 4487
rect 7093 4473 7107 4487
rect 7173 4473 7187 4487
rect 7193 4473 7207 4487
rect 7073 4453 7087 4467
rect 7113 4453 7127 4467
rect 7153 4453 7167 4467
rect 6833 4433 6847 4447
rect 6893 4433 6907 4447
rect 6853 4413 6867 4427
rect 6653 4273 6667 4287
rect 6613 4213 6627 4227
rect 6713 4253 6727 4267
rect 6753 4233 6767 4247
rect 6833 4233 6847 4247
rect 6793 4213 6807 4227
rect 6793 4193 6807 4207
rect 6553 4133 6567 4147
rect 6613 4173 6627 4187
rect 6633 4173 6647 4187
rect 6673 4173 6687 4187
rect 6733 4153 6747 4167
rect 6713 4133 6727 4147
rect 6553 4113 6567 4127
rect 6573 4113 6587 4127
rect 6533 4013 6547 4027
rect 6513 3993 6527 4007
rect 6593 4093 6607 4107
rect 6673 4093 6687 4107
rect 6533 3973 6547 3987
rect 6553 3973 6567 3987
rect 6573 3973 6587 3987
rect 7033 4433 7047 4447
rect 6993 4413 7007 4427
rect 6973 4233 6987 4247
rect 6873 4193 6887 4207
rect 6893 4153 6907 4167
rect 6853 4133 6867 4147
rect 6773 4053 6787 4067
rect 6873 4033 6887 4047
rect 6793 4013 6807 4027
rect 6773 3993 6787 4007
rect 6653 3973 6667 3987
rect 6693 3973 6707 3987
rect 6473 3953 6487 3967
rect 6273 3813 6287 3827
rect 6233 3753 6247 3767
rect 6353 3773 6367 3787
rect 6253 3713 6267 3727
rect 6533 3753 6547 3767
rect 6613 3753 6627 3767
rect 6393 3713 6407 3727
rect 6533 3733 6547 3747
rect 6573 3733 6587 3747
rect 6213 3693 6227 3707
rect 6333 3693 6347 3707
rect 6113 3673 6127 3687
rect 6093 3573 6107 3587
rect 6473 3693 6487 3707
rect 6553 3713 6567 3727
rect 6593 3713 6607 3727
rect 6513 3573 6527 3587
rect 6333 3533 6347 3547
rect 6373 3533 6387 3547
rect 6133 3513 6147 3527
rect 6173 3513 6187 3527
rect 6253 3513 6267 3527
rect 6113 3493 6127 3507
rect 6153 3493 6167 3507
rect 6153 3453 6167 3467
rect 6073 3253 6087 3267
rect 6113 3253 6127 3267
rect 6073 3233 6087 3247
rect 6053 3213 6067 3227
rect 6213 3493 6227 3507
rect 6173 3253 6187 3267
rect 6153 3233 6167 3247
rect 6293 3493 6307 3507
rect 6313 3493 6327 3507
rect 6353 3513 6367 3527
rect 6253 3433 6267 3447
rect 6593 3693 6607 3707
rect 6613 3573 6627 3587
rect 6493 3533 6507 3547
rect 6533 3533 6547 3547
rect 6553 3533 6567 3547
rect 6393 3493 6407 3507
rect 6573 3513 6587 3527
rect 6673 3733 6687 3747
rect 6693 3713 6707 3727
rect 6653 3693 6667 3707
rect 6633 3533 6647 3547
rect 6613 3473 6627 3487
rect 6693 3673 6707 3687
rect 6733 3653 6747 3667
rect 6713 3493 6727 3507
rect 6693 3473 6707 3487
rect 6513 3453 6527 3467
rect 6653 3453 6667 3467
rect 6733 3453 6747 3467
rect 6753 3313 6767 3327
rect 6413 3293 6427 3307
rect 6473 3293 6487 3307
rect 6273 3273 6287 3287
rect 6553 3273 6567 3287
rect 6673 3273 6687 3287
rect 6253 3253 6267 3267
rect 6233 3233 6247 3247
rect 6253 3233 6267 3247
rect 6033 3113 6047 3127
rect 6213 3113 6227 3127
rect 5993 3053 6007 3067
rect 5833 3013 5847 3027
rect 5873 3013 5887 3027
rect 5973 3013 5987 3027
rect 6153 3073 6167 3087
rect 6193 3073 6207 3087
rect 6053 3033 6067 3047
rect 6093 3013 6107 3027
rect 6193 3053 6207 3067
rect 6173 3033 6187 3047
rect 6173 3013 6187 3027
rect 5933 2993 5947 3007
rect 6153 2993 6167 3007
rect 6273 3213 6287 3227
rect 6313 3213 6327 3227
rect 6433 3253 6447 3267
rect 6473 3253 6487 3267
rect 6813 3973 6827 3987
rect 6973 4193 6987 4207
rect 7053 4413 7067 4427
rect 7073 4393 7087 4407
rect 6993 4173 7007 4187
rect 7053 4193 7067 4207
rect 7113 4313 7127 4327
rect 7093 4233 7107 4247
rect 7073 4173 7087 4187
rect 7093 4173 7107 4187
rect 7193 4413 7207 4427
rect 7153 4253 7167 4267
rect 7153 4213 7167 4227
rect 7193 4213 7207 4227
rect 7133 4193 7147 4207
rect 7173 4173 7187 4187
rect 7193 4173 7207 4187
rect 7013 4153 7027 4167
rect 6953 4113 6967 4127
rect 6913 4033 6927 4047
rect 7113 4153 7127 4167
rect 7093 4053 7107 4067
rect 7033 4033 7047 4047
rect 7033 4013 7047 4027
rect 7053 3993 7067 4007
rect 7133 3993 7147 4007
rect 6913 3973 6927 3987
rect 6953 3973 6967 3987
rect 6993 3973 7007 3987
rect 7033 3973 7047 3987
rect 7113 3973 7127 3987
rect 6793 3733 6807 3747
rect 6933 3733 6947 3747
rect 6833 3713 6847 3727
rect 6853 3693 6867 3707
rect 6813 3673 6827 3687
rect 6953 3713 6967 3727
rect 7013 3713 7027 3727
rect 6933 3693 6947 3707
rect 6913 3653 6927 3667
rect 6933 3653 6947 3667
rect 6833 3573 6847 3587
rect 6853 3553 6867 3567
rect 6833 3533 6847 3547
rect 6813 3493 6827 3507
rect 6913 3513 6927 3527
rect 6993 3653 7007 3667
rect 7013 3573 7027 3587
rect 6953 3533 6967 3547
rect 6973 3533 6987 3547
rect 6993 3533 7007 3547
rect 6793 3313 6807 3327
rect 6933 3473 6947 3487
rect 7133 3713 7147 3727
rect 7233 4513 7247 4527
rect 7273 4833 7287 4847
rect 7273 4733 7287 4747
rect 7293 4713 7307 4727
rect 7313 4693 7327 4707
rect 7453 5393 7467 5407
rect 7413 5373 7427 5387
rect 7533 5533 7547 5547
rect 7513 5453 7527 5467
rect 7613 5893 7627 5907
rect 7653 5893 7667 5907
rect 7713 5893 7727 5907
rect 7773 5853 7787 5867
rect 7693 5653 7707 5667
rect 7853 5653 7867 5667
rect 7633 5633 7647 5647
rect 7733 5633 7747 5647
rect 7793 5633 7807 5647
rect 7613 5613 7627 5627
rect 7593 5473 7607 5487
rect 7613 5453 7627 5467
rect 7573 5433 7587 5447
rect 7533 5413 7547 5427
rect 7373 5213 7387 5227
rect 7413 5213 7427 5227
rect 7473 5213 7487 5227
rect 7453 5193 7467 5207
rect 7553 5193 7567 5207
rect 7373 5153 7387 5167
rect 7413 5153 7427 5167
rect 7393 5113 7407 5127
rect 7433 5093 7447 5107
rect 7413 5013 7427 5027
rect 7353 4973 7367 4987
rect 7393 4973 7407 4987
rect 7373 4953 7387 4967
rect 7373 4933 7387 4947
rect 7493 5173 7507 5187
rect 7533 5173 7547 5187
rect 7633 5413 7647 5427
rect 7633 5393 7647 5407
rect 7593 5233 7607 5247
rect 7473 5153 7487 5167
rect 7513 5133 7527 5147
rect 7493 5113 7507 5127
rect 7513 5113 7527 5127
rect 7453 4993 7467 5007
rect 7453 4973 7467 4987
rect 7413 4953 7427 4967
rect 7493 4953 7507 4967
rect 7433 4933 7447 4947
rect 7453 4933 7467 4947
rect 7393 4913 7407 4927
rect 7473 4913 7487 4927
rect 7493 4913 7507 4927
rect 7373 4873 7387 4887
rect 7353 4853 7367 4867
rect 7453 4853 7467 4867
rect 7393 4693 7407 4707
rect 7433 4693 7447 4707
rect 7333 4673 7347 4687
rect 7373 4673 7387 4687
rect 7373 4653 7387 4667
rect 7353 4633 7367 4647
rect 7313 4533 7327 4547
rect 7253 4493 7267 4507
rect 7233 4473 7247 4487
rect 7313 4473 7327 4487
rect 7253 4453 7267 4467
rect 7293 4453 7307 4467
rect 7373 4573 7387 4587
rect 7353 4453 7367 4467
rect 7413 4553 7427 4567
rect 7413 4533 7427 4547
rect 7433 4513 7447 4527
rect 7413 4493 7427 4507
rect 7313 4433 7327 4447
rect 7353 4433 7367 4447
rect 7373 4373 7387 4387
rect 7273 4353 7287 4367
rect 7253 4233 7267 4247
rect 7233 4153 7247 4167
rect 7213 4013 7227 4027
rect 7253 3993 7267 4007
rect 7233 3973 7247 3987
rect 7333 4253 7347 4267
rect 7293 4213 7307 4227
rect 7273 3973 7287 3987
rect 7193 3753 7207 3767
rect 7253 3753 7267 3767
rect 7213 3733 7227 3747
rect 7253 3733 7267 3747
rect 7273 3733 7287 3747
rect 7233 3713 7247 3727
rect 7193 3693 7207 3707
rect 7113 3673 7127 3687
rect 7153 3673 7167 3687
rect 7073 3553 7087 3567
rect 7113 3553 7127 3567
rect 7033 3493 7047 3507
rect 7213 3553 7227 3567
rect 7253 3533 7267 3547
rect 7373 4193 7387 4207
rect 7353 4133 7367 4147
rect 7333 4013 7347 4027
rect 7313 3973 7327 3987
rect 7353 3973 7367 3987
rect 7353 3753 7367 3767
rect 7313 3733 7327 3747
rect 7153 3513 7167 3527
rect 7293 3493 7307 3507
rect 7133 3473 7147 3487
rect 6793 3293 6807 3307
rect 6893 3293 6907 3307
rect 7053 3293 7067 3307
rect 6773 3273 6787 3287
rect 6413 3233 6427 3247
rect 6373 3093 6387 3107
rect 6233 3053 6247 3067
rect 6333 3033 6347 3047
rect 6273 2993 6287 3007
rect 6233 2973 6247 2987
rect 5893 2793 5907 2807
rect 5933 2793 5947 2807
rect 6113 2793 6127 2807
rect 5853 2753 5867 2767
rect 6033 2773 6047 2787
rect 6233 2773 6247 2787
rect 6393 3053 6407 3067
rect 6673 3253 6687 3267
rect 6753 3253 6767 3267
rect 6513 3213 6527 3227
rect 6533 3213 6547 3227
rect 6493 3073 6507 3087
rect 6613 3213 6627 3227
rect 6613 3193 6627 3207
rect 6713 3233 6727 3247
rect 6893 3273 6907 3287
rect 6833 3253 6847 3267
rect 6873 3253 6887 3267
rect 6693 3213 6707 3227
rect 6733 3213 6747 3227
rect 6653 3173 6667 3187
rect 6573 3153 6587 3167
rect 6853 3153 6867 3167
rect 6573 3093 6587 3107
rect 6693 3093 6707 3107
rect 6533 3033 6547 3047
rect 6413 3013 6427 3027
rect 6453 3013 6467 3027
rect 6513 3013 6527 3027
rect 6593 3013 6607 3027
rect 6673 3013 6687 3027
rect 6633 2993 6647 3007
rect 6713 3033 6727 3047
rect 7013 3253 7027 3267
rect 7053 3253 7067 3267
rect 6973 3233 6987 3247
rect 6993 3213 7007 3227
rect 6953 3193 6967 3207
rect 7013 3193 7027 3207
rect 7073 3233 7087 3247
rect 7073 3193 7087 3207
rect 7033 3173 7047 3187
rect 7073 3053 7087 3067
rect 6753 3013 6767 3027
rect 6593 2973 6607 2987
rect 6373 2813 6387 2827
rect 6293 2773 6307 2787
rect 6353 2773 6367 2787
rect 6033 2753 6047 2767
rect 6093 2753 6107 2767
rect 6113 2753 6127 2767
rect 5673 2733 5687 2747
rect 5713 2733 5727 2747
rect 5873 2733 5887 2747
rect 5913 2733 5927 2747
rect 5233 2553 5247 2567
rect 5233 2533 5247 2547
rect 5153 2513 5167 2527
rect 5193 2493 5207 2507
rect 5253 2513 5267 2527
rect 5293 2713 5307 2727
rect 5353 2713 5367 2727
rect 5313 2633 5327 2647
rect 5293 2553 5307 2567
rect 5293 2493 5307 2507
rect 5273 2473 5287 2487
rect 5353 2573 5367 2587
rect 5633 2713 5647 2727
rect 5773 2713 5787 2727
rect 5953 2713 5967 2727
rect 5553 2633 5567 2647
rect 5493 2613 5507 2627
rect 5433 2573 5447 2587
rect 5373 2533 5387 2547
rect 5453 2553 5467 2567
rect 5573 2613 5587 2627
rect 5753 2613 5767 2627
rect 5953 2613 5967 2627
rect 5533 2553 5547 2567
rect 5913 2593 5927 2607
rect 5873 2573 5887 2587
rect 5633 2553 5647 2567
rect 5473 2533 5487 2547
rect 5653 2533 5667 2547
rect 5693 2533 5707 2547
rect 5333 2513 5347 2527
rect 5213 2453 5227 2467
rect 5313 2453 5327 2467
rect 5833 2553 5847 2567
rect 5773 2533 5787 2547
rect 5853 2533 5867 2547
rect 6173 2733 6187 2747
rect 6273 2753 6287 2767
rect 6353 2753 6367 2767
rect 6493 2773 6507 2787
rect 6013 2713 6027 2727
rect 6013 2693 6027 2707
rect 6073 2693 6087 2707
rect 5973 2573 5987 2587
rect 5953 2553 5967 2567
rect 5913 2513 5927 2527
rect 5133 2333 5147 2347
rect 5273 2333 5287 2347
rect 5713 2333 5727 2347
rect 5233 2313 5247 2327
rect 5133 2293 5147 2307
rect 5553 2293 5567 2307
rect 5653 2293 5667 2307
rect 5693 2293 5707 2307
rect 5733 2293 5747 2307
rect 5153 2273 5167 2287
rect 5193 2273 5207 2287
rect 5253 2273 5267 2287
rect 5173 2233 5187 2247
rect 5393 2253 5407 2267
rect 5133 2213 5147 2227
rect 5213 2213 5227 2227
rect 5113 2113 5127 2127
rect 5173 2113 5187 2127
rect 5093 2053 5107 2067
rect 5013 1953 5027 1967
rect 4973 1813 4987 1827
rect 5013 1813 5027 1827
rect 5053 1813 5067 1827
rect 4813 1773 4827 1787
rect 4853 1753 4867 1767
rect 4813 1633 4827 1647
rect 4713 1573 4727 1587
rect 4753 1573 4767 1587
rect 4833 1613 4847 1627
rect 4773 1453 4787 1467
rect 4953 1793 4967 1807
rect 4993 1793 5007 1807
rect 5013 1733 5027 1747
rect 4973 1573 4987 1587
rect 4873 1553 4887 1567
rect 4853 1453 4867 1467
rect 4813 1373 4827 1387
rect 4653 1333 4667 1347
rect 4613 1313 4627 1327
rect 4633 1313 4647 1327
rect 4573 1293 4587 1307
rect 4613 1273 4627 1287
rect 4733 1353 4747 1367
rect 4693 1333 4707 1347
rect 4813 1333 4827 1347
rect 4713 1313 4727 1327
rect 4853 1313 4867 1327
rect 4673 1273 4687 1287
rect 4613 1253 4627 1267
rect 4653 1253 4667 1267
rect 4553 1133 4567 1147
rect 4933 1553 4947 1567
rect 5133 2073 5147 2087
rect 5433 2093 5447 2107
rect 5213 2073 5227 2087
rect 5153 2053 5167 2067
rect 5193 2053 5207 2067
rect 5273 2053 5287 2067
rect 5213 2033 5227 2047
rect 5153 1973 5167 1987
rect 5073 1573 5087 1587
rect 5113 1573 5127 1587
rect 5293 2033 5307 2047
rect 5273 2013 5287 2027
rect 5173 1773 5187 1787
rect 5213 1773 5227 1787
rect 5253 1773 5267 1787
rect 5193 1573 5207 1587
rect 5073 1533 5087 1547
rect 5073 1473 5087 1487
rect 4933 1353 4947 1367
rect 5093 1433 5107 1447
rect 5173 1553 5187 1567
rect 5373 2053 5387 2067
rect 5333 1993 5347 2007
rect 5453 2053 5467 2067
rect 5473 2033 5487 2047
rect 5573 2273 5587 2287
rect 5613 2273 5627 2287
rect 5593 2253 5607 2267
rect 5713 2253 5727 2267
rect 5813 2293 5827 2307
rect 5873 2293 5887 2307
rect 5793 2273 5807 2287
rect 5573 2233 5587 2247
rect 5613 2233 5627 2247
rect 5633 2233 5647 2247
rect 5433 2013 5447 2027
rect 5573 1973 5587 1987
rect 5293 1813 5307 1827
rect 5373 1813 5387 1827
rect 5273 1653 5287 1667
rect 5413 1813 5427 1827
rect 5513 1813 5527 1827
rect 5553 1813 5567 1827
rect 5353 1793 5367 1807
rect 5393 1793 5407 1807
rect 5373 1773 5387 1787
rect 5333 1753 5347 1767
rect 5313 1733 5327 1747
rect 5293 1633 5307 1647
rect 5433 1793 5447 1807
rect 5473 1793 5487 1807
rect 5453 1773 5467 1787
rect 5573 1793 5587 1807
rect 5533 1753 5547 1767
rect 5593 1713 5607 1727
rect 5593 1693 5607 1707
rect 5513 1633 5527 1647
rect 5313 1613 5327 1627
rect 5393 1613 5407 1627
rect 5413 1613 5427 1627
rect 5293 1573 5307 1587
rect 5253 1553 5267 1567
rect 5333 1553 5347 1567
rect 5433 1573 5447 1587
rect 5413 1553 5427 1567
rect 5333 1533 5347 1547
rect 5393 1533 5407 1547
rect 5453 1533 5467 1547
rect 5453 1493 5467 1507
rect 5293 1473 5307 1487
rect 5173 1373 5187 1387
rect 5213 1373 5227 1387
rect 5133 1353 5147 1367
rect 4893 1313 4907 1327
rect 4953 1313 4967 1327
rect 4953 1293 4967 1307
rect 5073 1333 5087 1347
rect 5113 1333 5127 1347
rect 5113 1313 5127 1327
rect 4833 1273 4847 1287
rect 4873 1273 4887 1287
rect 4753 1193 4767 1207
rect 4793 1193 4807 1207
rect 4513 1073 4527 1087
rect 4573 1073 4587 1087
rect 4553 993 4567 1007
rect 4453 853 4467 867
rect 4473 813 4487 827
rect 4433 733 4447 747
rect 4333 653 4347 667
rect 4433 653 4447 667
rect 4453 653 4467 667
rect 4673 1113 4687 1127
rect 4713 1113 4727 1127
rect 4593 833 4607 847
rect 4953 1113 4967 1127
rect 5093 1273 5107 1287
rect 5153 1333 5167 1347
rect 5193 1333 5207 1347
rect 5253 1333 5267 1347
rect 5313 1333 5327 1347
rect 5373 1333 5387 1347
rect 5173 1313 5187 1327
rect 5233 1313 5247 1327
rect 5233 1273 5247 1287
rect 5133 1193 5147 1207
rect 5353 1193 5367 1207
rect 4993 1113 5007 1127
rect 5053 1113 5067 1127
rect 4873 1093 4887 1107
rect 4973 1093 4987 1107
rect 5113 1073 5127 1087
rect 5113 1033 5127 1047
rect 4813 853 4827 867
rect 4873 853 4887 867
rect 5233 1113 5247 1127
rect 5413 1313 5427 1327
rect 5393 1293 5407 1307
rect 5433 1293 5447 1307
rect 5553 1573 5567 1587
rect 5713 2093 5727 2107
rect 5753 2073 5767 2087
rect 5633 2033 5647 2047
rect 5873 2253 5887 2267
rect 5793 2233 5807 2247
rect 6353 2653 6367 2667
rect 6193 2613 6207 2627
rect 6133 2593 6147 2607
rect 6093 2573 6107 2587
rect 6153 2573 6167 2587
rect 6053 2533 6067 2547
rect 6033 2513 6047 2527
rect 6313 2553 6327 2567
rect 6453 2573 6467 2587
rect 6093 2493 6107 2507
rect 6513 2753 6527 2767
rect 6573 2733 6587 2747
rect 6793 2793 6807 2807
rect 6613 2773 6627 2787
rect 6633 2753 6647 2767
rect 6593 2713 6607 2727
rect 6713 2773 6727 2787
rect 6753 2773 6767 2787
rect 6773 2753 6787 2767
rect 6673 2733 6687 2747
rect 6913 3033 6927 3047
rect 6893 3013 6907 3027
rect 6933 2993 6947 3007
rect 6913 2793 6927 2807
rect 6873 2753 6887 2767
rect 6853 2733 6867 2747
rect 6973 2973 6987 2987
rect 6993 2793 7007 2807
rect 6953 2753 6967 2767
rect 7173 3253 7187 3267
rect 7473 4693 7487 4707
rect 7473 4653 7487 4667
rect 7473 4573 7487 4587
rect 7533 5013 7547 5027
rect 7593 5153 7607 5167
rect 7573 5133 7587 5147
rect 7633 5113 7647 5127
rect 7613 5093 7627 5107
rect 7593 5013 7607 5027
rect 7553 4973 7567 4987
rect 7633 4973 7647 4987
rect 7533 4953 7547 4967
rect 7573 4933 7587 4947
rect 7613 4933 7627 4947
rect 7513 4873 7527 4887
rect 7513 4833 7527 4847
rect 7673 5613 7687 5627
rect 7693 5593 7707 5607
rect 7773 5593 7787 5607
rect 7753 5573 7767 5587
rect 7773 5573 7787 5587
rect 7753 5473 7767 5487
rect 7713 5433 7727 5447
rect 7793 5513 7807 5527
rect 7833 5513 7847 5527
rect 7773 5453 7787 5467
rect 7753 5413 7767 5427
rect 7833 5453 7847 5467
rect 7793 5433 7807 5447
rect 7873 5433 7887 5447
rect 7813 5413 7827 5427
rect 7853 5413 7867 5427
rect 7773 5393 7787 5407
rect 7713 5193 7727 5207
rect 7753 5173 7767 5187
rect 7773 5173 7787 5187
rect 7733 5133 7747 5147
rect 7913 5433 7927 5447
rect 7793 5133 7807 5147
rect 7773 5113 7787 5127
rect 7773 5093 7787 5107
rect 7693 5073 7707 5087
rect 7733 5073 7747 5087
rect 7673 4993 7687 5007
rect 7693 4973 7707 4987
rect 7713 4953 7727 4967
rect 7593 4873 7607 4887
rect 7553 4853 7567 4867
rect 7533 4733 7547 4747
rect 7633 4733 7647 4747
rect 7533 4713 7547 4727
rect 7593 4713 7607 4727
rect 7573 4693 7587 4707
rect 7853 5153 7867 5167
rect 7893 5153 7907 5167
rect 7813 5093 7827 5107
rect 7873 5133 7887 5147
rect 7913 5133 7927 5147
rect 7873 5113 7887 5127
rect 7853 5073 7867 5087
rect 7813 4973 7827 4987
rect 7833 4973 7847 4987
rect 7793 4933 7807 4947
rect 7833 4933 7847 4947
rect 7893 4993 7907 5007
rect 7753 4873 7767 4887
rect 7753 4753 7767 4767
rect 7733 4733 7747 4747
rect 7673 4713 7687 4727
rect 7673 4693 7687 4707
rect 7713 4693 7727 4707
rect 7773 4733 7787 4747
rect 7593 4673 7607 4687
rect 7633 4673 7647 4687
rect 7573 4653 7587 4667
rect 7613 4633 7627 4647
rect 7633 4573 7647 4587
rect 7593 4553 7607 4567
rect 7553 4533 7567 4547
rect 7513 4513 7527 4527
rect 7553 4513 7567 4527
rect 7573 4513 7587 4527
rect 7453 4473 7467 4487
rect 7513 4473 7527 4487
rect 7533 4473 7547 4487
rect 7453 4453 7467 4467
rect 7433 4413 7447 4427
rect 7433 4253 7447 4267
rect 7413 4213 7427 4227
rect 7473 4433 7487 4447
rect 7493 4413 7507 4427
rect 7553 4393 7567 4407
rect 7473 4313 7487 4327
rect 7473 4293 7487 4307
rect 7513 4253 7527 4267
rect 7473 4213 7487 4227
rect 7413 4193 7427 4207
rect 7453 4193 7467 4207
rect 7493 4193 7507 4207
rect 7433 4173 7447 4187
rect 7413 4113 7427 4127
rect 7473 4153 7487 4167
rect 7453 4113 7467 4127
rect 7453 3993 7467 4007
rect 7453 3953 7467 3967
rect 7413 3933 7427 3947
rect 7453 3913 7467 3927
rect 7493 3993 7507 4007
rect 7493 3953 7507 3967
rect 7553 4353 7567 4367
rect 7733 4673 7747 4687
rect 7693 4653 7707 4667
rect 7713 4653 7727 4667
rect 7673 4633 7687 4647
rect 7653 4513 7667 4527
rect 7613 4453 7627 4467
rect 7633 4453 7647 4467
rect 7753 4533 7767 4547
rect 7733 4493 7747 4507
rect 7673 4453 7687 4467
rect 7693 4453 7707 4467
rect 7593 4373 7607 4387
rect 7673 4433 7687 4447
rect 7633 4413 7647 4427
rect 7693 4413 7707 4427
rect 7633 4393 7647 4407
rect 7613 4293 7627 4307
rect 7613 4233 7627 4247
rect 7533 4213 7547 4227
rect 7573 4213 7587 4227
rect 7553 4193 7567 4207
rect 7673 4273 7687 4287
rect 7673 4213 7687 4227
rect 7633 4193 7647 4207
rect 7653 4193 7667 4207
rect 7533 4173 7547 4187
rect 7593 4173 7607 4187
rect 7613 4173 7627 4187
rect 7633 4153 7647 4167
rect 7653 4153 7667 4167
rect 7613 4013 7627 4027
rect 7553 3993 7567 4007
rect 7573 3993 7587 4007
rect 7593 3993 7607 4007
rect 7533 3973 7547 3987
rect 7573 3973 7587 3987
rect 7613 3973 7627 3987
rect 7533 3933 7547 3947
rect 7593 3953 7607 3967
rect 7553 3913 7567 3927
rect 7533 3773 7547 3787
rect 7553 3773 7567 3787
rect 7513 3753 7527 3767
rect 7593 3753 7607 3767
rect 7613 3753 7627 3767
rect 7713 4253 7727 4267
rect 7713 4233 7727 4247
rect 7813 4913 7827 4927
rect 7853 4713 7867 4727
rect 7813 4693 7827 4707
rect 7773 4493 7787 4507
rect 7793 4493 7807 4507
rect 7833 4513 7847 4527
rect 7873 4513 7887 4527
rect 7853 4493 7867 4507
rect 7813 4473 7827 4487
rect 7753 4453 7767 4467
rect 7833 4453 7847 4467
rect 7773 4433 7787 4447
rect 7813 4433 7827 4447
rect 7753 4233 7767 4247
rect 7873 4393 7887 4407
rect 7913 4753 7927 4767
rect 7893 4273 7907 4287
rect 7773 4213 7787 4227
rect 7813 4213 7827 4227
rect 7833 4213 7847 4227
rect 7853 4213 7867 4227
rect 7893 4213 7907 4227
rect 7753 4193 7767 4207
rect 7793 4193 7807 4207
rect 7773 4173 7787 4187
rect 7733 4133 7747 4147
rect 7713 4053 7727 4067
rect 7713 4033 7727 4047
rect 7673 4013 7687 4027
rect 7693 4013 7707 4027
rect 7773 4153 7787 4167
rect 7753 4033 7767 4047
rect 7673 3993 7687 4007
rect 7833 4173 7847 4187
rect 7873 4173 7887 4187
rect 7813 4133 7827 4147
rect 7813 4093 7827 4107
rect 7853 4093 7867 4107
rect 7853 4053 7867 4067
rect 7833 4033 7847 4047
rect 7873 4033 7887 4047
rect 7793 4013 7807 4027
rect 7833 4013 7847 4027
rect 7853 4013 7867 4027
rect 7773 3993 7787 4007
rect 7653 3973 7667 3987
rect 7693 3973 7707 3987
rect 7713 3973 7727 3987
rect 7673 3953 7687 3967
rect 7693 3933 7707 3947
rect 7673 3873 7687 3887
rect 7653 3853 7667 3867
rect 7653 3833 7667 3847
rect 7373 3553 7387 3567
rect 7413 3553 7427 3567
rect 7433 3553 7447 3567
rect 7553 3733 7567 3747
rect 7593 3733 7607 3747
rect 7633 3733 7647 3747
rect 7573 3713 7587 3727
rect 7573 3693 7587 3707
rect 7393 3513 7407 3527
rect 7353 3493 7367 3507
rect 7193 3233 7207 3247
rect 7233 3233 7247 3247
rect 7313 3233 7327 3247
rect 7333 3233 7347 3247
rect 7133 3053 7147 3067
rect 7053 3013 7067 3027
rect 7113 3013 7127 3027
rect 7153 3033 7167 3047
rect 7213 3193 7227 3207
rect 7253 3213 7267 3227
rect 7373 3233 7387 3247
rect 7293 3193 7307 3207
rect 7313 3193 7327 3207
rect 7353 3193 7367 3207
rect 7273 3173 7287 3187
rect 7333 3093 7347 3107
rect 7253 3073 7267 3087
rect 7173 2993 7187 3007
rect 7053 2973 7067 2987
rect 7013 2773 7027 2787
rect 6933 2733 6947 2747
rect 6693 2713 6707 2727
rect 6813 2713 6827 2727
rect 6873 2713 6887 2727
rect 6653 2693 6667 2707
rect 6633 2653 6647 2667
rect 6573 2633 6587 2647
rect 6573 2573 6587 2587
rect 6513 2553 6527 2567
rect 6553 2553 6567 2567
rect 6433 2513 6447 2527
rect 6133 2293 6147 2307
rect 6193 2293 6207 2307
rect 6013 2273 6027 2287
rect 6113 2273 6127 2287
rect 6233 2273 6247 2287
rect 6273 2273 6287 2287
rect 6373 2293 6387 2307
rect 6333 2273 6347 2287
rect 6213 2233 6227 2247
rect 5993 2213 6007 2227
rect 6113 2173 6127 2187
rect 5953 2093 5967 2107
rect 5953 2073 5967 2087
rect 5873 2053 5887 2067
rect 5933 2053 5947 2067
rect 5973 2053 5987 2067
rect 6013 2053 6027 2067
rect 6073 2053 6087 2067
rect 5833 2033 5847 2047
rect 5773 2013 5787 2027
rect 5913 1973 5927 1987
rect 5633 1873 5647 1887
rect 5613 1593 5627 1607
rect 5753 1833 5767 1847
rect 5673 1813 5687 1827
rect 5713 1753 5727 1767
rect 5853 1793 5867 1807
rect 5833 1753 5847 1767
rect 5813 1733 5827 1747
rect 5753 1673 5767 1687
rect 5693 1653 5707 1667
rect 5893 1773 5907 1787
rect 5893 1733 5907 1747
rect 5773 1613 5787 1627
rect 5833 1613 5847 1627
rect 5873 1613 5887 1627
rect 5653 1593 5667 1607
rect 5793 1593 5807 1607
rect 5553 1533 5567 1547
rect 5573 1493 5587 1507
rect 5653 1553 5667 1567
rect 5633 1353 5647 1367
rect 5533 1333 5547 1347
rect 5573 1313 5587 1327
rect 5613 1313 5627 1327
rect 5593 1293 5607 1307
rect 5713 1573 5727 1587
rect 5753 1573 5767 1587
rect 5673 1473 5687 1487
rect 5693 1453 5707 1467
rect 5673 1333 5687 1347
rect 5733 1353 5747 1367
rect 5673 1293 5687 1307
rect 5693 1293 5707 1307
rect 5493 1273 5507 1287
rect 5613 1133 5627 1147
rect 5573 1113 5587 1127
rect 5653 1113 5667 1127
rect 5453 1093 5467 1107
rect 5353 1073 5367 1087
rect 5273 853 5287 867
rect 5313 853 5327 867
rect 5473 1073 5487 1087
rect 5633 1093 5647 1107
rect 5693 1093 5707 1107
rect 5593 1053 5607 1067
rect 5433 1033 5447 1047
rect 5473 1033 5487 1047
rect 5473 973 5487 987
rect 5553 973 5567 987
rect 5593 973 5607 987
rect 5433 933 5447 947
rect 5013 833 5027 847
rect 5213 833 5227 847
rect 5173 813 5187 827
rect 5333 833 5347 847
rect 5133 793 5147 807
rect 4513 773 4527 787
rect 4553 773 4567 787
rect 4593 773 4607 787
rect 4513 673 4527 687
rect 4033 633 4047 647
rect 4013 613 4027 627
rect 4053 613 4067 627
rect 4153 633 4167 647
rect 4233 633 4247 647
rect 4193 613 4207 627
rect 4233 613 4247 627
rect 4293 613 4307 627
rect 4333 613 4347 627
rect 4173 593 4187 607
rect 4093 573 4107 587
rect 4113 573 4127 587
rect 4093 553 4107 567
rect 4053 393 4067 407
rect 3993 373 4007 387
rect 4033 313 4047 327
rect 4073 313 4087 327
rect 4373 553 4387 567
rect 4353 493 4367 507
rect 4113 433 4127 447
rect 4133 433 4147 447
rect 4213 433 4227 447
rect 4113 393 4127 407
rect 4093 293 4107 307
rect 4053 273 4067 287
rect 3973 173 3987 187
rect 3953 153 3967 167
rect 3993 153 4007 167
rect 3973 133 3987 147
rect 4113 233 4127 247
rect 4093 153 4107 167
rect 4313 373 4327 387
rect 4253 353 4267 367
rect 4293 353 4307 367
rect 4193 313 4207 327
rect 4233 313 4247 327
rect 4273 213 4287 227
rect 4533 653 4547 667
rect 4993 713 5007 727
rect 4713 693 4727 707
rect 4833 693 4847 707
rect 4473 453 4487 467
rect 4413 433 4427 447
rect 4433 373 4447 387
rect 4553 633 4567 647
rect 4513 593 4527 607
rect 4493 393 4507 407
rect 4393 353 4407 367
rect 4433 353 4447 367
rect 4453 353 4467 367
rect 4313 273 4327 287
rect 4413 333 4427 347
rect 4373 273 4387 287
rect 4333 253 4347 267
rect 4173 193 4187 207
rect 4293 193 4307 207
rect 4313 193 4327 207
rect 4153 173 4167 187
rect 4153 153 4167 167
rect 4093 133 4107 147
rect 4133 133 4147 147
rect 4773 653 4787 667
rect 4613 613 4627 627
rect 4813 633 4827 647
rect 4773 533 4787 547
rect 4773 513 4787 527
rect 4693 493 4707 507
rect 4573 473 4587 487
rect 4633 433 4647 447
rect 4553 373 4567 387
rect 4573 353 4587 367
rect 4513 333 4527 347
rect 4533 253 4547 267
rect 4333 173 4347 187
rect 4433 173 4447 187
rect 4453 173 4467 187
rect 4033 113 4047 127
rect 4073 113 4087 127
rect 4273 93 4287 107
rect 4413 153 4427 167
rect 4493 153 4507 167
rect 4773 413 4787 427
rect 4653 373 4667 387
rect 4693 373 4707 387
rect 4713 373 4727 387
rect 4733 373 4747 387
rect 4593 333 4607 347
rect 4633 293 4647 307
rect 4553 233 4567 247
rect 4573 233 4587 247
rect 4513 133 4527 147
rect 4473 113 4487 127
rect 4593 133 4607 147
rect 4713 333 4727 347
rect 4753 313 4767 327
rect 4693 253 4707 267
rect 4713 253 4727 267
rect 4673 173 4687 187
rect 4693 133 4707 147
rect 4973 673 4987 687
rect 4933 633 4947 647
rect 5173 673 5187 687
rect 4993 653 5007 667
rect 5033 633 5047 647
rect 4813 573 4827 587
rect 4793 393 4807 407
rect 4893 573 4907 587
rect 4953 553 4967 567
rect 4893 533 4907 547
rect 4873 513 4887 527
rect 4833 473 4847 487
rect 4933 413 4947 427
rect 4853 353 4867 367
rect 4893 313 4907 327
rect 4813 293 4827 307
rect 4913 293 4927 307
rect 4993 453 5007 467
rect 4813 253 4827 267
rect 4953 253 4967 267
rect 4773 153 4787 167
rect 4953 213 4967 227
rect 4853 173 4867 187
rect 4793 133 4807 147
rect 4833 133 4847 147
rect 4913 133 4927 147
rect 4753 113 4767 127
rect 4893 113 4907 127
rect 4973 173 4987 187
rect 5053 613 5067 627
rect 5133 653 5147 667
rect 5113 613 5127 627
rect 5073 593 5087 607
rect 5073 433 5087 447
rect 5233 653 5247 667
rect 5393 713 5407 727
rect 5353 693 5367 707
rect 5253 633 5267 647
rect 5513 853 5527 867
rect 5513 833 5527 847
rect 5533 813 5547 827
rect 5453 793 5467 807
rect 5493 793 5507 807
rect 5433 633 5447 647
rect 5193 613 5207 627
rect 5253 533 5267 547
rect 5173 493 5187 507
rect 5133 413 5147 427
rect 5133 393 5147 407
rect 5033 373 5047 387
rect 5073 373 5087 387
rect 5093 353 5107 367
rect 5173 373 5187 387
rect 5113 313 5127 327
rect 5173 313 5187 327
rect 5153 273 5167 287
rect 5173 253 5187 267
rect 5013 213 5027 227
rect 5053 213 5067 227
rect 5133 193 5147 207
rect 5113 173 5127 187
rect 5133 153 5147 167
rect 5213 373 5227 387
rect 5373 613 5387 627
rect 5853 1593 5867 1607
rect 5893 1593 5907 1607
rect 5873 1573 5887 1587
rect 6293 2253 6307 2267
rect 6373 2233 6387 2247
rect 6253 2213 6267 2227
rect 6213 2113 6227 2127
rect 6173 2073 6187 2087
rect 6053 2013 6067 2027
rect 6193 2053 6207 2067
rect 6393 2113 6407 2127
rect 6353 2093 6367 2107
rect 6413 2093 6427 2107
rect 6293 2073 6307 2087
rect 6333 2073 6347 2087
rect 6373 2073 6387 2087
rect 6413 2073 6427 2087
rect 6313 2033 6327 2047
rect 6333 2033 6347 2047
rect 6233 1973 6247 1987
rect 6013 1873 6027 1887
rect 5993 1853 6007 1867
rect 6053 1853 6067 1867
rect 6193 1853 6207 1867
rect 6013 1833 6027 1847
rect 6053 1833 6067 1847
rect 6073 1793 6087 1807
rect 6113 1793 6127 1807
rect 6033 1773 6047 1787
rect 5953 1753 5967 1767
rect 5933 1673 5947 1687
rect 5973 1653 5987 1667
rect 5933 1633 5947 1647
rect 5953 1633 5967 1647
rect 6093 1773 6107 1787
rect 6133 1773 6147 1787
rect 6153 1673 6167 1687
rect 6073 1633 6087 1647
rect 6133 1633 6147 1647
rect 6073 1613 6087 1627
rect 5993 1593 6007 1607
rect 6393 1993 6407 2007
rect 6253 1813 6267 1827
rect 6233 1793 6247 1807
rect 6193 1773 6207 1787
rect 6313 1773 6327 1787
rect 6293 1753 6307 1767
rect 6273 1673 6287 1687
rect 6213 1653 6227 1667
rect 6173 1613 6187 1627
rect 6233 1613 6247 1627
rect 5933 1573 5947 1587
rect 6013 1573 6027 1587
rect 6053 1573 6067 1587
rect 5873 1553 5887 1567
rect 5913 1553 5927 1567
rect 5873 1473 5887 1487
rect 5793 1313 5807 1327
rect 5773 1293 5787 1307
rect 5813 1293 5827 1307
rect 6373 1813 6387 1827
rect 6373 1753 6387 1767
rect 6333 1653 6347 1667
rect 6593 2533 6607 2547
rect 6573 2493 6587 2507
rect 6493 2413 6507 2427
rect 6533 2413 6547 2427
rect 6453 2293 6467 2307
rect 6473 2273 6487 2287
rect 6513 2173 6527 2187
rect 6533 2113 6547 2127
rect 6433 1833 6447 1847
rect 6493 2033 6507 2047
rect 6473 1973 6487 1987
rect 6433 1793 6447 1807
rect 6453 1793 6467 1807
rect 6553 1833 6567 1847
rect 6513 1813 6527 1827
rect 6493 1793 6507 1807
rect 6533 1793 6547 1807
rect 6453 1753 6467 1767
rect 6493 1753 6507 1767
rect 6413 1713 6427 1727
rect 6833 2633 6847 2647
rect 6653 2613 6667 2627
rect 6733 2613 6747 2627
rect 6793 2613 6807 2627
rect 6693 2573 6707 2587
rect 6773 2573 6787 2587
rect 6673 2553 6687 2567
rect 6713 2553 6727 2567
rect 6753 2533 6767 2547
rect 6653 2493 6667 2507
rect 6673 2333 6687 2347
rect 6653 2253 6667 2267
rect 6633 2133 6647 2147
rect 6633 2113 6647 2127
rect 6593 2073 6607 2087
rect 6613 2053 6627 2067
rect 6813 2573 6827 2587
rect 6973 2733 6987 2747
rect 7013 2693 7027 2707
rect 6973 2653 6987 2667
rect 7013 2613 7027 2627
rect 6953 2533 6967 2547
rect 7233 3033 7247 3047
rect 7213 3013 7227 3027
rect 7293 3033 7307 3047
rect 7273 2993 7287 3007
rect 7273 2793 7287 2807
rect 7213 2733 7227 2747
rect 7193 2713 7207 2727
rect 7173 2653 7187 2667
rect 7213 2613 7227 2627
rect 7173 2593 7187 2607
rect 7133 2573 7147 2587
rect 7073 2513 7087 2527
rect 6893 2493 6907 2507
rect 6953 2333 6967 2347
rect 6853 2293 6867 2307
rect 7153 2553 7167 2567
rect 7313 2773 7327 2787
rect 7293 2593 7307 2607
rect 7293 2573 7307 2587
rect 7253 2553 7267 2567
rect 7193 2533 7207 2547
rect 7313 2553 7327 2567
rect 7473 3533 7487 3547
rect 7433 3513 7447 3527
rect 7453 3493 7467 3507
rect 7553 3553 7567 3567
rect 7513 3293 7527 3307
rect 7613 3713 7627 3727
rect 7673 3733 7687 3747
rect 7673 3693 7687 3707
rect 7673 3553 7687 3567
rect 7593 3533 7607 3547
rect 7633 3533 7647 3547
rect 7653 3533 7667 3547
rect 7573 3513 7587 3527
rect 7593 3513 7607 3527
rect 7573 3473 7587 3487
rect 7753 3973 7767 3987
rect 7733 3933 7747 3947
rect 7733 3853 7747 3867
rect 7713 3633 7727 3647
rect 7713 3553 7727 3567
rect 7813 3993 7827 4007
rect 7853 3993 7867 4007
rect 7793 3953 7807 3967
rect 7853 3953 7867 3967
rect 7793 3933 7807 3947
rect 7833 3933 7847 3947
rect 7773 3873 7787 3887
rect 7793 3813 7807 3827
rect 7753 3753 7767 3767
rect 7753 3733 7767 3747
rect 7813 3733 7827 3747
rect 7833 3733 7847 3747
rect 7773 3713 7787 3727
rect 7773 3693 7787 3707
rect 7733 3533 7747 3547
rect 7753 3533 7767 3547
rect 7833 3693 7847 3707
rect 7793 3653 7807 3667
rect 7793 3633 7807 3647
rect 7693 3513 7707 3527
rect 7793 3513 7807 3527
rect 7853 3553 7867 3567
rect 7913 3833 7927 3847
rect 7913 3813 7927 3827
rect 7893 3693 7907 3707
rect 7893 3673 7907 3687
rect 7673 3493 7687 3507
rect 7713 3493 7727 3507
rect 7753 3493 7767 3507
rect 7773 3493 7787 3507
rect 7813 3493 7827 3507
rect 7853 3493 7867 3507
rect 7553 3273 7567 3287
rect 7413 3253 7427 3267
rect 7473 3253 7487 3267
rect 7653 3453 7667 3467
rect 7593 3293 7607 3307
rect 7393 3073 7407 3087
rect 7373 3053 7387 3067
rect 7453 3173 7467 3187
rect 7493 3233 7507 3247
rect 7473 3093 7487 3107
rect 7433 3053 7447 3067
rect 7453 3053 7467 3067
rect 7373 3013 7387 3027
rect 7453 3013 7467 3027
rect 7533 3073 7547 3087
rect 7613 3253 7627 3267
rect 7633 3193 7647 3207
rect 7673 3273 7687 3287
rect 7733 3453 7747 3467
rect 7673 3253 7687 3267
rect 7713 3253 7727 3267
rect 7693 3213 7707 3227
rect 7713 3093 7727 3107
rect 7653 3073 7667 3087
rect 7693 3073 7707 3087
rect 7613 3053 7627 3067
rect 7653 3053 7667 3067
rect 7613 3033 7627 3047
rect 7533 3013 7547 3027
rect 7573 3013 7587 3027
rect 7513 2973 7527 2987
rect 7553 2993 7567 3007
rect 7593 2993 7607 3007
rect 7533 2913 7547 2927
rect 7533 2893 7547 2907
rect 7493 2793 7507 2807
rect 7513 2773 7527 2787
rect 7393 2733 7407 2747
rect 7353 2713 7367 2727
rect 7453 2733 7467 2747
rect 7433 2613 7447 2627
rect 7413 2593 7427 2607
rect 7393 2573 7407 2587
rect 7353 2553 7367 2567
rect 7373 2553 7387 2567
rect 7273 2513 7287 2527
rect 7333 2513 7347 2527
rect 7193 2493 7207 2507
rect 7233 2493 7247 2507
rect 7313 2493 7327 2507
rect 7153 2473 7167 2487
rect 6813 2273 6827 2287
rect 6753 2253 6767 2267
rect 6773 2253 6787 2267
rect 6813 2233 6827 2247
rect 6873 2233 6887 2247
rect 6713 2093 6727 2107
rect 6733 2093 6747 2107
rect 6753 2093 6767 2107
rect 6773 2093 6787 2107
rect 6793 2073 6807 2087
rect 6593 1973 6607 1987
rect 6653 1973 6667 1987
rect 6733 2053 6747 2067
rect 6713 2033 6727 2047
rect 6853 2213 6867 2227
rect 6973 2293 6987 2307
rect 6993 2293 7007 2307
rect 7033 2293 7047 2307
rect 7053 2293 7067 2307
rect 7133 2293 7147 2307
rect 6933 2273 6947 2287
rect 6973 2233 6987 2247
rect 7013 2233 7027 2247
rect 7033 2153 7047 2167
rect 6993 2133 7007 2147
rect 6893 2113 6907 2127
rect 6973 2093 6987 2107
rect 6873 2033 6887 2047
rect 6913 2033 6927 2047
rect 6593 1793 6607 1807
rect 6633 1793 6647 1807
rect 6653 1773 6667 1787
rect 6573 1693 6587 1707
rect 6653 1753 6667 1767
rect 6473 1653 6487 1667
rect 6493 1653 6507 1667
rect 6633 1653 6647 1667
rect 6653 1653 6667 1667
rect 6093 1373 6107 1387
rect 6213 1373 6227 1387
rect 6393 1593 6407 1607
rect 6593 1633 6607 1647
rect 6553 1613 6567 1627
rect 6613 1613 6627 1627
rect 6433 1573 6447 1587
rect 6693 1793 6707 1807
rect 6733 1873 6747 1887
rect 6713 1653 6727 1667
rect 6673 1633 6687 1647
rect 6713 1633 6727 1647
rect 6573 1573 6587 1587
rect 6793 1853 6807 1867
rect 6933 1853 6947 1867
rect 6753 1813 6767 1827
rect 6873 1833 6887 1847
rect 6833 1813 6847 1827
rect 6893 1813 6907 1827
rect 7173 2273 7187 2287
rect 7113 2253 7127 2267
rect 7153 2253 7167 2267
rect 7233 2473 7247 2487
rect 7253 2333 7267 2347
rect 7333 2313 7347 2327
rect 7313 2293 7327 2307
rect 7293 2273 7307 2287
rect 7133 2133 7147 2147
rect 7053 2073 7067 2087
rect 7053 2053 7067 2067
rect 7013 2033 7027 2047
rect 6773 1753 6787 1767
rect 6993 1793 7007 1807
rect 7053 1793 7067 1807
rect 7093 1793 7107 1807
rect 7073 1753 7087 1767
rect 7113 1753 7127 1767
rect 7033 1673 7047 1687
rect 7033 1633 7047 1647
rect 7053 1633 7067 1647
rect 6893 1613 6907 1627
rect 6953 1613 6967 1627
rect 6673 1553 6687 1567
rect 6733 1553 6747 1567
rect 6553 1533 6567 1547
rect 6693 1533 6707 1547
rect 6193 1313 6207 1327
rect 6233 1313 6247 1327
rect 6353 1333 6367 1347
rect 6373 1333 6387 1347
rect 6493 1333 6507 1347
rect 6513 1333 6527 1347
rect 6553 1333 6567 1347
rect 6613 1333 6627 1347
rect 5933 1273 5947 1287
rect 5773 1253 5787 1267
rect 5733 1133 5747 1147
rect 5893 1153 5907 1167
rect 5853 1113 5867 1127
rect 5833 1093 5847 1107
rect 5713 1053 5727 1067
rect 5793 1073 5807 1087
rect 5753 1033 5767 1047
rect 5653 953 5667 967
rect 5633 873 5647 887
rect 5593 853 5607 867
rect 5633 853 5647 867
rect 5853 1033 5867 1047
rect 5873 1033 5887 1047
rect 5793 933 5807 947
rect 5693 853 5707 867
rect 5753 853 5767 867
rect 5613 833 5627 847
rect 5673 833 5687 847
rect 5633 813 5647 827
rect 5573 633 5587 647
rect 5553 613 5567 627
rect 5413 593 5427 607
rect 5453 593 5467 607
rect 5333 573 5347 587
rect 5293 513 5307 527
rect 5313 413 5327 427
rect 5233 313 5247 327
rect 5253 233 5267 247
rect 5553 393 5567 407
rect 5373 373 5387 387
rect 5613 373 5627 387
rect 5353 353 5367 367
rect 5433 353 5447 367
rect 5473 353 5487 367
rect 5513 353 5527 367
rect 5273 173 5287 187
rect 5313 173 5327 187
rect 5173 133 5187 147
rect 5233 133 5247 147
rect 5533 333 5547 347
rect 5513 313 5527 327
rect 5553 313 5567 327
rect 5513 273 5527 287
rect 5493 253 5507 267
rect 5473 193 5487 207
rect 5333 133 5347 147
rect 5453 153 5467 167
rect 5573 233 5587 247
rect 5833 813 5847 827
rect 5673 793 5687 807
rect 5833 673 5847 687
rect 5753 653 5767 667
rect 5713 633 5727 647
rect 5733 613 5747 627
rect 5773 613 5787 627
rect 5813 613 5827 627
rect 5793 593 5807 607
rect 6093 1293 6107 1307
rect 6053 1233 6067 1247
rect 6073 1173 6087 1187
rect 6133 1173 6147 1187
rect 5993 1093 6007 1107
rect 6033 1093 6047 1107
rect 6093 1133 6107 1147
rect 6113 1133 6127 1147
rect 5953 1073 5967 1087
rect 5973 1073 5987 1087
rect 5993 1053 6007 1067
rect 5973 953 5987 967
rect 5933 873 5947 887
rect 5893 853 5907 867
rect 5873 813 5887 827
rect 5933 833 5947 847
rect 5953 573 5967 587
rect 6033 1053 6047 1067
rect 6153 1093 6167 1107
rect 6213 1293 6227 1307
rect 6253 1273 6267 1287
rect 6373 1313 6387 1327
rect 6373 1273 6387 1287
rect 6293 1253 6307 1267
rect 6333 1253 6347 1267
rect 6373 1253 6387 1267
rect 6413 1253 6427 1267
rect 6293 1173 6307 1187
rect 6353 1173 6367 1187
rect 6213 1153 6227 1167
rect 6433 1213 6447 1227
rect 6393 1173 6407 1187
rect 6373 1133 6387 1147
rect 6253 1113 6267 1127
rect 6293 1113 6307 1127
rect 6333 1113 6347 1127
rect 6453 1153 6467 1167
rect 6233 1093 6247 1107
rect 6273 1093 6287 1107
rect 6193 1053 6207 1067
rect 6313 1093 6327 1107
rect 6153 1033 6167 1047
rect 6253 1033 6267 1047
rect 6293 1033 6307 1047
rect 5993 893 6007 907
rect 6033 893 6047 907
rect 5993 833 6007 847
rect 6153 873 6167 887
rect 6013 813 6027 827
rect 6053 813 6067 827
rect 6093 813 6107 827
rect 6053 793 6067 807
rect 6013 613 6027 627
rect 6073 593 6087 607
rect 6173 793 6187 807
rect 6193 793 6207 807
rect 6173 753 6187 767
rect 6233 713 6247 727
rect 6133 653 6147 667
rect 6413 1073 6427 1087
rect 6433 853 6447 867
rect 6413 833 6427 847
rect 6533 1313 6547 1327
rect 6533 1293 6547 1307
rect 6613 1293 6627 1307
rect 6493 953 6507 967
rect 6513 873 6527 887
rect 6473 833 6487 847
rect 6373 813 6387 827
rect 6453 813 6467 827
rect 6493 813 6507 827
rect 6693 1273 6707 1287
rect 6653 1253 6667 1267
rect 6573 1093 6587 1107
rect 6693 1233 6707 1247
rect 6733 1213 6747 1227
rect 6553 1033 6567 1047
rect 6533 853 6547 867
rect 6633 1033 6647 1047
rect 6673 1033 6687 1047
rect 6593 993 6607 1007
rect 6533 813 6547 827
rect 6273 753 6287 767
rect 6313 793 6327 807
rect 6313 713 6327 727
rect 6493 713 6507 727
rect 6293 693 6307 707
rect 6133 613 6147 627
rect 6093 573 6107 587
rect 6033 553 6047 567
rect 5973 533 5987 547
rect 5853 473 5867 487
rect 5653 353 5667 367
rect 5753 373 5767 387
rect 5813 373 5827 387
rect 5853 373 5867 387
rect 5793 353 5807 367
rect 5673 293 5687 307
rect 5793 333 5807 347
rect 5853 353 5867 367
rect 6133 573 6147 587
rect 6113 533 6127 547
rect 6093 353 6107 367
rect 5953 333 5967 347
rect 5813 293 5827 307
rect 5733 253 5747 267
rect 5973 313 5987 327
rect 6013 313 6027 327
rect 5993 273 6007 287
rect 5833 233 5847 247
rect 6073 213 6087 227
rect 5633 193 5647 207
rect 5713 193 5727 207
rect 5973 193 5987 207
rect 5753 153 5767 167
rect 5933 153 5947 167
rect 6273 633 6287 647
rect 6193 553 6207 567
rect 6173 333 6187 347
rect 6213 333 6227 347
rect 6453 693 6467 707
rect 6373 653 6387 667
rect 6413 653 6427 667
rect 6433 653 6447 667
rect 6333 633 6347 647
rect 6313 613 6327 627
rect 6353 613 6367 627
rect 6393 613 6407 627
rect 6333 593 6347 607
rect 6473 653 6487 667
rect 6533 653 6547 667
rect 6433 613 6447 627
rect 6373 413 6387 427
rect 6333 373 6347 387
rect 6273 353 6287 367
rect 6353 353 6367 367
rect 6313 333 6327 347
rect 6233 293 6247 307
rect 6353 273 6367 287
rect 6193 193 6207 207
rect 6073 173 6087 187
rect 6093 173 6107 187
rect 6153 173 6167 187
rect 6187 173 6201 187
rect 6293 173 6307 187
rect 6573 593 6587 607
rect 6713 993 6727 1007
rect 6673 773 6687 787
rect 6773 1593 6787 1607
rect 6793 1353 6807 1367
rect 7013 1593 7027 1607
rect 6913 1373 6927 1387
rect 6853 1293 6867 1307
rect 6893 1293 6907 1307
rect 6793 1053 6807 1067
rect 6753 793 6767 807
rect 6693 673 6707 687
rect 6613 633 6627 647
rect 6753 653 6767 667
rect 6593 493 6607 507
rect 6553 433 6567 447
rect 6593 433 6607 447
rect 6453 393 6467 407
rect 6493 393 6507 407
rect 6553 393 6567 407
rect 6413 373 6427 387
rect 6473 373 6487 387
rect 6513 353 6527 367
rect 6433 313 6447 327
rect 6473 313 6487 327
rect 6493 313 6507 327
rect 6533 313 6547 327
rect 6473 273 6487 287
rect 6393 193 6407 207
rect 6213 153 6227 167
rect 6113 133 6127 147
rect 6193 133 6207 147
rect 6233 133 6247 147
rect 6313 153 6327 167
rect 6393 153 6407 167
rect 6553 253 6567 267
rect 6653 613 6667 627
rect 6773 613 6787 627
rect 6833 1113 6847 1127
rect 6833 1073 6847 1087
rect 6813 673 6827 687
rect 6633 593 6647 607
rect 6773 593 6787 607
rect 6693 573 6707 587
rect 6673 493 6687 507
rect 6613 373 6627 387
rect 6653 373 6667 387
rect 6953 1353 6967 1367
rect 6933 1273 6947 1287
rect 6973 1293 6987 1307
rect 7053 1333 7067 1347
rect 7033 1273 7047 1287
rect 6913 1093 6927 1107
rect 6993 1133 7007 1147
rect 7153 2033 7167 2047
rect 7233 2133 7247 2147
rect 7293 2113 7307 2127
rect 7273 2073 7287 2087
rect 7193 1873 7207 1887
rect 7213 1873 7227 1887
rect 7153 1753 7167 1767
rect 7173 1753 7187 1767
rect 7193 1733 7207 1747
rect 7133 1633 7147 1647
rect 7193 1573 7207 1587
rect 7133 1533 7147 1547
rect 7153 1533 7167 1547
rect 7133 1373 7147 1387
rect 7093 1333 7107 1347
rect 7233 1773 7247 1787
rect 7233 1753 7247 1767
rect 7253 1753 7267 1767
rect 7273 1753 7287 1767
rect 7473 2593 7487 2607
rect 7493 2593 7507 2607
rect 7473 2553 7487 2567
rect 7393 2513 7407 2527
rect 7373 2493 7387 2507
rect 7353 2253 7367 2267
rect 7453 2513 7467 2527
rect 7433 2313 7447 2327
rect 7493 2533 7507 2547
rect 7493 2513 7507 2527
rect 7473 2293 7487 2307
rect 7393 2213 7407 2227
rect 7453 2253 7467 2267
rect 7413 2153 7427 2167
rect 7373 2113 7387 2127
rect 7473 2093 7487 2107
rect 7433 2073 7447 2087
rect 7413 2053 7427 2067
rect 7453 2053 7467 2067
rect 7593 2913 7607 2927
rect 7553 2653 7567 2667
rect 7673 2973 7687 2987
rect 7653 2873 7667 2887
rect 7633 2773 7647 2787
rect 7813 3453 7827 3467
rect 7793 3273 7807 3287
rect 7813 3273 7827 3287
rect 7873 3473 7887 3487
rect 7853 3273 7867 3287
rect 7873 3253 7887 3267
rect 7853 3093 7867 3107
rect 7813 3073 7827 3087
rect 7853 3073 7867 3087
rect 7793 3053 7807 3067
rect 7833 3053 7847 3067
rect 7793 3033 7807 3047
rect 7733 2893 7747 2907
rect 7813 3013 7827 3027
rect 7853 3013 7867 3027
rect 7793 2993 7807 3007
rect 7733 2873 7747 2887
rect 7793 2793 7807 2807
rect 7833 2873 7847 2887
rect 7633 2733 7647 2747
rect 7753 2773 7767 2787
rect 7813 2773 7827 2787
rect 7533 2333 7547 2347
rect 7613 2553 7627 2567
rect 7793 2753 7807 2767
rect 7773 2733 7787 2747
rect 7813 2733 7827 2747
rect 7773 2713 7787 2727
rect 7813 2713 7827 2727
rect 7853 2713 7867 2727
rect 7673 2553 7687 2567
rect 7713 2553 7727 2567
rect 7753 2553 7767 2567
rect 7613 2513 7627 2527
rect 7633 2513 7647 2527
rect 7753 2513 7767 2527
rect 7573 2313 7587 2327
rect 7593 2313 7607 2327
rect 7513 2293 7527 2307
rect 7553 2293 7567 2307
rect 7653 2333 7667 2347
rect 7633 2313 7647 2327
rect 7533 2273 7547 2287
rect 7573 2253 7587 2267
rect 7513 2113 7527 2127
rect 7593 2113 7607 2127
rect 7493 2033 7507 2047
rect 7533 2033 7547 2047
rect 7413 1853 7427 1867
rect 7333 1833 7347 1847
rect 7313 1813 7327 1827
rect 7473 1833 7487 1847
rect 7453 1793 7467 1807
rect 7333 1773 7347 1787
rect 7313 1753 7327 1767
rect 7333 1753 7347 1767
rect 7293 1733 7307 1747
rect 7333 1733 7347 1747
rect 7233 1613 7247 1627
rect 7273 1593 7287 1607
rect 7253 1573 7267 1587
rect 7293 1573 7307 1587
rect 7333 1553 7347 1567
rect 7373 1733 7387 1747
rect 7393 1733 7407 1747
rect 7393 1653 7407 1667
rect 7373 1613 7387 1627
rect 7373 1573 7387 1587
rect 7373 1533 7387 1547
rect 7353 1373 7367 1387
rect 7333 1353 7347 1367
rect 7173 1333 7187 1347
rect 7213 1333 7227 1347
rect 7633 2053 7647 2067
rect 7573 1873 7587 1887
rect 7573 1853 7587 1867
rect 7533 1813 7547 1827
rect 7553 1793 7567 1807
rect 7533 1753 7547 1767
rect 7473 1653 7487 1667
rect 7453 1633 7467 1647
rect 7513 1633 7527 1647
rect 7433 1613 7447 1627
rect 7493 1613 7507 1627
rect 7413 1593 7427 1607
rect 7793 2293 7807 2307
rect 7733 2213 7747 2227
rect 7673 2133 7687 2147
rect 7773 2133 7787 2147
rect 7713 2113 7727 2127
rect 7773 2053 7787 2067
rect 7613 1813 7627 1827
rect 7653 1813 7667 1827
rect 7593 1733 7607 1747
rect 7573 1593 7587 1607
rect 7433 1573 7447 1587
rect 7473 1573 7487 1587
rect 7533 1573 7547 1587
rect 7573 1573 7587 1587
rect 7553 1553 7567 1567
rect 7493 1373 7507 1387
rect 7393 1353 7407 1367
rect 7073 1313 7087 1327
rect 7113 1313 7127 1327
rect 7113 1273 7127 1287
rect 7053 1133 7067 1147
rect 6953 1113 6967 1127
rect 7033 1113 7047 1127
rect 6933 1073 6947 1087
rect 7013 1093 7027 1107
rect 7033 1073 7047 1087
rect 7073 1073 7087 1087
rect 7133 1073 7147 1087
rect 6973 1053 6987 1067
rect 7113 1053 7127 1067
rect 6893 1033 6907 1047
rect 7193 1313 7207 1327
rect 7233 1313 7247 1327
rect 7213 1293 7227 1307
rect 7193 1273 7207 1287
rect 7253 1273 7267 1287
rect 7433 1313 7447 1327
rect 7413 1293 7427 1307
rect 7353 1273 7367 1287
rect 7393 1273 7407 1287
rect 7293 1253 7307 1267
rect 7253 1133 7267 1147
rect 6973 853 6987 867
rect 6853 813 6867 827
rect 6873 813 6887 827
rect 6913 813 6927 827
rect 6873 693 6887 707
rect 6933 653 6947 667
rect 6933 613 6947 627
rect 6853 593 6867 607
rect 6893 593 6907 607
rect 6953 593 6967 607
rect 6833 573 6847 587
rect 6913 573 6927 587
rect 6773 413 6787 427
rect 6733 393 6747 407
rect 6733 373 6747 387
rect 6633 333 6647 347
rect 6593 273 6607 287
rect 6613 273 6627 287
rect 6573 233 6587 247
rect 6553 193 6567 207
rect 6493 173 6507 187
rect 6613 213 6627 227
rect 6593 193 6607 207
rect 6593 173 6607 187
rect 6673 313 6687 327
rect 6673 293 6687 307
rect 6673 213 6687 227
rect 6633 173 6647 187
rect 6293 133 6307 147
rect 6333 133 6347 147
rect 6753 273 6767 287
rect 6693 173 6707 187
rect 6733 173 6747 187
rect 7033 833 7047 847
rect 6993 813 7007 827
rect 7013 813 7027 827
rect 7173 853 7187 867
rect 6993 673 7007 687
rect 6793 373 6807 387
rect 6913 373 6927 387
rect 6973 373 6987 387
rect 6813 333 6827 347
rect 6973 333 6987 347
rect 6873 313 6887 327
rect 6933 313 6947 327
rect 6953 313 6967 327
rect 6853 273 6867 287
rect 6833 253 6847 267
rect 7013 653 7027 667
rect 7153 713 7167 727
rect 7073 633 7087 647
rect 7053 613 7067 627
rect 7073 593 7087 607
rect 7113 593 7127 607
rect 7313 1113 7327 1127
rect 7213 813 7227 827
rect 7173 673 7187 687
rect 7193 673 7207 687
rect 7213 673 7227 687
rect 7113 393 7127 407
rect 7153 393 7167 407
rect 7053 373 7067 387
rect 7093 373 7107 387
rect 7013 353 7027 367
rect 7173 333 7187 347
rect 7233 633 7247 647
rect 7233 373 7247 387
rect 7293 353 7307 367
rect 7253 333 7267 347
rect 7373 1093 7387 1107
rect 7353 1073 7367 1087
rect 7333 853 7347 867
rect 7373 853 7387 867
rect 7353 813 7367 827
rect 7513 1353 7527 1367
rect 7493 1273 7507 1287
rect 7473 1253 7487 1267
rect 7473 1233 7487 1247
rect 7453 1193 7467 1207
rect 7433 1173 7447 1187
rect 7553 1333 7567 1347
rect 7653 1793 7667 1807
rect 7693 1793 7707 1807
rect 7753 1793 7767 1807
rect 7673 1733 7687 1747
rect 7633 1713 7647 1727
rect 7673 1713 7687 1727
rect 7653 1613 7667 1627
rect 7773 1753 7787 1767
rect 7693 1613 7707 1627
rect 7713 1613 7727 1627
rect 7733 1613 7747 1627
rect 7793 1633 7807 1647
rect 7633 1573 7647 1587
rect 7773 1573 7787 1587
rect 7793 1573 7807 1587
rect 7693 1553 7707 1567
rect 7753 1553 7767 1567
rect 7593 1353 7607 1367
rect 7613 1353 7627 1367
rect 7593 1333 7607 1347
rect 7673 1333 7687 1347
rect 7573 1293 7587 1307
rect 7533 1273 7547 1287
rect 7513 1213 7527 1227
rect 7493 1133 7507 1147
rect 7533 1133 7547 1147
rect 7613 1293 7627 1307
rect 7713 1353 7727 1367
rect 7693 1313 7707 1327
rect 7613 1213 7627 1227
rect 7613 1153 7627 1167
rect 7673 1173 7687 1187
rect 7473 1113 7487 1127
rect 7613 1133 7627 1147
rect 7473 1093 7487 1107
rect 7513 1093 7527 1107
rect 7613 1093 7627 1107
rect 7453 1073 7467 1087
rect 7573 1073 7587 1087
rect 7593 1073 7607 1087
rect 7433 893 7447 907
rect 7433 873 7447 887
rect 7413 853 7427 867
rect 7333 653 7347 667
rect 7393 653 7407 667
rect 7413 653 7427 667
rect 7373 633 7387 647
rect 7353 613 7367 627
rect 7393 613 7407 627
rect 7333 413 7347 427
rect 7393 413 7407 427
rect 7373 393 7387 407
rect 7333 373 7347 387
rect 7353 353 7367 367
rect 7033 313 7047 327
rect 7213 313 7227 327
rect 7313 313 7327 327
rect 7153 213 7167 227
rect 7473 893 7487 907
rect 7453 853 7467 867
rect 7513 873 7527 887
rect 7553 873 7567 887
rect 7573 853 7587 867
rect 7473 833 7487 847
rect 7453 813 7467 827
rect 7493 813 7507 827
rect 7533 813 7547 827
rect 7493 753 7507 767
rect 7473 713 7487 727
rect 7453 653 7467 667
rect 7573 733 7587 747
rect 7573 713 7587 727
rect 7513 613 7527 627
rect 7653 1153 7667 1167
rect 7653 1133 7667 1147
rect 7753 1333 7767 1347
rect 7833 2573 7847 2587
rect 7873 2573 7887 2587
rect 7853 2273 7867 2287
rect 7913 3653 7927 3667
rect 7913 2733 7927 2747
rect 7893 2293 7907 2307
rect 7893 2273 7907 2287
rect 7853 2213 7867 2227
rect 7873 2093 7887 2107
rect 7893 2073 7907 2087
rect 7833 2053 7847 2067
rect 7853 2033 7867 2047
rect 7893 2033 7907 2047
rect 7893 1933 7907 1947
rect 7893 1893 7907 1907
rect 7853 1793 7867 1807
rect 7873 1773 7887 1787
rect 7873 1753 7887 1767
rect 7853 1713 7867 1727
rect 7853 1613 7867 1627
rect 7833 1593 7847 1607
rect 7853 1573 7867 1587
rect 7833 1553 7847 1567
rect 7813 1313 7827 1327
rect 7733 1233 7747 1247
rect 7793 1193 7807 1207
rect 7693 1133 7707 1147
rect 7713 1133 7727 1147
rect 7653 1113 7667 1127
rect 7633 873 7647 887
rect 7773 1133 7787 1147
rect 7753 1113 7767 1127
rect 7773 1093 7787 1107
rect 7773 933 7787 947
rect 7613 833 7627 847
rect 7653 833 7667 847
rect 7673 813 7687 827
rect 7633 753 7647 767
rect 7653 733 7667 747
rect 7593 653 7607 667
rect 7633 653 7647 667
rect 7593 633 7607 647
rect 7673 673 7687 687
rect 7733 853 7747 867
rect 7753 813 7767 827
rect 7713 793 7727 807
rect 7713 773 7727 787
rect 7753 793 7767 807
rect 7793 853 7807 867
rect 7793 813 7807 827
rect 7793 793 7807 807
rect 7733 713 7747 727
rect 7773 713 7787 727
rect 7773 673 7787 687
rect 7693 653 7707 667
rect 7753 653 7767 667
rect 7673 633 7687 647
rect 7733 633 7747 647
rect 7533 593 7547 607
rect 7613 613 7627 627
rect 7713 613 7727 627
rect 7653 593 7667 607
rect 7673 573 7687 587
rect 7513 453 7527 467
rect 7553 453 7567 467
rect 7453 393 7467 407
rect 7413 373 7427 387
rect 7433 373 7447 387
rect 7473 333 7487 347
rect 7633 313 7647 327
rect 7653 313 7667 327
rect 7593 293 7607 307
rect 7473 213 7487 227
rect 7033 193 7047 207
rect 7393 193 7407 207
rect 7453 193 7467 207
rect 7593 193 7607 207
rect 6733 153 6747 167
rect 6773 153 6787 167
rect 6913 153 6927 167
rect 6993 153 7007 167
rect 7133 173 7147 187
rect 7393 173 7407 187
rect 7233 153 7247 167
rect 7273 153 7287 167
rect 7493 153 7507 167
rect 6673 133 6687 147
rect 6713 133 6727 147
rect 6753 133 6767 147
rect 6853 133 6867 147
rect 7413 133 7427 147
rect 7473 133 7487 147
rect 7513 133 7527 147
rect 5073 113 5087 127
rect 5393 113 5407 127
rect 6273 113 6287 127
rect 6433 113 6447 127
rect 7833 1273 7847 1287
rect 7833 1193 7847 1207
rect 7893 1553 7907 1567
rect 7873 1313 7887 1327
rect 7873 1273 7887 1287
rect 7853 1173 7867 1187
rect 7853 1153 7867 1167
rect 7893 1193 7907 1207
rect 7893 1173 7907 1187
rect 7873 1133 7887 1147
rect 7853 1093 7867 1107
rect 7873 1073 7887 1087
rect 7853 933 7867 947
rect 7833 853 7847 867
rect 7873 813 7887 827
rect 7853 773 7867 787
rect 7833 693 7847 707
rect 7853 693 7867 707
rect 7813 673 7827 687
rect 7833 673 7847 687
rect 7773 633 7787 647
rect 7813 633 7827 647
rect 7873 653 7887 667
rect 7793 493 7807 507
rect 7833 353 7847 367
rect 7873 613 7887 627
rect 7873 593 7887 607
rect 7893 493 7907 507
rect 7893 353 7907 367
rect 7713 333 7727 347
rect 7753 333 7767 347
rect 7813 333 7827 347
rect 7853 333 7867 347
rect 7773 313 7787 327
rect 7913 293 7927 307
rect 7833 213 7847 227
rect 7653 173 7667 187
rect 7673 173 7687 187
rect 7613 153 7627 167
rect 7593 133 7607 147
rect 7633 133 7647 147
rect 7673 133 7687 147
rect 7733 133 7747 147
rect 7733 113 7747 127
rect 7853 133 7867 147
rect 7553 93 7567 107
rect 7753 93 7767 107
<< metal3 >>
rect 4807 6176 5193 6184
rect 5207 6176 5313 6184
rect 7427 6176 7733 6184
rect -24 6156 13 6164
rect 1687 6156 1793 6164
rect 2107 6156 2173 6164
rect 3307 6156 3473 6164
rect 3607 6156 3673 6164
rect 3727 6156 3813 6164
rect 3827 6156 3853 6164
rect 4867 6156 4993 6164
rect 5487 6156 5533 6164
rect 5627 6156 6113 6164
rect 6127 6156 6173 6164
rect 6287 6156 6393 6164
rect 6896 6156 7033 6164
rect 47 6136 213 6144
rect 227 6136 233 6144
rect 327 6136 393 6144
rect 407 6136 413 6144
rect 427 6136 493 6144
rect 507 6136 553 6144
rect 576 6136 653 6144
rect 576 6124 584 6136
rect 1427 6136 1473 6144
rect 1847 6136 2164 6144
rect 387 6116 584 6124
rect 607 6116 693 6124
rect 1756 6124 1764 6133
rect 2156 6127 2164 6136
rect 2907 6136 4053 6144
rect 4067 6136 4513 6144
rect 4907 6136 4953 6144
rect 5027 6136 5213 6144
rect 5227 6136 5273 6144
rect 6027 6136 6784 6144
rect 1056 6116 1304 6124
rect 1756 6116 1893 6124
rect 1056 6107 1064 6116
rect -24 6096 53 6104
rect 627 6096 873 6104
rect 1187 6096 1273 6104
rect 1296 6104 1304 6116
rect 2027 6116 2093 6124
rect 2247 6116 2393 6124
rect 2447 6116 2693 6124
rect 3707 6116 3733 6124
rect 4227 6116 4373 6124
rect 4507 6116 4553 6124
rect 4607 6116 4633 6124
rect 4707 6116 4773 6124
rect 4827 6116 4873 6124
rect 4987 6116 5033 6124
rect 5496 6124 5504 6133
rect 6776 6127 6784 6136
rect 6896 6144 6904 6156
rect 7567 6156 7653 6164
rect 6887 6136 6904 6144
rect 6927 6136 7093 6144
rect 7107 6136 7513 6144
rect 7527 6136 7693 6144
rect 5307 6116 5504 6124
rect 5927 6116 5973 6124
rect 6047 6116 6073 6124
rect 6207 6116 6273 6124
rect 6327 6116 6353 6124
rect 6407 6116 6453 6124
rect 6527 6116 6573 6124
rect 6587 6116 6633 6124
rect 6787 6116 6893 6124
rect 6907 6116 6993 6124
rect 7287 6116 7333 6124
rect 7387 6116 7433 6124
rect 7487 6116 7593 6124
rect 7607 6116 7613 6124
rect 7647 6116 7664 6124
rect 1296 6096 1393 6104
rect 1447 6096 1493 6104
rect 1547 6096 1613 6104
rect 1976 6104 1984 6113
rect 1627 6096 2293 6104
rect 2387 6096 2513 6104
rect 2567 6096 2733 6104
rect 3047 6096 3233 6104
rect 3776 6104 3784 6113
rect 3667 6096 3784 6104
rect 3807 6096 3973 6104
rect 4287 6096 4973 6104
rect 5047 6096 5673 6104
rect 5756 6104 5764 6113
rect 5687 6096 5764 6104
rect 5787 6096 6013 6104
rect 6147 6096 6233 6104
rect 6347 6096 6593 6104
rect 6607 6096 6613 6104
rect 6667 6096 7044 6104
rect 647 6076 673 6084
rect 687 6076 733 6084
rect 847 6076 1093 6084
rect 1347 6076 1453 6084
rect 1487 6076 1513 6084
rect 1847 6076 1913 6084
rect 2007 6076 2073 6084
rect 2087 6076 2113 6084
rect 2287 6076 2353 6084
rect 3007 6076 3113 6084
rect 3467 6076 3513 6084
rect 3947 6076 4193 6084
rect 4347 6076 4633 6084
rect 4647 6076 4673 6084
rect 4727 6076 4853 6084
rect 4867 6076 4933 6084
rect 5407 6076 5473 6084
rect 5647 6076 5673 6084
rect 5707 6076 5953 6084
rect 5967 6076 6053 6084
rect 6307 6076 6433 6084
rect 6507 6076 6733 6084
rect 6747 6076 6853 6084
rect 6867 6076 7013 6084
rect 7036 6084 7044 6096
rect 7156 6104 7164 6113
rect 7067 6096 7164 6104
rect 7656 6087 7664 6116
rect 7727 6116 7813 6124
rect 7856 6104 7864 6113
rect 7687 6096 7864 6104
rect 7036 6076 7273 6084
rect 7527 6076 7613 6084
rect 7707 6076 7833 6084
rect 107 6056 653 6064
rect 1467 6056 2033 6064
rect 2047 6056 2253 6064
rect 3287 6056 3933 6064
rect 4487 6056 4573 6064
rect 4627 6056 4893 6064
rect 4907 6056 4913 6064
rect 4967 6056 5313 6064
rect 5327 6056 5713 6064
rect 5727 6056 5733 6064
rect 6067 6056 6353 6064
rect 6367 6056 6413 6064
rect 6567 6056 7573 6064
rect 7587 6056 7713 6064
rect 1247 6036 1693 6044
rect 1707 6036 1813 6044
rect 2107 6036 2153 6044
rect 2407 6036 3753 6044
rect 4547 6036 5013 6044
rect 5187 6036 5333 6044
rect 5347 6036 5413 6044
rect 5647 6036 5793 6044
rect 5807 6036 5853 6044
rect 5887 6036 6513 6044
rect 6547 6036 6753 6044
rect 6827 6036 7253 6044
rect 7267 6036 7353 6044
rect 1567 6016 1733 6024
rect 1827 6016 2873 6024
rect 3347 6016 3373 6024
rect 4127 6016 4153 6024
rect 4267 6016 4493 6024
rect 4507 6016 4733 6024
rect 4827 6016 5093 6024
rect 5127 6016 5673 6024
rect 5827 6016 6033 6024
rect 6047 6016 6293 6024
rect 6687 6016 6873 6024
rect 1527 5996 1853 6004
rect 3107 5996 3513 6004
rect 3527 5996 3653 6004
rect 4587 5996 4753 6004
rect 5527 5996 5773 6004
rect 5887 5996 7173 6004
rect 7187 5996 7233 6004
rect 7247 5996 7453 6004
rect 167 5976 313 5984
rect 867 5976 1633 5984
rect 1807 5976 2233 5984
rect 2347 5976 3173 5984
rect 5427 5976 5693 5984
rect 5707 5976 5793 5984
rect 5847 5976 6513 5984
rect 6527 5976 6613 5984
rect 7027 5976 7053 5984
rect 7067 5976 7133 5984
rect 7227 5976 7533 5984
rect 7587 5976 7833 5984
rect 227 5956 253 5964
rect 667 5956 713 5964
rect 927 5956 1253 5964
rect 1367 5956 1513 5964
rect 1667 5956 1673 5964
rect 1687 5956 2013 5964
rect 2027 5956 2553 5964
rect 2987 5956 3233 5964
rect 4287 5956 4573 5964
rect 4587 5956 4953 5964
rect 5107 5956 5293 5964
rect 5307 5956 5373 5964
rect 5547 5956 6033 5964
rect 6087 5956 6133 5964
rect 7047 5956 7073 5964
rect 7407 5956 7673 5964
rect 7687 5956 7693 5964
rect 267 5936 293 5944
rect 307 5936 524 5944
rect 87 5916 113 5924
rect 127 5916 273 5924
rect 367 5916 493 5924
rect 516 5924 524 5936
rect 547 5936 793 5944
rect 1027 5936 1313 5944
rect 1427 5936 1453 5944
rect 1467 5936 1473 5944
rect 1707 5936 1853 5944
rect 2547 5936 2593 5944
rect 2607 5936 2933 5944
rect 3007 5936 3033 5944
rect 3167 5936 3353 5944
rect 3367 5936 3413 5944
rect 3507 5936 3604 5944
rect 516 5916 613 5924
rect 1496 5924 1504 5933
rect 3596 5927 3604 5936
rect 3687 5936 3813 5944
rect 4667 5936 4753 5944
rect 4867 5936 4993 5944
rect 5167 5936 5413 5944
rect 5667 5936 5813 5944
rect 5867 5936 5933 5944
rect 5947 5936 6093 5944
rect 6247 5936 6373 5944
rect 6427 5936 7113 5944
rect 7127 5936 7153 5944
rect 7716 5936 7873 5944
rect 1307 5916 1504 5924
rect 1727 5916 1833 5924
rect 2287 5916 2313 5924
rect 2367 5916 2413 5924
rect 2587 5916 2693 5924
rect 2927 5916 3013 5924
rect 3127 5916 3193 5924
rect 3247 5916 3473 5924
rect 3667 5916 3704 5924
rect 247 5896 333 5904
rect 387 5896 513 5904
rect 1127 5896 1153 5904
rect 1256 5887 1264 5913
rect 3696 5907 3704 5916
rect 3847 5916 3933 5924
rect 4167 5916 4213 5924
rect 4447 5916 4513 5924
rect 4687 5916 4773 5924
rect 4787 5916 4813 5924
rect 4967 5916 5073 5924
rect 5367 5916 5384 5924
rect 1467 5896 1573 5904
rect 2067 5896 2473 5904
rect 2527 5896 2873 5904
rect 3087 5896 3164 5904
rect 27 5876 73 5884
rect 587 5876 1053 5884
rect 1067 5876 1093 5884
rect 1276 5864 1284 5893
rect 1347 5876 1713 5884
rect 1907 5876 1973 5884
rect 2107 5876 2133 5884
rect 2187 5876 2253 5884
rect 2267 5876 2273 5884
rect 2507 5876 2593 5884
rect 2827 5876 2853 5884
rect 2907 5876 2913 5884
rect 2927 5876 3133 5884
rect 3156 5884 3164 5896
rect 3267 5896 3313 5904
rect 3367 5896 3393 5904
rect 3407 5896 3633 5904
rect 3647 5896 3673 5904
rect 4027 5896 4093 5904
rect 4276 5904 4284 5913
rect 4147 5896 4284 5904
rect 4647 5896 4713 5904
rect 4856 5904 4864 5913
rect 4747 5896 4864 5904
rect 3156 5876 3693 5884
rect 4287 5876 4293 5884
rect 4307 5876 4413 5884
rect 4767 5876 4893 5884
rect 5256 5884 5264 5913
rect 5287 5896 5333 5904
rect 5376 5904 5384 5916
rect 5407 5916 5473 5924
rect 5507 5916 5653 5924
rect 5747 5916 6024 5924
rect 5376 5896 5713 5904
rect 5767 5896 5913 5904
rect 5927 5896 5993 5904
rect 6016 5904 6024 5916
rect 6047 5916 6153 5924
rect 6347 5916 6533 5924
rect 6667 5916 7064 5924
rect 6016 5896 6233 5904
rect 6267 5896 6353 5904
rect 6547 5896 6593 5904
rect 6727 5896 6753 5904
rect 6776 5896 6973 5904
rect 5256 5876 5424 5884
rect 687 5856 1284 5864
rect 2467 5856 2513 5864
rect 3227 5856 3333 5864
rect 3587 5856 3853 5864
rect 4387 5856 4953 5864
rect 5416 5864 5424 5876
rect 5447 5876 5513 5884
rect 5627 5876 5673 5884
rect 5687 5876 5693 5884
rect 5727 5876 5813 5884
rect 5967 5876 6013 5884
rect 6027 5876 6133 5884
rect 6256 5884 6264 5893
rect 6187 5876 6264 5884
rect 6776 5884 6784 5896
rect 6987 5896 7033 5904
rect 7056 5904 7064 5916
rect 7147 5916 7193 5924
rect 7267 5916 7293 5924
rect 7327 5916 7364 5924
rect 7356 5907 7364 5916
rect 7387 5916 7413 5924
rect 7427 5916 7453 5924
rect 7607 5916 7633 5924
rect 7716 5907 7724 5936
rect 7747 5916 7793 5924
rect 7056 5896 7093 5904
rect 7107 5896 7173 5904
rect 7367 5896 7393 5904
rect 7427 5896 7513 5904
rect 7527 5896 7613 5904
rect 7667 5896 7713 5904
rect 6287 5876 6784 5884
rect 6796 5876 6813 5884
rect 5416 5856 6373 5864
rect 6796 5864 6804 5876
rect 6827 5876 6993 5884
rect 7276 5884 7284 5893
rect 7007 5876 7284 5884
rect 6567 5856 6804 5864
rect 7316 5864 7324 5893
rect 7447 5876 7573 5884
rect 7247 5856 7324 5864
rect 7567 5856 7773 5864
rect 2307 5836 2553 5844
rect 2567 5836 3093 5844
rect 3687 5836 3993 5844
rect 5587 5836 5613 5844
rect 6067 5836 6493 5844
rect 6507 5836 6593 5844
rect 6607 5836 6773 5844
rect 7047 5836 7253 5844
rect 6207 5816 6393 5824
rect 4027 5796 4053 5804
rect 4787 5796 5453 5804
rect 5787 5796 6233 5804
rect 6247 5796 6733 5804
rect 4047 5776 4053 5784
rect 5067 5776 6573 5784
rect 4607 5756 4633 5764
rect 4947 5756 5713 5764
rect 5187 5736 5213 5744
rect 5227 5736 5373 5744
rect 6147 5736 6333 5744
rect 1167 5716 2153 5724
rect 2167 5716 2393 5724
rect 2427 5716 3273 5724
rect 4427 5716 5033 5724
rect 5387 5716 5993 5724
rect 6007 5716 6313 5724
rect 6327 5716 6473 5724
rect 6487 5716 6633 5724
rect 7127 5716 7473 5724
rect 1727 5696 2093 5704
rect 2707 5696 3113 5704
rect 3167 5696 3293 5704
rect 4627 5696 5113 5704
rect 5127 5696 5413 5704
rect 7067 5696 7133 5704
rect 7196 5696 7333 5704
rect 207 5676 353 5684
rect 1347 5676 1393 5684
rect 1767 5676 2213 5684
rect 2227 5676 2373 5684
rect 2387 5676 2813 5684
rect 2827 5676 2993 5684
rect 3767 5676 4113 5684
rect 4127 5676 4193 5684
rect 4207 5676 4333 5684
rect 4347 5676 4553 5684
rect 4567 5676 4613 5684
rect 4987 5676 5253 5684
rect 5267 5676 5793 5684
rect 5827 5676 6073 5684
rect 6087 5676 6213 5684
rect 6387 5676 6653 5684
rect 6667 5676 6693 5684
rect 6707 5676 6713 5684
rect 7047 5676 7153 5684
rect 67 5656 113 5664
rect 127 5656 133 5664
rect 307 5656 333 5664
rect 1007 5656 1193 5664
rect 1207 5656 1213 5664
rect 1327 5656 1373 5664
rect 2027 5656 2053 5664
rect 2667 5656 2753 5664
rect 2847 5656 2913 5664
rect 2967 5656 3053 5664
rect 3076 5656 3133 5664
rect 67 5636 173 5644
rect 307 5636 393 5644
rect 687 5636 713 5644
rect 1087 5636 1224 5644
rect 427 5616 553 5624
rect 707 5616 733 5624
rect 867 5616 1053 5624
rect 1107 5616 1193 5624
rect 1216 5624 1224 5636
rect 1387 5636 1533 5644
rect 1607 5636 1613 5644
rect 1627 5636 2033 5644
rect 2327 5636 2433 5644
rect 2627 5636 2773 5644
rect 2796 5644 2804 5653
rect 2796 5636 2933 5644
rect 3027 5636 3033 5644
rect 3076 5644 3084 5656
rect 3147 5656 3193 5664
rect 3247 5656 3353 5664
rect 3667 5656 3693 5664
rect 4067 5656 4213 5664
rect 4707 5656 4773 5664
rect 4967 5656 5013 5664
rect 5047 5656 5093 5664
rect 5127 5656 5144 5664
rect 3047 5636 3084 5644
rect 3107 5636 3113 5644
rect 3127 5636 3433 5644
rect 3647 5636 3713 5644
rect 4007 5636 4033 5644
rect 4047 5636 4073 5644
rect 4207 5636 4273 5644
rect 4287 5636 4293 5644
rect 4336 5636 4513 5644
rect 1216 5616 1413 5624
rect 1747 5616 1853 5624
rect 1927 5616 2113 5624
rect 2407 5616 2513 5624
rect 2527 5616 2853 5624
rect 3307 5616 3493 5624
rect 3747 5616 3873 5624
rect 4336 5624 4344 5636
rect 4567 5636 4713 5644
rect 4727 5636 4873 5644
rect 4927 5636 5053 5644
rect 5136 5644 5144 5656
rect 5167 5656 5673 5664
rect 5687 5656 5753 5664
rect 5856 5656 5873 5664
rect 5136 5636 5164 5644
rect 4327 5616 4344 5624
rect 4367 5616 4753 5624
rect 4807 5616 4833 5624
rect 4907 5616 4973 5624
rect 5156 5624 5164 5636
rect 5187 5636 5233 5644
rect 5327 5636 5444 5644
rect 5156 5616 5293 5624
rect 5316 5616 5393 5624
rect 327 5596 553 5604
rect 676 5604 684 5613
rect 567 5596 684 5604
rect 967 5596 1593 5604
rect 1987 5596 2273 5604
rect 2287 5596 2333 5604
rect 2607 5596 2713 5604
rect 2827 5596 2893 5604
rect 2907 5596 2993 5604
rect 3267 5596 3433 5604
rect 3707 5596 3773 5604
rect 3927 5596 4393 5604
rect 4407 5596 4644 5604
rect 607 5576 793 5584
rect 807 5576 813 5584
rect 1067 5576 1513 5584
rect 1907 5576 1913 5584
rect 1927 5576 1993 5584
rect 2247 5576 2393 5584
rect 2487 5576 2833 5584
rect 2847 5576 2873 5584
rect 3227 5576 3233 5584
rect 3247 5576 3313 5584
rect 4447 5576 4473 5584
rect 4547 5576 4593 5584
rect 4636 5584 4644 5596
rect 4667 5596 4733 5604
rect 4767 5596 4844 5604
rect 4636 5576 4653 5584
rect 4667 5576 4673 5584
rect 4747 5576 4813 5584
rect 4836 5584 4844 5596
rect 5316 5604 5324 5616
rect 5436 5624 5444 5636
rect 5467 5636 5573 5644
rect 5667 5636 5693 5644
rect 5747 5636 5833 5644
rect 5856 5627 5864 5656
rect 5896 5656 6013 5664
rect 5896 5644 5904 5656
rect 6027 5656 6193 5664
rect 6247 5656 6413 5664
rect 6467 5656 6853 5664
rect 6967 5656 6993 5664
rect 7016 5664 7024 5673
rect 7196 5667 7204 5696
rect 7267 5676 7413 5684
rect 7427 5676 7553 5684
rect 7016 5656 7084 5664
rect 5887 5636 5904 5644
rect 5947 5636 5973 5644
rect 5987 5636 6053 5644
rect 6447 5636 6513 5644
rect 6947 5636 7004 5644
rect 5436 5616 5593 5624
rect 6096 5624 6104 5633
rect 6096 5616 6233 5624
rect 6607 5616 6673 5624
rect 6747 5616 6773 5624
rect 6787 5616 6833 5624
rect 6996 5624 7004 5636
rect 7027 5636 7053 5644
rect 7076 5644 7084 5656
rect 7107 5656 7193 5664
rect 7247 5656 7284 5664
rect 7076 5636 7113 5644
rect 7127 5636 7213 5644
rect 7276 5644 7284 5656
rect 7307 5656 7373 5664
rect 7587 5656 7693 5664
rect 7707 5656 7853 5664
rect 7276 5636 7293 5644
rect 7387 5636 7453 5644
rect 7647 5636 7733 5644
rect 7756 5636 7793 5644
rect 6996 5616 7133 5624
rect 7147 5616 7173 5624
rect 7536 5624 7544 5633
rect 7447 5616 7613 5624
rect 7756 5624 7764 5636
rect 7687 5616 7764 5624
rect 4907 5596 5324 5604
rect 5347 5596 5473 5604
rect 5567 5596 5953 5604
rect 6007 5596 6033 5604
rect 6587 5596 6613 5604
rect 6627 5596 6793 5604
rect 6947 5596 7253 5604
rect 7267 5596 7273 5604
rect 7347 5596 7393 5604
rect 7707 5596 7773 5604
rect 4836 5576 4933 5584
rect 4967 5576 5013 5584
rect 5087 5576 5333 5584
rect 5407 5576 5513 5584
rect 5527 5576 5533 5584
rect 5767 5576 5773 5584
rect 5787 5576 5833 5584
rect 5847 5576 5913 5584
rect 6307 5576 6913 5584
rect 6927 5576 6973 5584
rect 6987 5576 7073 5584
rect 7367 5576 7493 5584
rect 7507 5576 7753 5584
rect 7767 5576 7773 5584
rect 867 5556 1273 5564
rect 1287 5556 1313 5564
rect 1487 5556 1573 5564
rect 1587 5556 1673 5564
rect 1907 5556 2013 5564
rect 2027 5556 2313 5564
rect 3127 5556 3353 5564
rect 4847 5556 4993 5564
rect 5067 5556 5153 5564
rect 5327 5556 5373 5564
rect 5447 5556 5733 5564
rect 5887 5556 6693 5564
rect 387 5536 433 5544
rect 627 5536 953 5544
rect 1047 5536 1913 5544
rect 2167 5536 2573 5544
rect 3187 5536 3293 5544
rect 4407 5536 4453 5544
rect 4467 5536 4573 5544
rect 4587 5536 4853 5544
rect 4967 5536 5073 5544
rect 5147 5536 5213 5544
rect 5747 5536 6173 5544
rect 7307 5536 7533 5544
rect 807 5516 1453 5524
rect 1467 5516 1553 5524
rect 1967 5516 2193 5524
rect 2207 5516 2233 5524
rect 2987 5516 3073 5524
rect 4527 5516 4693 5524
rect 4727 5516 4793 5524
rect 4827 5516 4913 5524
rect 4927 5516 4973 5524
rect 4987 5516 6253 5524
rect 6836 5516 7793 5524
rect 727 5496 1293 5504
rect 4267 5496 4853 5504
rect 4867 5496 5293 5504
rect 6836 5504 6844 5516
rect 7807 5516 7833 5524
rect 5347 5496 6844 5504
rect 7007 5496 7113 5504
rect 7127 5496 7173 5504
rect 7267 5496 7473 5504
rect 47 5476 93 5484
rect 147 5476 273 5484
rect 287 5476 513 5484
rect 527 5476 693 5484
rect 907 5476 1353 5484
rect 1687 5476 1713 5484
rect 1727 5476 1753 5484
rect 1876 5476 1973 5484
rect 107 5456 324 5464
rect 316 5447 324 5456
rect 607 5456 693 5464
rect 707 5456 733 5464
rect 767 5456 873 5464
rect 1027 5456 1473 5464
rect 1556 5456 1693 5464
rect 1556 5447 1564 5456
rect 1876 5464 1884 5476
rect 2087 5476 2473 5484
rect 2927 5476 2933 5484
rect 2947 5476 3253 5484
rect 3267 5476 3453 5484
rect 3467 5476 3493 5484
rect 3507 5476 3513 5484
rect 3527 5476 3933 5484
rect 3947 5476 4153 5484
rect 4367 5476 4873 5484
rect 4887 5476 5173 5484
rect 5187 5476 5193 5484
rect 5567 5476 5933 5484
rect 5947 5476 6053 5484
rect 6067 5476 6073 5484
rect 6887 5476 6953 5484
rect 7327 5476 7493 5484
rect 7607 5476 7753 5484
rect 1707 5456 1884 5464
rect 2127 5456 2173 5464
rect 2187 5456 2213 5464
rect 2327 5456 2433 5464
rect 2547 5456 2773 5464
rect 2787 5456 2953 5464
rect 3016 5456 3073 5464
rect 3016 5447 3024 5456
rect 3607 5456 3673 5464
rect 3887 5456 4173 5464
rect 4187 5456 4273 5464
rect 4287 5456 4353 5464
rect 4387 5456 4433 5464
rect 4467 5456 4493 5464
rect 4547 5456 4893 5464
rect 5667 5456 5693 5464
rect 5727 5456 6473 5464
rect 6487 5456 6553 5464
rect 6867 5456 6993 5464
rect 7167 5456 7313 5464
rect 7487 5456 7513 5464
rect 7527 5456 7613 5464
rect 7787 5456 7833 5464
rect 367 5436 393 5444
rect 447 5436 473 5444
rect 487 5436 573 5444
rect 907 5436 933 5444
rect 1327 5436 1493 5444
rect 1576 5436 1633 5444
rect -24 5416 173 5424
rect 687 5416 993 5424
rect 1207 5416 1253 5424
rect 1307 5416 1373 5424
rect 1576 5424 1584 5436
rect 1656 5436 1853 5444
rect 1467 5416 1584 5424
rect 1656 5424 1664 5436
rect 2507 5436 2664 5444
rect 1627 5416 1664 5424
rect 1787 5416 1833 5424
rect 1887 5416 1933 5424
rect 2007 5416 2093 5424
rect 2187 5416 2293 5424
rect 2387 5416 2413 5424
rect 2467 5416 2473 5424
rect 2487 5416 2633 5424
rect 2656 5424 2664 5436
rect 2767 5436 2793 5444
rect 2827 5436 2893 5444
rect 3227 5436 3733 5444
rect 3756 5436 3833 5444
rect 3756 5427 3764 5436
rect 3847 5436 4513 5444
rect 4587 5436 4673 5444
rect 4767 5436 4953 5444
rect 4996 5436 5033 5444
rect 2656 5416 3093 5424
rect 3587 5416 3713 5424
rect 3987 5416 4253 5424
rect 4327 5416 4384 5424
rect 1227 5396 1673 5404
rect 1687 5396 1793 5404
rect 2147 5396 2333 5404
rect 2347 5396 2353 5404
rect 2367 5396 2493 5404
rect 2567 5396 2573 5404
rect 2587 5396 3033 5404
rect 3347 5396 3853 5404
rect 3867 5396 3873 5404
rect 3947 5396 4053 5404
rect 4376 5387 4384 5416
rect 4536 5424 4544 5433
rect 4507 5416 4544 5424
rect 4996 5424 5004 5436
rect 5087 5436 5113 5444
rect 5267 5436 5313 5444
rect 5387 5436 5473 5444
rect 5527 5436 5624 5444
rect 4667 5416 4864 5424
rect 4527 5396 4553 5404
rect 4636 5404 4644 5413
rect 4856 5407 4864 5416
rect 4936 5416 5004 5424
rect 4587 5396 4644 5404
rect 4667 5396 4713 5404
rect 4936 5387 4944 5416
rect 5027 5416 5113 5424
rect 5227 5416 5353 5424
rect 5447 5416 5573 5424
rect 5587 5416 5593 5424
rect 5616 5424 5624 5436
rect 5647 5436 5673 5444
rect 5687 5436 5813 5444
rect 6387 5436 6413 5444
rect 6447 5436 6513 5444
rect 6527 5436 6633 5444
rect 6687 5436 6753 5444
rect 6827 5436 6884 5444
rect 5616 5416 5693 5424
rect 5807 5416 5893 5424
rect 5907 5416 5973 5424
rect 5987 5416 6033 5424
rect 6227 5416 6553 5424
rect 6607 5416 6793 5424
rect 6876 5424 6884 5436
rect 6907 5436 7013 5444
rect 7067 5436 7193 5444
rect 7287 5436 7353 5444
rect 7407 5436 7573 5444
rect 7587 5436 7713 5444
rect 7807 5436 7864 5444
rect 7856 5427 7864 5436
rect 7887 5436 7913 5444
rect 6876 5416 7033 5424
rect 7087 5416 7284 5424
rect 4987 5396 5033 5404
rect 5107 5396 5153 5404
rect 5247 5396 5293 5404
rect 5527 5396 5633 5404
rect 5647 5396 5773 5404
rect 5967 5396 6073 5404
rect 6547 5396 6593 5404
rect 6627 5396 6693 5404
rect 6927 5396 6973 5404
rect 7027 5396 7093 5404
rect 7276 5404 7284 5416
rect 7307 5416 7333 5424
rect 7356 5416 7433 5424
rect 7356 5407 7364 5416
rect 7547 5416 7633 5424
rect 7767 5416 7813 5424
rect 7276 5396 7333 5404
rect 7387 5396 7444 5404
rect 187 5376 1293 5384
rect 1667 5376 1773 5384
rect 1787 5376 2973 5384
rect 4007 5376 4033 5384
rect 4427 5376 4553 5384
rect 5147 5376 5253 5384
rect 5427 5376 5713 5384
rect 5747 5376 5813 5384
rect 7147 5376 7413 5384
rect 7436 5384 7444 5396
rect 7467 5396 7633 5404
rect 7656 5396 7773 5404
rect 7656 5384 7664 5396
rect 7436 5376 7664 5384
rect 627 5356 1813 5364
rect 1847 5356 1913 5364
rect 3987 5356 4333 5364
rect 4627 5356 4653 5364
rect 5247 5356 5393 5364
rect 5667 5356 5853 5364
rect 2047 5336 2633 5344
rect 2687 5336 2733 5344
rect 2747 5336 2933 5344
rect 2947 5336 3153 5344
rect 4267 5336 4453 5344
rect 4467 5336 4573 5344
rect 4867 5336 5113 5344
rect 5267 5336 6233 5344
rect 6247 5336 6293 5344
rect 4147 5316 4213 5324
rect 4247 5316 4333 5324
rect 4487 5316 5153 5324
rect 5727 5316 5893 5324
rect 4307 5296 4493 5304
rect 4507 5296 4673 5304
rect 4707 5296 6193 5304
rect 6207 5296 6273 5304
rect 4847 5276 6393 5284
rect 327 5256 413 5264
rect 4627 5256 5033 5264
rect 5047 5256 5073 5264
rect 5127 5256 5333 5264
rect 5367 5256 5913 5264
rect 2047 5236 2073 5244
rect 2087 5236 3613 5244
rect 4487 5236 4773 5244
rect 4787 5236 4933 5244
rect 4987 5236 5473 5244
rect 5707 5236 5733 5244
rect 5767 5236 5813 5244
rect 6967 5236 6993 5244
rect 7287 5236 7593 5244
rect 4427 5216 5253 5224
rect 5267 5216 5273 5224
rect 5407 5216 5533 5224
rect 5547 5216 5573 5224
rect 5847 5216 6293 5224
rect 6347 5216 6733 5224
rect 6867 5216 6953 5224
rect 7267 5216 7373 5224
rect 7427 5216 7473 5224
rect 2267 5196 2873 5204
rect 3327 5196 3393 5204
rect 4567 5196 4593 5204
rect 4607 5196 4713 5204
rect 4727 5196 5313 5204
rect 5327 5196 5453 5204
rect 5787 5196 5953 5204
rect 6007 5196 6193 5204
rect 6207 5196 6333 5204
rect 6347 5196 6433 5204
rect 6967 5196 7044 5204
rect 7036 5187 7044 5196
rect 7087 5196 7453 5204
rect 7567 5196 7713 5204
rect 2687 5176 2913 5184
rect 2967 5176 3133 5184
rect 3187 5176 3353 5184
rect 3627 5176 3673 5184
rect 3687 5176 4113 5184
rect 4527 5176 4613 5184
rect 4747 5176 4953 5184
rect 5067 5176 5273 5184
rect 5347 5176 5393 5184
rect 5427 5176 5473 5184
rect 5807 5176 5913 5184
rect 6127 5176 6164 5184
rect 267 5156 473 5164
rect 487 5156 753 5164
rect 867 5156 913 5164
rect 2167 5156 2213 5164
rect 2307 5156 2333 5164
rect 2356 5156 2373 5164
rect 287 5136 353 5144
rect 747 5136 913 5144
rect 1047 5136 1253 5144
rect 1507 5136 1553 5144
rect 2356 5144 2364 5156
rect 2387 5156 2433 5164
rect 2487 5156 2624 5164
rect 2616 5147 2624 5156
rect 2807 5156 2833 5164
rect 2947 5156 3064 5164
rect 3056 5147 3064 5156
rect 3387 5156 3573 5164
rect 3707 5156 3793 5164
rect 3847 5156 3893 5164
rect 3947 5156 4073 5164
rect 4167 5156 4253 5164
rect 2327 5136 2364 5144
rect 2827 5136 2853 5144
rect 3227 5136 3273 5144
rect 3307 5136 3353 5144
rect 3487 5136 3673 5144
rect 3827 5136 3953 5144
rect 4087 5136 4193 5144
rect 4327 5136 4353 5144
rect 4476 5144 4484 5173
rect 4576 5156 4733 5164
rect 4576 5147 4584 5156
rect 4747 5156 4773 5164
rect 4467 5136 4484 5144
rect 4647 5136 4653 5144
rect 4996 5144 5004 5173
rect 5107 5156 5193 5164
rect 5307 5156 5353 5164
rect 5496 5164 5504 5173
rect 5396 5156 5504 5164
rect 5576 5156 5673 5164
rect 4667 5136 5024 5144
rect 156 5124 164 5133
rect 5016 5127 5024 5136
rect 5187 5136 5233 5144
rect 5396 5144 5404 5156
rect 5387 5136 5404 5144
rect 5576 5144 5584 5156
rect 5787 5156 5953 5164
rect 6087 5156 6133 5164
rect 5427 5136 5584 5144
rect 5607 5136 5793 5144
rect 6076 5144 6084 5153
rect 5987 5136 6084 5144
rect 6107 5136 6113 5144
rect 6156 5144 6164 5176
rect 6287 5176 6313 5184
rect 6527 5176 6624 5184
rect 6616 5167 6624 5176
rect 6747 5176 6853 5184
rect 7007 5176 7024 5184
rect 7016 5167 7024 5176
rect 7127 5176 7153 5184
rect 7227 5176 7253 5184
rect 7267 5176 7493 5184
rect 7547 5176 7753 5184
rect 7767 5176 7773 5184
rect 6187 5156 6233 5164
rect 6267 5156 6293 5164
rect 6387 5156 6493 5164
rect 7096 5156 7273 5164
rect 6127 5136 6164 5144
rect 6576 5144 6584 5153
rect 6407 5136 6584 5144
rect 6607 5136 6933 5144
rect 7096 5144 7104 5156
rect 7387 5156 7404 5164
rect 6987 5136 7104 5144
rect 7127 5136 7233 5144
rect 7396 5144 7404 5156
rect 7427 5156 7473 5164
rect 7576 5156 7593 5164
rect 7576 5147 7584 5156
rect 7867 5156 7893 5164
rect 7396 5136 7513 5144
rect 7747 5136 7793 5144
rect 7887 5136 7913 5144
rect 156 5116 373 5124
rect 387 5116 393 5124
rect 787 5116 813 5124
rect 827 5116 993 5124
rect 1007 5116 1153 5124
rect 1167 5116 1333 5124
rect 2027 5116 2133 5124
rect 2367 5116 2413 5124
rect 2427 5116 2813 5124
rect 2827 5116 3013 5124
rect 3207 5116 3513 5124
rect 3527 5116 3993 5124
rect 4107 5116 4273 5124
rect 4767 5116 4953 5124
rect 5227 5116 5293 5124
rect 5507 5116 5513 5124
rect 5527 5116 5613 5124
rect 5707 5116 5813 5124
rect 5827 5116 5933 5124
rect 5967 5116 6033 5124
rect 6307 5116 6353 5124
rect 6367 5116 6473 5124
rect 6627 5116 6713 5124
rect 6727 5116 6833 5124
rect 7067 5116 7173 5124
rect 7407 5116 7493 5124
rect 7527 5116 7633 5124
rect 7787 5116 7873 5124
rect 987 5096 1213 5104
rect 1227 5096 1373 5104
rect 2347 5096 2353 5104
rect 2367 5096 2453 5104
rect 2467 5096 2953 5104
rect 2967 5096 3233 5104
rect 4227 5096 4393 5104
rect 4407 5096 4493 5104
rect 4687 5096 4993 5104
rect 6047 5096 6493 5104
rect 7147 5096 7213 5104
rect 7447 5096 7613 5104
rect 7787 5096 7813 5104
rect 1307 5076 1853 5084
rect 1867 5076 3273 5084
rect 4887 5076 5153 5084
rect 6167 5076 6673 5084
rect 6687 5076 6873 5084
rect 7707 5076 7733 5084
rect 7747 5076 7853 5084
rect 1707 5056 3453 5064
rect 3987 5056 4053 5064
rect 4447 5056 4533 5064
rect 4547 5056 4893 5064
rect 4987 5056 5233 5064
rect 5567 5056 5733 5064
rect 5747 5056 5793 5064
rect 6427 5056 6493 5064
rect 6687 5056 6773 5064
rect 1347 5036 1413 5044
rect 1807 5036 2473 5044
rect 4347 5036 4473 5044
rect 4707 5036 4913 5044
rect 4927 5036 5653 5044
rect 6067 5036 6633 5044
rect 6647 5036 6713 5044
rect 1807 5016 1993 5024
rect 2007 5016 2513 5024
rect 2527 5016 2613 5024
rect 4467 5016 4813 5024
rect 4967 5016 5073 5024
rect 5407 5016 7273 5024
rect 7287 5016 7413 5024
rect 7547 5016 7593 5024
rect 1967 4996 2153 5004
rect 2207 4996 2293 5004
rect 4387 4996 5033 5004
rect 5047 4996 5173 5004
rect 5227 4996 5413 5004
rect 5727 4996 5753 5004
rect 5867 4996 6213 5004
rect 6227 4996 6373 5004
rect 6387 4996 6413 5004
rect 6767 4996 6893 5004
rect 6947 4996 7093 5004
rect 7467 4996 7484 5004
rect 167 4976 384 4984
rect 376 4967 384 4976
rect 1607 4976 1793 4984
rect 2127 4976 2333 4984
rect 2647 4976 2713 4984
rect 2787 4976 2833 4984
rect 2907 4976 3233 4984
rect 3267 4976 3433 4984
rect 3627 4976 3653 4984
rect 3747 4976 3773 4984
rect 4027 4976 4204 4984
rect 67 4956 253 4964
rect 867 4956 953 4964
rect 1027 4956 1053 4964
rect 1387 4956 1453 4964
rect 1507 4956 1573 4964
rect 1647 4956 1873 4964
rect 1916 4964 1924 4973
rect 1887 4956 1924 4964
rect 2207 4956 2233 4964
rect 2707 4956 2793 4964
rect 2867 4956 2893 4964
rect 3087 4956 3393 4964
rect 3567 4956 3633 4964
rect 3647 4956 3704 4964
rect 87 4936 133 4944
rect 487 4936 593 4944
rect 947 4936 1653 4944
rect 1667 4936 1773 4944
rect 2047 4936 2133 4944
rect 2387 4936 2413 4944
rect 3467 4936 3533 4944
rect 3627 4936 3653 4944
rect 3696 4944 3704 4956
rect 3727 4956 3813 4964
rect 3847 4956 3873 4964
rect 3927 4956 4113 4964
rect 4196 4964 4204 4976
rect 4547 4976 4773 4984
rect 4787 4976 4813 4984
rect 4827 4976 5053 4984
rect 5067 4976 5113 4984
rect 5927 4976 5993 4984
rect 6007 4976 6253 4984
rect 6327 4976 6613 4984
rect 6627 4976 6753 4984
rect 6807 4976 7113 4984
rect 7127 4976 7153 4984
rect 7267 4976 7353 4984
rect 7407 4976 7453 4984
rect 4196 4956 4233 4964
rect 4427 4956 4553 4964
rect 4687 4956 4793 4964
rect 4867 4956 4924 4964
rect 3696 4936 3793 4944
rect 3947 4936 3993 4944
rect 4347 4936 4393 4944
rect 4447 4936 4733 4944
rect 4836 4944 4844 4953
rect 4916 4947 4924 4956
rect 4947 4956 4984 4964
rect 4976 4947 4984 4956
rect 5167 4956 5293 4964
rect 5307 4956 5353 4964
rect 5627 4956 5713 4964
rect 5767 4956 6013 4964
rect 6107 4956 6133 4964
rect 6176 4956 6453 4964
rect 4767 4936 4844 4944
rect 4927 4936 4933 4944
rect 4996 4927 5004 4953
rect 5247 4936 5373 4944
rect 5507 4936 5604 4944
rect 5596 4927 5604 4936
rect 5667 4936 5833 4944
rect 5987 4936 6053 4944
rect 6176 4944 6184 4956
rect 6567 4956 6593 4964
rect 6607 4956 6784 4964
rect 6776 4947 6784 4956
rect 6907 4956 7064 4964
rect 6067 4936 6184 4944
rect 6207 4936 6273 4944
rect 6287 4936 6353 4944
rect 6407 4936 6453 4944
rect 6567 4936 6693 4944
rect 6887 4936 6913 4944
rect 6987 4936 7013 4944
rect 7056 4944 7064 4956
rect 7087 4956 7133 4964
rect 7207 4956 7373 4964
rect 7427 4956 7464 4964
rect 7456 4947 7464 4956
rect 7056 4936 7093 4944
rect 7107 4936 7173 4944
rect 7387 4936 7433 4944
rect 387 4916 2073 4924
rect 2687 4916 2953 4924
rect 3907 4916 3933 4924
rect 4247 4916 4313 4924
rect 4747 4916 4893 4924
rect 5016 4916 5053 4924
rect 1367 4896 2873 4904
rect 3107 4896 3153 4904
rect 5016 4904 5024 4916
rect 5127 4916 5313 4924
rect 5327 4916 5393 4924
rect 5767 4916 5793 4924
rect 5876 4924 5884 4933
rect 7476 4927 7484 4996
rect 7687 4996 7893 5004
rect 7567 4976 7633 4984
rect 7707 4976 7813 4984
rect 7547 4956 7713 4964
rect 7836 4964 7844 4973
rect 7776 4956 7844 4964
rect 7496 4927 7504 4953
rect 7587 4936 7613 4944
rect 5827 4916 5884 4924
rect 6367 4916 6433 4924
rect 6667 4916 6853 4924
rect 6867 4916 6953 4924
rect 7176 4916 7393 4924
rect 4747 4896 5024 4904
rect 5087 4896 5213 4904
rect 5727 4896 5933 4904
rect 6047 4896 6153 4904
rect 7176 4904 7184 4916
rect 7407 4916 7464 4924
rect 6907 4896 7184 4904
rect 7456 4904 7464 4916
rect 7776 4924 7784 4956
rect 7807 4936 7833 4944
rect 7776 4916 7813 4924
rect 7456 4896 7564 4904
rect 1227 4876 1373 4884
rect 2027 4876 2493 4884
rect 3427 4876 4173 4884
rect 4987 4876 5273 4884
rect 5567 4876 5813 4884
rect 6587 4876 6613 4884
rect 7027 4876 7233 4884
rect 7387 4876 7513 4884
rect 7556 4884 7564 4896
rect 7556 4876 7593 4884
rect 7607 4876 7753 4884
rect 827 4856 3073 4864
rect 3847 4856 3913 4864
rect 4807 4856 5513 4864
rect 5527 4856 5653 4864
rect 5667 4856 5673 4864
rect 5807 4856 5833 4864
rect 6827 4856 7033 4864
rect 7367 4856 7453 4864
rect 7467 4856 7553 4864
rect 667 4836 1073 4844
rect 1087 4836 1573 4844
rect 3227 4836 3333 4844
rect 5107 4836 6533 4844
rect 6547 4836 6573 4844
rect 7287 4836 7513 4844
rect 1507 4816 2093 4824
rect 3547 4816 3713 4824
rect 3727 4816 3753 4824
rect 5267 4816 5853 4824
rect 5867 4816 5953 4824
rect 627 4796 1533 4804
rect 2707 4796 3173 4804
rect 3847 4796 3853 4804
rect 5147 4796 5273 4804
rect 247 4776 553 4784
rect 567 4776 1033 4784
rect 1347 4776 2313 4784
rect 3307 4776 3953 4784
rect 5207 4776 5233 4784
rect 5327 4776 5893 4784
rect 5907 4776 5913 4784
rect 967 4756 2393 4764
rect 3747 4756 3813 4764
rect 4367 4756 4693 4764
rect 5167 4756 5433 4764
rect 5447 4756 6613 4764
rect 7767 4756 7913 4764
rect 1036 4736 1133 4744
rect 1036 4724 1044 4736
rect 1207 4736 1233 4744
rect 1247 4736 1953 4744
rect 1967 4736 2373 4744
rect 4307 4736 4953 4744
rect 4967 4736 5253 4744
rect 5467 4736 5633 4744
rect 5647 4736 5713 4744
rect 5727 4736 5733 4744
rect 6307 4736 6413 4744
rect 6447 4736 6493 4744
rect 6927 4736 7273 4744
rect 7547 4736 7633 4744
rect 7747 4736 7773 4744
rect 996 4716 1044 4724
rect 807 4676 873 4684
rect 996 4684 1004 4716
rect 1067 4716 1213 4724
rect 1927 4716 1933 4724
rect 1947 4716 2173 4724
rect 2287 4716 2493 4724
rect 2947 4716 3193 4724
rect 3207 4716 3313 4724
rect 3807 4716 3873 4724
rect 3887 4716 3973 4724
rect 3987 4716 4013 4724
rect 4027 4716 4133 4724
rect 4567 4716 4673 4724
rect 4687 4716 5433 4724
rect 5487 4716 5604 4724
rect 5596 4707 5604 4716
rect 6007 4716 6173 4724
rect 6347 4716 6453 4724
rect 6487 4716 6504 4724
rect 6496 4707 6504 4716
rect 7096 4716 7133 4724
rect 7096 4707 7104 4716
rect 7227 4716 7293 4724
rect 7547 4716 7593 4724
rect 7687 4716 7853 4724
rect 1107 4696 1124 4704
rect 987 4676 1004 4684
rect 227 4656 253 4664
rect 467 4656 493 4664
rect 707 4656 753 4664
rect 956 4664 964 4673
rect 1116 4667 1124 4696
rect 1447 4696 1493 4704
rect 2047 4696 2133 4704
rect 2287 4696 2313 4704
rect 2607 4696 2624 4704
rect 1407 4676 1493 4684
rect 1516 4676 1713 4684
rect 907 4656 964 4664
rect 1516 4664 1524 4676
rect 1327 4656 1524 4664
rect 1647 4656 1693 4664
rect 1767 4656 1813 4664
rect 1827 4656 1853 4664
rect 1907 4656 1993 4664
rect 2196 4664 2204 4693
rect 2267 4676 2293 4684
rect 2347 4676 2433 4684
rect 2447 4676 2593 4684
rect 2616 4684 2624 4696
rect 2907 4696 2953 4704
rect 3187 4696 3213 4704
rect 3447 4696 3573 4704
rect 3987 4696 4073 4704
rect 4107 4696 4153 4704
rect 4167 4696 4233 4704
rect 5027 4696 5053 4704
rect 5207 4696 5233 4704
rect 5287 4696 5453 4704
rect 5467 4696 5473 4704
rect 5647 4696 6033 4704
rect 6087 4696 6264 4704
rect 2616 4676 2724 4684
rect 2196 4656 2353 4664
rect 2667 4656 2693 4664
rect 2716 4664 2724 4676
rect 2767 4676 3273 4684
rect 3327 4676 3413 4684
rect 3527 4676 3613 4684
rect 3807 4676 3993 4684
rect 4267 4676 4313 4684
rect 4467 4676 4693 4684
rect 4767 4676 4833 4684
rect 4956 4684 4964 4693
rect 4887 4676 4964 4684
rect 5276 4684 5284 4693
rect 5207 4676 5284 4684
rect 5307 4676 5413 4684
rect 5507 4676 5553 4684
rect 5567 4676 5613 4684
rect 5947 4676 5993 4684
rect 6007 4676 6013 4684
rect 6067 4676 6133 4684
rect 6256 4684 6264 4696
rect 6327 4696 6493 4704
rect 7327 4696 7393 4704
rect 7447 4696 7473 4704
rect 7587 4696 7673 4704
rect 7687 4696 7713 4704
rect 7756 4696 7813 4704
rect 6256 4676 6273 4684
rect 6287 4676 6333 4684
rect 6387 4676 6473 4684
rect 2716 4656 2753 4664
rect 3087 4656 3293 4664
rect 3307 4656 3313 4664
rect 3756 4664 3764 4673
rect 6576 4667 6584 4693
rect 6607 4676 6733 4684
rect 6867 4676 6933 4684
rect 7007 4676 7073 4684
rect 7087 4676 7173 4684
rect 7347 4676 7364 4684
rect 3647 4656 3764 4664
rect 4347 4656 4473 4664
rect 4527 4656 4613 4664
rect 4827 4656 4893 4664
rect 4947 4656 5173 4664
rect 5227 4656 5273 4664
rect 5447 4656 5533 4664
rect 5547 4656 5673 4664
rect 5747 4656 5833 4664
rect 6247 4656 6313 4664
rect 6327 4656 6364 4664
rect 6356 4647 6364 4656
rect 6467 4656 6513 4664
rect 6767 4656 6813 4664
rect 6967 4656 7013 4664
rect 7356 4647 7364 4676
rect 7387 4676 7504 4684
rect 7387 4656 7473 4664
rect 7496 4664 7504 4676
rect 7647 4676 7733 4684
rect 7496 4656 7573 4664
rect 7596 4664 7604 4673
rect 7596 4656 7693 4664
rect 7756 4664 7764 4696
rect 7727 4656 7764 4664
rect 147 4636 273 4644
rect 287 4636 373 4644
rect 387 4636 593 4644
rect 847 4636 873 4644
rect 887 4636 953 4644
rect 1027 4636 1253 4644
rect 1527 4636 1673 4644
rect 1747 4636 1773 4644
rect 2127 4636 2213 4644
rect 2327 4636 2413 4644
rect 2727 4636 2733 4644
rect 2747 4636 2953 4644
rect 3007 4636 3133 4644
rect 3207 4636 3233 4644
rect 3287 4636 3333 4644
rect 3647 4636 3813 4644
rect 3907 4636 3933 4644
rect 4787 4636 5533 4644
rect 5547 4636 5753 4644
rect 5767 4636 5773 4644
rect 6047 4636 6153 4644
rect 6407 4636 6593 4644
rect 6647 4636 6873 4644
rect 7107 4636 7193 4644
rect 7627 4636 7673 4644
rect 147 4616 473 4624
rect 567 4616 633 4624
rect 787 4616 1073 4624
rect 1107 4616 1173 4624
rect 2207 4616 2233 4624
rect 2387 4616 2773 4624
rect 3087 4616 3253 4624
rect 3267 4616 3373 4624
rect 3507 4616 3773 4624
rect 4747 4616 4853 4624
rect 4887 4616 5033 4624
rect 5287 4616 5573 4624
rect 5587 4616 5653 4624
rect 5827 4616 6053 4624
rect 6567 4616 6713 4624
rect 6727 4616 6773 4624
rect 6787 4616 6833 4624
rect 347 4596 373 4604
rect 467 4596 573 4604
rect 987 4596 1913 4604
rect 1927 4596 2433 4604
rect 3747 4596 3773 4604
rect 4187 4596 4213 4604
rect 4227 4596 4513 4604
rect 4687 4596 4993 4604
rect 5007 4596 5113 4604
rect 5127 4596 5233 4604
rect 6067 4596 6093 4604
rect 207 4576 253 4584
rect 267 4576 673 4584
rect 907 4576 984 4584
rect 507 4556 533 4564
rect 547 4556 773 4564
rect 827 4556 953 4564
rect 976 4564 984 4576
rect 1167 4576 2253 4584
rect 2707 4576 2793 4584
rect 4067 4576 4173 4584
rect 4507 4576 4853 4584
rect 6447 4576 6513 4584
rect 7047 4576 7373 4584
rect 7487 4576 7633 4584
rect 976 4556 1644 4564
rect 227 4536 313 4544
rect 587 4536 1053 4544
rect 1187 4536 1384 4544
rect 287 4516 344 4524
rect 336 4504 344 4516
rect 407 4516 453 4524
rect 507 4516 793 4524
rect 847 4516 1113 4524
rect 1376 4524 1384 4536
rect 1447 4536 1573 4544
rect 1587 4536 1613 4544
rect 1636 4544 1644 4556
rect 1707 4556 1813 4564
rect 2087 4556 3233 4564
rect 4127 4556 4153 4564
rect 4467 4556 4973 4564
rect 4987 4556 5093 4564
rect 5267 4556 5513 4564
rect 5527 4556 5553 4564
rect 6207 4556 6273 4564
rect 6507 4556 6693 4564
rect 7427 4556 7593 4564
rect 1636 4536 1753 4544
rect 2187 4536 2393 4544
rect 2427 4536 3153 4544
rect 3367 4536 4233 4544
rect 4327 4536 5193 4544
rect 5707 4536 6373 4544
rect 6387 4536 6473 4544
rect 6687 4536 7213 4544
rect 7327 4536 7413 4544
rect 7567 4536 7753 4544
rect 1376 4516 1593 4524
rect 2087 4516 2224 4524
rect 307 4496 324 4504
rect 336 4496 513 4504
rect 316 4484 324 4496
rect 647 4496 693 4504
rect 867 4496 973 4504
rect 1047 4496 1533 4504
rect 1567 4496 1633 4504
rect 1976 4496 2013 4504
rect 316 4476 353 4484
rect 396 4476 413 4484
rect 116 4464 124 4473
rect 116 4456 173 4464
rect 267 4456 373 4464
rect 396 4447 404 4476
rect 667 4476 773 4484
rect 847 4476 864 4484
rect 647 4456 753 4464
rect 807 4456 833 4464
rect 856 4464 864 4476
rect 907 4476 924 4484
rect 856 4456 884 4464
rect 416 4444 424 4453
rect 416 4436 473 4444
rect 527 4436 593 4444
rect 607 4436 853 4444
rect 876 4444 884 4456
rect 876 4436 893 4444
rect 916 4424 924 4476
rect 1007 4476 1073 4484
rect 1247 4476 1333 4484
rect 1587 4476 1653 4484
rect 1976 4484 1984 4496
rect 2047 4496 2113 4504
rect 2127 4496 2153 4504
rect 1856 4476 1984 4484
rect 936 4464 944 4473
rect 936 4456 973 4464
rect 1076 4456 1353 4464
rect 1076 4444 1084 4456
rect 1007 4436 1084 4444
rect 1107 4436 1193 4444
rect 1416 4444 1424 4473
rect 1607 4456 1713 4464
rect 1736 4464 1744 4473
rect 1856 4467 1864 4476
rect 2007 4476 2093 4484
rect 2216 4467 2224 4516
rect 2247 4516 2373 4524
rect 2387 4516 2733 4524
rect 2767 4516 2793 4524
rect 2867 4516 3033 4524
rect 3267 4516 3593 4524
rect 4207 4516 4313 4524
rect 4587 4516 5313 4524
rect 5487 4516 5713 4524
rect 5827 4516 5853 4524
rect 6227 4516 6753 4524
rect 6767 4516 6813 4524
rect 6827 4516 6913 4524
rect 7247 4516 7433 4524
rect 7527 4516 7553 4524
rect 7587 4516 7653 4524
rect 7847 4516 7873 4524
rect 2316 4496 2413 4504
rect 2267 4476 2293 4484
rect 1736 4456 1793 4464
rect 1887 4456 2053 4464
rect 2316 4464 2324 4496
rect 2756 4496 2813 4504
rect 2347 4476 2513 4484
rect 2607 4476 2673 4484
rect 2756 4467 2764 4496
rect 2847 4496 2913 4504
rect 3047 4496 3113 4504
rect 3527 4496 3573 4504
rect 3587 4496 3853 4504
rect 4087 4496 4253 4504
rect 4407 4496 4573 4504
rect 4967 4496 5133 4504
rect 5167 4496 5213 4504
rect 5227 4496 5293 4504
rect 5347 4496 5393 4504
rect 5667 4496 5753 4504
rect 5807 4496 6073 4504
rect 6207 4496 6253 4504
rect 6487 4496 6553 4504
rect 6947 4496 7053 4504
rect 7067 4496 7133 4504
rect 7267 4496 7413 4504
rect 7747 4496 7773 4504
rect 2887 4476 3053 4484
rect 3347 4476 3413 4484
rect 3447 4476 3493 4484
rect 3616 4476 3633 4484
rect 2316 4456 2424 4464
rect 2416 4447 2424 4456
rect 2436 4456 2473 4464
rect 1287 4436 1533 4444
rect 1567 4436 1744 4444
rect 547 4416 924 4424
rect 1047 4416 1133 4424
rect 1207 4416 1713 4424
rect 1736 4424 1744 4436
rect 1847 4436 1973 4444
rect 2187 4436 2313 4444
rect 2367 4436 2393 4444
rect 1736 4416 2253 4424
rect 2436 4424 2444 4456
rect 2507 4456 2713 4464
rect 2847 4456 2893 4464
rect 2947 4456 2993 4464
rect 3147 4456 3193 4464
rect 3287 4456 3313 4464
rect 3336 4456 3533 4464
rect 2467 4436 2913 4444
rect 3027 4436 3053 4444
rect 3067 4436 3173 4444
rect 3336 4444 3344 4456
rect 3616 4464 3624 4476
rect 3747 4476 3813 4484
rect 4507 4476 4533 4484
rect 4547 4476 4613 4484
rect 4647 4476 5013 4484
rect 5056 4476 5273 4484
rect 3547 4456 3624 4464
rect 3636 4456 3713 4464
rect 3227 4436 3344 4444
rect 3367 4436 3473 4444
rect 3636 4444 3644 4456
rect 3807 4456 3833 4464
rect 3947 4456 3993 4464
rect 4096 4447 4104 4473
rect 4387 4456 4433 4464
rect 4447 4456 4513 4464
rect 4667 4456 4713 4464
rect 4727 4456 4773 4464
rect 4827 4456 4913 4464
rect 3627 4436 3644 4444
rect 3707 4436 3813 4444
rect 3827 4436 3873 4444
rect 4467 4436 4553 4444
rect 4647 4436 4693 4444
rect 4716 4436 4793 4444
rect 2367 4416 2444 4424
rect 2487 4416 2533 4424
rect 2667 4416 3073 4424
rect 3167 4416 3593 4424
rect 4027 4416 4113 4424
rect 4247 4416 4473 4424
rect 4607 4416 4693 4424
rect 587 4396 653 4404
rect 667 4396 933 4404
rect 1407 4396 1473 4404
rect 1547 4396 2493 4404
rect 2827 4396 3093 4404
rect 3287 4396 3473 4404
rect 3527 4396 3853 4404
rect 4127 4396 4193 4404
rect 4716 4404 4724 4436
rect 5036 4427 5044 4453
rect 5056 4447 5064 4476
rect 5327 4476 5413 4484
rect 5447 4476 5564 4484
rect 5207 4456 5493 4464
rect 5556 4464 5564 4476
rect 5627 4476 5664 4484
rect 5556 4456 5604 4464
rect 5176 4444 5184 4453
rect 5176 4436 5253 4444
rect 5267 4436 5313 4444
rect 5347 4436 5393 4444
rect 5467 4436 5553 4444
rect 5567 4436 5573 4444
rect 5596 4444 5604 4456
rect 5596 4436 5613 4444
rect 5656 4444 5664 4476
rect 5676 4476 5713 4484
rect 5676 4467 5684 4476
rect 5847 4476 5904 4484
rect 5767 4456 5813 4464
rect 5896 4464 5904 4476
rect 5967 4476 6193 4484
rect 6267 4476 6313 4484
rect 6367 4476 6453 4484
rect 6507 4476 6584 4484
rect 6576 4467 6584 4476
rect 6927 4476 7073 4484
rect 7107 4476 7144 4484
rect 5896 4456 5933 4464
rect 5987 4456 6073 4464
rect 6247 4456 6273 4464
rect 6287 4456 6333 4464
rect 6467 4456 6533 4464
rect 6647 4456 6693 4464
rect 6707 4456 6793 4464
rect 6816 4456 6933 4464
rect 5656 4436 5813 4444
rect 5827 4436 5833 4444
rect 4747 4416 4773 4424
rect 5127 4416 5453 4424
rect 5747 4416 5833 4424
rect 5856 4424 5864 4453
rect 5887 4436 5933 4444
rect 6027 4436 6093 4444
rect 6116 4424 6124 4453
rect 6427 4436 6473 4444
rect 6816 4444 6824 4456
rect 6967 4456 6993 4464
rect 7087 4456 7113 4464
rect 7136 4464 7144 4476
rect 7207 4476 7233 4484
rect 7327 4476 7453 4484
rect 7476 4476 7513 4484
rect 7136 4456 7153 4464
rect 7176 4464 7184 4473
rect 7176 4456 7253 4464
rect 7367 4456 7444 4464
rect 6756 4436 6824 4444
rect 5847 4416 6124 4424
rect 6756 4424 6764 4436
rect 6847 4436 6893 4444
rect 7296 4444 7304 4453
rect 7047 4436 7304 4444
rect 7327 4436 7353 4444
rect 7436 4444 7444 4456
rect 7476 4464 7484 4476
rect 7796 4484 7804 4493
rect 7547 4476 7564 4484
rect 7467 4456 7484 4464
rect 7556 4464 7564 4476
rect 7756 4476 7804 4484
rect 7756 4467 7764 4476
rect 7827 4476 7844 4484
rect 7836 4467 7844 4476
rect 7556 4456 7613 4464
rect 7647 4456 7673 4464
rect 7436 4436 7473 4444
rect 7487 4436 7673 4444
rect 7696 4444 7704 4453
rect 7696 4436 7773 4444
rect 7856 4444 7864 4493
rect 7827 4436 7864 4444
rect 6447 4416 6764 4424
rect 6867 4416 6993 4424
rect 7067 4416 7193 4424
rect 7447 4416 7493 4424
rect 7647 4416 7693 4424
rect 4547 4396 4724 4404
rect 5027 4396 5184 4404
rect 647 4376 813 4384
rect 847 4376 1053 4384
rect 1087 4376 1233 4384
rect 1267 4376 1433 4384
rect 1507 4376 1553 4384
rect 1747 4376 1973 4384
rect 2027 4376 2113 4384
rect 2127 4376 2213 4384
rect 2307 4376 2653 4384
rect 2687 4376 3193 4384
rect 3287 4376 4053 4384
rect 4567 4376 4593 4384
rect 4627 4376 4953 4384
rect 5176 4384 5184 4396
rect 5307 4396 5593 4404
rect 5827 4396 5893 4404
rect 7087 4396 7553 4404
rect 7647 4396 7873 4404
rect 5176 4376 5433 4384
rect 7387 4376 7593 4384
rect 607 4356 713 4364
rect 1187 4356 1313 4364
rect 1967 4356 2033 4364
rect 2067 4356 2833 4364
rect 2887 4356 3113 4364
rect 3567 4356 3653 4364
rect 3807 4356 4173 4364
rect 4187 4356 4773 4364
rect 4847 4356 6173 4364
rect 7287 4356 7553 4364
rect 27 4336 53 4344
rect 327 4336 833 4344
rect 907 4336 1213 4344
rect 1247 4336 2233 4344
rect 2347 4336 2813 4344
rect 2827 4336 3033 4344
rect 3367 4336 3493 4344
rect 3507 4336 3753 4344
rect 3767 4336 3913 4344
rect 4507 4336 4673 4344
rect 4867 4336 5013 4344
rect 5047 4336 5293 4344
rect 5307 4336 5633 4344
rect 587 4316 993 4324
rect 1067 4316 1173 4324
rect 1227 4316 2084 4324
rect 127 4296 453 4304
rect 467 4296 824 4304
rect 387 4276 553 4284
rect 816 4284 824 4296
rect 847 4296 1293 4304
rect 1327 4296 1533 4304
rect 1667 4296 1853 4304
rect 2007 4296 2053 4304
rect 2076 4304 2084 4316
rect 2107 4316 2293 4324
rect 2527 4316 2753 4324
rect 2787 4316 3733 4324
rect 3987 4316 4173 4324
rect 4467 4316 5253 4324
rect 5276 4316 5613 4324
rect 2076 4296 2133 4304
rect 2507 4296 2733 4304
rect 2847 4296 3173 4304
rect 4307 4296 4553 4304
rect 4567 4296 4753 4304
rect 4907 4296 4993 4304
rect 5276 4304 5284 4316
rect 7127 4316 7473 4324
rect 5167 4296 5284 4304
rect 7487 4296 7613 4304
rect 816 4276 933 4284
rect 987 4276 1553 4284
rect 1927 4276 2073 4284
rect 2267 4276 3133 4284
rect 4427 4276 4673 4284
rect 4707 4276 5073 4284
rect 5427 4276 5793 4284
rect 5807 4276 6013 4284
rect 6147 4276 6293 4284
rect 6607 4276 6653 4284
rect 7687 4276 7893 4284
rect 107 4256 453 4264
rect 527 4256 613 4264
rect 867 4256 993 4264
rect 1027 4256 1273 4264
rect 1367 4256 1733 4264
rect 1827 4256 1844 4264
rect 67 4236 153 4244
rect 247 4236 344 4244
rect 207 4216 313 4224
rect 36 4184 44 4213
rect 67 4196 84 4204
rect -4 4176 44 4184
rect 76 4184 84 4196
rect 107 4196 153 4204
rect 167 4196 273 4204
rect 296 4196 313 4204
rect 76 4176 93 4184
rect -4 4144 4 4176
rect 127 4176 213 4184
rect 296 4184 304 4196
rect 336 4187 344 4236
rect 427 4236 493 4244
rect 727 4236 1033 4244
rect 1056 4236 1413 4244
rect 407 4216 424 4224
rect 287 4176 304 4184
rect 27 4156 53 4164
rect 87 4156 353 4164
rect 416 4164 424 4216
rect 636 4216 773 4224
rect 436 4187 444 4213
rect 456 4196 533 4204
rect 456 4167 464 4196
rect 636 4204 644 4216
rect 1056 4224 1064 4236
rect 1607 4236 1633 4244
rect 1836 4244 1844 4256
rect 1867 4256 2093 4264
rect 2147 4256 2273 4264
rect 2287 4256 2533 4264
rect 2727 4256 2953 4264
rect 3087 4256 3813 4264
rect 4167 4256 4633 4264
rect 4727 4256 4893 4264
rect 4947 4256 4973 4264
rect 5047 4256 5073 4264
rect 5367 4256 6373 4264
rect 6547 4256 6713 4264
rect 6727 4256 7153 4264
rect 7347 4256 7433 4264
rect 7527 4256 7713 4264
rect 1787 4236 1824 4244
rect 1836 4236 1964 4244
rect 807 4216 1064 4224
rect 1107 4216 1153 4224
rect 1176 4216 1193 4224
rect 616 4196 644 4204
rect 616 4184 624 4196
rect 787 4196 793 4204
rect 807 4196 913 4204
rect 947 4196 1084 4204
rect 567 4176 624 4184
rect 967 4176 1013 4184
rect 1076 4184 1084 4196
rect 1147 4196 1153 4204
rect 1176 4204 1184 4216
rect 1496 4216 1513 4224
rect 1167 4196 1184 4204
rect 1207 4196 1313 4204
rect 1367 4196 1453 4204
rect 1076 4176 1284 4184
rect 416 4156 433 4164
rect 516 4164 524 4173
rect 516 4156 613 4164
rect 687 4156 693 4164
rect 707 4156 793 4164
rect 827 4156 853 4164
rect 927 4156 933 4164
rect 947 4156 973 4164
rect 1047 4156 1113 4164
rect 1276 4164 1284 4176
rect 1307 4176 1473 4184
rect 1276 4156 1353 4164
rect 1496 4164 1504 4216
rect 1627 4216 1704 4224
rect 1547 4196 1593 4204
rect 1647 4196 1673 4204
rect 1696 4187 1704 4216
rect 1767 4216 1804 4224
rect 1727 4196 1773 4204
rect 1587 4176 1653 4184
rect 1387 4156 1504 4164
rect 1607 4156 1753 4164
rect 1796 4164 1804 4216
rect 1816 4167 1824 4236
rect 1867 4216 1893 4224
rect 1916 4216 1933 4224
rect 1836 4167 1844 4213
rect 1787 4156 1804 4164
rect -4 4136 173 4144
rect 307 4136 393 4144
rect 547 4136 593 4144
rect 647 4136 733 4144
rect 747 4136 873 4144
rect 887 4136 913 4144
rect 1007 4136 1173 4144
rect 1347 4136 1393 4144
rect 1427 4136 1493 4144
rect 1876 4144 1884 4173
rect 1896 4167 1904 4193
rect 1916 4187 1924 4216
rect 1956 4204 1964 4236
rect 2047 4236 2093 4244
rect 2196 4236 2433 4244
rect 2196 4224 2204 4236
rect 2456 4236 2833 4244
rect 1987 4216 2204 4224
rect 1947 4196 2033 4204
rect 2076 4204 2084 4216
rect 2227 4216 2244 4224
rect 2047 4196 2064 4204
rect 2076 4196 2104 4204
rect 1936 4164 1944 4193
rect 1987 4176 2033 4184
rect 2056 4184 2064 4196
rect 2096 4184 2104 4196
rect 2127 4196 2173 4204
rect 2236 4204 2244 4216
rect 2456 4224 2464 4236
rect 2967 4236 3093 4244
rect 3107 4236 3153 4244
rect 3347 4236 3364 4244
rect 3356 4227 3364 4236
rect 3427 4236 3553 4244
rect 3567 4236 3693 4244
rect 4416 4236 5113 4244
rect 2327 4216 2464 4224
rect 2687 4216 2713 4224
rect 2787 4216 2853 4224
rect 2867 4216 3053 4224
rect 3267 4216 3304 4224
rect 2236 4196 2253 4204
rect 2307 4196 2473 4204
rect 2496 4204 2504 4213
rect 3296 4207 3304 4216
rect 3547 4216 3613 4224
rect 4376 4224 4384 4233
rect 4416 4227 4424 4236
rect 5156 4236 5253 4244
rect 5156 4227 5164 4236
rect 5407 4236 5693 4244
rect 6147 4236 6753 4244
rect 6847 4236 6973 4244
rect 6987 4236 7093 4244
rect 7267 4236 7613 4244
rect 7727 4236 7753 4244
rect 4376 4216 4404 4224
rect 2496 4196 2553 4204
rect 2587 4196 2653 4204
rect 2727 4196 2793 4204
rect 2816 4196 2873 4204
rect 2056 4176 2084 4184
rect 2096 4176 2193 4184
rect 2076 4164 2084 4176
rect 2216 4184 2224 4193
rect 2216 4176 2273 4184
rect 2287 4176 2333 4184
rect 2387 4176 2473 4184
rect 2487 4176 2613 4184
rect 2816 4184 2824 4196
rect 2947 4196 2973 4204
rect 2987 4196 3284 4204
rect 2767 4176 2824 4184
rect 2967 4176 3073 4184
rect 3276 4184 3284 4196
rect 3347 4196 3453 4204
rect 3467 4196 3833 4204
rect 3887 4196 4093 4204
rect 4396 4204 4404 4216
rect 4687 4216 4724 4224
rect 4396 4196 4513 4204
rect 4716 4204 4724 4216
rect 4747 4216 4813 4224
rect 4967 4216 4984 4224
rect 4716 4196 4804 4204
rect 3276 4176 3333 4184
rect 3447 4176 3653 4184
rect 3687 4176 3893 4184
rect 4207 4176 4273 4184
rect 4347 4176 4433 4184
rect 4507 4176 4573 4184
rect 4687 4176 4713 4184
rect 4796 4184 4804 4196
rect 4976 4204 4984 4216
rect 5007 4216 5073 4224
rect 5207 4216 5233 4224
rect 5487 4216 5553 4224
rect 6187 4216 6233 4224
rect 6807 4216 7153 4224
rect 7307 4216 7413 4224
rect 7436 4216 7473 4224
rect 4827 4196 5153 4204
rect 5187 4196 5213 4204
rect 5236 4196 5293 4204
rect 4796 4176 4873 4184
rect 4987 4176 5073 4184
rect 5236 4184 5244 4196
rect 5447 4196 5753 4204
rect 5767 4196 5873 4204
rect 5896 4196 5913 4204
rect 5147 4176 5244 4184
rect 5427 4176 5513 4184
rect 5527 4176 5613 4184
rect 5647 4176 5764 4184
rect 1927 4156 1944 4164
rect 1956 4156 2064 4164
rect 2076 4156 2173 4164
rect 1687 4136 1884 4144
rect 1956 4144 1964 4156
rect 1947 4136 1964 4144
rect 2007 4136 2033 4144
rect 2056 4144 2064 4156
rect 2207 4156 2393 4164
rect 2567 4156 2653 4164
rect 2927 4156 2973 4164
rect 3007 4156 3044 4164
rect 2056 4136 2493 4144
rect 2607 4136 2753 4144
rect 2787 4136 2893 4144
rect 2907 4136 3013 4144
rect 3036 4144 3044 4156
rect 3327 4156 3393 4164
rect 3587 4156 3613 4164
rect 3707 4156 3713 4164
rect 3727 4156 3873 4164
rect 3887 4156 4073 4164
rect 4087 4156 4113 4164
rect 4227 4156 4273 4164
rect 4647 4156 4753 4164
rect 4847 4156 5053 4164
rect 5227 4156 5273 4164
rect 5327 4156 5553 4164
rect 5607 4156 5733 4164
rect 5756 4164 5764 4176
rect 5896 4184 5904 4196
rect 5927 4196 6013 4204
rect 6067 4196 6333 4204
rect 5787 4176 5904 4184
rect 6127 4176 6193 4184
rect 6436 4184 6444 4193
rect 6616 4187 6624 4213
rect 6887 4196 6973 4204
rect 7067 4196 7133 4204
rect 6367 4176 6444 4184
rect 6467 4176 6533 4184
rect 6627 4176 6633 4184
rect 6796 4184 6804 4193
rect 7196 4187 7204 4213
rect 7387 4196 7413 4204
rect 7436 4187 7444 4216
rect 7587 4216 7673 4224
rect 7867 4216 7893 4224
rect 7467 4196 7493 4204
rect 7536 4187 7544 4213
rect 7667 4196 7753 4204
rect 6687 4176 6804 4184
rect 7007 4176 7073 4184
rect 7107 4176 7173 4184
rect 7447 4176 7524 4184
rect 5756 4156 5893 4164
rect 5907 4156 5993 4164
rect 6387 4156 6733 4164
rect 6907 4156 7013 4164
rect 7127 4156 7233 4164
rect 7247 4156 7473 4164
rect 7516 4164 7524 4176
rect 7556 4184 7564 4193
rect 7556 4176 7593 4184
rect 7636 4184 7644 4193
rect 7776 4187 7784 4213
rect 7627 4176 7644 4184
rect 7516 4156 7633 4164
rect 7647 4156 7653 4164
rect 7796 4164 7804 4193
rect 7816 4184 7824 4213
rect 7836 4204 7844 4213
rect 7836 4196 7884 4204
rect 7876 4187 7884 4196
rect 7816 4176 7833 4184
rect 7787 4156 7804 4164
rect 3036 4136 3113 4144
rect 3127 4136 3453 4144
rect 3467 4136 3533 4144
rect 4047 4136 4233 4144
rect 4547 4136 4793 4144
rect 5067 4136 5353 4144
rect 5516 4136 5653 4144
rect 67 4116 233 4124
rect 267 4116 293 4124
rect 1127 4116 1293 4124
rect 1347 4116 1353 4124
rect 1367 4116 1513 4124
rect 1967 4116 2053 4124
rect 2067 4116 2193 4124
rect 2227 4116 2313 4124
rect 2327 4116 2413 4124
rect 2447 4116 3464 4124
rect 47 4096 613 4104
rect 1187 4096 1433 4104
rect 1527 4096 1704 4104
rect 287 4076 313 4084
rect 407 4076 593 4084
rect 667 4076 713 4084
rect 747 4076 793 4084
rect 1067 4076 1393 4084
rect 1696 4084 1704 4096
rect 1727 4096 2013 4104
rect 2047 4096 2073 4104
rect 2147 4096 2353 4104
rect 2567 4096 2853 4104
rect 2867 4096 3073 4104
rect 3187 4096 3273 4104
rect 3456 4104 3464 4116
rect 3487 4116 3593 4124
rect 5516 4124 5524 4136
rect 5667 4136 6113 4144
rect 6167 4136 6413 4144
rect 6427 4136 6453 4144
rect 6567 4136 6713 4144
rect 6727 4136 6853 4144
rect 7367 4136 7733 4144
rect 7747 4136 7813 4144
rect 4867 4116 5524 4124
rect 5587 4116 6073 4124
rect 6087 4116 6133 4124
rect 6267 4116 6553 4124
rect 6587 4116 6953 4124
rect 7427 4116 7453 4124
rect 3456 4096 4353 4104
rect 5107 4096 5213 4104
rect 5247 4096 5913 4104
rect 5947 4096 6593 4104
rect 6607 4096 6673 4104
rect 7827 4096 7853 4104
rect 1696 4076 1993 4084
rect 2067 4076 2213 4084
rect 2267 4076 2473 4084
rect 2507 4076 2813 4084
rect 3007 4076 3033 4084
rect 3227 4076 3393 4084
rect 3627 4076 3733 4084
rect 4387 4076 4533 4084
rect 4547 4076 4753 4084
rect 4767 4076 5333 4084
rect 5347 4076 5493 4084
rect 5507 4076 5933 4084
rect 6047 4076 6353 4084
rect 27 4056 333 4064
rect 347 4056 473 4064
rect 496 4056 853 4064
rect 96 4036 204 4044
rect 96 4007 104 4036
rect 147 4016 173 4024
rect 196 4024 204 4036
rect 247 4036 253 4044
rect 496 4044 504 4056
rect 1247 4056 1273 4064
rect 1367 4056 1653 4064
rect 1667 4056 1693 4064
rect 1887 4056 1973 4064
rect 2027 4056 2253 4064
rect 2287 4056 2333 4064
rect 2427 4056 2593 4064
rect 2687 4056 2773 4064
rect 2887 4056 2913 4064
rect 2936 4056 3053 4064
rect 267 4036 504 4044
rect 627 4036 904 4044
rect 196 4016 353 4024
rect 387 4016 413 4024
rect 447 4016 564 4024
rect 376 3996 513 4004
rect 136 3964 144 3993
rect 167 3976 233 3984
rect 316 3984 324 3993
rect 376 3987 384 3996
rect 556 4004 564 4016
rect 587 4016 633 4024
rect 667 4016 693 4024
rect 707 4016 753 4024
rect 767 4016 793 4024
rect 896 4024 904 4036
rect 1207 4036 1293 4044
rect 1487 4036 1513 4044
rect 1587 4036 2073 4044
rect 2187 4036 2733 4044
rect 2936 4044 2944 4056
rect 3207 4056 3233 4064
rect 3267 4056 3313 4064
rect 5007 4056 5073 4064
rect 5127 4056 5473 4064
rect 5567 4056 5633 4064
rect 5656 4056 5853 4064
rect 2767 4036 2944 4044
rect 2987 4036 3013 4044
rect 3167 4036 3284 4044
rect 847 4016 884 4024
rect 896 4016 1253 4024
rect 556 3996 604 4004
rect 596 3987 604 3996
rect 287 3976 324 3984
rect 447 3976 533 3984
rect 616 3984 624 3993
rect 616 3976 773 3984
rect 136 3956 153 3964
rect 467 3956 493 3964
rect 507 3956 513 3964
rect 647 3956 853 3964
rect 876 3964 884 4016
rect 1327 4016 1533 4024
rect 1567 4016 1613 4024
rect 1627 4016 1753 4024
rect 1787 4016 1953 4024
rect 1976 4016 2013 4024
rect 1976 4007 1984 4016
rect 2127 4016 2144 4024
rect 916 3996 1124 4004
rect 916 3984 924 3996
rect 907 3976 924 3984
rect 947 3976 973 3984
rect 1047 3976 1073 3984
rect 1116 3984 1124 3996
rect 1147 3996 1184 4004
rect 1116 3976 1153 3984
rect 1176 3967 1184 3996
rect 1287 3996 1693 4004
rect 1867 3996 1953 4004
rect 1987 3996 2004 4004
rect 876 3956 1153 3964
rect 1216 3964 1224 3993
rect 1996 3987 2004 3996
rect 1267 3976 1773 3984
rect 1796 3976 1924 3984
rect 1216 3956 1413 3964
rect 1796 3964 1804 3976
rect 1447 3956 1804 3964
rect 1827 3956 1833 3964
rect 1847 3956 1893 3964
rect 1916 3964 1924 3976
rect 2016 3964 2024 3993
rect 2076 3987 2084 4013
rect 2136 4007 2144 4016
rect 2196 4016 2313 4024
rect 2196 3987 2204 4016
rect 2407 4016 2493 4024
rect 2647 4016 2793 4024
rect 2827 4016 2933 4024
rect 2947 4016 3033 4024
rect 3107 4016 3133 4024
rect 3187 4016 3253 4024
rect 3276 4024 3284 4036
rect 3307 4036 3353 4044
rect 4447 4036 4744 4044
rect 3276 4016 3593 4024
rect 3776 4016 3833 4024
rect 3776 4007 3784 4016
rect 3867 4016 3913 4024
rect 3967 4016 4073 4024
rect 4567 4016 4653 4024
rect 4736 4024 4744 4036
rect 4787 4036 4953 4044
rect 4967 4036 4993 4044
rect 5027 4036 5193 4044
rect 5227 4036 5313 4044
rect 5367 4036 5413 4044
rect 5656 4044 5664 4056
rect 5927 4056 6233 4064
rect 6247 4056 6313 4064
rect 6327 4056 6373 4064
rect 6787 4056 7093 4064
rect 7727 4056 7853 4064
rect 5467 4036 5664 4044
rect 5687 4036 6873 4044
rect 6887 4036 6913 4044
rect 6927 4036 7033 4044
rect 7727 4036 7753 4044
rect 7847 4036 7873 4044
rect 4736 4016 4773 4024
rect 4807 4016 4933 4024
rect 4947 4016 4973 4024
rect 4987 4016 5104 4024
rect 2227 3996 2253 4004
rect 2336 3996 2393 4004
rect 2276 3984 2284 3993
rect 2267 3976 2284 3984
rect 1916 3956 1964 3964
rect 2016 3956 2113 3964
rect 567 3936 733 3944
rect 827 3936 833 3944
rect 847 3936 1613 3944
rect 1727 3936 1933 3944
rect 1956 3944 1964 3956
rect 2127 3956 2293 3964
rect 2316 3964 2324 3993
rect 2336 3987 2344 3996
rect 2727 3996 2764 4004
rect 2347 3976 2364 3984
rect 2316 3956 2333 3964
rect 2356 3944 2364 3976
rect 2436 3964 2444 3993
rect 2467 3976 2693 3984
rect 2756 3967 2764 3996
rect 2776 3996 3013 4004
rect 2776 3967 2784 3996
rect 3027 3996 3044 4004
rect 2816 3976 2873 3984
rect 2436 3956 2493 3964
rect 2567 3956 2613 3964
rect 2727 3956 2744 3964
rect 1956 3936 2364 3944
rect 2407 3936 2713 3944
rect 2736 3944 2744 3956
rect 2816 3964 2824 3976
rect 3036 3984 3044 3996
rect 3067 3996 3233 4004
rect 3956 3996 3973 4004
rect 3036 3976 3124 3984
rect 3116 3967 3124 3976
rect 3247 3976 3304 3984
rect 2796 3956 2824 3964
rect 2796 3947 2804 3956
rect 2907 3956 2973 3964
rect 2987 3956 3013 3964
rect 3187 3956 3253 3964
rect 3296 3964 3304 3976
rect 3336 3984 3344 3993
rect 3327 3976 3344 3984
rect 3936 3984 3944 3993
rect 3956 3987 3964 3996
rect 4127 3996 4224 4004
rect 3867 3976 3944 3984
rect 4216 3984 4224 3996
rect 4607 3996 4733 4004
rect 5096 4004 5104 4016
rect 5307 4016 5373 4024
rect 5447 4016 5553 4024
rect 5567 4016 5793 4024
rect 5967 4016 6093 4024
rect 6107 4016 6153 4024
rect 6167 4016 6253 4024
rect 6367 4016 6493 4024
rect 6547 4016 6793 4024
rect 7227 4016 7333 4024
rect 7627 4016 7673 4024
rect 7807 4016 7833 4024
rect 7867 4016 7884 4024
rect 5096 3996 5604 4004
rect 4216 3976 4313 3984
rect 4327 3976 4433 3984
rect 4556 3976 4613 3984
rect 4556 3967 4564 3976
rect 5247 3976 5433 3984
rect 5596 3984 5604 3996
rect 5627 3996 5713 4004
rect 5727 3996 5753 4004
rect 5867 3996 5953 4004
rect 6276 3996 6353 4004
rect 5596 3976 5673 3984
rect 3296 3956 3553 3964
rect 4067 3956 4453 3964
rect 4467 3956 4473 3964
rect 4587 3956 4673 3964
rect 5007 3956 5253 3964
rect 5367 3956 5393 3964
rect 5447 3956 5533 3964
rect 5576 3956 5593 3964
rect 5576 3947 5584 3956
rect 2736 3936 2773 3944
rect 2827 3936 2853 3944
rect 2867 3936 2913 3944
rect 3027 3936 3213 3944
rect 4107 3936 4933 3944
rect 5027 3936 5573 3944
rect 5636 3944 5644 3976
rect 5727 3976 5773 3984
rect 5847 3976 5873 3984
rect 6067 3976 6173 3984
rect 6187 3976 6213 3984
rect 6276 3984 6284 3996
rect 6527 3996 6773 4004
rect 7036 3987 7044 4013
rect 7067 3996 7124 4004
rect 7116 3987 7124 3996
rect 7147 3996 7253 4004
rect 7467 3996 7493 4004
rect 7567 3996 7573 4004
rect 7607 3996 7673 4004
rect 7696 4004 7704 4013
rect 7696 3996 7724 4004
rect 7716 3987 7724 3996
rect 7787 3996 7813 4004
rect 6227 3976 6284 3984
rect 6307 3976 6393 3984
rect 6447 3976 6473 3984
rect 6487 3976 6533 3984
rect 6547 3976 6553 3984
rect 6587 3976 6653 3984
rect 6707 3976 6813 3984
rect 6927 3976 6953 3984
rect 6967 3976 6993 3984
rect 7247 3976 7273 3984
rect 7327 3976 7344 3984
rect 5667 3956 5693 3964
rect 5747 3956 5813 3964
rect 5907 3956 5973 3964
rect 6007 3956 6013 3964
rect 6027 3956 6073 3964
rect 6247 3956 6273 3964
rect 6327 3956 6473 3964
rect 7336 3964 7344 3976
rect 7367 3976 7404 3984
rect 7396 3964 7404 3976
rect 7547 3976 7573 3984
rect 7667 3976 7693 3984
rect 7856 3984 7864 3993
rect 7767 3976 7864 3984
rect 7336 3956 7384 3964
rect 7396 3956 7453 3964
rect 5636 3936 5673 3944
rect 7376 3944 7384 3956
rect 7507 3956 7593 3964
rect 7616 3964 7624 3973
rect 7616 3956 7673 3964
rect 7687 3956 7704 3964
rect 7807 3956 7853 3964
rect 7376 3936 7413 3944
rect 7547 3936 7693 3944
rect 7747 3936 7793 3944
rect 7876 3944 7884 4016
rect 7847 3936 7884 3944
rect 787 3916 1173 3924
rect 1187 3916 1433 3924
rect 1487 3916 1513 3924
rect 1587 3916 1853 3924
rect 1907 3916 2193 3924
rect 2347 3916 2473 3924
rect 2507 3916 3133 3924
rect 3307 3916 3413 3924
rect 4227 3916 4273 3924
rect 5067 3916 5133 3924
rect 5407 3916 5773 3924
rect 7467 3916 7553 3924
rect 327 3896 1013 3904
rect 1147 3896 1533 3904
rect 1547 3896 1633 3904
rect 1747 3896 1933 3904
rect 2167 3896 2413 3904
rect 2447 3896 2793 3904
rect 2816 3896 2833 3904
rect 347 3876 433 3884
rect 447 3876 473 3884
rect 947 3876 1293 3884
rect 1327 3876 1353 3884
rect 1387 3876 1473 3884
rect 1927 3876 2233 3884
rect 2307 3876 2453 3884
rect 2567 3876 2673 3884
rect 2707 3876 2733 3884
rect 2816 3884 2824 3896
rect 2847 3896 3293 3904
rect 4687 3896 5333 3904
rect 5647 3896 5873 3904
rect 2787 3876 2824 3884
rect 2947 3876 4033 3884
rect 4647 3876 5104 3884
rect 307 3856 393 3864
rect 847 3856 1133 3864
rect 1187 3856 1353 3864
rect 1387 3856 1673 3864
rect 1787 3856 2393 3864
rect 2487 3856 2513 3864
rect 2527 3856 2853 3864
rect 2987 3856 3053 3864
rect 3127 3856 3713 3864
rect 4547 3856 4813 3864
rect 4847 3856 4993 3864
rect 5096 3864 5104 3876
rect 7687 3876 7773 3884
rect 5096 3856 5213 3864
rect 7667 3856 7733 3864
rect 267 3836 593 3844
rect 767 3836 1393 3844
rect 1447 3836 1973 3844
rect 2087 3836 2213 3844
rect 2347 3836 2533 3844
rect 2667 3836 2933 3844
rect 3067 3836 3193 3844
rect 5127 3836 5273 3844
rect 5287 3836 5493 3844
rect 5527 3836 5553 3844
rect 7667 3836 7913 3844
rect 367 3816 753 3824
rect 907 3816 1113 3824
rect 1567 3816 1713 3824
rect 1947 3816 2393 3824
rect 2427 3816 2433 3824
rect 2447 3816 2524 3824
rect 587 3796 713 3804
rect 1207 3796 1373 3804
rect 1507 3796 1824 3804
rect 87 3776 213 3784
rect 227 3776 593 3784
rect 627 3776 713 3784
rect 967 3776 1133 3784
rect 1267 3776 1593 3784
rect 1767 3776 1793 3784
rect 1816 3784 1824 3796
rect 1847 3796 2053 3804
rect 2067 3796 2493 3804
rect 2516 3804 2524 3816
rect 2587 3816 3313 3824
rect 3427 3816 3453 3824
rect 4527 3816 4633 3824
rect 4647 3816 5293 3824
rect 5307 3816 5393 3824
rect 5487 3816 5893 3824
rect 5907 3816 6013 3824
rect 6027 3816 6273 3824
rect 7807 3816 7913 3824
rect 2516 3796 2593 3804
rect 2627 3796 3033 3804
rect 3047 3796 3153 3804
rect 4567 3796 4653 3804
rect 4987 3796 5433 3804
rect 5767 3796 5833 3804
rect 5987 3796 6113 3804
rect 1816 3776 2073 3784
rect 2107 3776 2113 3784
rect 2127 3776 2293 3784
rect 2407 3776 2533 3784
rect 2567 3776 2633 3784
rect 2687 3776 2973 3784
rect 3007 3776 3073 3784
rect 3087 3776 3353 3784
rect 3567 3776 3873 3784
rect 4707 3776 4793 3784
rect 4827 3776 4853 3784
rect 4867 3776 5653 3784
rect 5667 3776 5773 3784
rect 5967 3776 6353 3784
rect 7547 3776 7553 3784
rect 476 3756 693 3764
rect 396 3716 453 3724
rect 147 3696 153 3704
rect 167 3696 373 3704
rect 327 3676 353 3684
rect 396 3684 404 3716
rect 476 3704 484 3756
rect 927 3756 993 3764
rect 1127 3756 1204 3764
rect 736 3736 753 3744
rect 567 3716 653 3724
rect 467 3696 484 3704
rect 547 3696 613 3704
rect 676 3704 684 3733
rect 736 3704 744 3736
rect 1196 3744 1204 3756
rect 1307 3756 1333 3764
rect 1427 3756 1493 3764
rect 1507 3756 1613 3764
rect 1667 3756 1913 3764
rect 1967 3756 2453 3764
rect 2507 3756 2653 3764
rect 2727 3756 2753 3764
rect 3107 3756 3173 3764
rect 3227 3756 3993 3764
rect 4187 3756 4253 3764
rect 4907 3756 4973 3764
rect 5007 3756 5053 3764
rect 5187 3756 5253 3764
rect 5267 3756 5353 3764
rect 5367 3756 5633 3764
rect 5867 3756 6113 3764
rect 6127 3756 6233 3764
rect 6547 3756 6613 3764
rect 7207 3756 7244 3764
rect 1027 3736 1124 3744
rect 1196 3736 1224 3744
rect 776 3724 784 3733
rect 767 3716 784 3724
rect 976 3724 984 3733
rect 907 3716 964 3724
rect 976 3716 1004 3724
rect 647 3696 684 3704
rect 696 3696 744 3704
rect 796 3704 804 3713
rect 796 3696 813 3704
rect 387 3676 404 3684
rect 507 3676 653 3684
rect 696 3684 704 3696
rect 956 3704 964 3716
rect 956 3696 973 3704
rect 687 3676 704 3684
rect 727 3676 793 3684
rect 996 3684 1004 3716
rect 1047 3716 1073 3724
rect 1116 3707 1124 3736
rect 1216 3724 1224 3736
rect 1247 3736 1333 3744
rect 1367 3736 1933 3744
rect 2007 3736 2033 3744
rect 2087 3736 2273 3744
rect 1216 3716 1244 3724
rect 1236 3707 1244 3716
rect 1307 3716 1724 3724
rect 1287 3696 1413 3704
rect 1487 3696 1693 3704
rect 1716 3687 1724 3716
rect 1907 3716 1953 3724
rect 1976 3724 1984 3733
rect 1976 3716 2004 3724
rect 1856 3704 1864 3713
rect 1747 3696 1864 3704
rect 1927 3696 1973 3704
rect 996 3676 1033 3684
rect 1067 3676 1253 3684
rect 1287 3676 1453 3684
rect 1487 3676 1513 3684
rect 1527 3676 1633 3684
rect 1807 3676 1853 3684
rect 1996 3684 2004 3716
rect 1947 3676 2004 3684
rect 2096 3684 2104 3736
rect 2387 3736 2413 3744
rect 2487 3736 2633 3744
rect 2656 3736 2693 3744
rect 2227 3716 2284 3724
rect 2276 3704 2284 3716
rect 2307 3716 2353 3724
rect 2427 3716 2464 3724
rect 2276 3696 2353 3704
rect 2456 3687 2464 3716
rect 2527 3716 2533 3724
rect 2547 3716 2613 3724
rect 2656 3724 2664 3736
rect 2747 3736 2773 3744
rect 2787 3736 2813 3744
rect 2836 3736 2853 3744
rect 2647 3716 2664 3724
rect 2836 3724 2844 3736
rect 3267 3736 3813 3744
rect 3867 3736 4053 3744
rect 4107 3736 4233 3744
rect 4347 3736 4593 3744
rect 4607 3736 4873 3744
rect 4887 3736 4933 3744
rect 5036 3736 5133 3744
rect 2727 3716 2844 3724
rect 2947 3716 3013 3724
rect 3087 3716 3113 3724
rect 3167 3716 3204 3724
rect 3196 3707 3204 3716
rect 3367 3716 3393 3724
rect 3536 3716 3613 3724
rect 2667 3696 2733 3704
rect 3216 3687 3224 3713
rect 3247 3696 3293 3704
rect 2096 3676 2113 3684
rect 2207 3676 2213 3684
rect 2227 3676 2433 3684
rect 2827 3676 2973 3684
rect 2987 3676 3213 3684
rect 3336 3684 3344 3713
rect 3536 3687 3544 3716
rect 3676 3716 3753 3724
rect 3676 3707 3684 3716
rect 3827 3716 4013 3724
rect 4087 3716 4253 3724
rect 4727 3716 4893 3724
rect 4956 3707 4964 3733
rect 5036 3727 5044 3736
rect 5227 3736 5493 3744
rect 5507 3736 5513 3744
rect 5687 3736 5733 3744
rect 5927 3736 6053 3744
rect 6067 3736 6153 3744
rect 6207 3736 6524 3744
rect 5247 3716 5293 3724
rect 5307 3716 5333 3724
rect 5487 3716 5653 3724
rect 5767 3716 5833 3724
rect 6027 3716 6173 3724
rect 6267 3716 6393 3724
rect 6516 3724 6524 3736
rect 6547 3736 6573 3744
rect 6587 3736 6673 3744
rect 6687 3736 6793 3744
rect 6947 3736 7213 3744
rect 7236 3727 7244 3756
rect 7267 3756 7353 3764
rect 7527 3756 7564 3764
rect 7556 3747 7564 3756
rect 7576 3756 7593 3764
rect 7267 3736 7273 3744
rect 7287 3736 7313 3744
rect 7576 3727 7584 3756
rect 7627 3756 7724 3764
rect 7607 3736 7633 3744
rect 6516 3716 6553 3724
rect 6607 3716 6693 3724
rect 6916 3716 6953 3724
rect 3727 3696 3953 3704
rect 3967 3696 4113 3704
rect 4287 3696 4413 3704
rect 4967 3696 5093 3704
rect 5267 3696 5313 3704
rect 5387 3696 5453 3704
rect 5547 3696 5793 3704
rect 5807 3696 5813 3704
rect 5976 3687 5984 3713
rect 5996 3687 6004 3713
rect 6227 3696 6333 3704
rect 6487 3696 6593 3704
rect 6836 3704 6844 3713
rect 6667 3696 6844 3704
rect 6916 3704 6924 3716
rect 7027 3716 7133 3724
rect 6867 3696 6924 3704
rect 6947 3696 7193 3704
rect 7616 3704 7624 3713
rect 7676 3707 7684 3733
rect 7587 3696 7624 3704
rect 7716 3704 7724 3756
rect 7736 3756 7753 3764
rect 7736 3724 7744 3756
rect 7767 3736 7813 3744
rect 7736 3716 7773 3724
rect 7836 3724 7844 3733
rect 7816 3716 7844 3724
rect 7716 3696 7773 3704
rect 3327 3676 3344 3684
rect 3667 3676 3693 3684
rect 4247 3676 4313 3684
rect 4887 3676 4973 3684
rect 5167 3676 5353 3684
rect 5367 3676 5453 3684
rect 6047 3676 6113 3684
rect 6707 3676 6813 3684
rect 7127 3676 7153 3684
rect 7816 3684 7824 3716
rect 7847 3696 7893 3704
rect 7816 3676 7893 3684
rect 167 3656 393 3664
rect 607 3656 773 3664
rect 787 3656 833 3664
rect 847 3656 893 3664
rect 1107 3656 1193 3664
rect 1267 3656 1353 3664
rect 1567 3656 1593 3664
rect 1687 3656 2073 3664
rect 2187 3656 2273 3664
rect 2367 3656 2393 3664
rect 2487 3656 2533 3664
rect 2647 3656 2713 3664
rect 2747 3656 3024 3664
rect 107 3636 1013 3644
rect 1047 3636 1524 3644
rect 307 3616 473 3624
rect 487 3616 553 3624
rect 647 3616 1193 3624
rect 1516 3624 1524 3636
rect 1547 3636 1833 3644
rect 2147 3636 2233 3644
rect 2247 3636 2293 3644
rect 2336 3636 2833 3644
rect 2336 3627 2344 3636
rect 3016 3644 3024 3656
rect 3156 3656 3333 3664
rect 3016 3636 3093 3644
rect 3156 3644 3164 3656
rect 3347 3656 3473 3664
rect 3507 3656 3793 3664
rect 4227 3656 4273 3664
rect 4907 3656 5253 3664
rect 5307 3656 5433 3664
rect 6747 3656 6913 3664
rect 6927 3656 6933 3664
rect 6947 3656 6993 3664
rect 7807 3656 7913 3664
rect 3116 3636 3164 3644
rect 1516 3616 1684 3624
rect 127 3596 413 3604
rect 527 3596 713 3604
rect 747 3596 793 3604
rect 867 3596 1013 3604
rect 1087 3596 1153 3604
rect 1227 3596 1293 3604
rect 1676 3604 1684 3616
rect 1707 3616 1873 3624
rect 1907 3616 2173 3624
rect 2367 3616 2433 3624
rect 2567 3616 2653 3624
rect 2667 3616 2753 3624
rect 2767 3616 2773 3624
rect 3116 3624 3124 3636
rect 3207 3636 3253 3644
rect 3287 3636 4413 3644
rect 4787 3636 4953 3644
rect 5047 3636 5493 3644
rect 7727 3636 7793 3644
rect 2927 3616 3124 3624
rect 3147 3616 3293 3624
rect 3407 3616 3833 3624
rect 3847 3616 4033 3624
rect 4847 3616 5113 3624
rect 5127 3616 5593 3624
rect 1676 3596 1953 3604
rect 1987 3596 2133 3604
rect 2167 3596 2213 3604
rect 2487 3596 2753 3604
rect 2767 3596 2793 3604
rect 2907 3596 3053 3604
rect 3087 3596 3253 3604
rect 3267 3596 3313 3604
rect 3327 3596 3593 3604
rect 4267 3596 4333 3604
rect 5007 3596 5053 3604
rect 5087 3596 5344 3604
rect 107 3576 473 3584
rect 547 3576 613 3584
rect 687 3576 753 3584
rect 967 3576 1093 3584
rect 1247 3576 1273 3584
rect 1447 3576 1613 3584
rect 1636 3576 1853 3584
rect 87 3556 253 3564
rect 327 3556 493 3564
rect 567 3556 633 3564
rect 667 3556 753 3564
rect 767 3556 933 3564
rect 1127 3556 1253 3564
rect 1287 3556 1353 3564
rect 1407 3556 1533 3564
rect 1636 3564 1644 3576
rect 1986 3576 2033 3584
rect 1627 3556 1644 3564
rect 1787 3556 1833 3564
rect 1986 3564 1994 3576
rect 2047 3576 2193 3584
rect 2327 3576 2633 3584
rect 2647 3576 2693 3584
rect 2967 3576 3053 3584
rect 3107 3576 3193 3584
rect 3647 3576 3993 3584
rect 4027 3576 4313 3584
rect 4927 3576 5053 3584
rect 5107 3576 5253 3584
rect 5267 3576 5293 3584
rect 5336 3584 5344 3596
rect 5336 3576 5353 3584
rect 5667 3576 6093 3584
rect 6527 3576 6613 3584
rect 6847 3576 7013 3584
rect 1867 3556 1994 3564
rect 2107 3556 2153 3564
rect 2167 3556 2233 3564
rect 2407 3556 2553 3564
rect 2947 3556 3033 3564
rect 3207 3556 3233 3564
rect 3387 3556 3493 3564
rect 3527 3556 3713 3564
rect 4407 3556 4513 3564
rect 4527 3556 4613 3564
rect 4627 3556 4913 3564
rect 4927 3556 5033 3564
rect 5047 3556 5173 3564
rect 5207 3556 5753 3564
rect 5867 3556 6853 3564
rect 6867 3556 7073 3564
rect 7087 3556 7113 3564
rect 7127 3556 7213 3564
rect 7387 3556 7413 3564
rect 7447 3556 7553 3564
rect 7687 3556 7713 3564
rect 116 3536 153 3544
rect 116 3507 124 3536
rect 267 3536 293 3544
rect 316 3536 353 3544
rect 316 3524 324 3536
rect 587 3536 624 3544
rect 376 3524 384 3533
rect 227 3516 324 3524
rect 356 3516 384 3524
rect 356 3507 364 3516
rect 516 3507 524 3533
rect 616 3507 624 3536
rect 847 3536 973 3544
rect 1007 3536 1033 3544
rect 1047 3536 1513 3544
rect 1527 3536 1573 3544
rect 1807 3536 1893 3544
rect 2013 3544 2027 3547
rect 2013 3536 2164 3544
rect 816 3524 824 3533
rect 687 3516 824 3524
rect 907 3516 953 3524
rect 987 3516 1113 3524
rect 1167 3516 1384 3524
rect 1376 3507 1384 3516
rect 1487 3516 1653 3524
rect 1827 3516 1893 3524
rect 1916 3524 1924 3533
rect 1916 3516 2004 3524
rect 387 3496 433 3504
rect 827 3496 1164 3504
rect 247 3476 673 3484
rect 27 3456 464 3464
rect 27 3436 113 3444
rect 267 3436 373 3444
rect 456 3444 464 3456
rect 696 3464 704 3493
rect 747 3476 1133 3484
rect 1156 3484 1164 3496
rect 1187 3496 1273 3504
rect 1487 3496 1773 3504
rect 1807 3496 1833 3504
rect 1996 3487 2004 3516
rect 1156 3476 1384 3484
rect 487 3456 704 3464
rect 887 3456 1073 3464
rect 1147 3456 1173 3464
rect 1207 3456 1233 3464
rect 1247 3456 1353 3464
rect 1376 3464 1384 3476
rect 1427 3476 1513 3484
rect 1547 3476 1673 3484
rect 1696 3476 1993 3484
rect 1696 3464 1704 3476
rect 2016 3484 2024 3513
rect 2036 3504 2044 3536
rect 2067 3516 2104 3524
rect 2036 3496 2073 3504
rect 2096 3487 2104 3516
rect 2016 3476 2053 3484
rect 2156 3484 2164 3536
rect 2207 3536 2253 3544
rect 2407 3536 2473 3544
rect 2507 3536 2793 3544
rect 2867 3536 2944 3544
rect 2176 3516 2213 3524
rect 2176 3507 2184 3516
rect 2247 3516 2293 3524
rect 2316 3507 2324 3533
rect 2547 3516 2553 3524
rect 2567 3516 2733 3524
rect 2936 3524 2944 3536
rect 3027 3536 3144 3544
rect 2767 3516 2904 3524
rect 2936 3516 2964 3524
rect 2336 3484 2344 3513
rect 2376 3504 2384 3513
rect 2376 3496 2484 3504
rect 2156 3476 2344 3484
rect 2387 3476 2453 3484
rect 2476 3484 2484 3496
rect 2547 3496 2613 3504
rect 2687 3496 2813 3504
rect 2827 3496 2833 3504
rect 2896 3487 2904 3516
rect 2956 3507 2964 3516
rect 2987 3516 3113 3524
rect 3136 3504 3144 3536
rect 3547 3536 3573 3544
rect 3627 3536 3973 3544
rect 4007 3536 4073 3544
rect 4207 3536 4333 3544
rect 4547 3536 4613 3544
rect 4767 3536 4844 3544
rect 3316 3524 3324 3533
rect 4836 3527 4844 3536
rect 5427 3536 5773 3544
rect 5827 3536 6053 3544
rect 6347 3536 6373 3544
rect 6387 3536 6493 3544
rect 6507 3536 6533 3544
rect 6547 3536 6553 3544
rect 6647 3536 6833 3544
rect 6967 3536 6973 3544
rect 6987 3536 6993 3544
rect 7007 3536 7253 3544
rect 7487 3536 7593 3544
rect 7607 3536 7633 3544
rect 7667 3536 7733 3544
rect 7767 3536 7824 3544
rect 3247 3516 3324 3524
rect 3416 3516 3553 3524
rect 3136 3496 3333 3504
rect 3347 3496 3393 3504
rect 3416 3487 3424 3516
rect 4216 3516 4253 3524
rect 3447 3496 3533 3504
rect 3696 3487 3704 3513
rect 4216 3507 4224 3516
rect 4467 3516 4513 3524
rect 4587 3516 4713 3524
rect 4847 3516 4973 3524
rect 5027 3516 5144 3524
rect 3827 3496 4013 3504
rect 4127 3496 4173 3504
rect 4527 3496 4553 3504
rect 4607 3496 4633 3504
rect 2476 3476 2504 3484
rect 1376 3456 1704 3464
rect 1747 3456 1833 3464
rect 1887 3456 2033 3464
rect 2047 3456 2193 3464
rect 2207 3456 2473 3464
rect 456 3436 773 3444
rect 787 3436 973 3444
rect 1767 3436 1973 3444
rect 2496 3444 2504 3476
rect 2527 3476 2553 3484
rect 2596 3476 2673 3484
rect 2596 3464 2604 3476
rect 3007 3476 3393 3484
rect 3507 3476 3624 3484
rect 2547 3456 2604 3464
rect 2756 3464 2764 3473
rect 2627 3456 2764 3464
rect 2887 3456 3273 3464
rect 3367 3456 3513 3464
rect 3616 3464 3624 3476
rect 3887 3476 3913 3484
rect 4627 3476 4653 3484
rect 5136 3484 5144 3516
rect 5187 3516 5313 3524
rect 5427 3516 5524 3524
rect 5167 3496 5213 3504
rect 5347 3496 5393 3504
rect 5416 3496 5433 3504
rect 5136 3476 5153 3484
rect 5287 3476 5333 3484
rect 5416 3484 5424 3496
rect 5516 3504 5524 3516
rect 5547 3516 5713 3524
rect 5827 3516 5853 3524
rect 6147 3516 6173 3524
rect 6267 3516 6353 3524
rect 6587 3516 6913 3524
rect 6927 3516 7153 3524
rect 7336 3516 7393 3524
rect 5516 3496 5673 3504
rect 5767 3496 5793 3504
rect 5847 3496 5913 3504
rect 5976 3496 6013 3504
rect 5407 3476 5424 3484
rect 5507 3476 5553 3484
rect 5627 3476 5693 3484
rect 5747 3476 5893 3484
rect 5976 3484 5984 3496
rect 6067 3496 6113 3504
rect 6227 3496 6293 3504
rect 6327 3496 6393 3504
rect 6727 3496 6813 3504
rect 6827 3496 7033 3504
rect 7336 3504 7344 3516
rect 7407 3516 7433 3524
rect 7607 3516 7693 3524
rect 7716 3516 7793 3524
rect 7307 3496 7344 3504
rect 7367 3496 7453 3504
rect 5947 3476 5984 3484
rect 6156 3484 6164 3493
rect 7576 3487 7584 3513
rect 7716 3507 7724 3516
rect 7816 3507 7824 3536
rect 7856 3507 7864 3553
rect 7656 3496 7673 3504
rect 6007 3476 6164 3484
rect 6627 3476 6693 3484
rect 6947 3476 7133 3484
rect 3616 3456 3773 3464
rect 5087 3456 5473 3464
rect 5996 3464 6004 3473
rect 7656 3467 7664 3496
rect 7767 3496 7773 3504
rect 7776 3484 7784 3493
rect 7776 3476 7873 3484
rect 5907 3456 6004 3464
rect 6167 3456 6513 3464
rect 6527 3456 6653 3464
rect 6667 3456 6733 3464
rect 7747 3456 7813 3464
rect 2267 3436 3253 3444
rect 3487 3436 3553 3444
rect 5267 3436 5513 3444
rect 6047 3436 6253 3444
rect 47 3416 113 3424
rect 747 3416 1793 3424
rect 1967 3416 2073 3424
rect 2447 3416 2633 3424
rect 2687 3416 3253 3424
rect 3447 3416 3633 3424
rect 5207 3416 5933 3424
rect 47 3396 293 3404
rect 307 3396 813 3404
rect 867 3396 993 3404
rect 1007 3396 1473 3404
rect 1527 3396 1673 3404
rect 1707 3396 1873 3404
rect 2427 3396 2613 3404
rect 2807 3396 3353 3404
rect 3407 3396 3893 3404
rect 147 3376 153 3384
rect 167 3376 1033 3384
rect 1147 3376 1453 3384
rect 1496 3376 1793 3384
rect 347 3356 853 3364
rect 1496 3364 1504 3376
rect 1827 3376 2013 3384
rect 2047 3376 2053 3384
rect 2067 3376 2353 3384
rect 2487 3376 2873 3384
rect 2927 3376 3113 3384
rect 3187 3376 3433 3384
rect 987 3356 1504 3364
rect 1627 3356 1733 3364
rect 1907 3356 1973 3364
rect 1996 3356 2273 3364
rect 1287 3336 1413 3344
rect 1507 3336 1553 3344
rect 1596 3336 1693 3344
rect 167 3316 393 3324
rect 527 3316 573 3324
rect 1047 3316 1213 3324
rect 1267 3316 1533 3324
rect 1596 3324 1604 3336
rect 1996 3344 2004 3356
rect 2567 3356 2773 3364
rect 2827 3356 2993 3364
rect 3327 3356 3493 3364
rect 3527 3356 3793 3364
rect 3807 3356 4433 3364
rect 1727 3336 2004 3344
rect 2087 3336 2213 3344
rect 2247 3336 2333 3344
rect 2347 3336 3193 3344
rect 3207 3336 3673 3344
rect 5027 3336 5133 3344
rect 1556 3316 1604 3324
rect 347 3296 873 3304
rect 927 3296 1193 3304
rect 1556 3304 1564 3316
rect 1687 3316 2093 3324
rect 2127 3316 2153 3324
rect 2307 3316 2513 3324
rect 2627 3316 2653 3324
rect 2667 3316 3193 3324
rect 3207 3316 3333 3324
rect 3367 3316 3553 3324
rect 3567 3316 3993 3324
rect 6767 3316 6793 3324
rect 1207 3296 1564 3304
rect 1587 3296 1593 3304
rect 1607 3296 1813 3304
rect 1947 3296 2173 3304
rect 2207 3296 2233 3304
rect 2407 3296 2453 3304
rect 2567 3296 2753 3304
rect 2987 3296 3653 3304
rect 4807 3296 5273 3304
rect 5827 3296 5853 3304
rect 6427 3296 6473 3304
rect 6807 3296 6893 3304
rect 7036 3296 7053 3304
rect 287 3276 293 3284
rect 307 3276 613 3284
rect 887 3276 1073 3284
rect 1787 3276 1933 3284
rect 2107 3276 2253 3284
rect 2287 3276 2493 3284
rect 2607 3276 2673 3284
rect 2887 3276 2913 3284
rect 3027 3276 3133 3284
rect 3307 3276 3373 3284
rect 3507 3276 3573 3284
rect 3687 3276 3713 3284
rect 4567 3276 4713 3284
rect 4727 3276 4773 3284
rect 5047 3276 5313 3284
rect 5327 3276 5573 3284
rect 5867 3276 5873 3284
rect 5887 3276 6013 3284
rect 6256 3276 6273 3284
rect 6256 3267 6264 3276
rect 6287 3276 6553 3284
rect 6567 3276 6673 3284
rect 6787 3276 6893 3284
rect 267 3256 413 3264
rect 576 3256 753 3264
rect 136 3227 144 3253
rect 227 3236 304 3244
rect 227 3216 273 3224
rect 296 3224 304 3236
rect 327 3236 393 3244
rect 527 3236 544 3244
rect 296 3216 313 3224
rect 436 3207 444 3233
rect 107 3196 413 3204
rect 476 3204 484 3233
rect 536 3227 544 3236
rect 576 3227 584 3256
rect 856 3256 913 3264
rect 607 3236 733 3244
rect 747 3236 793 3244
rect 856 3227 864 3256
rect 1387 3256 1713 3264
rect 1747 3256 2124 3264
rect 2116 3247 2124 3256
rect 2147 3256 2313 3264
rect 2327 3256 2473 3264
rect 876 3236 933 3244
rect 476 3196 573 3204
rect 876 3204 884 3236
rect 987 3236 1053 3244
rect 1127 3236 1253 3244
rect 1527 3236 1564 3244
rect 1556 3227 1564 3236
rect 1627 3236 1653 3244
rect 1676 3236 1693 3244
rect 1676 3227 1684 3236
rect 1787 3236 1833 3244
rect 1887 3236 1913 3244
rect 2147 3236 2173 3244
rect 2307 3236 2353 3244
rect 2416 3227 2424 3256
rect 2647 3256 2693 3264
rect 2787 3256 2873 3264
rect 2967 3256 3053 3264
rect 3127 3256 3144 3264
rect 2747 3236 2833 3244
rect 907 3216 953 3224
rect 1087 3216 1133 3224
rect 1187 3216 1253 3224
rect 1807 3216 1864 3224
rect 847 3196 884 3204
rect 1107 3196 1213 3204
rect 1316 3204 1324 3213
rect 1856 3207 1864 3216
rect 2027 3216 2093 3224
rect 2107 3216 2273 3224
rect 2507 3216 2533 3224
rect 2616 3224 2624 3233
rect 2616 3216 2693 3224
rect 2767 3216 2793 3224
rect 2867 3216 3013 3224
rect 3036 3224 3044 3233
rect 3036 3216 3064 3224
rect 1316 3196 1433 3204
rect 1447 3196 1493 3204
rect 1507 3196 1533 3204
rect 1647 3196 1693 3204
rect 1767 3196 1793 3204
rect 1887 3196 1913 3204
rect 1927 3196 2173 3204
rect 2387 3196 2573 3204
rect 2627 3196 2653 3204
rect 2787 3196 2993 3204
rect 3007 3196 3033 3204
rect 507 3176 813 3184
rect 827 3176 1133 3184
rect 1207 3176 1593 3184
rect 1667 3176 1813 3184
rect 1836 3176 2333 3184
rect 447 3156 513 3164
rect 727 3156 913 3164
rect 1267 3156 1313 3164
rect 1836 3164 1844 3176
rect 2367 3176 2393 3184
rect 2487 3176 2593 3184
rect 2667 3176 2933 3184
rect 3056 3184 3064 3216
rect 3136 3207 3144 3256
rect 3176 3256 3233 3264
rect 3176 3227 3184 3256
rect 3276 3256 3353 3264
rect 3256 3244 3264 3253
rect 3276 3247 3284 3256
rect 3516 3256 3533 3264
rect 3247 3236 3264 3244
rect 3307 3236 3393 3244
rect 3416 3224 3424 3253
rect 3516 3244 3524 3256
rect 3556 3256 3593 3264
rect 3556 3244 3564 3256
rect 3607 3256 3773 3264
rect 4067 3256 4113 3264
rect 4427 3256 4593 3264
rect 4647 3256 4733 3264
rect 4927 3256 5093 3264
rect 5147 3256 5273 3264
rect 5396 3256 5444 3264
rect 3447 3236 3464 3244
rect 3396 3216 3424 3224
rect 3396 3207 3404 3216
rect 3456 3207 3464 3236
rect 3496 3236 3524 3244
rect 3536 3236 3564 3244
rect 3596 3236 3633 3244
rect 3496 3227 3504 3236
rect 3187 3196 3393 3204
rect 3027 3176 3064 3184
rect 3516 3184 3524 3213
rect 3536 3207 3544 3236
rect 3596 3227 3604 3236
rect 3756 3236 3853 3244
rect 3756 3227 3764 3236
rect 4307 3236 4353 3244
rect 4427 3236 4453 3244
rect 4467 3236 4473 3244
rect 4627 3236 4653 3244
rect 5396 3244 5404 3256
rect 5307 3236 5404 3244
rect 5436 3244 5444 3256
rect 5467 3256 5533 3264
rect 5647 3256 5693 3264
rect 5707 3256 5773 3264
rect 5827 3256 5944 3264
rect 5936 3247 5944 3256
rect 5967 3256 5993 3264
rect 6087 3256 6113 3264
rect 6187 3256 6244 3264
rect 6236 3247 6244 3256
rect 6447 3256 6473 3264
rect 6687 3256 6704 3264
rect 5436 3236 5473 3244
rect 5727 3236 5833 3244
rect 6087 3236 6153 3244
rect 6267 3236 6413 3244
rect 3667 3216 3693 3224
rect 3887 3216 3933 3224
rect 4187 3216 4233 3224
rect 4747 3216 4813 3224
rect 4907 3216 5193 3224
rect 5416 3224 5424 3233
rect 6696 3227 6704 3256
rect 6767 3256 6833 3264
rect 6887 3256 7013 3264
rect 7036 3244 7044 3296
rect 7527 3296 7593 3304
rect 7567 3276 7604 3284
rect 7067 3256 7173 3264
rect 7427 3256 7473 3264
rect 7596 3264 7604 3276
rect 7687 3276 7793 3284
rect 7827 3276 7853 3284
rect 7596 3256 7613 3264
rect 7627 3256 7673 3264
rect 7727 3256 7873 3264
rect 7036 3236 7073 3244
rect 7247 3236 7313 3244
rect 7347 3236 7373 3244
rect 7387 3236 7493 3244
rect 5416 3216 5493 3224
rect 5507 3216 5673 3224
rect 6067 3216 6273 3224
rect 6327 3216 6513 3224
rect 6527 3216 6533 3224
rect 6547 3216 6613 3224
rect 3627 3196 3873 3204
rect 4027 3196 4273 3204
rect 4287 3196 4393 3204
rect 4407 3196 4713 3204
rect 4727 3196 4953 3204
rect 5207 3196 5353 3204
rect 5467 3196 5573 3204
rect 6716 3204 6724 3233
rect 6976 3224 6984 3233
rect 6747 3216 6984 3224
rect 7196 3224 7204 3233
rect 7007 3216 7253 3224
rect 7267 3216 7693 3224
rect 6627 3196 6724 3204
rect 6967 3196 7013 3204
rect 7027 3196 7073 3204
rect 7227 3196 7293 3204
rect 7307 3196 7313 3204
rect 7327 3196 7353 3204
rect 7367 3196 7633 3204
rect 3267 3176 3524 3184
rect 3807 3176 3833 3184
rect 3907 3176 4353 3184
rect 4607 3176 4753 3184
rect 4787 3176 4913 3184
rect 5047 3176 5433 3184
rect 5487 3176 5553 3184
rect 5567 3176 5593 3184
rect 6667 3176 7033 3184
rect 7287 3176 7453 3184
rect 1327 3156 1844 3164
rect 2067 3156 2153 3164
rect 2267 3156 2573 3164
rect 3147 3156 3213 3164
rect 3227 3156 3333 3164
rect 3367 3156 3773 3164
rect 3787 3156 3813 3164
rect 3827 3156 3833 3164
rect 5527 3156 5913 3164
rect 6587 3156 6853 3164
rect 467 3136 613 3144
rect 1027 3136 1393 3144
rect 1487 3136 1533 3144
rect 1707 3136 1873 3144
rect 1907 3136 2073 3144
rect 2087 3136 2113 3144
rect 2567 3136 2833 3144
rect 3127 3136 3473 3144
rect 3567 3136 4053 3144
rect 87 3116 333 3124
rect 407 3116 693 3124
rect 727 3116 813 3124
rect 887 3116 1124 3124
rect 167 3096 213 3104
rect 1116 3104 1124 3116
rect 1207 3116 1393 3124
rect 1607 3116 1713 3124
rect 1767 3116 1873 3124
rect 1887 3116 1953 3124
rect 2187 3116 2193 3124
rect 2207 3116 2713 3124
rect 2727 3116 3053 3124
rect 3087 3116 3193 3124
rect 3587 3116 3633 3124
rect 3687 3116 3753 3124
rect 3947 3116 4013 3124
rect 4327 3116 4733 3124
rect 5767 3116 6033 3124
rect 6047 3116 6213 3124
rect 1116 3096 1204 3104
rect 187 3076 413 3084
rect 447 3076 533 3084
rect 547 3076 673 3084
rect 847 3076 913 3084
rect 1196 3084 1204 3096
rect 1247 3096 1373 3104
rect 1827 3096 2253 3104
rect 2447 3096 2913 3104
rect 3167 3096 3933 3104
rect 5227 3096 5753 3104
rect 5767 3096 5853 3104
rect 6387 3096 6573 3104
rect 6587 3096 6693 3104
rect 7347 3096 7473 3104
rect 7727 3096 7853 3104
rect 1196 3076 1344 3084
rect -24 3056 173 3064
rect 207 3056 253 3064
rect 307 3056 444 3064
rect 47 3036 93 3044
rect 167 3036 393 3044
rect 436 3044 444 3056
rect 467 3056 633 3064
rect 647 3056 813 3064
rect 827 3056 1113 3064
rect 1147 3056 1173 3064
rect 1196 3056 1233 3064
rect 436 3036 513 3044
rect 767 3036 1113 3044
rect 1196 3044 1204 3056
rect 1296 3056 1313 3064
rect 1127 3036 1204 3044
rect 1247 3036 1273 3044
rect 67 3016 133 3024
rect 187 3016 273 3024
rect 636 3024 644 3033
rect 1296 3027 1304 3056
rect 1336 3044 1344 3076
rect 1407 3076 1853 3084
rect 1867 3076 1933 3084
rect 2107 3076 2133 3084
rect 2207 3076 2293 3084
rect 2307 3076 2513 3084
rect 2547 3076 2613 3084
rect 2687 3076 2753 3084
rect 2807 3076 2844 3084
rect 1387 3056 1433 3064
rect 1487 3056 1613 3064
rect 1736 3056 1813 3064
rect 1736 3047 1744 3056
rect 1927 3056 1953 3064
rect 1976 3056 1993 3064
rect 1327 3036 1344 3044
rect 1367 3036 1413 3044
rect 1527 3036 1553 3044
rect 636 3016 753 3024
rect 807 3016 853 3024
rect 987 3016 1033 3024
rect 1107 3016 1253 3024
rect 1267 3016 1284 3024
rect -24 2996 33 3004
rect 87 2996 153 3004
rect 167 2996 253 3004
rect 327 2996 633 3004
rect 1027 2996 1113 3004
rect 1276 3004 1284 3016
rect 1316 3024 1324 3033
rect 1976 3027 1984 3056
rect 2267 3056 2604 3064
rect 2007 3036 2253 3044
rect 2387 3036 2473 3044
rect 2596 3044 2604 3056
rect 2627 3056 2813 3064
rect 2836 3064 2844 3076
rect 2967 3076 3073 3084
rect 3427 3076 3613 3084
rect 4047 3076 4053 3084
rect 4067 3076 4173 3084
rect 4347 3076 4573 3084
rect 4587 3076 4693 3084
rect 4967 3076 5333 3084
rect 5347 3076 5713 3084
rect 5907 3076 6153 3084
rect 6207 3076 6493 3084
rect 7267 3076 7393 3084
rect 7407 3076 7533 3084
rect 7667 3076 7693 3084
rect 7827 3076 7853 3084
rect 2836 3056 3133 3064
rect 3167 3056 3233 3064
rect 2596 3036 2653 3044
rect 2707 3036 2824 3044
rect 2816 3027 2824 3036
rect 2836 3036 2873 3044
rect 1316 3016 1753 3024
rect 2127 3016 2144 3024
rect 1276 2996 1464 3004
rect 767 2976 1013 2984
rect 1227 2976 1433 2984
rect 1456 2984 1464 2996
rect 1487 2996 1533 3004
rect 1567 2996 1833 3004
rect 2047 2996 2093 3004
rect 2136 3004 2144 3016
rect 2167 3016 2373 3024
rect 2136 2996 2293 3004
rect 2507 2996 2533 3004
rect 2647 2996 2713 3004
rect 2836 3004 2844 3036
rect 3036 3036 3273 3044
rect 2867 3016 2953 3024
rect 2996 3024 3004 3033
rect 2987 3016 3004 3024
rect 3036 3024 3044 3036
rect 3027 3016 3044 3024
rect 3067 3016 3213 3024
rect 3296 3024 3304 3073
rect 3327 3056 3373 3064
rect 3407 3056 3464 3064
rect 3347 3036 3413 3044
rect 3456 3044 3464 3056
rect 3487 3056 4073 3064
rect 4487 3056 4653 3064
rect 4667 3056 4713 3064
rect 5207 3056 5733 3064
rect 5827 3056 5984 3064
rect 3456 3036 3473 3044
rect 3567 3036 3584 3044
rect 3267 3016 3304 3024
rect 3327 3016 3393 3024
rect 2747 2996 3093 3004
rect 3147 2996 3353 3004
rect 3516 3004 3524 3033
rect 3576 3027 3584 3036
rect 3687 3036 3704 3044
rect 3516 2996 3613 3004
rect 3696 3004 3704 3036
rect 3907 3036 4093 3044
rect 3716 3024 3724 3033
rect 3716 3016 3793 3024
rect 4116 3024 4124 3053
rect 4147 3036 4433 3044
rect 4687 3036 4933 3044
rect 5307 3036 5573 3044
rect 5976 3044 5984 3056
rect 6007 3056 6193 3064
rect 6247 3056 6393 3064
rect 7087 3056 7133 3064
rect 7596 3056 7613 3064
rect 5747 3036 5884 3044
rect 5976 3036 6053 3044
rect 3847 3016 4124 3024
rect 4167 3016 4313 3024
rect 4976 3024 4984 3033
rect 5876 3027 5884 3036
rect 6187 3036 6333 3044
rect 6547 3036 6713 3044
rect 6927 3036 7153 3044
rect 7056 3027 7064 3036
rect 7247 3036 7293 3044
rect 7376 3027 7384 3053
rect 4867 3016 4993 3024
rect 5087 3016 5173 3024
rect 5487 3016 5513 3024
rect 5607 3016 5673 3024
rect 5787 3016 5833 3024
rect 5987 3016 6093 3024
rect 6107 3016 6173 3024
rect 6427 3016 6453 3024
rect 6527 3016 6593 3024
rect 6607 3016 6673 3024
rect 6767 3016 6893 3024
rect 7127 3016 7213 3024
rect 3696 2996 3953 3004
rect 5647 2996 5933 3004
rect 6167 2996 6273 3004
rect 6647 2996 6933 3004
rect 7187 2996 7273 3004
rect 7436 3004 7444 3053
rect 7456 3027 7464 3053
rect 7547 3016 7573 3024
rect 7596 3007 7604 3056
rect 7627 3056 7653 3064
rect 7676 3056 7793 3064
rect 7676 3044 7684 3056
rect 7807 3056 7833 3064
rect 7627 3036 7684 3044
rect 7796 3007 7804 3033
rect 7827 3016 7853 3024
rect 7436 2996 7553 3004
rect 1456 2976 1493 2984
rect 1527 2976 1673 2984
rect 1687 2976 2193 2984
rect 2907 2976 3013 2984
rect 3027 2976 3253 2984
rect 3547 2976 3593 2984
rect 5707 2976 6233 2984
rect 6247 2976 6593 2984
rect 6607 2976 6973 2984
rect 6987 2976 7053 2984
rect 7527 2976 7673 2984
rect 767 2956 893 2964
rect 907 2956 1053 2964
rect 1247 2956 1453 2964
rect 1476 2956 2753 2964
rect 247 2936 373 2944
rect 727 2936 773 2944
rect 947 2936 1133 2944
rect 1476 2944 1484 2956
rect 3327 2956 3473 2964
rect 3487 2956 3693 2964
rect 4187 2956 4353 2964
rect 1427 2936 1484 2944
rect 1787 2936 1913 2944
rect 2127 2936 2513 2944
rect 3587 2936 3933 2944
rect 667 2916 833 2924
rect 1007 2916 1113 2924
rect 1267 2916 1833 2924
rect 1867 2916 2024 2924
rect 287 2896 1293 2904
rect 1427 2896 1513 2904
rect 2016 2904 2024 2916
rect 2287 2916 2693 2924
rect 3407 2916 3653 2924
rect 3887 2916 3913 2924
rect 4507 2916 4533 2924
rect 7547 2916 7593 2924
rect 2016 2896 2193 2904
rect 2227 2896 2353 2904
rect 2607 2896 2633 2904
rect 2667 2896 3893 2904
rect 4007 2896 4033 2904
rect 7547 2896 7733 2904
rect 807 2876 1093 2884
rect 1116 2876 1844 2884
rect 567 2856 613 2864
rect 1116 2864 1124 2876
rect 927 2856 1124 2864
rect 1187 2856 1813 2864
rect 1836 2864 1844 2876
rect 1887 2876 2133 2884
rect 2147 2876 3413 2884
rect 3547 2876 3773 2884
rect 4007 2876 4213 2884
rect 4807 2876 4833 2884
rect 5567 2876 5653 2884
rect 7667 2876 7733 2884
rect 7747 2876 7833 2884
rect 1836 2856 1953 2864
rect 1967 2856 2233 2864
rect 2296 2856 2673 2864
rect 87 2836 333 2844
rect 1147 2836 1233 2844
rect 1507 2836 2033 2844
rect 2296 2844 2304 2856
rect 2867 2856 3313 2864
rect 3507 2856 4413 2864
rect 2167 2836 2304 2844
rect 2327 2836 2853 2844
rect 2927 2836 3664 2844
rect 127 2816 353 2824
rect 407 2816 513 2824
rect 587 2816 1453 2824
rect 1727 2816 1784 2824
rect 247 2796 453 2804
rect 507 2796 1173 2804
rect 1536 2796 1593 2804
rect 1536 2787 1544 2796
rect 1776 2804 1784 2816
rect 1807 2816 1993 2824
rect 2047 2816 2173 2824
rect 2207 2816 2313 2824
rect 2327 2816 2433 2824
rect 2447 2816 2973 2824
rect 2987 2816 3613 2824
rect 3627 2816 3633 2824
rect 3656 2824 3664 2836
rect 3687 2836 3833 2844
rect 3847 2836 4693 2844
rect 4867 2836 5093 2844
rect 3656 2816 3693 2824
rect 3727 2816 3753 2824
rect 3827 2816 3953 2824
rect 4467 2816 6373 2824
rect 1707 2796 1764 2804
rect 1776 2796 1793 2804
rect 47 2776 93 2784
rect 127 2776 273 2784
rect 347 2776 433 2784
rect 487 2776 593 2784
rect 607 2776 793 2784
rect 887 2776 953 2784
rect 976 2776 1033 2784
rect 187 2756 213 2764
rect 327 2756 473 2764
rect 496 2756 813 2764
rect 496 2747 504 2756
rect 827 2756 904 2764
rect 896 2747 904 2756
rect 227 2736 253 2744
rect 307 2736 333 2744
rect 576 2736 593 2744
rect 147 2716 293 2724
rect 576 2724 584 2736
rect 976 2744 984 2776
rect 1056 2776 1133 2784
rect 1056 2764 1064 2776
rect 1167 2776 1293 2784
rect 1467 2776 1524 2784
rect 1007 2756 1064 2764
rect 1207 2756 1273 2764
rect 1407 2756 1473 2764
rect 1516 2764 1524 2776
rect 1687 2776 1713 2784
rect 1516 2756 1733 2764
rect 1756 2764 1764 2796
rect 1867 2796 2153 2804
rect 2247 2796 2293 2804
rect 2427 2796 2464 2804
rect 1847 2776 1913 2784
rect 1947 2776 2113 2784
rect 2287 2776 2333 2784
rect 2367 2776 2393 2784
rect 2456 2784 2464 2796
rect 2527 2796 2544 2804
rect 2456 2776 2473 2784
rect 2496 2776 2513 2784
rect 1756 2756 1773 2764
rect 1787 2756 2004 2764
rect 947 2736 984 2744
rect 1067 2736 1133 2744
rect 1356 2744 1364 2753
rect 1227 2736 1573 2744
rect 1607 2736 1653 2744
rect 1676 2736 1733 2744
rect 467 2716 584 2724
rect 607 2716 673 2724
rect 747 2716 793 2724
rect 827 2716 833 2724
rect 847 2716 973 2724
rect 1307 2716 1333 2724
rect 1467 2716 1493 2724
rect 1676 2724 1684 2736
rect 1747 2736 1753 2744
rect 1867 2736 1973 2744
rect 1996 2744 2004 2756
rect 2067 2756 2253 2764
rect 2307 2756 2373 2764
rect 2496 2764 2504 2776
rect 2536 2767 2544 2796
rect 2587 2796 2953 2804
rect 2967 2796 3053 2804
rect 3367 2796 3453 2804
rect 3747 2796 3913 2804
rect 4767 2796 5253 2804
rect 5907 2796 5933 2804
rect 5956 2796 6113 2804
rect 2687 2776 2913 2784
rect 2987 2776 3073 2784
rect 3387 2776 3413 2784
rect 3447 2776 3733 2784
rect 3787 2776 3813 2784
rect 3827 2776 4273 2784
rect 4907 2776 5033 2784
rect 5047 2776 5053 2784
rect 5956 2784 5964 2796
rect 6807 2796 6913 2804
rect 6927 2796 6993 2804
rect 7287 2796 7493 2804
rect 7736 2796 7793 2804
rect 5856 2776 5964 2784
rect 5856 2767 5864 2776
rect 6047 2776 6233 2784
rect 6307 2776 6353 2784
rect 6507 2776 6613 2784
rect 6727 2776 6753 2784
rect 7027 2776 7313 2784
rect 7527 2776 7633 2784
rect 2427 2756 2504 2764
rect 2587 2756 2793 2764
rect 2907 2756 2953 2764
rect 3076 2756 3113 2764
rect 1996 2736 2193 2744
rect 2467 2736 2673 2744
rect 3016 2744 3024 2753
rect 3076 2747 3084 2756
rect 3227 2756 3353 2764
rect 3367 2756 3413 2764
rect 3467 2756 3533 2764
rect 3567 2756 3604 2764
rect 2887 2736 3024 2744
rect 3367 2736 3513 2744
rect 1547 2716 1684 2724
rect 1707 2716 1893 2724
rect 1987 2716 2033 2724
rect 2087 2716 2253 2724
rect 2527 2716 2893 2724
rect 3047 2716 3233 2724
rect 3287 2716 3493 2724
rect 3596 2724 3604 2756
rect 3616 2756 3633 2764
rect 3616 2747 3624 2756
rect 3836 2756 4013 2764
rect 3596 2716 3613 2724
rect 3776 2724 3784 2753
rect 3836 2747 3844 2756
rect 4947 2756 5173 2764
rect 5327 2756 5484 2764
rect 5476 2747 5484 2756
rect 5916 2756 6033 2764
rect 5916 2747 5924 2756
rect 6127 2756 6273 2764
rect 6367 2756 6513 2764
rect 6647 2756 6773 2764
rect 6887 2756 6953 2764
rect 7736 2764 7744 2796
rect 7767 2776 7813 2784
rect 7736 2756 7784 2764
rect 3996 2736 4073 2744
rect 3996 2727 4004 2736
rect 4267 2736 4313 2744
rect 4387 2736 4553 2744
rect 4687 2736 4813 2744
rect 4987 2736 5113 2744
rect 5687 2736 5713 2744
rect 5736 2736 5873 2744
rect 3647 2716 3784 2724
rect 4167 2716 4393 2724
rect 4407 2716 4633 2724
rect 4847 2716 4873 2724
rect 5107 2716 5153 2724
rect 5167 2716 5193 2724
rect 5307 2716 5353 2724
rect 5736 2724 5744 2736
rect 6096 2744 6104 2753
rect 7776 2747 7784 2756
rect 6096 2736 6173 2744
rect 6587 2736 6673 2744
rect 6867 2736 6933 2744
rect 6947 2736 6973 2744
rect 7227 2736 7393 2744
rect 7467 2736 7633 2744
rect 5647 2716 5744 2724
rect 5787 2716 5953 2724
rect 5967 2716 6013 2724
rect 6607 2716 6693 2724
rect 6827 2716 6873 2724
rect 7207 2716 7353 2724
rect 7796 2724 7804 2753
rect 7827 2736 7913 2744
rect 7787 2716 7804 2724
rect 7827 2716 7853 2724
rect 307 2696 533 2704
rect 547 2696 633 2704
rect 647 2696 713 2704
rect 967 2696 1013 2704
rect 1107 2696 1213 2704
rect 1367 2696 1413 2704
rect 1547 2696 1553 2704
rect 1567 2696 1933 2704
rect 2167 2696 2453 2704
rect 2727 2696 3033 2704
rect 3047 2696 3273 2704
rect 3447 2696 3753 2704
rect 3807 2696 4193 2704
rect 4647 2696 4773 2704
rect 6027 2696 6073 2704
rect 6667 2696 7013 2704
rect 427 2676 533 2684
rect 787 2676 913 2684
rect 1167 2676 1373 2684
rect 1387 2676 1413 2684
rect 1427 2676 1513 2684
rect 1847 2676 1873 2684
rect 1927 2676 1993 2684
rect 2047 2676 2173 2684
rect 2187 2676 2213 2684
rect 2227 2676 2553 2684
rect 2887 2676 2993 2684
rect 3167 2676 3273 2684
rect 3287 2676 3573 2684
rect 4147 2676 4433 2684
rect 807 2656 1093 2664
rect 1247 2656 1893 2664
rect 2007 2656 2493 2664
rect 3087 2656 3093 2664
rect 3107 2656 3513 2664
rect 4247 2656 4513 2664
rect 6367 2656 6633 2664
rect 6647 2656 6973 2664
rect 6987 2656 7173 2664
rect 7187 2656 7553 2664
rect 187 2636 493 2644
rect 667 2636 733 2644
rect 1007 2636 1253 2644
rect 1667 2636 1793 2644
rect 1827 2636 2333 2644
rect 2347 2636 2373 2644
rect 2447 2636 2733 2644
rect 2767 2636 2853 2644
rect 3507 2636 3773 2644
rect 4747 2636 4793 2644
rect 5327 2636 5553 2644
rect 6587 2636 6833 2644
rect 107 2616 173 2624
rect 287 2616 573 2624
rect 947 2616 1353 2624
rect 1367 2616 1513 2624
rect 1647 2616 2233 2624
rect 2487 2616 2573 2624
rect 2627 2616 2933 2624
rect 3027 2616 3233 2624
rect 3447 2616 3553 2624
rect 3567 2616 3993 2624
rect 4007 2616 4053 2624
rect 5507 2616 5573 2624
rect 5587 2616 5753 2624
rect 5967 2616 6193 2624
rect 6667 2616 6733 2624
rect 6747 2616 6793 2624
rect 7027 2616 7213 2624
rect 47 2596 133 2604
rect 467 2596 513 2604
rect 527 2596 1053 2604
rect 1447 2596 1853 2604
rect 1876 2596 2153 2604
rect 107 2576 153 2584
rect 167 2576 213 2584
rect 567 2576 613 2584
rect 627 2576 653 2584
rect 1567 2576 1613 2584
rect 1727 2576 1793 2584
rect 1876 2584 1884 2596
rect 2207 2596 2253 2604
rect 2567 2596 2633 2604
rect 2676 2596 2693 2604
rect 1827 2576 1884 2584
rect 1907 2576 2473 2584
rect 87 2556 184 2564
rect 67 2536 153 2544
rect -24 2516 33 2524
rect 176 2524 184 2556
rect 527 2556 604 2564
rect 207 2536 253 2544
rect 287 2536 293 2544
rect 307 2536 333 2544
rect 407 2536 473 2544
rect 596 2544 604 2556
rect 627 2556 673 2564
rect 727 2556 933 2564
rect 987 2556 1173 2564
rect 1207 2556 1233 2564
rect 1267 2556 1293 2564
rect 1347 2556 1384 2564
rect 596 2536 853 2544
rect 716 2527 724 2536
rect 867 2536 993 2544
rect 1087 2536 1353 2544
rect 1376 2544 1384 2556
rect 1527 2556 1613 2564
rect 1627 2556 1753 2564
rect 1827 2556 2093 2564
rect 2207 2556 2293 2564
rect 2327 2556 2384 2564
rect 1376 2536 1913 2544
rect 176 2516 253 2524
rect 1376 2524 1384 2536
rect 1947 2536 2013 2544
rect 2127 2536 2153 2544
rect 2267 2536 2353 2544
rect 2376 2544 2384 2556
rect 2427 2556 2453 2564
rect 2376 2536 2393 2544
rect 1247 2516 1384 2524
rect 1507 2516 1733 2524
rect 1747 2516 1793 2524
rect 1807 2516 1913 2524
rect 1927 2516 1944 2524
rect 27 2496 33 2504
rect 47 2496 693 2504
rect 1147 2496 1253 2504
rect 1287 2496 1653 2504
rect 1787 2496 1893 2504
rect 1936 2504 1944 2516
rect 2076 2524 2084 2533
rect 1967 2516 2084 2524
rect 2107 2516 2193 2524
rect 2216 2524 2224 2533
rect 2516 2527 2524 2593
rect 2656 2584 2664 2593
rect 2567 2576 2664 2584
rect 2536 2556 2593 2564
rect 2216 2516 2313 2524
rect 2356 2516 2393 2524
rect 1936 2496 2033 2504
rect 2356 2504 2364 2516
rect 2187 2496 2364 2504
rect 2536 2504 2544 2556
rect 2676 2564 2684 2596
rect 2767 2596 2993 2604
rect 3647 2596 3953 2604
rect 4407 2596 4733 2604
rect 4747 2596 4813 2604
rect 5087 2596 5913 2604
rect 5927 2596 6133 2604
rect 7187 2596 7293 2604
rect 7307 2596 7413 2604
rect 7436 2604 7444 2613
rect 7436 2596 7473 2604
rect 7507 2596 7584 2604
rect 2707 2576 2893 2584
rect 2947 2576 3013 2584
rect 3067 2576 3253 2584
rect 3307 2576 3333 2584
rect 3347 2576 3373 2584
rect 3396 2576 3473 2584
rect 2676 2556 2784 2564
rect 2776 2547 2784 2556
rect 2807 2556 2824 2564
rect 2816 2544 2824 2556
rect 2907 2556 3013 2564
rect 3276 2564 3284 2573
rect 3396 2564 3404 2576
rect 3627 2576 3653 2584
rect 3807 2576 4013 2584
rect 4187 2576 4253 2584
rect 4347 2576 4373 2584
rect 4447 2576 4473 2584
rect 4667 2576 4764 2584
rect 3127 2556 3284 2564
rect 3296 2556 3404 2564
rect 3296 2547 3304 2556
rect 3427 2556 3504 2564
rect 3496 2547 3504 2556
rect 3527 2556 3733 2564
rect 3867 2556 3953 2564
rect 3987 2556 4033 2564
rect 4476 2556 4633 2564
rect 2816 2536 3113 2544
rect 3127 2536 3173 2544
rect 3307 2536 3424 2544
rect 3416 2527 3424 2536
rect 3547 2536 3613 2544
rect 4476 2544 4484 2556
rect 4756 2564 4764 2576
rect 4787 2576 5064 2584
rect 4756 2556 4773 2564
rect 4787 2556 4833 2564
rect 4887 2556 4913 2564
rect 4956 2556 5033 2564
rect 4327 2536 4484 2544
rect 4676 2544 4684 2553
rect 4956 2544 4964 2556
rect 5056 2547 5064 2576
rect 5127 2576 5173 2584
rect 5367 2576 5433 2584
rect 5447 2576 5664 2584
rect 5107 2556 5133 2564
rect 5147 2556 5233 2564
rect 5307 2556 5453 2564
rect 5547 2556 5633 2564
rect 5656 2564 5664 2576
rect 5887 2576 5973 2584
rect 5987 2576 6093 2584
rect 6107 2576 6153 2584
rect 6467 2576 6573 2584
rect 6707 2576 6773 2584
rect 6827 2576 7133 2584
rect 7307 2576 7393 2584
rect 7576 2584 7584 2596
rect 7576 2576 7604 2584
rect 5656 2556 5833 2564
rect 4507 2536 4964 2544
rect 5156 2536 5233 2544
rect 2647 2516 2933 2524
rect 3887 2516 3973 2524
rect 4107 2516 4213 2524
rect 4327 2516 4353 2524
rect 4827 2516 4853 2524
rect 4976 2507 4984 2533
rect 5156 2527 5164 2536
rect 5387 2536 5473 2544
rect 5536 2544 5544 2553
rect 5656 2547 5664 2556
rect 5856 2556 5953 2564
rect 5856 2547 5864 2556
rect 6327 2556 6513 2564
rect 6567 2556 6673 2564
rect 7167 2556 7253 2564
rect 7327 2556 7353 2564
rect 7387 2556 7473 2564
rect 5487 2536 5544 2544
rect 5707 2536 5773 2544
rect 6556 2544 6564 2553
rect 6067 2536 6104 2544
rect 6556 2536 6593 2544
rect 5267 2516 5333 2524
rect 5927 2516 6033 2524
rect 6096 2507 6104 2536
rect 6716 2544 6724 2553
rect 6716 2536 6753 2544
rect 6967 2536 7193 2544
rect 7436 2536 7493 2544
rect 6447 2516 7073 2524
rect 7087 2516 7273 2524
rect 7347 2516 7393 2524
rect 2387 2496 2593 2504
rect 3407 2496 3433 2504
rect 5207 2496 5293 2504
rect 6587 2496 6653 2504
rect 6907 2496 7193 2504
rect 7247 2496 7313 2504
rect 7436 2504 7444 2536
rect 7596 2544 7604 2576
rect 7847 2576 7873 2584
rect 7627 2556 7673 2564
rect 7727 2556 7753 2564
rect 7596 2536 7624 2544
rect 7616 2527 7624 2536
rect 7467 2516 7493 2524
rect 7647 2516 7753 2524
rect 7387 2496 7444 2504
rect 347 2476 953 2484
rect 1587 2476 1753 2484
rect 1767 2476 2353 2484
rect 2367 2476 2433 2484
rect 2467 2476 2733 2484
rect 2767 2476 3313 2484
rect 3687 2476 4493 2484
rect 5027 2476 5273 2484
rect 7167 2476 7233 2484
rect 27 2456 393 2464
rect 907 2456 953 2464
rect 1227 2456 1733 2464
rect 1867 2456 2173 2464
rect 2287 2456 2613 2464
rect 3247 2456 3413 2464
rect 3587 2456 4193 2464
rect 5227 2456 5313 2464
rect 167 2436 753 2444
rect 827 2436 853 2444
rect 1347 2436 1773 2444
rect 1927 2436 2453 2444
rect 2496 2436 2573 2444
rect 227 2416 993 2424
rect 1067 2416 1704 2424
rect 367 2396 473 2404
rect 507 2396 1093 2404
rect 1127 2396 1393 2404
rect 1696 2404 1704 2416
rect 1727 2416 2053 2424
rect 2496 2424 2504 2436
rect 2607 2436 2873 2444
rect 2947 2436 3453 2444
rect 4087 2436 4113 2444
rect 4627 2436 4653 2444
rect 2407 2416 2504 2424
rect 2527 2416 2713 2424
rect 2787 2416 3073 2424
rect 3187 2416 3453 2424
rect 3507 2416 3593 2424
rect 4267 2416 4333 2424
rect 6507 2416 6533 2424
rect 1696 2396 1913 2404
rect 2047 2396 2293 2404
rect 2327 2396 2413 2404
rect 2467 2396 2593 2404
rect 2627 2396 2833 2404
rect 3067 2396 3313 2404
rect 3347 2396 3593 2404
rect 3687 2396 4053 2404
rect 407 2376 593 2384
rect 607 2376 1253 2384
rect 1276 2376 1633 2384
rect 747 2356 813 2364
rect 1276 2364 1284 2376
rect 1687 2376 1873 2384
rect 1987 2376 2053 2384
rect 2347 2376 2813 2384
rect 2827 2376 3053 2384
rect 3367 2376 4353 2384
rect 1167 2356 1284 2364
rect 1887 2356 1993 2364
rect 2027 2356 2173 2364
rect 2347 2356 2833 2364
rect 3087 2356 3113 2364
rect 3427 2356 3613 2364
rect 3807 2356 3833 2364
rect 3907 2356 3953 2364
rect 887 2336 973 2344
rect 1127 2336 1193 2344
rect 1387 2336 1533 2344
rect 1907 2336 2024 2344
rect 467 2316 553 2324
rect 576 2316 653 2324
rect 87 2296 133 2304
rect 187 2296 233 2304
rect 407 2296 524 2304
rect 516 2287 524 2296
rect 156 2276 273 2284
rect 156 2264 164 2276
rect 307 2276 384 2284
rect 376 2267 384 2276
rect 147 2256 164 2264
rect 227 2256 253 2264
rect 436 2264 444 2273
rect 436 2256 533 2264
rect 107 2236 413 2244
rect 556 2244 564 2273
rect 576 2247 584 2316
rect 847 2316 1033 2324
rect 1107 2316 1644 2324
rect 647 2296 773 2304
rect 807 2296 984 2304
rect 667 2276 813 2284
rect 867 2276 884 2284
rect 607 2256 713 2264
rect 727 2256 824 2264
rect 816 2247 824 2256
rect 876 2247 884 2276
rect 976 2264 984 2296
rect 1087 2296 1173 2304
rect 1487 2296 1564 2304
rect 996 2267 1004 2293
rect 1556 2287 1564 2296
rect 1636 2287 1644 2316
rect 1687 2316 1713 2324
rect 1807 2316 2004 2324
rect 1996 2307 2004 2316
rect 1656 2296 1693 2304
rect 1027 2276 1093 2284
rect 1207 2276 1413 2284
rect 1447 2276 1493 2284
rect 947 2256 984 2264
rect 1007 2256 1073 2264
rect 1327 2256 1373 2264
rect 1467 2256 1513 2264
rect 1656 2264 1664 2296
rect 1827 2296 1853 2304
rect 1867 2296 1913 2304
rect 1687 2276 1893 2284
rect 1587 2256 1664 2264
rect 1767 2256 1893 2264
rect 1956 2264 1964 2293
rect 2016 2287 2024 2336
rect 2147 2336 2433 2344
rect 2507 2336 2533 2344
rect 2547 2336 2793 2344
rect 2887 2336 3273 2344
rect 3307 2336 3793 2344
rect 5147 2336 5273 2344
rect 5727 2336 6673 2344
rect 6687 2336 6953 2344
rect 6967 2336 7253 2344
rect 7547 2336 7653 2344
rect 2167 2316 2473 2324
rect 2607 2316 3113 2324
rect 3127 2316 3133 2324
rect 3227 2316 3333 2324
rect 3387 2316 3873 2324
rect 4007 2316 4413 2324
rect 4567 2316 4573 2324
rect 4587 2316 4633 2324
rect 4707 2316 4733 2324
rect 4927 2316 5233 2324
rect 7347 2316 7433 2324
rect 7536 2316 7573 2324
rect 2047 2296 2093 2304
rect 2116 2296 2193 2304
rect 2116 2287 2124 2296
rect 2247 2296 2293 2304
rect 2387 2296 2404 2304
rect 2067 2276 2104 2284
rect 1956 2256 2053 2264
rect 2096 2264 2104 2276
rect 2187 2276 2213 2284
rect 2396 2284 2404 2296
rect 2427 2296 2493 2304
rect 2567 2296 2753 2304
rect 3127 2296 3253 2304
rect 3327 2296 3473 2304
rect 3556 2296 3913 2304
rect 2396 2276 2473 2284
rect 2527 2276 2593 2284
rect 2767 2276 2813 2284
rect 2847 2276 3153 2284
rect 3167 2276 3233 2284
rect 3276 2276 3373 2284
rect 2096 2256 2233 2264
rect 2267 2256 2293 2264
rect 2676 2264 2684 2273
rect 2587 2256 2684 2264
rect 2707 2256 2993 2264
rect 3067 2256 3093 2264
rect 3276 2264 3284 2276
rect 3556 2284 3564 2296
rect 4267 2296 4693 2304
rect 4707 2296 5053 2304
rect 5107 2296 5133 2304
rect 5567 2296 5653 2304
rect 5667 2296 5693 2304
rect 5827 2296 5873 2304
rect 6147 2296 6193 2304
rect 6387 2296 6453 2304
rect 6867 2296 6973 2304
rect 7067 2296 7133 2304
rect 7327 2296 7473 2304
rect 7487 2296 7513 2304
rect 3467 2276 3564 2284
rect 3556 2267 3564 2276
rect 3627 2276 3913 2284
rect 3936 2276 4013 2284
rect 3936 2267 3944 2276
rect 4067 2276 4113 2284
rect 4136 2267 4144 2293
rect 4287 2276 4593 2284
rect 5087 2276 5153 2284
rect 5207 2276 5253 2284
rect 5587 2276 5613 2284
rect 5736 2284 5744 2293
rect 5736 2276 5793 2284
rect 5856 2276 6013 2284
rect 3147 2256 3284 2264
rect 3307 2256 3393 2264
rect 3436 2256 3513 2264
rect 547 2236 564 2244
rect 627 2236 793 2244
rect 1287 2236 1613 2244
rect 1627 2236 1964 2244
rect 167 2216 293 2224
rect 347 2216 413 2224
rect 447 2216 613 2224
rect 647 2216 773 2224
rect 867 2216 933 2224
rect 947 2216 1133 2224
rect 1247 2216 1273 2224
rect 1467 2216 1684 2224
rect 247 2196 273 2204
rect 507 2196 633 2204
rect 687 2196 713 2204
rect 747 2196 873 2204
rect 907 2196 1084 2204
rect 227 2176 393 2184
rect 407 2176 493 2184
rect 556 2176 693 2184
rect 127 2156 233 2164
rect 556 2164 564 2176
rect 767 2176 793 2184
rect 847 2176 973 2184
rect 1076 2184 1084 2196
rect 1167 2196 1193 2204
rect 1267 2196 1453 2204
rect 1507 2196 1653 2204
rect 1676 2204 1684 2216
rect 1827 2216 1873 2224
rect 1956 2224 1964 2236
rect 1987 2236 2393 2244
rect 2447 2236 2473 2244
rect 2547 2236 2573 2244
rect 2587 2236 2633 2244
rect 2656 2236 2933 2244
rect 1956 2216 2373 2224
rect 2656 2224 2664 2236
rect 2967 2236 3113 2244
rect 3247 2236 3353 2244
rect 3436 2244 3444 2256
rect 3747 2256 3793 2264
rect 3976 2256 4093 2264
rect 3387 2236 3444 2244
rect 3616 2244 3624 2253
rect 3467 2236 3624 2244
rect 3976 2244 3984 2256
rect 3827 2236 3984 2244
rect 4007 2236 4193 2244
rect 4216 2227 4224 2273
rect 4287 2256 4353 2264
rect 4967 2256 5033 2264
rect 5407 2256 5593 2264
rect 5856 2264 5864 2276
rect 6127 2276 6233 2284
rect 6287 2276 6333 2284
rect 6487 2276 6813 2284
rect 6996 2284 7004 2293
rect 6947 2276 7004 2284
rect 7036 2284 7044 2293
rect 7536 2287 7544 2316
rect 7607 2316 7633 2324
rect 7567 2296 7584 2304
rect 7036 2276 7144 2284
rect 5727 2256 5864 2264
rect 5887 2256 6293 2264
rect 6667 2256 6753 2264
rect 6787 2256 7113 2264
rect 7136 2264 7144 2276
rect 7187 2276 7293 2284
rect 7576 2267 7584 2296
rect 7807 2296 7893 2304
rect 7867 2276 7893 2284
rect 7136 2256 7153 2264
rect 7367 2256 7453 2264
rect 4307 2236 4553 2244
rect 4827 2236 5173 2244
rect 5587 2236 5613 2244
rect 5647 2236 5793 2244
rect 6227 2236 6373 2244
rect 6387 2236 6813 2244
rect 6827 2236 6873 2244
rect 6987 2236 7013 2244
rect 2407 2216 2664 2224
rect 2687 2216 3173 2224
rect 3187 2216 3253 2224
rect 3327 2216 3433 2224
rect 3547 2216 3853 2224
rect 3907 2216 4204 2224
rect 1676 2196 1853 2204
rect 1947 2196 2073 2204
rect 2107 2196 2533 2204
rect 2667 2196 2873 2204
rect 2887 2196 3373 2204
rect 3447 2196 3604 2204
rect 1076 2176 1113 2184
rect 1127 2176 1333 2184
rect 1607 2176 1793 2184
rect 1927 2176 2373 2184
rect 2427 2176 2953 2184
rect 2976 2176 3393 2184
rect 287 2156 564 2164
rect 587 2156 664 2164
rect -4 2136 73 2144
rect -4 2044 4 2136
rect 167 2136 593 2144
rect 656 2144 664 2156
rect 687 2156 953 2164
rect 1007 2156 1393 2164
rect 1707 2156 1753 2164
rect 1807 2156 1993 2164
rect 2087 2156 2193 2164
rect 2267 2156 2293 2164
rect 2367 2156 2453 2164
rect 2467 2156 2653 2164
rect 2707 2156 2744 2164
rect 656 2136 853 2144
rect 1027 2136 1213 2144
rect 1307 2136 1353 2144
rect 1627 2136 1833 2144
rect 1867 2136 2053 2144
rect 2147 2136 2173 2144
rect 2247 2136 2313 2144
rect 2736 2144 2744 2156
rect 2827 2156 2913 2164
rect 2976 2164 2984 2176
rect 3547 2176 3573 2184
rect 3596 2184 3604 2196
rect 3627 2196 4113 2204
rect 4196 2204 4204 2216
rect 5007 2216 5133 2224
rect 5147 2216 5213 2224
rect 6007 2216 6253 2224
rect 6867 2216 7393 2224
rect 7747 2216 7853 2224
rect 4196 2196 4333 2204
rect 3596 2176 3853 2184
rect 3927 2176 4333 2184
rect 4387 2176 4513 2184
rect 6127 2176 6513 2184
rect 2967 2156 2984 2164
rect 3167 2156 3193 2164
rect 3487 2156 3713 2164
rect 3956 2156 4293 2164
rect 2736 2136 3053 2144
rect 3127 2136 3693 2144
rect 3707 2136 3833 2144
rect 3956 2144 3964 2156
rect 4527 2156 4573 2164
rect 7047 2156 7413 2164
rect 3847 2136 3964 2144
rect 3987 2136 4093 2144
rect 4307 2136 4433 2144
rect 6647 2136 6993 2144
rect 7007 2136 7133 2144
rect 7147 2136 7233 2144
rect 7247 2136 7673 2144
rect 7687 2136 7773 2144
rect 16 2116 73 2124
rect 16 2064 24 2116
rect 127 2116 173 2124
rect 367 2116 493 2124
rect 596 2116 653 2124
rect 67 2096 84 2104
rect 36 2084 44 2093
rect 36 2076 64 2084
rect 56 2067 64 2076
rect 16 2056 33 2064
rect 76 2047 84 2096
rect 136 2096 253 2104
rect 136 2067 144 2096
rect 287 2096 304 2104
rect 296 2087 304 2096
rect 387 2096 484 2104
rect 476 2087 484 2096
rect 247 2076 284 2084
rect 276 2067 284 2076
rect 447 2076 464 2084
rect 456 2067 464 2076
rect 476 2064 484 2073
rect 596 2067 604 2116
rect 767 2116 833 2124
rect 947 2116 1093 2124
rect 1127 2116 1153 2124
rect 1307 2116 1413 2124
rect 1447 2116 1593 2124
rect 1647 2116 2253 2124
rect 2676 2116 2853 2124
rect 2676 2107 2684 2116
rect 2867 2116 3013 2124
rect 3087 2116 3233 2124
rect 3287 2116 3433 2124
rect 3476 2116 3573 2124
rect 627 2096 793 2104
rect 887 2096 973 2104
rect 1047 2096 1073 2104
rect 1127 2096 1344 2104
rect 627 2076 684 2084
rect 476 2056 544 2064
rect -4 2036 64 2044
rect 56 2024 64 2036
rect 236 2044 244 2053
rect 107 2036 293 2044
rect 307 2036 313 2044
rect 336 2044 344 2053
rect 336 2036 513 2044
rect 56 2016 253 2024
rect 367 2016 453 2024
rect 536 2024 544 2056
rect 676 2047 684 2076
rect 996 2084 1004 2093
rect 1336 2087 1344 2096
rect 1587 2096 1653 2104
rect 1667 2096 1713 2104
rect 1776 2096 1813 2104
rect 707 2076 1004 2084
rect 1487 2076 1513 2084
rect 707 2056 733 2064
rect 967 2056 993 2064
rect 1056 2064 1064 2073
rect 1056 2056 1093 2064
rect 867 2036 913 2044
rect 1256 2044 1264 2073
rect 1396 2047 1404 2073
rect 1567 2056 1633 2064
rect 1676 2064 1684 2073
rect 1676 2056 1693 2064
rect 1227 2036 1264 2044
rect 1716 2044 1724 2073
rect 1547 2036 1744 2044
rect 536 2016 773 2024
rect 847 2016 973 2024
rect 1007 2016 1693 2024
rect 1736 2024 1744 2036
rect 1776 2044 1784 2096
rect 1947 2096 2033 2104
rect 2047 2096 2413 2104
rect 2447 2096 2553 2104
rect 2747 2096 2904 2104
rect 1856 2084 1864 2093
rect 1856 2076 2013 2084
rect 2027 2076 2113 2084
rect 2136 2076 2273 2084
rect 1836 2064 1844 2073
rect 1836 2056 1873 2064
rect 2136 2064 2144 2076
rect 2436 2076 2473 2084
rect 1896 2056 2144 2064
rect 1767 2036 1784 2044
rect 1896 2044 1904 2056
rect 2436 2064 2444 2076
rect 2527 2076 2604 2084
rect 2247 2056 2444 2064
rect 2467 2056 2564 2064
rect 2556 2047 2564 2056
rect 1807 2036 1904 2044
rect 2187 2036 2513 2044
rect 2596 2044 2604 2076
rect 2896 2084 2904 2096
rect 2927 2096 3073 2104
rect 3287 2096 3413 2104
rect 3476 2104 3484 2116
rect 3607 2116 3973 2124
rect 3987 2116 4013 2124
rect 4047 2116 4153 2124
rect 5127 2116 5173 2124
rect 6227 2116 6393 2124
rect 6547 2116 6633 2124
rect 6647 2116 6893 2124
rect 6776 2107 6784 2116
rect 7307 2116 7373 2124
rect 7387 2116 7513 2124
rect 7607 2116 7713 2124
rect 3447 2096 3484 2104
rect 3507 2096 3593 2104
rect 3667 2096 3713 2104
rect 3747 2096 3993 2104
rect 4507 2096 4613 2104
rect 4647 2096 4773 2104
rect 4787 2096 4993 2104
rect 5007 2096 5433 2104
rect 5447 2096 5713 2104
rect 5727 2096 5953 2104
rect 6367 2096 6413 2104
rect 6727 2096 6733 2104
rect 6747 2096 6753 2104
rect 6987 2096 7473 2104
rect 7856 2096 7873 2104
rect 2647 2076 2884 2084
rect 2896 2076 2944 2084
rect 2627 2056 2673 2064
rect 2816 2056 2853 2064
rect 2816 2044 2824 2056
rect 2876 2064 2884 2076
rect 2936 2067 2944 2076
rect 3027 2076 3193 2084
rect 3216 2076 3313 2084
rect 2876 2056 2924 2064
rect 2596 2036 2824 2044
rect 2847 2036 2893 2044
rect 2916 2044 2924 2056
rect 3216 2064 3224 2076
rect 3467 2076 3513 2084
rect 4036 2076 4193 2084
rect 3027 2056 3224 2064
rect 3407 2056 3453 2064
rect 3656 2064 3664 2073
rect 3567 2056 3664 2064
rect 3776 2064 3784 2073
rect 3707 2056 3784 2064
rect 3956 2047 3964 2073
rect 4036 2067 4044 2076
rect 4207 2076 4413 2084
rect 4447 2076 4673 2084
rect 5147 2076 5213 2084
rect 5767 2076 5953 2084
rect 5976 2076 6173 2084
rect 5976 2067 5984 2076
rect 6196 2076 6293 2084
rect 6196 2067 6204 2076
rect 6347 2076 6373 2084
rect 6427 2076 6593 2084
rect 6807 2076 7053 2084
rect 7287 2076 7433 2084
rect 4187 2056 4233 2064
rect 4407 2056 4493 2064
rect 5107 2056 5153 2064
rect 5207 2056 5273 2064
rect 5387 2056 5453 2064
rect 5887 2056 5933 2064
rect 6027 2056 6073 2064
rect 6627 2056 6733 2064
rect 7067 2056 7413 2064
rect 7467 2056 7633 2064
rect 7787 2056 7833 2064
rect 7856 2047 7864 2096
rect 7896 2047 7904 2073
rect 2916 2036 2993 2044
rect 3127 2036 3793 2044
rect 3807 2036 3933 2044
rect 4027 2036 4053 2044
rect 4227 2036 4273 2044
rect 4527 2036 4853 2044
rect 5227 2036 5293 2044
rect 5487 2036 5633 2044
rect 5647 2036 5833 2044
rect 6327 2036 6333 2044
rect 6347 2036 6493 2044
rect 6727 2036 6873 2044
rect 6887 2036 6913 2044
rect 7027 2036 7153 2044
rect 7507 2036 7533 2044
rect 1736 2016 2133 2024
rect 2507 2016 2813 2024
rect 3007 2016 3353 2024
rect 3527 2016 3593 2024
rect 3607 2016 3633 2024
rect 3867 2016 4033 2024
rect 5287 2016 5433 2024
rect 5447 2016 5773 2024
rect 5787 2016 6053 2024
rect 467 1996 833 2004
rect 947 1996 1253 2004
rect 1447 1996 1733 2004
rect 1747 1996 1993 2004
rect 2127 1996 2413 2004
rect 2447 1996 2613 2004
rect 2787 1996 2833 2004
rect 2867 1996 3444 2004
rect 287 1976 653 1984
rect 727 1976 1033 1984
rect 1176 1976 1373 1984
rect 1176 1967 1184 1976
rect 1476 1976 1493 1984
rect 387 1956 533 1964
rect 707 1956 1153 1964
rect 1476 1964 1484 1976
rect 1607 1976 1773 1984
rect 1827 1976 2053 1984
rect 2067 1976 2333 1984
rect 2547 1976 2733 1984
rect 3247 1976 3293 1984
rect 3436 1984 3444 1996
rect 3467 1996 3733 2004
rect 4047 1996 4073 2004
rect 4327 1996 4393 2004
rect 4407 1996 5333 2004
rect 5347 1996 6393 2004
rect 3436 1976 3613 1984
rect 3667 1976 3953 1984
rect 4027 1976 4353 1984
rect 5167 1976 5573 1984
rect 5927 1976 6233 1984
rect 6487 1976 6593 1984
rect 6607 1976 6653 1984
rect 1327 1956 1484 1964
rect 1507 1956 1913 1964
rect 1967 1956 2653 1964
rect 2687 1956 2753 1964
rect 3747 1956 3893 1964
rect 4947 1956 5013 1964
rect 227 1936 1473 1944
rect 1487 1936 1553 1944
rect 1827 1936 2153 1944
rect 2167 1936 2713 1944
rect 3567 1936 3833 1944
rect 87 1916 213 1924
rect 307 1916 733 1924
rect 747 1916 1013 1924
rect 1267 1916 1573 1924
rect 1707 1916 1953 1924
rect 2007 1916 2173 1924
rect 2387 1916 2473 1924
rect 2487 1916 2793 1924
rect 2807 1916 3113 1924
rect 3187 1916 3333 1924
rect 7896 1907 7904 1933
rect 207 1896 273 1904
rect 487 1896 593 1904
rect 727 1896 3913 1904
rect 547 1876 1413 1884
rect 1527 1876 1893 1884
rect 1947 1876 2073 1884
rect 2127 1876 2453 1884
rect 2527 1876 3513 1884
rect 4367 1876 4653 1884
rect 5647 1876 6013 1884
rect 6747 1876 7193 1884
rect 7227 1876 7573 1884
rect 527 1856 613 1864
rect 887 1856 1473 1864
rect 1587 1856 1853 1864
rect 1907 1856 2013 1864
rect 2067 1856 2153 1864
rect 2227 1856 2373 1864
rect 2427 1856 3573 1864
rect 3807 1856 4133 1864
rect 4247 1856 4453 1864
rect 6007 1856 6053 1864
rect 6207 1856 6793 1864
rect 6947 1856 7413 1864
rect 7427 1856 7573 1864
rect 487 1836 513 1844
rect 787 1836 993 1844
rect 1147 1836 1313 1844
rect 1387 1836 1593 1844
rect 1707 1836 1753 1844
rect 2187 1836 2313 1844
rect 2327 1836 2813 1844
rect 2827 1836 3253 1844
rect 3347 1836 3713 1844
rect 4176 1836 4293 1844
rect 47 1816 453 1824
rect 567 1816 793 1824
rect 827 1816 913 1824
rect 936 1816 1133 1824
rect 507 1796 573 1804
rect 667 1796 693 1804
rect 936 1804 944 1816
rect 1476 1816 1513 1824
rect 827 1796 944 1804
rect 1007 1796 1093 1804
rect 1156 1796 1233 1804
rect 107 1776 173 1784
rect 327 1776 493 1784
rect 567 1776 584 1784
rect 147 1756 373 1764
rect 387 1756 553 1764
rect 576 1764 584 1776
rect 576 1756 753 1764
rect 816 1764 824 1793
rect 847 1776 884 1784
rect 816 1756 833 1764
rect 876 1764 884 1776
rect 907 1776 1013 1784
rect 1047 1776 1073 1784
rect 1136 1784 1144 1793
rect 1156 1787 1164 1796
rect 1336 1787 1344 1813
rect 1116 1776 1144 1784
rect 876 1756 953 1764
rect 1116 1764 1124 1776
rect 1476 1767 1484 1816
rect 1536 1816 1553 1824
rect 1536 1784 1544 1816
rect 1627 1816 1653 1824
rect 1807 1816 1833 1824
rect 2067 1816 2213 1824
rect 2227 1816 2473 1824
rect 2527 1816 2633 1824
rect 2907 1816 2993 1824
rect 3007 1816 3113 1824
rect 3267 1816 3433 1824
rect 3647 1816 3673 1824
rect 3707 1816 3753 1824
rect 3907 1816 3973 1824
rect 1576 1804 1584 1813
rect 4176 1807 4184 1836
rect 4427 1836 4593 1844
rect 4676 1836 4813 1844
rect 4327 1816 4653 1824
rect 1567 1796 1584 1804
rect 1627 1796 1724 1804
rect 1716 1787 1724 1796
rect 1776 1796 1913 1804
rect 1776 1787 1784 1796
rect 2007 1796 2313 1804
rect 2347 1796 2444 1804
rect 1536 1776 1573 1784
rect 1647 1776 1673 1784
rect 2047 1776 2253 1784
rect 1107 1756 1124 1764
rect 1227 1756 1293 1764
rect 1307 1756 1393 1764
rect 1527 1756 1593 1764
rect 1647 1756 1813 1764
rect 1947 1756 2033 1764
rect 2047 1756 2133 1764
rect 2307 1756 2353 1764
rect 2367 1756 2393 1764
rect 2436 1764 2444 1796
rect 2567 1796 2584 1804
rect 2576 1787 2584 1796
rect 2727 1796 2773 1804
rect 2867 1796 2933 1804
rect 3327 1796 3353 1804
rect 3427 1796 3464 1804
rect 2467 1776 2493 1784
rect 2587 1776 2693 1784
rect 2887 1776 3013 1784
rect 3136 1784 3144 1793
rect 3047 1776 3144 1784
rect 3287 1776 3393 1784
rect 3456 1784 3464 1796
rect 3487 1796 3513 1804
rect 3547 1796 3564 1804
rect 3456 1776 3473 1784
rect 2436 1756 2493 1764
rect 2547 1756 2833 1764
rect 2927 1756 3213 1764
rect 3227 1756 3253 1764
rect 3556 1764 3564 1796
rect 3716 1796 3733 1804
rect 3587 1776 3673 1784
rect 3556 1756 3573 1764
rect 3716 1764 3724 1796
rect 3767 1796 3853 1804
rect 3867 1796 3953 1804
rect 4196 1804 4204 1813
rect 4676 1807 4684 1836
rect 5767 1836 6013 1844
rect 6067 1836 6433 1844
rect 6567 1836 6873 1844
rect 7347 1836 7473 1844
rect 4707 1816 4913 1824
rect 4927 1816 4973 1824
rect 5027 1816 5053 1824
rect 5067 1816 5293 1824
rect 5387 1816 5413 1824
rect 5527 1816 5553 1824
rect 5567 1816 5673 1824
rect 5687 1816 6253 1824
rect 6387 1816 6513 1824
rect 6527 1816 6753 1824
rect 6847 1816 6893 1824
rect 7327 1816 7533 1824
rect 7627 1816 7653 1824
rect 4196 1796 4273 1804
rect 4527 1796 4573 1804
rect 4696 1796 4733 1804
rect 3987 1776 4013 1784
rect 4476 1784 4484 1793
rect 4087 1776 4484 1784
rect 4696 1784 4704 1796
rect 4967 1796 4993 1804
rect 5407 1796 5433 1804
rect 5487 1796 5573 1804
rect 5587 1796 5853 1804
rect 6087 1796 6113 1804
rect 6247 1796 6324 1804
rect 4607 1776 4704 1784
rect 4787 1776 4813 1784
rect 4827 1776 5173 1784
rect 5227 1776 5253 1784
rect 3667 1756 3724 1764
rect 3747 1756 3833 1764
rect 3847 1756 3893 1764
rect 3907 1756 3933 1764
rect 3967 1756 4053 1764
rect 4507 1756 4673 1764
rect 4867 1756 5333 1764
rect 5356 1764 5364 1793
rect 6316 1787 6324 1796
rect 6467 1796 6493 1804
rect 6547 1796 6593 1804
rect 6647 1796 6693 1804
rect 7007 1796 7053 1804
rect 7107 1796 7244 1804
rect 5387 1776 5453 1784
rect 5907 1776 6033 1784
rect 6047 1776 6093 1784
rect 6147 1776 6193 1784
rect 6436 1784 6444 1793
rect 7236 1787 7244 1796
rect 7467 1796 7553 1804
rect 7567 1796 7653 1804
rect 7707 1796 7753 1804
rect 7867 1796 7884 1804
rect 7876 1787 7884 1796
rect 6436 1776 6653 1784
rect 7256 1776 7333 1784
rect 7256 1767 7264 1776
rect 5356 1756 5533 1764
rect 5727 1756 5833 1764
rect 5847 1756 5953 1764
rect 6307 1756 6373 1764
rect 6467 1756 6493 1764
rect 6667 1756 6773 1764
rect 7087 1756 7113 1764
rect 7127 1756 7153 1764
rect 7187 1756 7233 1764
rect 7287 1756 7313 1764
rect 7347 1756 7533 1764
rect 7787 1756 7873 1764
rect 227 1736 333 1744
rect 407 1736 513 1744
rect 667 1736 753 1744
rect 787 1736 913 1744
rect 1087 1736 1333 1744
rect 1667 1736 1733 1744
rect 1787 1736 2013 1744
rect 2067 1736 2193 1744
rect 2207 1736 2273 1744
rect 2347 1736 2544 1744
rect 167 1716 473 1724
rect 487 1716 893 1724
rect 1127 1716 1273 1724
rect 1307 1716 1793 1724
rect 1887 1716 1893 1724
rect 1907 1716 2213 1724
rect 2307 1716 2373 1724
rect 2407 1716 2513 1724
rect 2536 1724 2544 1736
rect 2587 1736 3153 1744
rect 3207 1736 3533 1744
rect 3607 1736 3633 1744
rect 3767 1736 3793 1744
rect 3887 1736 4093 1744
rect 4307 1736 4413 1744
rect 5027 1736 5313 1744
rect 5827 1736 5893 1744
rect 7207 1736 7293 1744
rect 7347 1736 7373 1744
rect 7387 1736 7393 1744
rect 7607 1736 7673 1744
rect 2536 1716 2713 1724
rect 2787 1716 2873 1724
rect 2887 1716 2893 1724
rect 2947 1716 3473 1724
rect 3547 1716 3613 1724
rect 3787 1716 4033 1724
rect 4267 1716 4633 1724
rect 5607 1716 6413 1724
rect 7647 1716 7673 1724
rect 7687 1716 7853 1724
rect 307 1696 413 1704
rect 687 1696 853 1704
rect 867 1696 913 1704
rect 947 1696 1053 1704
rect 1107 1696 1133 1704
rect 1207 1696 1293 1704
rect 1427 1696 1973 1704
rect 1987 1696 2113 1704
rect 2127 1696 2153 1704
rect 2507 1696 2793 1704
rect 2967 1696 3313 1704
rect 3567 1696 3613 1704
rect 3887 1696 4033 1704
rect 4047 1696 4073 1704
rect 4107 1696 4353 1704
rect 4727 1696 4753 1704
rect 5607 1696 6573 1704
rect 87 1676 453 1684
rect 707 1676 953 1684
rect 1167 1676 1313 1684
rect 1336 1676 1653 1684
rect 267 1656 413 1664
rect 727 1656 813 1664
rect 1336 1664 1344 1676
rect 1667 1676 1993 1684
rect 2447 1676 2533 1684
rect 2607 1676 2753 1684
rect 2867 1676 3033 1684
rect 3047 1676 3633 1684
rect 4087 1676 4233 1684
rect 4647 1676 5753 1684
rect 5767 1676 5933 1684
rect 6167 1676 6273 1684
rect 6287 1676 7033 1684
rect 987 1656 1344 1664
rect 1607 1656 1753 1664
rect 1807 1656 2073 1664
rect 2087 1656 2233 1664
rect 2267 1656 2553 1664
rect 2667 1656 2993 1664
rect 3127 1656 3153 1664
rect 3227 1656 3553 1664
rect 4147 1656 4193 1664
rect 4207 1656 4453 1664
rect 4567 1656 5273 1664
rect 5707 1656 5973 1664
rect 5987 1656 6213 1664
rect 6347 1656 6473 1664
rect 6507 1656 6633 1664
rect 6667 1656 6713 1664
rect 7407 1656 7473 1664
rect 87 1636 533 1644
rect 547 1636 733 1644
rect 767 1636 1073 1644
rect 1087 1636 1384 1644
rect 67 1616 93 1624
rect 247 1616 313 1624
rect 327 1616 333 1624
rect 367 1616 433 1624
rect 847 1616 873 1624
rect 947 1616 1013 1624
rect 1207 1616 1353 1624
rect 1376 1624 1384 1636
rect 1407 1636 1693 1644
rect 2007 1636 2473 1644
rect 2547 1636 2673 1644
rect 2747 1636 2793 1644
rect 3027 1636 3233 1644
rect 3287 1636 3673 1644
rect 4167 1636 4273 1644
rect 4367 1636 4813 1644
rect 5307 1636 5513 1644
rect 5947 1636 5953 1644
rect 5967 1636 6073 1644
rect 6087 1636 6133 1644
rect 6607 1636 6673 1644
rect 6687 1636 6713 1644
rect 7047 1636 7053 1644
rect 7067 1636 7133 1644
rect 7467 1636 7513 1644
rect 7807 1636 7884 1644
rect 1376 1616 1413 1624
rect 1427 1616 1533 1624
rect 1547 1616 1664 1624
rect 267 1596 373 1604
rect 527 1596 593 1604
rect 647 1596 693 1604
rect 736 1596 873 1604
rect 176 1584 184 1593
rect 147 1576 184 1584
rect 207 1576 393 1584
rect 507 1576 633 1584
rect 187 1556 293 1564
rect 367 1556 453 1564
rect 107 1536 233 1544
rect 716 1544 724 1573
rect 736 1567 744 1596
rect 1227 1596 1433 1604
rect 1656 1604 1664 1616
rect 1687 1616 1713 1624
rect 1847 1616 1933 1624
rect 2227 1616 2453 1624
rect 2487 1616 2573 1624
rect 2607 1616 2813 1624
rect 2847 1616 3053 1624
rect 3147 1616 3264 1624
rect 1547 1596 1584 1604
rect 1656 1596 1693 1604
rect 907 1576 953 1584
rect 816 1564 824 1573
rect 796 1556 824 1564
rect 796 1544 804 1556
rect 716 1536 804 1544
rect 827 1536 853 1544
rect 976 1544 984 1593
rect 1367 1576 1413 1584
rect 1467 1576 1553 1584
rect 1576 1584 1584 1596
rect 1707 1596 1753 1604
rect 1827 1596 2013 1604
rect 2047 1596 2133 1604
rect 2307 1596 2444 1604
rect 1576 1576 1673 1584
rect 1727 1576 1793 1584
rect 2347 1576 2413 1584
rect 2436 1584 2444 1596
rect 2747 1596 2893 1604
rect 2907 1596 2933 1604
rect 3067 1596 3084 1604
rect 3076 1587 3084 1596
rect 3256 1587 3264 1616
rect 3387 1616 3433 1624
rect 3447 1616 3493 1624
rect 3707 1616 3853 1624
rect 4127 1616 4533 1624
rect 4547 1616 4833 1624
rect 5327 1616 5393 1624
rect 5407 1616 5413 1624
rect 5787 1616 5833 1624
rect 5847 1616 5873 1624
rect 6087 1616 6173 1624
rect 6187 1616 6233 1624
rect 6567 1616 6613 1624
rect 6907 1616 6953 1624
rect 6967 1616 7233 1624
rect 7247 1616 7373 1624
rect 7447 1616 7493 1624
rect 3407 1596 3433 1604
rect 3447 1596 3453 1604
rect 3507 1596 3553 1604
rect 3847 1596 3893 1604
rect 4127 1596 4273 1604
rect 4327 1596 4353 1604
rect 4527 1596 4613 1604
rect 4636 1596 4673 1604
rect 2436 1576 2873 1584
rect 3007 1576 3064 1584
rect 1007 1556 1613 1564
rect 1627 1556 1813 1564
rect 2276 1564 2284 1573
rect 1847 1556 2353 1564
rect 2547 1556 2573 1564
rect 2596 1556 3033 1564
rect 976 1536 1033 1544
rect 1067 1536 1353 1544
rect 1476 1536 2173 1544
rect 787 1516 833 1524
rect 1476 1524 1484 1536
rect 2596 1544 2604 1556
rect 3056 1564 3064 1576
rect 3307 1576 3593 1584
rect 3636 1584 3644 1593
rect 3636 1576 3913 1584
rect 4027 1576 4033 1584
rect 4047 1576 4133 1584
rect 4347 1576 4573 1584
rect 4636 1584 4644 1596
rect 5416 1596 5613 1604
rect 4587 1576 4644 1584
rect 4656 1576 4713 1584
rect 4656 1567 4664 1576
rect 4767 1576 4973 1584
rect 5087 1576 5113 1584
rect 5136 1576 5193 1584
rect 3056 1556 3293 1564
rect 2327 1536 2604 1544
rect 3056 1544 3064 1556
rect 3487 1556 3533 1564
rect 4147 1556 4213 1564
rect 4407 1556 4433 1564
rect 4487 1556 4513 1564
rect 4527 1556 4533 1564
rect 4887 1556 4933 1564
rect 5136 1564 5144 1576
rect 5416 1584 5424 1596
rect 5807 1596 5853 1604
rect 5907 1596 5993 1604
rect 6407 1596 6773 1604
rect 7027 1596 7273 1604
rect 7296 1596 7413 1604
rect 5307 1576 5424 1584
rect 5447 1576 5553 1584
rect 5656 1567 5664 1593
rect 7296 1587 7304 1596
rect 7476 1587 7484 1616
rect 7667 1616 7693 1624
rect 7727 1616 7733 1624
rect 7747 1616 7853 1624
rect 7587 1596 7784 1604
rect 7776 1587 7784 1596
rect 7876 1604 7884 1636
rect 7856 1596 7884 1604
rect 5727 1576 5753 1584
rect 5887 1576 5933 1584
rect 6027 1576 6053 1584
rect 6447 1576 6573 1584
rect 7207 1576 7253 1584
rect 7387 1576 7433 1584
rect 7547 1576 7573 1584
rect 7587 1576 7633 1584
rect 7836 1584 7844 1593
rect 7856 1587 7864 1596
rect 7807 1576 7844 1584
rect 4947 1556 5144 1564
rect 5187 1556 5253 1564
rect 5347 1556 5413 1564
rect 5887 1556 5913 1564
rect 6687 1556 6733 1564
rect 7347 1556 7553 1564
rect 7707 1556 7753 1564
rect 7847 1556 7893 1564
rect 2627 1536 3064 1544
rect 5087 1536 5333 1544
rect 5407 1536 5453 1544
rect 5567 1536 6553 1544
rect 6567 1536 6693 1544
rect 7147 1536 7153 1544
rect 7167 1536 7373 1544
rect 1147 1516 1484 1524
rect 1827 1516 2333 1524
rect 2367 1516 2613 1524
rect 2667 1516 2693 1524
rect 2767 1516 3073 1524
rect 227 1496 533 1504
rect 547 1496 873 1504
rect 1376 1496 1833 1504
rect 1376 1484 1384 1496
rect 2207 1496 2573 1504
rect 2827 1496 3213 1504
rect 5467 1496 5573 1504
rect 207 1476 1384 1484
rect 1607 1476 1953 1484
rect 1987 1476 2413 1484
rect 2587 1476 3413 1484
rect 3427 1476 3513 1484
rect 5087 1476 5293 1484
rect 5687 1476 5873 1484
rect 407 1456 793 1464
rect 867 1456 1293 1464
rect 1347 1456 1493 1464
rect 1947 1456 2033 1464
rect 2047 1456 2253 1464
rect 2347 1456 2373 1464
rect 2667 1456 2864 1464
rect 2856 1447 2864 1456
rect 3127 1456 4773 1464
rect 4867 1456 5693 1464
rect 587 1436 893 1444
rect 1187 1436 1333 1444
rect 1367 1436 1973 1444
rect 2207 1436 2233 1444
rect 2247 1436 2313 1444
rect 2607 1436 2833 1444
rect 2867 1436 4093 1444
rect 4247 1436 5093 1444
rect 167 1416 433 1424
rect 1147 1416 1933 1424
rect 2367 1416 2753 1424
rect 2807 1416 2913 1424
rect 2987 1416 3673 1424
rect 267 1396 853 1404
rect 1867 1396 2373 1404
rect 2656 1396 4253 1404
rect 467 1376 593 1384
rect 607 1376 693 1384
rect 727 1376 1613 1384
rect 1747 1376 1933 1384
rect 2656 1384 2664 1396
rect 4447 1396 4593 1404
rect 2247 1376 2664 1384
rect 2687 1376 2733 1384
rect 2767 1376 3113 1384
rect 3187 1376 3253 1384
rect 4607 1376 4813 1384
rect 5187 1376 5213 1384
rect 5616 1376 6093 1384
rect 576 1356 624 1364
rect 576 1344 584 1356
rect 556 1336 584 1344
rect 556 1327 564 1336
rect 487 1316 513 1324
rect 87 1296 213 1304
rect 347 1296 533 1304
rect 596 1304 604 1333
rect 616 1327 624 1356
rect 947 1356 973 1364
rect 1067 1356 1233 1364
rect 1327 1356 1453 1364
rect 1687 1356 2173 1364
rect 2427 1356 2513 1364
rect 2596 1356 3453 1364
rect 887 1336 933 1344
rect 1027 1336 1084 1344
rect 787 1316 1053 1324
rect 1076 1324 1084 1336
rect 1247 1336 1373 1344
rect 1667 1336 1713 1344
rect 1787 1336 1813 1344
rect 2596 1344 2604 1356
rect 3547 1356 3953 1364
rect 4527 1356 4733 1364
rect 4747 1356 4933 1364
rect 4947 1356 5133 1364
rect 5616 1364 5624 1376
rect 6107 1376 6213 1384
rect 6927 1376 7133 1384
rect 7367 1376 7493 1384
rect 5176 1356 5624 1364
rect 2087 1336 2604 1344
rect 2616 1336 2693 1344
rect 1076 1316 1313 1324
rect 1427 1316 1684 1324
rect 596 1296 693 1304
rect 1087 1296 1173 1304
rect 1367 1296 1413 1304
rect 1527 1296 1633 1304
rect 1676 1304 1684 1316
rect 1707 1316 1853 1324
rect 1876 1316 1913 1324
rect 1876 1307 1884 1316
rect 1927 1316 1973 1324
rect 2076 1324 2084 1333
rect 2616 1327 2624 1336
rect 2707 1336 2813 1344
rect 2947 1336 2953 1344
rect 2967 1336 3233 1344
rect 3567 1336 3693 1344
rect 3807 1336 3853 1344
rect 4327 1336 4473 1344
rect 4667 1336 4693 1344
rect 4827 1336 5073 1344
rect 5127 1336 5153 1344
rect 5176 1327 5184 1356
rect 5647 1356 5733 1364
rect 6807 1356 6953 1364
rect 6967 1356 7333 1364
rect 7407 1356 7424 1364
rect 5267 1336 5313 1344
rect 5327 1336 5373 1344
rect 5547 1336 5673 1344
rect 6387 1336 6493 1344
rect 6507 1336 6513 1344
rect 6567 1336 6613 1344
rect 7067 1336 7093 1344
rect 7187 1336 7213 1344
rect 2076 1316 2124 1324
rect 2116 1307 2124 1316
rect 2487 1316 2553 1324
rect 2727 1316 2773 1324
rect 2796 1316 2873 1324
rect 1676 1296 1753 1304
rect 2007 1296 2093 1304
rect 2367 1296 2393 1304
rect 127 1276 133 1284
rect 147 1276 373 1284
rect 767 1276 793 1284
rect 867 1276 893 1284
rect 996 1284 1004 1293
rect 996 1276 1093 1284
rect 1127 1276 1273 1284
rect 1307 1276 1853 1284
rect 1967 1276 1973 1284
rect 1987 1276 2073 1284
rect 2227 1276 2313 1284
rect 2416 1284 2424 1313
rect 2507 1296 2573 1304
rect 2796 1304 2804 1316
rect 2927 1316 2944 1324
rect 2627 1296 2804 1304
rect 2887 1296 2913 1304
rect 2407 1276 2424 1284
rect 2487 1276 2533 1284
rect 2936 1284 2944 1316
rect 3067 1316 3173 1324
rect 3196 1316 3313 1324
rect 3196 1304 3204 1316
rect 3327 1316 3393 1324
rect 3687 1316 3813 1324
rect 3927 1316 3973 1324
rect 4087 1316 4193 1324
rect 4207 1316 4453 1324
rect 4507 1316 4613 1324
rect 4627 1316 4633 1324
rect 4727 1316 4853 1324
rect 4867 1316 4893 1324
rect 4967 1316 5113 1324
rect 5196 1324 5204 1333
rect 5196 1316 5233 1324
rect 5427 1316 5573 1324
rect 5627 1316 5793 1324
rect 6076 1316 6193 1324
rect 2987 1296 3204 1304
rect 3227 1296 3573 1304
rect 3787 1296 3833 1304
rect 3907 1296 4013 1304
rect 4267 1296 4313 1304
rect 4387 1296 4573 1304
rect 4967 1296 5393 1304
rect 5447 1296 5593 1304
rect 5687 1296 5693 1304
rect 5707 1296 5773 1304
rect 6076 1304 6084 1316
rect 6207 1316 6233 1324
rect 6356 1324 6364 1333
rect 6356 1316 6373 1324
rect 6387 1316 6533 1324
rect 7087 1316 7113 1324
rect 7207 1316 7233 1324
rect 7416 1307 7424 1356
rect 7527 1356 7593 1364
rect 7627 1356 7713 1364
rect 7567 1336 7593 1344
rect 7607 1336 7673 1344
rect 7687 1336 7753 1344
rect 7447 1316 7693 1324
rect 7827 1316 7873 1324
rect 5827 1296 6084 1304
rect 6107 1296 6213 1304
rect 6547 1296 6613 1304
rect 6867 1296 6893 1304
rect 6987 1296 7213 1304
rect 7587 1296 7613 1304
rect 2567 1276 2944 1284
rect 3227 1276 3293 1284
rect 3427 1276 3633 1284
rect 3667 1276 4033 1284
rect 4627 1276 4673 1284
rect 4847 1276 4873 1284
rect 5107 1276 5233 1284
rect 5507 1276 5933 1284
rect 6267 1276 6373 1284
rect 6707 1276 6933 1284
rect 6947 1276 7033 1284
rect 7127 1276 7193 1284
rect 7267 1276 7353 1284
rect 7367 1276 7393 1284
rect 7507 1276 7533 1284
rect 7847 1276 7873 1284
rect 407 1256 533 1264
rect 847 1256 1553 1264
rect 1567 1256 1653 1264
rect 1767 1256 1893 1264
rect 1967 1256 2033 1264
rect 2347 1256 3053 1264
rect 3307 1256 3333 1264
rect 3407 1256 3433 1264
rect 3467 1256 3533 1264
rect 3587 1256 3753 1264
rect 3807 1256 3933 1264
rect 4627 1256 4653 1264
rect 5787 1256 6293 1264
rect 6347 1256 6373 1264
rect 6387 1256 6413 1264
rect 6667 1256 7293 1264
rect 7307 1256 7473 1264
rect 107 1236 953 1244
rect 1167 1236 1233 1244
rect 1267 1236 1393 1244
rect 1456 1236 1513 1244
rect 387 1216 413 1224
rect 1456 1224 1464 1236
rect 1547 1236 1833 1244
rect 2007 1236 2153 1244
rect 2427 1236 2753 1244
rect 2807 1236 3693 1244
rect 3727 1236 3873 1244
rect 6067 1236 6693 1244
rect 7487 1236 7733 1244
rect 536 1216 1464 1224
rect 536 1204 544 1216
rect 1627 1216 2273 1224
rect 2487 1216 3273 1224
rect 3767 1216 3953 1224
rect 3967 1216 3993 1224
rect 6447 1216 6733 1224
rect 7527 1216 7613 1224
rect 327 1196 544 1204
rect 567 1196 653 1204
rect 927 1196 1073 1204
rect 1256 1196 1573 1204
rect 247 1176 753 1184
rect 1256 1184 1264 1196
rect 1747 1196 2073 1204
rect 2087 1196 2113 1204
rect 2167 1196 2353 1204
rect 2407 1196 2433 1204
rect 2447 1196 2613 1204
rect 2647 1196 2713 1204
rect 2807 1196 3073 1204
rect 3927 1196 3973 1204
rect 4767 1196 4793 1204
rect 5147 1196 5353 1204
rect 7467 1196 7793 1204
rect 7847 1196 7893 1204
rect 907 1176 1264 1184
rect 1547 1176 1693 1184
rect 1727 1176 1753 1184
rect 1856 1176 1973 1184
rect 427 1156 473 1164
rect 667 1156 733 1164
rect 1187 1156 1524 1164
rect 407 1136 613 1144
rect 647 1136 753 1144
rect 867 1136 913 1144
rect 1067 1136 1233 1144
rect 1427 1136 1453 1144
rect 1476 1136 1493 1144
rect 127 1116 253 1124
rect 287 1116 473 1124
rect 547 1116 593 1124
rect 627 1116 673 1124
rect 787 1116 813 1124
rect 887 1116 973 1124
rect 1087 1116 1113 1124
rect 147 1096 173 1104
rect 487 1096 504 1104
rect 267 1076 313 1084
rect 496 1084 504 1096
rect 527 1096 573 1104
rect 727 1096 793 1104
rect 1007 1096 1033 1104
rect 1107 1096 1133 1104
rect 1387 1096 1433 1104
rect 496 1076 613 1084
rect 667 1076 693 1084
rect 767 1076 833 1084
rect 1476 1084 1484 1136
rect 1516 1124 1524 1156
rect 1556 1156 1613 1164
rect 1556 1144 1564 1156
rect 1856 1164 1864 1176
rect 2287 1176 2373 1184
rect 2387 1176 2424 1184
rect 1687 1156 1864 1164
rect 1967 1156 2053 1164
rect 2107 1156 2133 1164
rect 2147 1156 2213 1164
rect 2416 1164 2424 1176
rect 2447 1176 2613 1184
rect 2687 1176 2793 1184
rect 2827 1176 2873 1184
rect 2927 1176 3173 1184
rect 3347 1176 3373 1184
rect 3387 1176 3433 1184
rect 3447 1176 3473 1184
rect 3487 1176 3513 1184
rect 6087 1176 6133 1184
rect 6147 1176 6293 1184
rect 6367 1176 6393 1184
rect 7447 1176 7673 1184
rect 7867 1176 7893 1184
rect 2416 1156 2653 1164
rect 2667 1156 2693 1164
rect 2847 1156 2973 1164
rect 3067 1156 3253 1164
rect 3527 1156 3613 1164
rect 5907 1156 6213 1164
rect 6227 1156 6453 1164
rect 7627 1156 7644 1164
rect 1507 1116 1524 1124
rect 1536 1136 1564 1144
rect 1536 1104 1544 1136
rect 1607 1136 1693 1144
rect 1716 1136 1773 1144
rect 1716 1124 1724 1136
rect 1796 1136 1913 1144
rect 1587 1116 1724 1124
rect 1796 1124 1804 1136
rect 2147 1136 2344 1144
rect 2336 1127 2344 1136
rect 2447 1136 2453 1144
rect 2467 1136 2813 1144
rect 2836 1136 2853 1144
rect 1747 1116 1804 1124
rect 1847 1116 1933 1124
rect 1947 1116 2153 1124
rect 2267 1116 2324 1124
rect 1527 1096 1544 1104
rect 2316 1104 2324 1116
rect 2287 1096 2304 1104
rect 2316 1096 2353 1104
rect 1476 1076 1493 1084
rect 1736 1084 1744 1093
rect 1627 1076 1744 1084
rect 1867 1076 2033 1084
rect 2296 1084 2304 1096
rect 2296 1076 2373 1084
rect 207 1056 1133 1064
rect 1527 1056 1553 1064
rect 1647 1056 1753 1064
rect 2396 1064 2404 1133
rect 2687 1116 2713 1124
rect 2416 1104 2424 1113
rect 2836 1107 2844 1136
rect 2887 1136 3093 1144
rect 3116 1136 3133 1144
rect 2867 1116 2964 1124
rect 2416 1096 2773 1104
rect 2956 1104 2964 1116
rect 3116 1124 3124 1136
rect 3167 1136 3353 1144
rect 3647 1136 3673 1144
rect 3736 1136 3873 1144
rect 2987 1116 3124 1124
rect 3667 1116 3684 1124
rect 2956 1096 2993 1104
rect 3156 1104 3164 1113
rect 3676 1107 3684 1116
rect 3156 1096 3173 1104
rect 3207 1096 3253 1104
rect 3267 1096 3493 1104
rect 3567 1096 3613 1104
rect 2427 1076 2453 1084
rect 2507 1076 2513 1084
rect 2527 1076 2573 1084
rect 2876 1084 2884 1093
rect 2667 1076 3033 1084
rect 3536 1084 3544 1093
rect 3107 1076 3544 1084
rect 3656 1067 3664 1093
rect 3736 1084 3744 1136
rect 4007 1136 4033 1144
rect 4047 1136 4233 1144
rect 4387 1136 4553 1144
rect 5627 1136 5733 1144
rect 5836 1136 6093 1144
rect 3807 1116 3833 1124
rect 3896 1124 3904 1133
rect 3856 1116 3904 1124
rect 3856 1107 3864 1116
rect 4107 1116 4173 1124
rect 4347 1116 4673 1124
rect 4687 1116 4713 1124
rect 4727 1116 4953 1124
rect 5007 1116 5053 1124
rect 5247 1116 5573 1124
rect 5836 1124 5844 1136
rect 6127 1136 6373 1144
rect 7007 1136 7053 1144
rect 7267 1136 7493 1144
rect 7547 1136 7613 1144
rect 7636 1144 7644 1156
rect 7667 1156 7853 1164
rect 7636 1136 7653 1144
rect 7707 1136 7713 1144
rect 7727 1136 7773 1144
rect 5667 1116 5844 1124
rect 5867 1116 5984 1124
rect 3767 1096 3844 1104
rect 3836 1084 3844 1096
rect 4227 1096 4393 1104
rect 4407 1096 4873 1104
rect 4887 1096 4973 1104
rect 5467 1096 5633 1104
rect 5707 1096 5833 1104
rect 5976 1087 5984 1116
rect 6307 1116 6333 1124
rect 6847 1116 6953 1124
rect 7047 1116 7313 1124
rect 7487 1116 7524 1124
rect 6007 1096 6033 1104
rect 6167 1096 6233 1104
rect 3736 1076 3784 1084
rect 3836 1076 3853 1084
rect 3776 1067 3784 1076
rect 4027 1076 4193 1084
rect 4207 1076 4513 1084
rect 4587 1076 5113 1084
rect 5367 1076 5473 1084
rect 5807 1076 5953 1084
rect 6256 1084 6264 1113
rect 7516 1107 7524 1116
rect 7596 1116 7653 1124
rect 6287 1096 6313 1104
rect 6587 1096 6913 1104
rect 6927 1096 7013 1104
rect 7387 1096 7473 1104
rect 7596 1087 7604 1116
rect 7767 1116 7804 1124
rect 7627 1096 7773 1104
rect 6256 1076 6413 1084
rect 6847 1076 6933 1084
rect 6947 1076 7033 1084
rect 7087 1076 7133 1084
rect 7147 1076 7353 1084
rect 7467 1076 7573 1084
rect 7796 1084 7804 1116
rect 7876 1104 7884 1133
rect 7867 1096 7884 1104
rect 7796 1076 7873 1084
rect 1996 1056 2513 1064
rect 247 1036 313 1044
rect 567 1036 653 1044
rect 1447 1036 1693 1044
rect 1996 1044 2004 1056
rect 2547 1056 2593 1064
rect 2687 1056 2793 1064
rect 3667 1056 3733 1064
rect 5607 1056 5713 1064
rect 6007 1056 6033 1064
rect 6207 1056 6793 1064
rect 6807 1056 6973 1064
rect 6987 1056 7113 1064
rect 1947 1036 2004 1044
rect 2347 1036 2453 1044
rect 2467 1036 2553 1044
rect 2707 1036 2933 1044
rect 3287 1036 3453 1044
rect 3527 1036 3573 1044
rect 3727 1036 3753 1044
rect 3987 1036 4073 1044
rect 4087 1036 4193 1044
rect 4207 1036 4313 1044
rect 5127 1036 5433 1044
rect 5487 1036 5753 1044
rect 5767 1036 5853 1044
rect 5887 1036 6153 1044
rect 6267 1036 6293 1044
rect 6567 1036 6633 1044
rect 6687 1036 6893 1044
rect 347 1016 2193 1024
rect 2327 1016 2633 1024
rect 2747 1016 3173 1024
rect 1227 996 2493 1004
rect 2567 996 3313 1004
rect 3507 996 3593 1004
rect 4567 996 6593 1004
rect 6607 996 6713 1004
rect 987 976 1733 984
rect 1767 976 2233 984
rect 2247 976 2833 984
rect 5487 976 5553 984
rect 5567 976 5593 984
rect 487 956 1873 964
rect 2007 956 2413 964
rect 2507 956 2813 964
rect 5667 956 5973 964
rect 5987 956 6493 964
rect 447 936 533 944
rect 547 936 1213 944
rect 1227 936 1413 944
rect 1487 936 1573 944
rect 1587 936 1773 944
rect 1847 936 1953 944
rect 2407 936 2713 944
rect 2887 936 2913 944
rect 3067 936 4293 944
rect 5447 936 5793 944
rect 7787 936 7853 944
rect 747 916 993 924
rect 1007 916 1993 924
rect 2067 916 2473 924
rect 2527 916 2713 924
rect 3547 916 3693 924
rect 3987 916 4133 924
rect 807 896 1393 904
rect 1427 896 1533 904
rect 1587 896 1753 904
rect 1787 896 2373 904
rect 2587 896 2733 904
rect 3307 896 3633 904
rect 6007 896 6033 904
rect 7447 896 7473 904
rect 267 876 373 884
rect 787 876 853 884
rect 1287 876 1313 884
rect 1407 876 1473 884
rect 1487 876 1973 884
rect 2087 876 2133 884
rect 2527 876 3013 884
rect 3027 876 3413 884
rect 3576 876 3793 884
rect 276 856 293 864
rect 276 847 284 856
rect 387 856 513 864
rect 587 856 713 864
rect 727 856 773 864
rect 787 856 893 864
rect 947 856 1933 864
rect 1967 856 2013 864
rect 2087 856 2553 864
rect 2607 856 2893 864
rect 2947 856 2973 864
rect 3147 856 3353 864
rect 3376 856 3553 864
rect 327 836 404 844
rect 147 816 173 824
rect 247 816 273 824
rect 287 816 373 824
rect 396 824 404 836
rect 587 836 613 844
rect 627 836 753 844
rect 767 836 953 844
rect 1156 836 1313 844
rect 1156 827 1164 836
rect 1347 836 1373 844
rect 1467 836 1613 844
rect 1656 836 1693 844
rect 396 816 493 824
rect 1287 816 1353 824
rect 1656 824 1664 836
rect 1747 836 2093 844
rect 2707 836 2833 844
rect 3007 836 3093 844
rect 3247 836 3293 844
rect 3376 844 3384 856
rect 3576 847 3584 876
rect 3807 876 3824 884
rect 3816 867 3824 876
rect 4107 876 4393 884
rect 5616 876 5633 884
rect 3607 856 3633 864
rect 3656 856 3773 864
rect 3327 836 3384 844
rect 3656 844 3664 856
rect 4356 856 4424 864
rect 3627 836 3664 844
rect 3707 836 3793 844
rect 4147 836 4293 844
rect 4356 827 4364 856
rect 4416 844 4424 856
rect 4467 856 4813 864
rect 4827 856 4873 864
rect 5287 856 5313 864
rect 5527 856 5593 864
rect 5616 847 5624 876
rect 5947 876 6153 884
rect 6167 876 6513 884
rect 7447 876 7513 884
rect 7567 876 7633 884
rect 5707 856 5753 864
rect 5767 856 5893 864
rect 6447 856 6533 864
rect 6987 856 7173 864
rect 7387 856 7413 864
rect 7587 856 7733 864
rect 7807 856 7833 864
rect 4416 836 4593 844
rect 5027 836 5213 844
rect 1607 816 1664 824
rect 1787 816 2133 824
rect 2407 816 2433 824
rect 2567 816 2593 824
rect 2667 816 2693 824
rect 2727 816 2773 824
rect 3127 816 3413 824
rect 3547 816 3673 824
rect 3747 816 3853 824
rect 4227 816 4313 824
rect 4396 824 4404 833
rect 5176 827 5184 836
rect 5347 836 5513 844
rect 5636 844 5644 853
rect 5636 836 5673 844
rect 5947 836 5993 844
rect 6427 836 6473 844
rect 7336 844 7344 853
rect 7047 836 7344 844
rect 7456 827 7464 853
rect 7487 836 7613 844
rect 4396 816 4473 824
rect 5187 816 5533 824
rect 5547 816 5633 824
rect 5647 816 5833 824
rect 5887 816 6013 824
rect 6067 816 6093 824
rect 6107 816 6373 824
rect 6467 816 6493 824
rect 6547 816 6853 824
rect 6867 816 6873 824
rect 6927 816 6993 824
rect 7007 816 7013 824
rect 7227 816 7353 824
rect 7507 816 7533 824
rect 107 796 293 804
rect 347 796 393 804
rect 547 796 593 804
rect 607 796 1373 804
rect 1676 804 1684 813
rect 1587 796 1684 804
rect 1727 796 1793 804
rect 1927 796 2013 804
rect 2027 796 2053 804
rect 2167 796 2193 804
rect 2207 796 2733 804
rect 2827 796 3353 804
rect 3387 796 3533 804
rect 3967 796 4033 804
rect 4047 796 4333 804
rect 4387 796 4413 804
rect 5147 796 5453 804
rect 5507 796 5673 804
rect 6067 796 6173 804
rect 6207 796 6313 804
rect 6327 796 6753 804
rect 7656 804 7664 833
rect 7687 816 7753 824
rect 7807 816 7873 824
rect 7656 796 7713 804
rect 7767 796 7793 804
rect 367 776 533 784
rect 547 776 693 784
rect 967 776 1693 784
rect 1727 776 1933 784
rect 2156 776 2673 784
rect 147 756 913 764
rect 927 756 1053 764
rect 1207 756 1253 764
rect 1267 756 1353 764
rect 2156 764 2164 776
rect 3467 776 3713 784
rect 4007 776 4113 784
rect 4127 776 4513 784
rect 4527 776 4553 784
rect 4607 776 6673 784
rect 7727 776 7853 784
rect 1387 756 2164 764
rect 3347 756 3393 764
rect 3407 756 3853 764
rect 6187 756 6273 764
rect 7507 756 7633 764
rect 427 736 453 744
rect 467 736 933 744
rect 1076 736 1513 744
rect 1076 724 1084 736
rect 1567 736 1733 744
rect 1787 736 1913 744
rect 1947 736 2613 744
rect 2747 736 4433 744
rect 7587 736 7653 744
rect 767 716 1084 724
rect 1247 716 1333 724
rect 1347 716 1873 724
rect 1887 716 2033 724
rect 2727 716 3253 724
rect 5007 716 5393 724
rect 6247 716 6313 724
rect 6327 716 6493 724
rect 7167 716 7473 724
rect 7587 716 7733 724
rect 7787 716 7884 724
rect 387 696 433 704
rect 467 696 613 704
rect 1167 696 1313 704
rect 1367 696 1713 704
rect 1867 696 1893 704
rect 2227 696 2433 704
rect 2807 696 3113 704
rect 4727 696 4833 704
rect 4847 696 5353 704
rect 6307 696 6453 704
rect 6887 696 7833 704
rect 7847 696 7853 704
rect 167 676 293 684
rect 307 676 473 684
rect 647 676 733 684
rect 847 676 1033 684
rect 1067 676 1193 684
rect 1207 676 1233 684
rect 1307 676 1413 684
rect 1507 676 1913 684
rect 1927 676 2273 684
rect 2287 676 2353 684
rect 2367 676 2473 684
rect 2487 676 2953 684
rect 2967 676 3153 684
rect 3167 676 3173 684
rect 3187 676 3493 684
rect 3587 676 3633 684
rect 4527 676 4973 684
rect 4987 676 5173 684
rect 5847 676 6693 684
rect 6707 676 6813 684
rect 6827 676 6993 684
rect 7007 676 7173 684
rect 7187 676 7193 684
rect 7227 676 7673 684
rect 7787 676 7813 684
rect 7876 684 7884 716
rect 7847 676 7884 684
rect 107 656 413 664
rect 436 656 493 664
rect 47 636 133 644
rect 436 627 444 656
rect 527 656 673 664
rect 727 656 853 664
rect 1076 656 1113 664
rect 587 636 753 644
rect 776 636 793 644
rect 347 616 393 624
rect 567 616 633 624
rect 776 624 784 636
rect 887 636 933 644
rect 736 616 784 624
rect 327 596 613 604
rect 656 604 664 613
rect 736 607 744 616
rect 1027 616 1053 624
rect 1076 624 1084 656
rect 1287 656 1433 664
rect 1527 656 1553 664
rect 1747 656 1953 664
rect 2067 656 2093 664
rect 2187 656 2293 664
rect 2347 656 2524 664
rect 1107 636 1233 644
rect 1307 636 1324 644
rect 1316 627 1324 636
rect 1427 636 1453 644
rect 1496 636 1513 644
rect 1076 616 1113 624
rect 1347 616 1393 624
rect 627 596 664 604
rect 967 596 1073 604
rect 1307 596 1353 604
rect 1496 587 1504 636
rect 1607 636 1793 644
rect 1887 636 1933 644
rect 2107 636 2173 644
rect 2516 644 2524 656
rect 2907 656 3133 664
rect 3147 656 3264 664
rect 3256 647 3264 656
rect 3307 656 3333 664
rect 3447 656 3473 664
rect 3507 656 3653 664
rect 4136 656 4293 664
rect 2516 636 2553 644
rect 2647 636 2753 644
rect 3027 636 3153 644
rect 3167 636 3193 644
rect 3587 636 3613 644
rect 3707 636 4033 644
rect 1667 616 1693 624
rect 1767 616 1853 624
rect 2127 616 2233 624
rect 2256 624 2264 633
rect 4056 627 4064 653
rect 2256 616 2313 624
rect 2427 616 2653 624
rect 2667 616 2713 624
rect 2747 616 2773 624
rect 3047 616 3293 624
rect 3347 616 3393 624
rect 3487 616 3733 624
rect 3907 616 4013 624
rect 4136 624 4144 656
rect 4347 656 4433 664
rect 4467 656 4533 664
rect 4787 656 4993 664
rect 5147 656 5233 664
rect 5767 656 6133 664
rect 6387 656 6413 664
rect 6447 656 6473 664
rect 6487 656 6533 664
rect 6767 656 6933 664
rect 7027 656 7333 664
rect 7347 656 7393 664
rect 7407 656 7413 664
rect 7467 656 7593 664
rect 7607 656 7633 664
rect 7656 656 7693 664
rect 4167 636 4233 644
rect 4827 636 4933 644
rect 4956 636 5033 644
rect 4136 616 4184 624
rect 4176 607 4184 616
rect 4247 616 4293 624
rect 4556 624 4564 633
rect 4347 616 4613 624
rect 4956 624 4964 636
rect 5267 636 5433 644
rect 5376 627 5384 636
rect 5587 636 5713 644
rect 6287 636 6333 644
rect 6627 636 7073 644
rect 7247 636 7373 644
rect 7536 636 7593 644
rect 4636 616 4964 624
rect 1687 596 1713 604
rect 1767 596 1813 604
rect 2107 596 2493 604
rect 3127 596 3493 604
rect 3507 596 3633 604
rect 3687 596 3713 604
rect 3807 596 3833 604
rect 287 576 333 584
rect 607 576 773 584
rect 787 576 1484 584
rect 227 556 353 564
rect 367 556 693 564
rect 707 556 873 564
rect 1476 564 1484 576
rect 1527 576 1533 584
rect 1547 576 1644 584
rect 1476 556 1613 564
rect 1636 564 1644 576
rect 1727 576 1793 584
rect 2207 576 2293 584
rect 2607 576 2813 584
rect 2827 576 3053 584
rect 3767 576 3873 584
rect 3927 576 4093 584
rect 4196 584 4204 613
rect 4636 604 4644 616
rect 5067 616 5113 624
rect 5127 616 5193 624
rect 5567 616 5733 624
rect 5787 616 5813 624
rect 5827 616 6013 624
rect 6076 616 6133 624
rect 6076 607 6084 616
rect 6327 616 6353 624
rect 6407 616 6433 624
rect 6667 616 6773 624
rect 6896 616 6933 624
rect 6896 607 6904 616
rect 7067 616 7353 624
rect 7407 616 7513 624
rect 7536 607 7544 636
rect 7656 644 7664 656
rect 7767 656 7873 664
rect 7616 636 7664 644
rect 7616 627 7624 636
rect 7696 636 7733 644
rect 4527 596 4644 604
rect 5087 596 5413 604
rect 5427 596 5453 604
rect 5467 596 5793 604
rect 6347 596 6573 604
rect 6587 596 6633 604
rect 6787 596 6853 604
rect 6967 596 7073 604
rect 7087 596 7113 604
rect 7547 596 7653 604
rect 7676 587 7684 633
rect 7696 604 7704 636
rect 7756 636 7773 644
rect 7756 624 7764 636
rect 7727 616 7764 624
rect 7816 624 7824 633
rect 7816 616 7873 624
rect 7696 596 7873 604
rect 4127 576 4204 584
rect 4827 576 4893 584
rect 5347 576 5953 584
rect 5967 576 6093 584
rect 6107 576 6133 584
rect 6707 576 6833 584
rect 6847 576 6913 584
rect 1636 556 2073 564
rect 2087 556 2413 564
rect 2867 556 2933 564
rect 3627 556 3773 564
rect 4107 556 4373 564
rect 4387 556 4953 564
rect 6047 556 6193 564
rect 307 536 453 544
rect 547 536 1433 544
rect 1587 536 1933 544
rect 1967 536 2073 544
rect 2247 536 2593 544
rect 2807 536 3273 544
rect 4787 536 4893 544
rect 5267 536 5973 544
rect 5987 536 6113 544
rect 427 516 1693 524
rect 1747 516 1813 524
rect 4787 516 4873 524
rect 4887 516 5293 524
rect 1467 496 3973 504
rect 4367 496 4693 504
rect 5187 496 6593 504
rect 6607 496 6673 504
rect 7807 496 7893 504
rect 367 476 753 484
rect 1047 476 3513 484
rect 3887 476 4573 484
rect 4847 476 5853 484
rect 567 456 673 464
rect 687 456 853 464
rect 1227 456 1813 464
rect 3427 456 3793 464
rect 4487 456 4993 464
rect 7527 456 7553 464
rect 627 436 873 444
rect 887 436 993 444
rect 1267 436 1673 444
rect 2827 436 2913 444
rect 3547 436 3693 444
rect 3847 436 4113 444
rect 4147 436 4213 444
rect 4227 436 4413 444
rect 4647 436 5073 444
rect 6567 436 6593 444
rect 687 416 813 424
rect 1347 416 1613 424
rect 2027 416 2353 424
rect 2367 416 2573 424
rect 2767 416 2973 424
rect 3807 416 4773 424
rect 4947 416 5133 424
rect 5327 416 6373 424
rect 6387 416 6773 424
rect 7347 416 7393 424
rect 127 396 213 404
rect 1507 396 1533 404
rect 1587 396 1893 404
rect 2227 396 2573 404
rect 2927 396 3033 404
rect 3307 396 3593 404
rect 3947 396 3973 404
rect 4067 396 4113 404
rect 4127 396 4493 404
rect 4516 396 4793 404
rect 107 376 233 384
rect 927 376 1233 384
rect 1327 376 1353 384
rect 1487 376 1653 384
rect 1667 376 2233 384
rect 2267 376 2473 384
rect 2907 376 2933 384
rect 2987 376 3033 384
rect 3056 376 3073 384
rect 76 364 84 373
rect 76 356 144 364
rect 136 347 144 356
rect 327 356 373 364
rect 667 356 733 364
rect 787 356 893 364
rect 1027 356 1153 364
rect 1467 356 1553 364
rect 1567 356 1653 364
rect 1707 356 1853 364
rect 1907 356 1953 364
rect 2247 356 2373 364
rect 2507 356 2613 364
rect 2927 356 2953 364
rect 3056 364 3064 376
rect 3327 376 3373 384
rect 3967 376 3993 384
rect 4327 376 4433 384
rect 4516 384 4524 396
rect 5147 396 5553 404
rect 6467 396 6493 404
rect 6567 396 6733 404
rect 7127 396 7153 404
rect 7387 396 7453 404
rect 4447 376 4524 384
rect 4536 376 4553 384
rect 3007 356 3064 364
rect 3107 356 3153 364
rect 3767 356 3933 364
rect 4267 356 4293 364
rect 4407 356 4433 364
rect 4536 364 4544 376
rect 4707 376 4713 384
rect 4727 376 4733 384
rect 5087 376 5173 384
rect 5227 376 5373 384
rect 5387 376 5613 384
rect 5767 376 5813 384
rect 5867 376 6333 384
rect 6487 376 6613 384
rect 6667 376 6733 384
rect 6807 376 6913 384
rect 6927 376 6973 384
rect 6996 376 7053 384
rect 4467 356 4544 364
rect 4656 364 4664 373
rect 4587 356 4664 364
rect 5036 364 5044 373
rect 4867 356 5093 364
rect 5367 356 5433 364
rect 5487 356 5513 364
rect 5536 356 5653 364
rect 87 336 104 344
rect 96 327 104 336
rect 147 336 613 344
rect 647 336 713 344
rect 867 336 1073 344
rect 1196 344 1204 353
rect 5536 347 5544 356
rect 5807 356 5853 364
rect 6107 356 6184 364
rect 6176 347 6184 356
rect 6216 356 6273 364
rect 6216 347 6224 356
rect 6416 364 6424 373
rect 6367 356 6513 364
rect 1167 336 1204 344
rect 1227 336 1253 344
rect 1287 336 1373 344
rect 1447 336 1513 344
rect 1707 336 1793 344
rect 1807 336 2013 344
rect 2067 336 2133 344
rect 2167 336 2293 344
rect 2607 336 2793 344
rect 2867 336 2993 344
rect 3007 336 3233 344
rect 3156 327 3164 336
rect 3747 336 3833 344
rect 4427 336 4513 344
rect 4607 336 4713 344
rect 5807 336 5953 344
rect 6327 336 6633 344
rect 6827 336 6973 344
rect 6996 344 7004 376
rect 7107 376 7233 384
rect 7347 376 7413 384
rect 7427 376 7433 384
rect 7027 356 7284 364
rect 6987 336 7004 344
rect 127 316 153 324
rect 307 316 533 324
rect 627 316 1313 324
rect 1487 316 1593 324
rect 1727 316 1833 324
rect 1847 316 2433 324
rect 3267 316 3313 324
rect 3707 316 3873 324
rect 3887 316 4033 324
rect 4087 316 4193 324
rect 4207 316 4233 324
rect 4767 316 4893 324
rect 5127 316 5173 324
rect 5187 316 5233 324
rect 5527 316 5553 324
rect 5987 316 6013 324
rect 6447 316 6473 324
rect 6507 316 6533 324
rect 6547 316 6673 324
rect 6887 316 6933 324
rect 7016 324 7024 353
rect 7187 336 7253 344
rect 7276 344 7284 356
rect 7307 356 7353 364
rect 7847 356 7893 364
rect 7276 336 7473 344
rect 7727 336 7753 344
rect 7827 336 7853 344
rect 6967 316 7024 324
rect 7047 316 7213 324
rect 7327 316 7633 324
rect 7667 316 7773 324
rect 367 296 393 304
rect 607 296 653 304
rect 707 296 813 304
rect 827 296 973 304
rect 1107 296 1153 304
rect 1307 296 1333 304
rect 1387 296 2153 304
rect 3607 296 3773 304
rect 4107 296 4633 304
rect 4656 296 4813 304
rect 1067 276 1773 284
rect 1787 276 2113 284
rect 2127 276 2253 284
rect 3067 276 3233 284
rect 3907 276 3933 284
rect 3947 276 4053 284
rect 4067 276 4313 284
rect 4656 284 4664 296
rect 4827 296 4913 304
rect 5687 296 5813 304
rect 5827 296 6233 304
rect 6247 296 6673 304
rect 7607 296 7913 304
rect 4387 276 4664 284
rect 5167 276 5513 284
rect 6007 276 6353 284
rect 6367 276 6473 284
rect 6487 276 6593 284
rect 6627 276 6753 284
rect 6767 276 6853 284
rect 487 256 1413 264
rect 1807 256 1933 264
rect 2007 256 2073 264
rect 2147 256 2193 264
rect 3827 256 4333 264
rect 4347 256 4533 264
rect 4547 256 4693 264
rect 4727 256 4813 264
rect 4967 256 5173 264
rect 5507 256 5733 264
rect 6567 256 6833 264
rect 327 236 533 244
rect 547 236 853 244
rect 1127 236 1693 244
rect 4127 236 4553 244
rect 4587 236 5253 244
rect 5587 236 5833 244
rect 5847 236 6573 244
rect 427 216 673 224
rect 1187 216 1613 224
rect 1647 216 1913 224
rect 1987 216 2293 224
rect 4287 216 4953 224
rect 4967 216 5013 224
rect 5067 216 6073 224
rect 6087 216 6613 224
rect 6687 216 7153 224
rect 7487 216 7833 224
rect 227 196 313 204
rect 447 196 473 204
rect 1167 196 1453 204
rect 1607 196 1813 204
rect 1827 196 1993 204
rect 2607 196 2813 204
rect 2907 196 2933 204
rect 3207 196 3293 204
rect 3307 196 3533 204
rect 4187 196 4293 204
rect 4307 196 4313 204
rect 4327 196 5133 204
rect 5487 196 5633 204
rect 5647 196 5713 204
rect 5727 196 5973 204
rect 6207 196 6393 204
rect 6407 196 6553 204
rect 6607 196 7033 204
rect 7407 196 7453 204
rect 7467 196 7593 204
rect 147 176 713 184
rect 727 176 953 184
rect 967 176 1193 184
rect 1327 176 1353 184
rect 1667 176 1953 184
rect 1967 176 2273 184
rect 2287 176 2733 184
rect 2747 176 2773 184
rect 2787 176 3053 184
rect 3247 176 3373 184
rect 3687 176 3713 184
rect 3927 176 3973 184
rect 4167 176 4333 184
rect 4347 176 4433 184
rect 4447 176 4453 184
rect 4687 176 4853 184
rect 4987 176 5113 184
rect 5287 176 5313 184
rect 6087 176 6093 184
rect 6107 176 6153 184
rect 6201 176 6293 184
rect 6607 176 6633 184
rect 6647 176 6693 184
rect 6747 176 7133 184
rect 7147 176 7393 184
rect 47 156 133 164
rect 187 156 333 164
rect 467 156 493 164
rect 587 156 693 164
rect 767 156 913 164
rect 1047 156 1233 164
rect 1287 156 1353 164
rect 1507 156 1533 164
rect 1747 156 1773 164
rect 2007 156 2033 164
rect 2167 156 2193 164
rect 2407 156 2453 164
rect 2507 156 2693 164
rect 2867 156 3253 164
rect 3447 156 3493 164
rect 3867 156 3953 164
rect 4007 156 4093 164
rect 4107 156 4144 164
rect 4136 147 4144 156
rect 4427 156 4493 164
rect 4516 156 4773 164
rect 227 136 353 144
rect 367 136 1133 144
rect 1347 136 1393 144
rect 1447 136 1553 144
rect 1687 136 1793 144
rect 2067 136 2113 144
rect 2347 136 2473 144
rect 2907 136 2993 144
rect 3287 136 3413 144
rect 3747 136 3973 144
rect 4107 136 4124 144
rect 87 116 293 124
rect 347 116 553 124
rect 567 116 1753 124
rect 1767 116 2133 124
rect 2387 116 2513 124
rect 3147 116 3393 124
rect 3407 116 3473 124
rect 3567 116 3613 124
rect 3687 116 4033 124
rect 4116 124 4124 136
rect 4156 124 4164 153
rect 4516 147 4524 156
rect 5147 156 5264 164
rect 4536 136 4593 144
rect 4116 116 4164 124
rect 4536 124 4544 136
rect 4707 136 4793 144
rect 4847 136 4913 144
rect 5187 136 5233 144
rect 5256 144 5264 156
rect 5467 156 5753 164
rect 5947 156 6213 164
rect 6236 156 6313 164
rect 6236 147 6244 156
rect 6496 164 6504 173
rect 6407 156 6733 164
rect 6787 156 6913 164
rect 7007 156 7233 164
rect 7287 156 7493 164
rect 7516 156 7613 164
rect 7516 147 7524 156
rect 5256 136 5333 144
rect 6127 136 6193 144
rect 6307 136 6333 144
rect 6687 136 6713 144
rect 6767 136 6853 144
rect 7427 136 7473 144
rect 7607 136 7633 144
rect 4487 116 4544 124
rect 4767 116 4893 124
rect 4907 116 5073 124
rect 5087 116 5393 124
rect 6287 116 6433 124
rect 7656 124 7664 173
rect 7676 147 7684 173
rect 7747 136 7853 144
rect 7656 116 7733 124
rect 387 96 513 104
rect 867 96 2053 104
rect 4076 104 4084 113
rect 4076 96 4273 104
rect 7567 96 7753 104
use NAND2X1  _1434_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304996
transform -1 0 4630 0 1 730
box -12 -8 92 252
use NAND2X1  _1435_
timestamp 1728304996
transform -1 0 4250 0 1 730
box -12 -8 92 252
use NOR2X1  _1436_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305106
transform -1 0 4370 0 1 730
box -12 -8 92 252
use INVX1  _1437_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304789
transform 1 0 5270 0 -1 730
box -12 -8 72 252
use INVX1  _1438_
timestamp 1728304789
transform 1 0 4110 0 1 730
box -12 -8 72 252
use INVX1  _1439_
timestamp 1728304789
transform 1 0 4590 0 -1 730
box -12 -8 72 252
use AND2X2  _1440_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304163
transform -1 0 4610 0 -1 1210
box -12 -8 112 252
use AND2X2  _1441_
timestamp 1728304163
transform 1 0 4030 0 -1 1210
box -12 -8 112 252
use NAND3X1  _1442_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305047
transform -1 0 4230 0 -1 1210
box -12 -8 112 252
use AOI21X1  _1443_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304211
transform 1 0 4290 0 -1 730
box -12 -8 112 252
use INVX1  _1444_
timestamp 1728304789
transform 1 0 5310 0 -1 250
box -12 -8 72 252
use NOR2X1  _1445_
timestamp 1728305106
transform 1 0 5090 0 -1 250
box -12 -8 92 252
use INVX1  _1446_
timestamp 1728304789
transform 1 0 5090 0 -1 730
box -12 -8 72 252
use NOR2X1  _1447_
timestamp 1728305106
transform -1 0 5270 0 -1 730
box -12 -8 92 252
use AND2X2  _1448_
timestamp 1728304163
transform -1 0 4990 0 1 250
box -12 -8 112 252
use OAI21X1  _1449_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305162
transform -1 0 4990 0 -1 730
box -12 -8 112 252
use AOI21X1  _1450_
timestamp 1728304211
transform -1 0 5430 0 -1 730
box -12 -8 112 252
use NAND3X1  _1451_
timestamp 1728305047
transform -1 0 4870 0 -1 730
box -12 -8 112 252
use AOI21X1  _1452_
timestamp 1728304211
transform -1 0 4030 0 -1 1210
box -12 -8 112 252
use OAI21X1  _1453_
timestamp 1728305162
transform -1 0 3970 0 1 730
box -12 -8 112 252
use INVX1  _1454_
timestamp 1728304789
transform -1 0 4150 0 -1 730
box -12 -8 72 252
use NOR2X1  _1455_
timestamp 1728305106
transform -1 0 4090 0 1 730
box -12 -8 92 252
use OAI21X1  _1456_
timestamp 1728305162
transform -1 0 4090 0 -1 730
box -12 -8 112 252
use NAND2X1  _1457_
timestamp 1728304996
transform 1 0 4170 0 -1 730
box -12 -8 92 252
use INVX1  _1458_
timestamp 1728304789
transform 1 0 4370 0 1 730
box -12 -8 72 252
use NOR2X1  _1459_
timestamp 1728305106
transform -1 0 4530 0 1 730
box -12 -8 92 252
use NOR2X1  _1460_
timestamp 1728305106
transform 1 0 4510 0 -1 730
box -12 -8 92 252
use NAND3X1  _1461_
timestamp 1728305047
transform -1 0 4490 0 -1 730
box -12 -8 112 252
use AOI21X1  _1462_
timestamp 1728304211
transform 1 0 4010 0 1 250
box -12 -8 112 252
use NAND2X1  _1463_
timestamp 1728304996
transform -1 0 4190 0 1 250
box -12 -8 92 252
use INVX1  _1464_
timestamp 1728304789
transform -1 0 4730 0 -1 730
box -12 -8 72 252
use AOI21X1  _1465_
timestamp 1728304211
transform -1 0 4410 0 1 250
box -12 -8 112 252
use NAND2X1  _1466_
timestamp 1728304996
transform -1 0 3970 0 1 250
box -12 -8 92 252
use AOI22X1  _1467_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304278
transform 1 0 3730 0 1 250
box -14 -8 132 252
use OR2X2  _1468_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305284
transform -1 0 3730 0 1 250
box -12 -8 112 252
use INVX1  _1469_
timestamp 1728304789
transform 1 0 3710 0 -1 250
box -12 -8 72 252
use OAI21X1  _1470_
timestamp 1728305162
transform -1 0 4010 0 -1 250
box -12 -8 112 252
use NAND2X1  _1471_
timestamp 1728304996
transform 1 0 4570 0 -1 250
box -12 -8 92 252
use AOI22X1  _1472_
timestamp 1728304278
transform 1 0 4450 0 -1 250
box -14 -8 132 252
use OAI21X1  _1473_
timestamp 1728305162
transform 1 0 4110 0 -1 250
box -12 -8 112 252
use OR2X2  _1474_
timestamp 1728305284
transform -1 0 4350 0 -1 250
box -12 -8 112 252
use NAND3X1  _1475_
timestamp 1728305047
transform -1 0 4110 0 -1 250
box -12 -8 112 252
use INVX1  _1476_
timestamp 1728304789
transform -1 0 4770 0 1 250
box -12 -8 72 252
use OAI21X1  _1477_
timestamp 1728305162
transform 1 0 5210 0 -1 250
box -12 -8 112 252
use NAND2X1  _1478_
timestamp 1728304996
transform -1 0 4710 0 1 250
box -12 -8 92 252
use AOI21X1  _1479_
timestamp 1728304211
transform 1 0 4210 0 1 250
box -12 -8 112 252
use NAND2X1  _1480_
timestamp 1728304996
transform 1 0 4890 0 -1 250
box -12 -8 92 252
use AOI22X1  _1481_
timestamp 1728304278
transform 1 0 4770 0 -1 250
box -14 -8 132 252
use OAI21X1  _1482_
timestamp 1728305162
transform 1 0 4990 0 -1 730
box -12 -8 112 252
use NAND3X1  _1483_
timestamp 1728305047
transform -1 0 4630 0 1 250
box -12 -8 112 252
use NAND3X1  _1484_
timestamp 1728305047
transform 1 0 4410 0 1 250
box -12 -8 112 252
use NAND2X1  _1485_
timestamp 1728304996
transform -1 0 2950 0 1 4570
box -12 -8 92 252
use NAND2X1  _1486_
timestamp 1728304996
transform 1 0 2970 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1487_
timestamp 1728305162
transform 1 0 2870 0 -1 4570
box -12 -8 112 252
use INVX1  _1488_
timestamp 1728304789
transform 1 0 2730 0 -1 5050
box -12 -8 72 252
use NAND2X1  _1489_
timestamp 1728304996
transform 1 0 3390 0 1 4570
box -12 -8 92 252
use OAI21X1  _1490_
timestamp 1728305162
transform 1 0 3250 0 1 4570
box -12 -8 112 252
use INVX1  _1491_
timestamp 1728304789
transform 1 0 2790 0 -1 4570
box -12 -8 72 252
use NAND2X1  _1492_
timestamp 1728304996
transform 1 0 3170 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1493_
timestamp 1728305162
transform 1 0 3070 0 -1 4570
box -12 -8 112 252
use INVX1  _1494_
timestamp 1728304789
transform 1 0 3270 0 -1 4570
box -12 -8 72 252
use NAND2X1  _1495_
timestamp 1728304996
transform 1 0 3470 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1496_
timestamp 1728305162
transform 1 0 3370 0 -1 4570
box -12 -8 112 252
use AND2X2  _1497_
timestamp 1728304163
transform 1 0 2730 0 1 4570
box -12 -8 112 252
use AND2X2  _1498_
timestamp 1728304163
transform 1 0 2970 0 1 4570
box -12 -8 112 252
use AND2X2  _1499_
timestamp 1728304163
transform 1 0 2630 0 -1 5050
box -12 -8 112 252
use INVX1  _1500_
timestamp 1728304789
transform -1 0 110 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1501_
timestamp 1728304996
transform 1 0 230 0 1 6010
box -12 -8 92 252
use OAI21X1  _1502_
timestamp 1728305162
transform 1 0 150 0 1 5530
box -12 -8 112 252
use INVX1  _1503_
timestamp 1728304789
transform -1 0 170 0 -1 5050
box -12 -8 72 252
use NAND2X1  _1504_
timestamp 1728304996
transform -1 0 130 0 1 5530
box -12 -8 92 252
use OAI21X1  _1505_
timestamp 1728305162
transform -1 0 110 0 -1 5050
box -12 -8 112 252
use INVX1  _1506_
timestamp 1728304789
transform -1 0 270 0 -1 6010
box -12 -8 72 252
use NAND2X1  _1507_
timestamp 1728304996
transform 1 0 490 0 1 6010
box -12 -8 92 252
use OAI21X1  _1508_
timestamp 1728305162
transform 1 0 310 0 -1 6010
box -12 -8 112 252
use INVX1  _1509_
timestamp 1728304789
transform -1 0 290 0 -1 2650
box -12 -8 72 252
use NAND2X1  _1510_
timestamp 1728304996
transform -1 0 90 0 -1 2650
box -12 -8 92 252
use OAI21X1  _1511_
timestamp 1728305162
transform -1 0 230 0 -1 2650
box -12 -8 112 252
use INVX1  _1512_
timestamp 1728304789
transform 1 0 670 0 1 6010
box -12 -8 72 252
use NAND2X1  _1513_
timestamp 1728304996
transform -1 0 410 0 1 6010
box -12 -8 92 252
use OAI21X1  _1514_
timestamp 1728305162
transform 1 0 570 0 1 6010
box -12 -8 112 252
use INVX1  _1515_
timestamp 1728304789
transform -1 0 310 0 -1 3130
box -12 -8 72 252
use NAND2X1  _1516_
timestamp 1728304996
transform -1 0 90 0 -1 3130
box -12 -8 92 252
use OAI21X1  _1517_
timestamp 1728305162
transform -1 0 210 0 -1 3130
box -12 -8 112 252
use INVX1  _1518_
timestamp 1728304789
transform 1 0 370 0 1 5050
box -12 -8 72 252
use NAND2X1  _1519_
timestamp 1728304996
transform -1 0 230 0 1 6010
box -12 -8 92 252
use OAI21X1  _1520_
timestamp 1728305162
transform -1 0 450 0 -1 5530
box -12 -8 112 252
use INVX1  _1521_
timestamp 1728304789
transform -1 0 330 0 1 5530
box -12 -8 72 252
use NAND2X1  _1522_
timestamp 1728304996
transform 1 0 410 0 1 6010
box -12 -8 92 252
use OAI21X1  _1523_
timestamp 1728305162
transform 1 0 370 0 1 5530
box -12 -8 112 252
use INVX1  _1524_
timestamp 1728304789
transform -1 0 1870 0 1 5050
box -12 -8 72 252
use INVX1  _1525_
timestamp 1728304789
transform 1 0 650 0 -1 6010
box -12 -8 72 252
use NOR2X1  _1526_
timestamp 1728305106
transform 1 0 1470 0 -1 6010
box -12 -8 92 252
use INVX1  _1527_
timestamp 1728304789
transform 1 0 950 0 1 5530
box -12 -8 72 252
use NOR2X1  _1528_
timestamp 1728305106
transform -1 0 1050 0 -1 6010
box -12 -8 92 252
use NAND3X1  _1529_
timestamp 1728305047
transform 1 0 1270 0 -1 6010
box -12 -8 112 252
use NOR2X1  _1530_
timestamp 1728305106
transform 1 0 570 0 -1 5530
box -12 -8 92 252
use INVX1  _1531_
timestamp 1728304789
transform -1 0 1430 0 -1 6010
box -12 -8 72 252
use NOR2X1  _1532_
timestamp 1728305106
transform -1 0 910 0 -1 5530
box -12 -8 92 252
use NAND3X1  _1533_
timestamp 1728305047
transform 1 0 710 0 -1 5530
box -12 -8 112 252
use NAND2X1  _1534_
timestamp 1728304996
transform 1 0 1390 0 1 5530
box -12 -8 92 252
use INVX1  _1535_
timestamp 1728304789
transform -1 0 710 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1536_
timestamp 1728304996
transform -1 0 1150 0 -1 6010
box -12 -8 92 252
use NAND3X1  _1537_
timestamp 1728305047
transform -1 0 1350 0 1 5530
box -12 -8 112 252
use OAI21X1  _1538_
timestamp 1728305162
transform -1 0 1250 0 1 5530
box -12 -8 112 252
use OAI21X1  _1539_
timestamp 1728305162
transform -1 0 1110 0 1 5530
box -12 -8 112 252
use OAI21X1  _1540_
timestamp 1728305162
transform 1 0 2070 0 1 5530
box -12 -8 112 252
use AND2X2  _1541_
timestamp 1728304163
transform -1 0 1930 0 1 5530
box -12 -8 112 252
use NAND3X1  _1542_
timestamp 1728305047
transform -1 0 2050 0 1 5530
box -12 -8 112 252
use NOR2X1  _1543_
timestamp 1728305106
transform -1 0 1890 0 -1 6010
box -12 -8 92 252
use INVX1  _1544_
timestamp 1728304789
transform -1 0 1930 0 1 6010
box -12 -8 72 252
use NOR2X1  _1545_
timestamp 1728305106
transform -1 0 1270 0 -1 6010
box -12 -8 92 252
use NAND2X1  _1546_
timestamp 1728304996
transform -1 0 1770 0 1 6010
box -12 -8 92 252
use AOI21X1  _1547_
timestamp 1728304211
transform -1 0 1590 0 1 5530
box -12 -8 112 252
use NAND3X1  _1548_
timestamp 1728305047
transform -1 0 1870 0 1 6010
box -12 -8 112 252
use NOR2X1  _1549_
timestamp 1728305106
transform 1 0 1610 0 1 6010
box -12 -8 92 252
use INVX1  _1550_
timestamp 1728304789
transform 1 0 3570 0 1 6010
box -12 -8 72 252
use NAND2X1  _1551_
timestamp 1728304996
transform -1 0 3730 0 1 6010
box -12 -8 92 252
use AOI21X1  _1552_
timestamp 1728304211
transform 1 0 3730 0 1 6010
box -12 -8 112 252
use INVX1  _1553_
timestamp 1728304789
transform -1 0 1230 0 1 5050
box -12 -8 72 252
use NAND2X1  _1554_
timestamp 1728304996
transform -1 0 1230 0 -1 5530
box -12 -8 92 252
use AOI21X1  _1555_
timestamp 1728304211
transform 1 0 1250 0 -1 5530
box -12 -8 112 252
use DFFPOSX1  _1556_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728340458
transform -1 0 950 0 1 5530
box -13 -8 253 252
use DFFPOSX1  _1557_
timestamp 1728340458
transform -1 0 1830 0 1 5530
box -13 -8 253 252
use DFFPOSX1  _1558_
timestamp 1728340458
transform -1 0 1790 0 -1 6010
box -13 -8 253 252
use DFFPOSX1  _1559_
timestamp 1728340458
transform -1 0 1150 0 -1 5530
box -13 -8 253 252
use DFFPOSX1  _1560_
timestamp 1728340458
transform -1 0 950 0 -1 6010
box -13 -8 253 252
use DFFPOSX1  _1561_
timestamp 1728340458
transform -1 0 4070 0 1 6010
box -13 -8 253 252
use DFFPOSX1  _1562_
timestamp 1728340458
transform 1 0 1470 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _1563_
timestamp 1728340458
transform 1 0 110 0 -1 5530
box -13 -8 253 252
use DFFPOSX1  _1564_
timestamp 1728340458
transform 1 0 170 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _1565_
timestamp 1728340458
transform 1 0 410 0 -1 6010
box -13 -8 253 252
use DFFPOSX1  _1566_
timestamp 1728340458
transform 1 0 10 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _1567_
timestamp 1728340458
transform -1 0 970 0 1 6010
box -13 -8 253 252
use DFFPOSX1  _1568_
timestamp 1728340458
transform 1 0 310 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _1569_
timestamp 1728340458
transform -1 0 370 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _1570_
timestamp 1728340458
transform 1 0 470 0 1 5530
box -13 -8 253 252
use INVX1  _1571_
timestamp 1728304789
transform 1 0 3870 0 -1 1210
box -12 -8 72 252
use NOR2X1  _1572_
timestamp 1728305106
transform -1 0 3890 0 -1 1690
box -12 -8 92 252
use INVX2  _1573_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304826
transform -1 0 3870 0 -1 1210
box -12 -8 72 252
use NAND2X1  _1574_
timestamp 1728304996
transform 1 0 3730 0 -1 1210
box -12 -8 92 252
use INVX1  _1575_
timestamp 1728304789
transform 1 0 3890 0 1 2650
box -12 -8 72 252
use NAND2X1  _1576_
timestamp 1728304996
transform 1 0 3070 0 1 250
box -12 -8 92 252
use INVX1  _1577_
timestamp 1728304789
transform -1 0 3550 0 1 1690
box -12 -8 72 252
use NAND2X1  _1578_
timestamp 1728304996
transform 1 0 3770 0 1 730
box -12 -8 92 252
use AND2X2  _1579_
timestamp 1728304163
transform -1 0 3450 0 -1 250
box -12 -8 112 252
use NOR2X1  _1580_
timestamp 1728305106
transform -1 0 3290 0 1 250
box -12 -8 92 252
use NAND3X1  _1581_
timestamp 1728305047
transform -1 0 3410 0 1 250
box -12 -8 112 252
use INVX1  _1582_
timestamp 1728304789
transform 1 0 3670 0 -1 1210
box -12 -8 72 252
use NOR2X1  _1583_
timestamp 1728305106
transform -1 0 3390 0 1 730
box -12 -8 92 252
use INVX4  _1584_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304878
transform -1 0 4590 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1585_
timestamp 1728304996
transform 1 0 4550 0 1 1690
box -12 -8 92 252
use NAND2X1  _1586_
timestamp 1728304996
transform -1 0 4710 0 1 1690
box -12 -8 92 252
use NAND2X1  _1587_
timestamp 1728304996
transform 1 0 4810 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1588_
timestamp 1728304996
transform 1 0 4430 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1589_
timestamp 1728304996
transform -1 0 4310 0 1 1690
box -12 -8 92 252
use NAND2X1  _1590_
timestamp 1728304996
transform -1 0 4210 0 1 1690
box -12 -8 92 252
use NAND2X1  _1591_
timestamp 1728304996
transform 1 0 5530 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1592_
timestamp 1728304996
transform 1 0 5770 0 1 2170
box -12 -8 92 252
use NAND2X1  _1593_
timestamp 1728304996
transform -1 0 5750 0 1 2170
box -12 -8 92 252
use NAND2X1  _1594_
timestamp 1728304996
transform 1 0 4690 0 1 1210
box -12 -8 92 252
use NAND2X1  _1595_
timestamp 1728304996
transform 1 0 5170 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1596_
timestamp 1728304996
transform -1 0 4950 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1597_
timestamp 1728304996
transform 1 0 5430 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1598_
timestamp 1728304996
transform 1 0 6050 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1599_
timestamp 1728304996
transform -1 0 5630 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1600_
timestamp 1728304996
transform 1 0 5090 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1601_
timestamp 1728304996
transform 1 0 5430 0 -1 2170
box -12 -8 92 252
use NAND2X1  _1602_
timestamp 1728304996
transform -1 0 5470 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1603_
timestamp 1728304996
transform 1 0 4470 0 1 1210
box -12 -8 92 252
use NAND2X1  _1604_
timestamp 1728304996
transform 1 0 4690 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1605_
timestamp 1728304996
transform -1 0 4670 0 -1 1690
box -12 -8 92 252
use NAND2X1  _1606_
timestamp 1728304996
transform -1 0 4990 0 1 1210
box -12 -8 92 252
use NAND2X1  _1607_
timestamp 1728304996
transform 1 0 5210 0 1 1210
box -12 -8 92 252
use NAND2X1  _1608_
timestamp 1728304996
transform -1 0 5210 0 1 1210
box -12 -8 92 252
use NAND2X1  _1609_
timestamp 1728304996
transform -1 0 6610 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1610_
timestamp 1728304996
transform 1 0 7030 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1611_
timestamp 1728304996
transform 1 0 7090 0 1 1210
box -12 -8 92 252
use NAND2X1  _1612_
timestamp 1728304996
transform -1 0 6690 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1613_
timestamp 1728304996
transform 1 0 7330 0 1 1210
box -12 -8 92 252
use NAND2X1  _1614_
timestamp 1728304996
transform 1 0 7410 0 1 1210
box -12 -8 92 252
use NAND2X1  _1615_
timestamp 1728304996
transform -1 0 6690 0 -1 730
box -12 -8 92 252
use NAND2X1  _1616_
timestamp 1728304996
transform 1 0 6910 0 -1 730
box -12 -8 92 252
use NAND2X1  _1617_
timestamp 1728304996
transform -1 0 6910 0 -1 730
box -12 -8 92 252
use NAND2X1  _1618_
timestamp 1728304996
transform -1 0 6390 0 1 250
box -12 -8 92 252
use NAND2X1  _1619_
timestamp 1728304996
transform -1 0 6710 0 1 250
box -12 -8 92 252
use NAND2X1  _1620_
timestamp 1728304996
transform -1 0 6470 0 1 250
box -12 -8 92 252
use NAND2X1  _1621_
timestamp 1728304996
transform -1 0 4890 0 1 250
box -12 -8 92 252
use NAND2X1  _1622_
timestamp 1728304996
transform -1 0 5270 0 1 250
box -12 -8 92 252
use NAND2X1  _1623_
timestamp 1728304996
transform -1 0 5090 0 1 250
box -12 -8 92 252
use NAND2X1  _1624_
timestamp 1728304996
transform 1 0 5790 0 -1 730
box -12 -8 92 252
use NAND2X1  _1625_
timestamp 1728304996
transform 1 0 6110 0 -1 730
box -12 -8 92 252
use NAND2X1  _1626_
timestamp 1728304996
transform -1 0 6090 0 -1 730
box -12 -8 92 252
use NAND2X1  _1627_
timestamp 1728304996
transform -1 0 5810 0 -1 1210
box -12 -8 92 252
use NAND2X1  _1628_
timestamp 1728304996
transform 1 0 6510 0 1 1210
box -12 -8 92 252
use NAND2X1  _1629_
timestamp 1728304996
transform -1 0 6370 0 1 1210
box -12 -8 92 252
use NAND2X1  _1630_
timestamp 1728304996
transform 1 0 5310 0 1 730
box -12 -8 92 252
use NAND2X1  _1631_
timestamp 1728304996
transform 1 0 5650 0 1 730
box -12 -8 92 252
use NAND2X1  _1632_
timestamp 1728304996
transform -1 0 5650 0 1 730
box -12 -8 92 252
use INVX1  _1633_
timestamp 1728304789
transform 1 0 4230 0 -1 4090
box -12 -8 72 252
use INVX1  _1634_
timestamp 1728304789
transform 1 0 3830 0 -1 4090
box -12 -8 72 252
use INVX1  _1635_
timestamp 1728304789
transform -1 0 3790 0 1 3610
box -12 -8 72 252
use OR2X2  _1636_
timestamp 1728305284
transform 1 0 1250 0 1 6010
box -12 -8 112 252
use NAND3X1  _1637_
timestamp 1728305047
transform 1 0 3610 0 -1 730
box -12 -8 112 252
use NAND3X1  _1638_
timestamp 1728305047
transform 1 0 3810 0 -1 730
box -12 -8 112 252
use NAND2X1  _1639_
timestamp 1728304996
transform 1 0 3710 0 -1 730
box -12 -8 92 252
use OAI21X1  _1640_
timestamp 1728305162
transform 1 0 3670 0 1 730
box -12 -8 112 252
use NAND3X1  _1641_
timestamp 1728305047
transform -1 0 3670 0 -1 1210
box -12 -8 112 252
use AND2X2  _1642_
timestamp 1728304163
transform -1 0 3490 0 1 730
box -12 -8 112 252
use NAND3X1  _1643_
timestamp 1728305047
transform -1 0 3630 0 1 730
box -12 -8 112 252
use NOR2X1  _1644_
timestamp 1728305106
transform -1 0 3370 0 -1 730
box -12 -8 92 252
use MUX2X1  _1645_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304958
transform -1 0 3050 0 -1 730
box -12 -8 131 252
use INVX1  _1646_
timestamp 1728304789
transform 1 0 3150 0 1 250
box -12 -8 72 252
use OAI21X1  _1647_
timestamp 1728305162
transform -1 0 3310 0 -1 250
box -12 -8 112 252
use INVX1  _1648_
timestamp 1728304789
transform -1 0 3070 0 1 250
box -12 -8 72 252
use NAND3X1  _1649_
timestamp 1728305047
transform -1 0 3010 0 1 250
box -12 -8 112 252
use NAND2X1  _1650_
timestamp 1728304996
transform -1 0 2930 0 -1 250
box -12 -8 92 252
use AOI21X1  _1651_
timestamp 1728304211
transform -1 0 4530 0 1 1690
box -12 -8 112 252
use AOI21X1  _1652_
timestamp 1728304211
transform -1 0 4190 0 -1 1690
box -12 -8 112 252
use AOI21X1  _1653_
timestamp 1728304211
transform -1 0 5670 0 1 2170
box -12 -8 112 252
use AOI21X1  _1654_
timestamp 1728304211
transform -1 0 4870 0 1 1210
box -12 -8 112 252
use AOI21X1  _1655_
timestamp 1728304211
transform -1 0 5650 0 -1 1210
box -12 -8 112 252
use AOI21X1  _1656_
timestamp 1728304211
transform -1 0 5350 0 -1 1690
box -12 -8 112 252
use AOI21X1  _1657_
timestamp 1728304211
transform -1 0 4650 0 1 1210
box -12 -8 112 252
use AOI21X1  _1658_
timestamp 1728304211
transform -1 0 5130 0 1 1210
box -12 -8 112 252
use AOI21X1  _1659_
timestamp 1728304211
transform -1 0 7030 0 -1 1210
box -12 -8 112 252
use AOI21X1  _1660_
timestamp 1728304211
transform -1 0 7290 0 1 1210
box -12 -8 112 252
use AOI21X1  _1661_
timestamp 1728304211
transform -1 0 6790 0 -1 730
box -12 -8 112 252
use AOI21X1  _1662_
timestamp 1728304211
transform 1 0 6510 0 1 250
box -12 -8 112 252
use AOI21X1  _1663_
timestamp 1728304211
transform 1 0 5090 0 1 250
box -12 -8 112 252
use AOI21X1  _1664_
timestamp 1728304211
transform -1 0 5790 0 -1 730
box -12 -8 112 252
use AOI21X1  _1665_
timestamp 1728304211
transform -1 0 6290 0 1 1210
box -12 -8 112 252
use AOI21X1  _1666_
timestamp 1728304211
transform -1 0 5530 0 1 730
box -12 -8 112 252
use NOR2X1  _1667_
timestamp 1728305106
transform 1 0 4110 0 1 3610
box -12 -8 92 252
use NOR2X1  _1668_
timestamp 1728305106
transform -1 0 3990 0 -1 4090
box -12 -8 92 252
use OAI21X1  _1669_
timestamp 1728305162
transform 1 0 3890 0 1 1210
box -12 -8 112 252
use NAND3X1  _1670_
timestamp 1728305047
transform 1 0 3490 0 -1 250
box -12 -8 112 252
use OAI21X1  _1671_
timestamp 1728305162
transform -1 0 3890 0 1 1210
box -12 -8 112 252
use NOR2X1  _1672_
timestamp 1728305106
transform -1 0 3950 0 -1 3610
box -12 -8 92 252
use NOR2X1  _1673_
timestamp 1728305106
transform -1 0 3730 0 1 3610
box -12 -8 92 252
use NOR2X1  _1674_
timestamp 1728305106
transform 1 0 1490 0 1 6010
box -12 -8 92 252
use AND2X2  _1675_
timestamp 1728304163
transform -1 0 1470 0 1 6010
box -12 -8 112 252
use DFFPOSX1  _1676_
timestamp 1728340458
transform 1 0 3370 0 -1 730
box -13 -8 253 252
use DFFPOSX1  _1677_
timestamp 1728340458
transform 1 0 3030 0 1 730
box -13 -8 253 252
use DFFPOSX1  _1678_
timestamp 1728340458
transform 1 0 2650 0 1 250
box -13 -8 253 252
use DFFPOSX1  _1679_
timestamp 1728340458
transform 1 0 2930 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _1680_
timestamp 1728340458
transform 1 0 650 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _1681_
timestamp 1728340458
transform -1 0 1470 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _1682_
timestamp 1728340458
transform -1 0 1130 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _1683_
timestamp 1728340458
transform -1 0 4770 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _1684_
timestamp 1728340458
transform 1 0 4190 0 -1 1690
box -13 -8 253 252
use DFFPOSX1  _1685_
timestamp 1728340458
transform 1 0 5310 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _1686_
timestamp 1728340458
transform -1 0 4850 0 -1 1210
box -13 -8 253 252
use DFFPOSX1  _1687_
timestamp 1728340458
transform -1 0 5330 0 -1 1210
box -13 -8 253 252
use DFFPOSX1  _1688_
timestamp 1728340458
transform -1 0 4470 0 -1 1210
box -13 -8 253 252
use DFFPOSX1  _1689_
timestamp 1728340458
transform -1 0 4470 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _1690_
timestamp 1728340458
transform -1 0 5090 0 -1 1210
box -13 -8 253 252
use DFFPOSX1  _1691_
timestamp 1728340458
transform -1 0 6930 0 -1 1210
box -13 -8 253 252
use DFFPOSX1  _1692_
timestamp 1728340458
transform -1 0 7070 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _1693_
timestamp 1728340458
transform -1 0 6830 0 1 730
box -13 -8 253 252
use DFFPOSX1  _1694_
timestamp 1728340458
transform -1 0 7130 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _1695_
timestamp 1728340458
transform -1 0 5610 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _1696_
timestamp 1728340458
transform -1 0 5670 0 -1 730
box -13 -8 253 252
use DFFPOSX1  _1697_
timestamp 1728340458
transform -1 0 6190 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _1698_
timestamp 1728340458
transform 1 0 5050 0 1 730
box -13 -8 253 252
use DFFPOSX1  _1699_
timestamp 1728340458
transform 1 0 4150 0 1 3130
box -13 -8 253 252
use DFFPOSX1  _1700_
timestamp 1728340458
transform 1 0 3990 0 -1 4090
box -13 -8 253 252
use DFFPOSX1  _1701_
timestamp 1728340458
transform -1 0 4030 0 1 3610
box -13 -8 253 252
use DFFPOSX1  _1702_
timestamp 1728340458
transform 1 0 3570 0 -1 4090
box -13 -8 253 252
use DFFPOSX1  _1703_
timestamp 1728340458
transform 1 0 970 0 1 6010
box -13 -8 253 252
use INVX2  _1704_
timestamp 1728304826
transform 1 0 3530 0 -1 5050
box -12 -8 72 252
use NAND2X1  _1705_
timestamp 1728304996
transform 1 0 4090 0 1 4570
box -12 -8 92 252
use INVX1  _1706_
timestamp 1728304789
transform -1 0 3590 0 1 4090
box -12 -8 72 252
use INVX1  _1707_
timestamp 1728304789
transform -1 0 3530 0 1 4090
box -12 -8 72 252
use OAI21X1  _1708_
timestamp 1728305162
transform -1 0 3450 0 1 4090
box -12 -8 112 252
use INVX1  _1709_
timestamp 1728304789
transform -1 0 3570 0 1 4570
box -12 -8 72 252
use OAI21X1  _1710_
timestamp 1728305162
transform -1 0 3650 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1711_
timestamp 1728305047
transform -1 0 3350 0 1 4090
box -12 -8 112 252
use NAND2X1  _1712_
timestamp 1728304996
transform -1 0 4110 0 -1 4570
box -12 -8 92 252
use NAND2X1  _1713_
timestamp 1728304996
transform 1 0 3970 0 1 4570
box -12 -8 92 252
use NAND2X1  _1714_
timestamp 1728304996
transform 1 0 3650 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1715_
timestamp 1728305162
transform 1 0 3590 0 1 4570
box -12 -8 112 252
use OAI21X1  _1716_
timestamp 1728305162
transform 1 0 3730 0 -1 4570
box -12 -8 112 252
use OAI21X1  _1717_
timestamp 1728305162
transform 1 0 3730 0 1 4570
box -12 -8 112 252
use INVX1  _1718_
timestamp 1728304789
transform -1 0 4030 0 -1 5050
box -12 -8 72 252
use AOI21X1  _1719_
timestamp 1728304211
transform 1 0 3830 0 1 4570
box -12 -8 112 252
use NAND2X1  _1720_
timestamp 1728304996
transform 1 0 3870 0 -1 4570
box -12 -8 92 252
use AOI22X1  _1721_
timestamp 1728304278
transform -1 0 3970 0 -1 5050
box -14 -8 132 252
use INVX1  _1722_
timestamp 1728304789
transform -1 0 3690 0 -1 5530
box -12 -8 72 252
use AOI21X1  _1723_
timestamp 1728304211
transform 1 0 3750 0 -1 5050
box -12 -8 112 252
use AOI22X1  _1724_
timestamp 1728304278
transform 1 0 3630 0 -1 5050
box -14 -8 132 252
use DFFPOSX1  _1725_
timestamp 1728340458
transform -1 0 4350 0 -1 4570
box -13 -8 253 252
use DFFPOSX1  _1726_
timestamp 1728340458
transform 1 0 3410 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _1727_
timestamp 1728340458
transform 1 0 4030 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _1728_
timestamp 1728340458
transform 1 0 3370 0 -1 5530
box -13 -8 253 252
use INVX1  _1729_
timestamp 1728304789
transform 1 0 2030 0 1 6010
box -12 -8 72 252
use INVX1  _1730_
timestamp 1728304789
transform 1 0 2230 0 -1 6010
box -12 -8 72 252
use NAND2X1  _1731_
timestamp 1728304996
transform 1 0 2130 0 -1 6010
box -12 -8 92 252
use NAND2X1  _1732_
timestamp 1728304996
transform 1 0 2130 0 1 6010
box -12 -8 92 252
use INVX1  _1733_
timestamp 1728304789
transform 1 0 2670 0 1 6010
box -12 -8 72 252
use NOR2X1  _1734_
timestamp 1728305106
transform 1 0 2310 0 -1 6010
box -12 -8 92 252
use AOI21X1  _1735_
timestamp 1728304211
transform -1 0 2030 0 1 6010
box -12 -8 112 252
use NOR2X1  _1736_
timestamp 1728305106
transform 1 0 2250 0 1 6010
box -12 -8 92 252
use OAI21X1  _1737_
timestamp 1728305162
transform -1 0 2430 0 1 6010
box -12 -8 112 252
use DFFPOSX1  _1738_
timestamp 1728340458
transform 1 0 1890 0 -1 6010
box -13 -8 253 252
use DFFPOSX1  _1739_
timestamp 1728340458
transform 1 0 2430 0 1 6010
box -13 -8 253 252
use INVX1  _1740_
timestamp 1728304789
transform -1 0 4970 0 -1 4090
box -12 -8 72 252
use NAND2X1  _1741_
timestamp 1728304996
transform -1 0 4030 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1742_
timestamp 1728305162
transform 1 0 3850 0 1 4090
box -12 -8 112 252
use INVX2  _1743_
timestamp 1728304826
transform -1 0 4710 0 1 4570
box -12 -8 72 252
use NAND2X1  _1744_
timestamp 1728304996
transform -1 0 4190 0 1 5050
box -12 -8 92 252
use OAI21X1  _1745_
timestamp 1728305162
transform -1 0 4330 0 1 5050
box -12 -8 112 252
use INVX2  _1746_
timestamp 1728304826
transform 1 0 4730 0 1 5050
box -12 -8 72 252
use NAND2X1  _1747_
timestamp 1728304996
transform -1 0 4370 0 -1 5050
box -12 -8 92 252
use OAI21X1  _1748_
timestamp 1728305162
transform -1 0 4470 0 -1 5050
box -12 -8 112 252
use INVX2  _1749_
timestamp 1728304826
transform -1 0 4430 0 1 5050
box -12 -8 72 252
use NAND2X1  _1750_
timestamp 1728304996
transform -1 0 4050 0 -1 6010
box -12 -8 92 252
use OAI21X1  _1751_
timestamp 1728305162
transform -1 0 4170 0 -1 6010
box -12 -8 112 252
use INVX2  _1752_
timestamp 1728304826
transform -1 0 4730 0 1 5050
box -12 -8 72 252
use NAND2X1  _1753_
timestamp 1728304996
transform -1 0 4290 0 1 4570
box -12 -8 92 252
use OAI21X1  _1754_
timestamp 1728305162
transform -1 0 4390 0 1 4570
box -12 -8 112 252
use INVX2  _1755_
timestamp 1728304826
transform -1 0 3950 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1756_
timestamp 1728304996
transform -1 0 3730 0 1 5050
box -12 -8 92 252
use OAI21X1  _1757_
timestamp 1728305162
transform -1 0 3870 0 1 5050
box -12 -8 112 252
use INVX1  _1758_
timestamp 1728304789
transform -1 0 4550 0 -1 4090
box -12 -8 72 252
use NAND2X1  _1759_
timestamp 1728304996
transform -1 0 4270 0 -1 2650
box -12 -8 92 252
use OAI21X1  _1760_
timestamp 1728305162
transform -1 0 4630 0 -1 3610
box -12 -8 112 252
use INVX1  _1761_
timestamp 1728304789
transform -1 0 4630 0 1 3610
box -12 -8 72 252
use NAND2X1  _1762_
timestamp 1728304996
transform -1 0 4150 0 -1 3610
box -12 -8 92 252
use OAI21X1  _1763_
timestamp 1728305162
transform -1 0 4250 0 -1 3610
box -12 -8 112 252
use INVX2  _1764_
timestamp 1728304826
transform -1 0 4810 0 1 4570
box -12 -8 72 252
use NAND2X1  _1765_
timestamp 1728304996
transform -1 0 4610 0 -1 2650
box -12 -8 92 252
use OAI21X1  _1766_
timestamp 1728305162
transform -1 0 4830 0 1 3130
box -12 -8 112 252
use INVX1  _1767_
timestamp 1728304789
transform 1 0 4570 0 -1 4570
box -12 -8 72 252
use NAND2X1  _1768_
timestamp 1728304996
transform 1 0 4630 0 1 3130
box -12 -8 92 252
use OAI21X1  _1769_
timestamp 1728305162
transform 1 0 4550 0 -1 4090
box -12 -8 112 252
use INVX1  _1770_
timestamp 1728304789
transform -1 0 4790 0 -1 5050
box -12 -8 72 252
use NAND2X1  _1771_
timestamp 1728304996
transform -1 0 4110 0 1 3610
box -12 -8 92 252
use OAI21X1  _1772_
timestamp 1728305162
transform -1 0 4330 0 1 3610
box -12 -8 112 252
use INVX2  _1773_
timestamp 1728304826
transform -1 0 4490 0 1 5050
box -12 -8 72 252
use NAND2X1  _1774_
timestamp 1728304996
transform 1 0 4210 0 -1 3130
box -12 -8 92 252
use OAI21X1  _1775_
timestamp 1728305162
transform -1 0 4290 0 1 4090
box -12 -8 112 252
use INVX2  _1776_
timestamp 1728304826
transform -1 0 3870 0 -1 5530
box -12 -8 72 252
use NAND2X1  _1777_
timestamp 1728304996
transform -1 0 3410 0 1 5050
box -12 -8 92 252
use OAI21X1  _1778_
timestamp 1728305162
transform -1 0 3790 0 -1 5530
box -12 -8 112 252
use INVX2  _1779_
timestamp 1728304826
transform 1 0 4070 0 1 5530
box -12 -8 72 252
use NAND2X1  _1780_
timestamp 1728304996
transform -1 0 3670 0 1 5530
box -12 -8 92 252
use OAI21X1  _1781_
timestamp 1728305162
transform -1 0 3790 0 1 5530
box -12 -8 112 252
use INVX1  _1782_
timestamp 1728304789
transform 1 0 4830 0 -1 3130
box -12 -8 72 252
use NAND3X1  _1783_
timestamp 1728305047
transform -1 0 5010 0 -1 3610
box -12 -8 112 252
use OAI21X1  _1784_
timestamp 1728305162
transform -1 0 4990 0 -1 3130
box -12 -8 112 252
use INVX1  _1785_
timestamp 1728304789
transform -1 0 4350 0 -1 2650
box -12 -8 72 252
use NAND2X1  _1786_
timestamp 1728304996
transform -1 0 5150 0 1 3130
box -12 -8 92 252
use NAND2X1  _1787_
timestamp 1728304996
transform -1 0 4750 0 1 3610
box -12 -8 92 252
use NOR2X1  _1788_
timestamp 1728305106
transform 1 0 5150 0 1 3130
box -12 -8 92 252
use INVX1  _1789_
timestamp 1728304789
transform -1 0 5210 0 -1 3130
box -12 -8 72 252
use OAI21X1  _1790_
timestamp 1728305162
transform -1 0 4970 0 1 3610
box -12 -8 112 252
use NAND3X1  _1791_
timestamp 1728305047
transform 1 0 5030 0 -1 3130
box -12 -8 112 252
use OAI21X1  _1792_
timestamp 1728305162
transform 1 0 4770 0 1 2650
box -12 -8 112 252
use INVX1  _1793_
timestamp 1728304789
transform 1 0 6010 0 1 2650
box -12 -8 72 252
use NAND2X1  _1794_
timestamp 1728304996
transform 1 0 5270 0 1 3130
box -12 -8 92 252
use NAND2X1  _1795_
timestamp 1728304996
transform -1 0 5270 0 1 3610
box -12 -8 92 252
use NAND2X1  _1796_
timestamp 1728304996
transform -1 0 5690 0 1 3610
box -12 -8 92 252
use OAI21X1  _1797_
timestamp 1728305162
transform 1 0 5410 0 1 3610
box -12 -8 112 252
use OAI21X1  _1798_
timestamp 1728305162
transform 1 0 5310 0 1 3610
box -12 -8 112 252
use OR2X2  _1799_
timestamp 1728305284
transform 1 0 5570 0 1 3130
box -12 -8 112 252
use OAI21X1  _1800_
timestamp 1728305162
transform 1 0 5090 0 1 3610
box -12 -8 112 252
use NAND3X1  _1801_
timestamp 1728305047
transform 1 0 5730 0 -1 3130
box -12 -8 112 252
use INVX1  _1802_
timestamp 1728304789
transform 1 0 6070 0 -1 3130
box -12 -8 72 252
use AOI21X1  _1803_
timestamp 1728304211
transform 1 0 5830 0 -1 3130
box -12 -8 112 252
use NOR2X1  _1804_
timestamp 1728305106
transform 1 0 6290 0 -1 3130
box -12 -8 92 252
use NAND2X1  _1805_
timestamp 1728304996
transform 1 0 6250 0 1 2650
box -12 -8 92 252
use OAI21X1  _1806_
timestamp 1728305162
transform -1 0 5930 0 1 2650
box -12 -8 112 252
use INVX1  _1807_
timestamp 1728304789
transform 1 0 5450 0 -1 3130
box -12 -8 72 252
use OR2X2  _1808_
timestamp 1728305284
transform 1 0 5350 0 1 3130
box -12 -8 112 252
use NAND2X1  _1809_
timestamp 1728304996
transform -1 0 4870 0 1 3610
box -12 -8 92 252
use INVX1  _1810_
timestamp 1728304789
transform 1 0 5590 0 -1 3610
box -12 -8 72 252
use AND2X2  _1811_
timestamp 1728304163
transform 1 0 5030 0 -1 3610
box -12 -8 112 252
use AND2X2  _1812_
timestamp 1728304163
transform 1 0 4970 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1813_
timestamp 1728304996
transform 1 0 5510 0 -1 3610
box -12 -8 92 252
use OAI21X1  _1814_
timestamp 1728305162
transform 1 0 5370 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1815_
timestamp 1728305047
transform 1 0 5670 0 -1 3610
box -12 -8 112 252
use OAI21X1  _1816_
timestamp 1728305162
transform 1 0 4970 0 1 3610
box -12 -8 112 252
use OAI21X1  _1817_
timestamp 1728305162
transform -1 0 5370 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1818_
timestamp 1728305047
transform 1 0 5130 0 -1 3610
box -12 -8 112 252
use NAND2X1  _1819_
timestamp 1728304996
transform 1 0 5890 0 -1 3610
box -12 -8 92 252
use OAI21X1  _1820_
timestamp 1728305162
transform 1 0 5770 0 -1 3610
box -12 -8 112 252
use AND2X2  _1821_
timestamp 1728304163
transform 1 0 5930 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1822_
timestamp 1728305047
transform 1 0 5970 0 -1 3610
box -12 -8 112 252
use NAND2X1  _1823_
timestamp 1728304996
transform -1 0 5870 0 1 3130
box -12 -8 92 252
use NAND3X1  _1824_
timestamp 1728305047
transform 1 0 5670 0 1 3130
box -12 -8 112 252
use OAI21X1  _1825_
timestamp 1728305162
transform -1 0 5570 0 1 3130
box -12 -8 112 252
use NAND3X1  _1826_
timestamp 1728305047
transform 1 0 5890 0 1 3130
box -12 -8 112 252
use AOI21X1  _1827_
timestamp 1728304211
transform -1 0 6030 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1828_
timestamp 1728305047
transform 1 0 6170 0 -1 3130
box -12 -8 112 252
use NAND2X1  _1829_
timestamp 1728304996
transform 1 0 5650 0 -1 3130
box -12 -8 92 252
use OAI22X1  _1830_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728305200
transform 1 0 5530 0 -1 3130
box -12 -8 132 252
use INVX1  _1831_
timestamp 1728304789
transform 1 0 6570 0 -1 2650
box -12 -8 72 252
use INVX1  _1832_
timestamp 1728304789
transform 1 0 6490 0 -1 3130
box -12 -8 72 252
use NAND2X1  _1833_
timestamp 1728304996
transform 1 0 5510 0 1 3610
box -12 -8 92 252
use OAI21X1  _1834_
timestamp 1728305162
transform 1 0 6090 0 -1 3610
box -12 -8 112 252
use INVX1  _1835_
timestamp 1728304789
transform -1 0 6250 0 -1 3610
box -12 -8 72 252
use NAND2X1  _1836_
timestamp 1728304996
transform -1 0 5270 0 -1 4090
box -12 -8 92 252
use INVX1  _1837_
timestamp 1728304789
transform -1 0 5570 0 -1 4090
box -12 -8 72 252
use AND2X2  _1838_
timestamp 1728304163
transform 1 0 4610 0 1 4090
box -12 -8 112 252
use NAND2X1  _1839_
timestamp 1728304996
transform -1 0 5150 0 -1 4090
box -12 -8 92 252
use OAI21X1  _1840_
timestamp 1728305162
transform 1 0 5310 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1841_
timestamp 1728305047
transform 1 0 5410 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1842_
timestamp 1728305047
transform 1 0 5670 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1843_
timestamp 1728304996
transform 1 0 5730 0 1 3610
box -12 -8 92 252
use NAND3X1  _1844_
timestamp 1728305047
transform 1 0 5570 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1845_
timestamp 1728305047
transform 1 0 5790 0 -1 4090
box -12 -8 112 252
use AND2X2  _1846_
timestamp 1728304163
transform 1 0 5510 0 1 4090
box -12 -8 112 252
use AOI22X1  _1847_
timestamp 1728304278
transform -1 0 5510 0 1 4090
box -14 -8 132 252
use AOI21X1  _1848_
timestamp 1728304211
transform -1 0 6010 0 1 3610
box -12 -8 112 252
use NAND3X1  _1849_
timestamp 1728305047
transform 1 0 6130 0 1 3610
box -12 -8 112 252
use NAND2X1  _1850_
timestamp 1728304996
transform 1 0 6230 0 1 3610
box -12 -8 92 252
use NAND2X1  _1851_
timestamp 1728304996
transform 1 0 6070 0 -1 4090
box -12 -8 92 252
use INVX1  _1852_
timestamp 1728304789
transform 1 0 6150 0 -1 4090
box -12 -8 72 252
use OAI21X1  _1853_
timestamp 1728305162
transform 1 0 6330 0 1 3610
box -12 -8 112 252
use NAND3X1  _1854_
timestamp 1728305047
transform -1 0 6350 0 -1 3610
box -12 -8 112 252
use INVX1  _1855_
timestamp 1728304789
transform 1 0 6490 0 -1 3610
box -12 -8 72 252
use AOI21X1  _1856_
timestamp 1728304211
transform 1 0 6010 0 1 3610
box -12 -8 112 252
use OAI21X1  _1857_
timestamp 1728305162
transform -1 0 6110 0 1 3130
box -12 -8 112 252
use NAND3X1  _1858_
timestamp 1728305047
transform 1 0 6230 0 1 3130
box -12 -8 112 252
use INVX1  _1859_
timestamp 1728304789
transform 1 0 6390 0 -1 3130
box -12 -8 72 252
use OAI21X1  _1860_
timestamp 1728305162
transform 1 0 6130 0 1 3130
box -12 -8 112 252
use NAND3X1  _1861_
timestamp 1728305047
transform 1 0 6350 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1862_
timestamp 1728305047
transform -1 0 6470 0 1 3130
box -12 -8 112 252
use AOI21X1  _1863_
timestamp 1728304211
transform 1 0 6550 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1864_
timestamp 1728305047
transform 1 0 6670 0 -1 3130
box -12 -8 112 252
use INVX1  _1865_
timestamp 1728304789
transform 1 0 6770 0 -1 3130
box -12 -8 72 252
use OAI21X1  _1866_
timestamp 1728305162
transform 1 0 6970 0 1 2650
box -12 -8 112 252
use INVX1  _1867_
timestamp 1728304789
transform 1 0 6690 0 1 2650
box -12 -8 72 252
use NOR2X1  _1868_
timestamp 1728305106
transform 1 0 6850 0 1 2650
box -12 -8 92 252
use NAND2X1  _1869_
timestamp 1728304996
transform 1 0 6750 0 1 2650
box -12 -8 92 252
use NAND3X1  _1870_
timestamp 1728305047
transform -1 0 6690 0 1 2650
box -12 -8 112 252
use OAI21X1  _1871_
timestamp 1728305162
transform -1 0 6570 0 -1 2650
box -12 -8 112 252
use INVX8  _1872_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304916
transform 1 0 6470 0 1 730
box -12 -8 133 252
use NAND2X1  _1873_
timestamp 1728304996
transform -1 0 6890 0 -1 2170
box -12 -8 92 252
use OAI21X1  _1874_
timestamp 1728305162
transform -1 0 6970 0 -1 3130
box -12 -8 112 252
use NAND2X1  _1875_
timestamp 1728304996
transform -1 0 6690 0 1 3130
box -12 -8 92 252
use OAI21X1  _1876_
timestamp 1728305162
transform 1 0 5810 0 1 3610
box -12 -8 112 252
use NAND2X1  _1877_
timestamp 1728304996
transform -1 0 4750 0 -1 4570
box -12 -8 92 252
use INVX1  _1878_
timestamp 1728304789
transform -1 0 4770 0 1 4090
box -12 -8 72 252
use AND2X2  _1879_
timestamp 1728304163
transform 1 0 4910 0 1 4090
box -12 -8 112 252
use NAND2X1  _1880_
timestamp 1728304996
transform -1 0 5090 0 1 4090
box -12 -8 92 252
use NAND2X1  _1881_
timestamp 1728304996
transform -1 0 4470 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1882_
timestamp 1728305162
transform -1 0 4590 0 1 4090
box -12 -8 112 252
use NAND3X1  _1883_
timestamp 1728305047
transform 1 0 4790 0 1 4090
box -12 -8 112 252
use NAND3X1  _1884_
timestamp 1728305047
transform 1 0 4470 0 -1 4570
box -12 -8 112 252
use NAND2X1  _1885_
timestamp 1728304996
transform 1 0 5270 0 -1 5050
box -12 -8 92 252
use NAND2X1  _1886_
timestamp 1728304996
transform -1 0 4950 0 -1 4570
box -12 -8 92 252
use NAND3X1  _1887_
timestamp 1728305047
transform 1 0 4770 0 -1 4570
box -12 -8 112 252
use AND2X2  _1888_
timestamp 1728304163
transform 1 0 6190 0 1 4090
box -12 -8 112 252
use NAND2X1  _1889_
timestamp 1728304996
transform -1 0 5070 0 -1 4570
box -12 -8 92 252
use INVX1  _1890_
timestamp 1728304789
transform 1 0 5750 0 -1 4570
box -12 -8 72 252
use AND2X2  _1891_
timestamp 1728304163
transform 1 0 5550 0 -1 4570
box -12 -8 112 252
use AND2X2  _1892_
timestamp 1728304163
transform 1 0 5670 0 1 4570
box -12 -8 112 252
use NAND2X1  _1893_
timestamp 1728304996
transform 1 0 5830 0 -1 4570
box -12 -8 92 252
use NAND2X1  _1894_
timestamp 1728304996
transform -1 0 5170 0 -1 4570
box -12 -8 92 252
use OAI21X1  _1895_
timestamp 1728305162
transform -1 0 5370 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1896_
timestamp 1728305047
transform 1 0 6070 0 -1 4570
box -12 -8 112 252
use NAND2X1  _1897_
timestamp 1728304996
transform -1 0 4370 0 1 4090
box -12 -8 92 252
use NAND3X1  _1898_
timestamp 1728305047
transform 1 0 4390 0 1 4090
box -12 -8 112 252
use NAND3X1  _1899_
timestamp 1728305047
transform 1 0 5170 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1900_
timestamp 1728305047
transform 1 0 5130 0 1 4090
box -12 -8 112 252
use NAND3X1  _1901_
timestamp 1728305047
transform 1 0 6350 0 -1 4090
box -12 -8 112 252
use AOI21X1  _1902_
timestamp 1728304211
transform 1 0 5250 0 1 4090
box -12 -8 112 252
use AOI22X1  _1903_
timestamp 1728304278
transform 1 0 5730 0 1 4090
box -14 -8 132 252
use OAI21X1  _1904_
timestamp 1728305162
transform 1 0 5890 0 1 4090
box -12 -8 112 252
use NAND3X1  _1905_
timestamp 1728305047
transform 1 0 6550 0 -1 4090
box -12 -8 112 252
use NAND2X1  _1906_
timestamp 1728304996
transform -1 0 6190 0 1 4090
box -12 -8 92 252
use OAI21X1  _1907_
timestamp 1728305162
transform 1 0 5990 0 1 4090
box -12 -8 112 252
use NAND3X1  _1908_
timestamp 1728305047
transform 1 0 6250 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1909_
timestamp 1728305047
transform 1 0 6450 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1910_
timestamp 1728305047
transform 1 0 6650 0 1 3610
box -12 -8 112 252
use NAND2X1  _1911_
timestamp 1728304996
transform -1 0 6550 0 1 3610
box -12 -8 92 252
use NAND2X1  _1912_
timestamp 1728304996
transform 1 0 6550 0 -1 3610
box -12 -8 92 252
use NAND3X1  _1913_
timestamp 1728305047
transform 1 0 7110 0 -1 3610
box -12 -8 112 252
use INVX1  _1914_
timestamp 1728304789
transform 1 0 7210 0 -1 3610
box -12 -8 72 252
use NAND2X1  _1915_
timestamp 1728304996
transform -1 0 6750 0 -1 3610
box -12 -8 92 252
use NAND3X1  _1916_
timestamp 1728305047
transform 1 0 6550 0 1 3610
box -12 -8 112 252
use NAND3X1  _1917_
timestamp 1728305047
transform 1 0 6990 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1918_
timestamp 1728305047
transform 1 0 7030 0 1 3130
box -12 -8 112 252
use AND2X2  _1919_
timestamp 1728304163
transform 1 0 6510 0 1 3130
box -12 -8 112 252
use NAND3X1  _1920_
timestamp 1728305047
transform -1 0 6970 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1921_
timestamp 1728305047
transform -1 0 6870 0 -1 3610
box -12 -8 112 252
use NAND3X1  _1922_
timestamp 1728305047
transform 1 0 6810 0 1 3130
box -12 -8 112 252
use AOI21X1  _1923_
timestamp 1728304211
transform -1 0 7110 0 -1 3130
box -12 -8 112 252
use NAND3X1  _1924_
timestamp 1728305047
transform 1 0 7110 0 -1 3130
box -12 -8 112 252
use NAND2X1  _1925_
timestamp 1728304996
transform 1 0 7450 0 1 2650
box -12 -8 92 252
use OAI21X1  _1926_
timestamp 1728305162
transform -1 0 7470 0 1 2170
box -12 -8 112 252
use NAND2X1  _1927_
timestamp 1728304996
transform 1 0 7270 0 -1 2650
box -12 -8 92 252
use NAND2X1  _1928_
timestamp 1728304996
transform 1 0 7230 0 -1 3130
box -12 -8 92 252
use INVX1  _1929_
timestamp 1728304789
transform 1 0 6990 0 1 3610
box -12 -8 72 252
use AOI21X1  _1930_
timestamp 1728304211
transform 1 0 7090 0 1 3610
box -12 -8 112 252
use AOI21X1  _1931_
timestamp 1728304211
transform 1 0 6290 0 1 4090
box -12 -8 112 252
use OAI21X1  _1932_
timestamp 1728305162
transform 1 0 6410 0 1 4090
box -12 -8 112 252
use NAND2X1  _1933_
timestamp 1728304996
transform -1 0 4350 0 -1 5530
box -12 -8 92 252
use INVX1  _1934_
timestamp 1728304789
transform 1 0 5170 0 -1 5050
box -12 -8 72 252
use AND2X2  _1935_
timestamp 1728304163
transform 1 0 4790 0 -1 5050
box -12 -8 112 252
use AND2X2  _1936_
timestamp 1728304163
transform -1 0 5110 0 1 4570
box -12 -8 112 252
use NAND2X1  _1937_
timestamp 1728304996
transform 1 0 4910 0 1 4570
box -12 -8 92 252
use NAND2X1  _1938_
timestamp 1728304996
transform -1 0 5450 0 1 4570
box -12 -8 92 252
use OAI21X1  _1939_
timestamp 1728305162
transform 1 0 5230 0 1 4570
box -12 -8 112 252
use NAND3X1  _1940_
timestamp 1728305047
transform -1 0 5230 0 1 4570
box -12 -8 112 252
use OAI21X1  _1941_
timestamp 1728305162
transform 1 0 4810 0 1 4570
box -12 -8 112 252
use OAI21X1  _1942_
timestamp 1728305162
transform -1 0 5010 0 -1 5050
box -12 -8 112 252
use NAND3X1  _1943_
timestamp 1728305047
transform 1 0 5030 0 -1 5050
box -12 -8 112 252
use NAND2X1  _1944_
timestamp 1728304996
transform -1 0 6590 0 -1 5050
box -12 -8 92 252
use AOI22X1  _1945_
timestamp 1728304278
transform -1 0 5530 0 -1 4570
box -14 -8 132 252
use OAI21X1  _1946_
timestamp 1728305162
transform 1 0 5650 0 -1 4570
box -12 -8 112 252
use NAND2X1  _1947_
timestamp 1728304996
transform -1 0 5970 0 1 4570
box -12 -8 92 252
use NAND2X1  _1948_
timestamp 1728304996
transform -1 0 5530 0 1 4570
box -12 -8 92 252
use NAND3X1  _1949_
timestamp 1728305047
transform 1 0 5570 0 1 4570
box -12 -8 112 252
use OAI21X1  _1950_
timestamp 1728305162
transform 1 0 5770 0 1 4570
box -12 -8 112 252
use AOI21X1  _1951_
timestamp 1728304211
transform 1 0 6130 0 1 4570
box -12 -8 112 252
use INVX1  _1952_
timestamp 1728304789
transform 1 0 6250 0 -1 5050
box -12 -8 72 252
use AND2X2  _1953_
timestamp 1728304163
transform 1 0 5690 0 -1 5050
box -12 -8 112 252
use NAND2X1  _1954_
timestamp 1728304996
transform -1 0 6090 0 -1 5050
box -12 -8 92 252
use OAI21X1  _1955_
timestamp 1728305162
transform 1 0 5810 0 -1 5050
box -12 -8 112 252
use AOI21X1  _1956_
timestamp 1728304211
transform -1 0 6410 0 -1 5050
box -12 -8 112 252
use OAI21X1  _1957_
timestamp 1728305162
transform 1 0 6310 0 -1 4570
box -12 -8 112 252
use AOI22X1  _1958_
timestamp 1728304278
transform 1 0 5910 0 -1 4570
box -14 -8 132 252
use NAND3X1  _1959_
timestamp 1728305047
transform 1 0 6410 0 -1 5050
box -12 -8 112 252
use NAND3X1  _1960_
timestamp 1728305047
transform 1 0 6010 0 1 4570
box -12 -8 112 252
use NAND3X1  _1961_
timestamp 1728305047
transform 1 0 6230 0 1 4570
box -12 -8 112 252
use AOI21X1  _1962_
timestamp 1728304211
transform 1 0 6530 0 -1 4570
box -12 -8 112 252
use AND2X2  _1963_
timestamp 1728304163
transform 1 0 6570 0 1 4570
box -12 -8 112 252
use NAND3X1  _1964_
timestamp 1728305047
transform 1 0 6470 0 1 4570
box -12 -8 112 252
use OAI21X1  _1965_
timestamp 1728305162
transform -1 0 6270 0 -1 4570
box -12 -8 112 252
use AOI21X1  _1966_
timestamp 1728304211
transform -1 0 6750 0 -1 4570
box -12 -8 112 252
use OAI21X1  _1967_
timestamp 1728305162
transform 1 0 6630 0 1 4090
box -12 -8 112 252
use INVX1  _1968_
timestamp 1728304789
transform 1 0 6790 0 -1 4090
box -12 -8 72 252
use AOI21X1  _1969_
timestamp 1728304211
transform 1 0 6650 0 -1 4090
box -12 -8 112 252
use NAND3X1  _1970_
timestamp 1728305047
transform 1 0 6770 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1971_
timestamp 1728305047
transform -1 0 6510 0 -1 4570
box -12 -8 112 252
use NAND3X1  _1972_
timestamp 1728305047
transform 1 0 6910 0 -1 4570
box -12 -8 112 252
use AOI22X1  _1973_
timestamp 1728304278
transform 1 0 6730 0 1 4090
box -14 -8 132 252
use OAI21X1  _1974_
timestamp 1728305162
transform -1 0 5730 0 1 4090
box -12 -8 112 252
use NAND3X1  _1975_
timestamp 1728305047
transform -1 0 7110 0 -1 4570
box -12 -8 112 252
use OAI21X1  _1976_
timestamp 1728305162
transform -1 0 6630 0 1 4090
box -12 -8 112 252
use AOI21X1  _1977_
timestamp 1728304211
transform 1 0 6990 0 -1 4090
box -12 -8 112 252
use OAI21X1  _1978_
timestamp 1728305162
transform 1 0 7090 0 -1 4090
box -12 -8 112 252
use AOI21X1  _1979_
timestamp 1728304211
transform 1 0 6790 0 1 3610
box -12 -8 112 252
use OAI21X1  _1980_
timestamp 1728305162
transform -1 0 6990 0 1 3610
box -12 -8 112 252
use NAND3X1  _1981_
timestamp 1728305047
transform 1 0 6870 0 -1 4090
box -12 -8 112 252
use INVX1  _1982_
timestamp 1728304789
transform 1 0 7030 0 1 4090
box -12 -8 72 252
use NAND3X1  _1983_
timestamp 1728305047
transform 1 0 7130 0 1 4090
box -12 -8 112 252
use NAND3X1  _1984_
timestamp 1728305047
transform 1 0 7190 0 1 3610
box -12 -8 112 252
use NAND2X1  _1985_
timestamp 1728304996
transform 1 0 7310 0 1 3610
box -12 -8 92 252
use INVX1  _1986_
timestamp 1728304789
transform 1 0 7310 0 1 3130
box -12 -8 72 252
use NOR2X1  _1987_
timestamp 1728305106
transform 1 0 7350 0 -1 3130
box -12 -8 92 252
use AOI22X1  _1988_
timestamp 1728304278
transform 1 0 6690 0 1 3130
box -14 -8 132 252
use AOI21X1  _1989_
timestamp 1728304211
transform 1 0 6930 0 1 3130
box -12 -8 112 252
use OAI21X1  _1990_
timestamp 1728305162
transform -1 0 7230 0 1 3130
box -12 -8 112 252
use OAI21X1  _1991_
timestamp 1728305162
transform 1 0 7350 0 1 2650
box -12 -8 112 252
use INVX1  _1992_
timestamp 1728304789
transform 1 0 7270 0 -1 3610
box -12 -8 72 252
use NOR2X1  _1993_
timestamp 1728305106
transform -1 0 7310 0 1 3130
box -12 -8 92 252
use NOR2X1  _1994_
timestamp 1728305106
transform 1 0 7410 0 1 3130
box -12 -8 92 252
use INVX1  _1995_
timestamp 1728304789
transform -1 0 6910 0 1 4090
box -12 -8 72 252
use AOI21X1  _1996_
timestamp 1728304211
transform 1 0 6930 0 1 4090
box -12 -8 112 252
use AND2X2  _1997_
timestamp 1728304163
transform 1 0 4570 0 1 5050
box -12 -8 112 252
use INVX1  _1998_
timestamp 1728304789
transform -1 0 5030 0 1 5050
box -12 -8 72 252
use OAI21X1  _1999_
timestamp 1728305162
transform 1 0 5350 0 -1 5050
box -12 -8 112 252
use INVX1  _2000_
timestamp 1728304789
transform 1 0 7270 0 -1 5050
box -12 -8 72 252
use AOI21X1  _2001_
timestamp 1728304211
transform 1 0 6330 0 1 4570
box -12 -8 112 252
use OAI21X1  _2002_
timestamp 1728305162
transform 1 0 6710 0 1 4570
box -12 -8 112 252
use NAND2X1  _2003_
timestamp 1728304996
transform 1 0 3950 0 -1 5530
box -12 -8 92 252
use INVX1  _2004_
timestamp 1728304789
transform -1 0 4510 0 -1 5530
box -12 -8 72 252
use AND2X2  _2005_
timestamp 1728304163
transform 1 0 4850 0 -1 5530
box -12 -8 112 252
use NAND2X1  _2006_
timestamp 1728304996
transform 1 0 4990 0 -1 5530
box -12 -8 92 252
use NAND2X1  _2007_
timestamp 1728304996
transform -1 0 5250 0 -1 5530
box -12 -8 92 252
use OAI21X1  _2008_
timestamp 1728305162
transform 1 0 5070 0 1 5530
box -12 -8 112 252
use NAND3X1  _2009_
timestamp 1728305047
transform 1 0 5070 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2010_
timestamp 1728305162
transform 1 0 4750 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2011_
timestamp 1728305162
transform 1 0 4530 0 -1 5530
box -12 -8 112 252
use NAND3X1  _2012_
timestamp 1728305047
transform 1 0 4630 0 -1 5530
box -12 -8 112 252
use NAND2X1  _2013_
timestamp 1728304996
transform -1 0 6250 0 -1 5530
box -12 -8 92 252
use NAND2X1  _2014_
timestamp 1728304996
transform -1 0 5530 0 -1 5050
box -12 -8 92 252
use AND2X2  _2015_
timestamp 1728304163
transform 1 0 5550 0 -1 5050
box -12 -8 112 252
use OAI21X1  _2016_
timestamp 1728305162
transform 1 0 5910 0 -1 5050
box -12 -8 112 252
use NAND2X1  _2017_
timestamp 1728304996
transform -1 0 5810 0 1 5530
box -12 -8 92 252
use AND2X2  _2018_
timestamp 1728304163
transform 1 0 5430 0 1 5050
box -12 -8 112 252
use OAI21X1  _2019_
timestamp 1728305162
transform 1 0 5550 0 1 5050
box -12 -8 112 252
use OAI21X1  _2020_
timestamp 1728305162
transform 1 0 5650 0 1 5050
box -12 -8 112 252
use AOI21X1  _2021_
timestamp 1728304211
transform 1 0 5910 0 1 5050
box -12 -8 112 252
use INVX1  _2022_
timestamp 1728304789
transform 1 0 5910 0 1 5530
box -12 -8 72 252
use NAND2X1  _2023_
timestamp 1728304996
transform -1 0 5830 0 -1 5530
box -12 -8 92 252
use NAND2X1  _2024_
timestamp 1728304996
transform -1 0 5470 0 -1 5530
box -12 -8 92 252
use OAI21X1  _2025_
timestamp 1728305162
transform 1 0 5510 0 -1 5530
box -12 -8 112 252
use AOI21X1  _2026_
timestamp 1728304211
transform 1 0 6030 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2027_
timestamp 1728305162
transform -1 0 6110 0 1 5050
box -12 -8 112 252
use AOI22X1  _2028_
timestamp 1728304278
transform 1 0 6130 0 -1 5050
box -14 -8 132 252
use NAND3X1  _2029_
timestamp 1728305047
transform 1 0 5930 0 -1 5530
box -12 -8 112 252
use NAND3X1  _2030_
timestamp 1728305047
transform 1 0 5770 0 1 5050
box -12 -8 112 252
use NAND3X1  _2031_
timestamp 1728305047
transform 1 0 6210 0 1 5050
box -12 -8 112 252
use AOI21X1  _2032_
timestamp 1728304211
transform 1 0 6730 0 -1 5050
box -12 -8 112 252
use AND2X2  _2033_
timestamp 1728304163
transform 1 0 6250 0 -1 5530
box -12 -8 112 252
use NAND3X1  _2034_
timestamp 1728305047
transform 1 0 6450 0 1 5050
box -12 -8 112 252
use OAI21X1  _2035_
timestamp 1728305162
transform 1 0 6110 0 1 5050
box -12 -8 112 252
use AOI21X1  _2036_
timestamp 1728304211
transform 1 0 6690 0 1 5050
box -12 -8 112 252
use OAI21X1  _2037_
timestamp 1728305162
transform -1 0 7130 0 -1 5050
box -12 -8 112 252
use INVX1  _2038_
timestamp 1728304789
transform 1 0 6830 0 1 4570
box -12 -8 72 252
use AOI21X1  _2039_
timestamp 1728304211
transform 1 0 6890 0 1 4570
box -12 -8 112 252
use NAND3X1  _2040_
timestamp 1728305047
transform 1 0 6830 0 1 5050
box -12 -8 112 252
use NAND3X1  _2041_
timestamp 1728305047
transform 1 0 6590 0 -1 5050
box -12 -8 112 252
use NAND3X1  _2042_
timestamp 1728305047
transform 1 0 6930 0 -1 5050
box -12 -8 112 252
use AOI21X1  _2043_
timestamp 1728304211
transform 1 0 7170 0 1 4570
box -12 -8 112 252
use NAND3X1  _2044_
timestamp 1728305047
transform 1 0 6830 0 -1 5050
box -12 -8 112 252
use OAI21X1  _2045_
timestamp 1728305162
transform 1 0 7150 0 -1 5050
box -12 -8 112 252
use AOI21X1  _2046_
timestamp 1728304211
transform 1 0 7430 0 -1 5050
box -12 -8 112 252
use OAI21X1  _2047_
timestamp 1728305162
transform 1 0 7470 0 -1 4570
box -12 -8 112 252
use AOI21X1  _2048_
timestamp 1728304211
transform 1 0 7110 0 -1 4570
box -12 -8 112 252
use OAI21X1  _2049_
timestamp 1728305162
transform 1 0 7230 0 -1 4570
box -12 -8 112 252
use NAND3X1  _2050_
timestamp 1728305047
transform -1 0 7430 0 -1 5050
box -12 -8 112 252
use NAND3X1  _2051_
timestamp 1728305047
transform -1 0 7130 0 1 4570
box -12 -8 112 252
use NAND3X1  _2052_
timestamp 1728305047
transform 1 0 7330 0 -1 4570
box -12 -8 112 252
use NAND2X1  _2053_
timestamp 1728304996
transform 1 0 7410 0 1 3610
box -12 -8 92 252
use NAND2X1  _2054_
timestamp 1728304996
transform -1 0 7610 0 -1 3130
box -12 -8 92 252
use INVX1  _2055_
timestamp 1728304789
transform 1 0 7650 0 -1 3130
box -12 -8 72 252
use OAI21X1  _2056_
timestamp 1728305162
transform 1 0 7430 0 -1 3130
box -12 -8 112 252
use NAND2X1  _2057_
timestamp 1728304996
transform 1 0 7550 0 1 2650
box -12 -8 92 252
use NAND2X1  _2058_
timestamp 1728304996
transform -1 0 7030 0 1 1690
box -12 -8 92 252
use OAI21X1  _2059_
timestamp 1728305162
transform -1 0 7490 0 -1 2170
box -12 -8 112 252
use INVX1  _2060_
timestamp 1728304789
transform 1 0 7510 0 -1 2170
box -12 -8 72 252
use INVX1  _2061_
timestamp 1728304789
transform -1 0 7390 0 -1 3610
box -12 -8 72 252
use OAI21X1  _2062_
timestamp 1728305162
transform 1 0 7430 0 -1 3610
box -12 -8 112 252
use NAND3X1  _2063_
timestamp 1728305047
transform 1 0 7490 0 1 3130
box -12 -8 112 252
use NAND2X1  _2064_
timestamp 1728304996
transform -1 0 7630 0 -1 3610
box -12 -8 92 252
use AND2X2  _2065_
timestamp 1728304163
transform 1 0 7710 0 -1 5050
box -12 -8 112 252
use OAI21X1  _2066_
timestamp 1728305162
transform -1 0 5390 0 -1 5530
box -12 -8 112 252
use INVX1  _2067_
timestamp 1728304789
transform 1 0 7830 0 1 5530
box -12 -8 72 252
use AOI21X1  _2068_
timestamp 1728304211
transform 1 0 6330 0 1 5050
box -12 -8 112 252
use OAI21X1  _2069_
timestamp 1728305162
transform 1 0 6550 0 1 5050
box -12 -8 112 252
use OAI22X1  _2070_
timestamp 1728305200
transform 1 0 5390 0 1 5530
box -12 -8 132 252
use NOR2X1  _2071_
timestamp 1728305106
transform -1 0 5350 0 1 5530
box -12 -8 92 252
use INVX1  _2072_
timestamp 1728304789
transform -1 0 6050 0 1 5530
box -12 -8 72 252
use OAI21X1  _2073_
timestamp 1728305162
transform -1 0 5910 0 1 5530
box -12 -8 112 252
use NOR2X1  _2074_
timestamp 1728305106
transform -1 0 5730 0 -1 5530
box -12 -8 92 252
use OAI21X1  _2075_
timestamp 1728305162
transform 1 0 5830 0 -1 5530
box -12 -8 112 252
use NOR2X1  _2076_
timestamp 1728305106
transform -1 0 5730 0 1 6010
box -12 -8 92 252
use INVX1  _2077_
timestamp 1728304789
transform 1 0 5950 0 1 6010
box -12 -8 72 252
use NAND2X1  _2078_
timestamp 1728304996
transform -1 0 5690 0 1 5530
box -12 -8 92 252
use NAND2X1  _2079_
timestamp 1728304996
transform -1 0 5330 0 1 5050
box -12 -8 92 252
use OAI21X1  _2080_
timestamp 1728305162
transform -1 0 5430 0 1 5050
box -12 -8 112 252
use OAI21X1  _2081_
timestamp 1728305162
transform 1 0 5590 0 -1 6010
box -12 -8 112 252
use NOR2X1  _2082_
timestamp 1728305106
transform -1 0 5910 0 1 6010
box -12 -8 92 252
use INVX1  _2083_
timestamp 1728304789
transform -1 0 5650 0 1 6010
box -12 -8 72 252
use NAND2X1  _2084_
timestamp 1728304996
transform -1 0 6230 0 1 6010
box -12 -8 92 252
use AOI21X1  _2085_
timestamp 1728304211
transform 1 0 6270 0 1 6010
box -12 -8 112 252
use OAI21X1  _2086_
timestamp 1728305162
transform 1 0 6610 0 1 6010
box -12 -8 112 252
use AND2X2  _2087_
timestamp 1728304163
transform 1 0 6170 0 1 5530
box -12 -8 112 252
use AOI21X1  _2088_
timestamp 1728304211
transform 1 0 6050 0 1 5530
box -12 -8 112 252
use NAND3X1  _2089_
timestamp 1728305047
transform 1 0 6410 0 1 6010
box -12 -8 112 252
use OAI21X1  _2090_
timestamp 1728305162
transform 1 0 5730 0 1 6010
box -12 -8 112 252
use NAND3X1  _2091_
timestamp 1728305047
transform 1 0 6730 0 1 6010
box -12 -8 112 252
use AOI21X1  _2092_
timestamp 1728304211
transform 1 0 7330 0 1 6010
box -12 -8 112 252
use INVX1  _2093_
timestamp 1728304789
transform 1 0 7450 0 1 6010
box -12 -8 72 252
use NAND3X1  _2094_
timestamp 1728305047
transform 1 0 6850 0 1 6010
box -12 -8 112 252
use OAI21X1  _2095_
timestamp 1728305162
transform -1 0 6610 0 1 6010
box -12 -8 112 252
use AOI21X1  _2096_
timestamp 1728304211
transform 1 0 7810 0 1 6010
box -12 -8 112 252
use OAI21X1  _2097_
timestamp 1728305162
transform 1 0 7690 0 -1 6010
box -12 -8 112 252
use INVX1  _2098_
timestamp 1728304789
transform -1 0 7550 0 -1 6010
box -12 -8 72 252
use NAND3X1  _2099_
timestamp 1728305047
transform 1 0 7670 0 1 6010
box -12 -8 112 252
use NAND3X1  _2100_
timestamp 1728305047
transform 1 0 7230 0 1 6010
box -12 -8 112 252
use NAND3X1  _2101_
timestamp 1728305047
transform 1 0 7370 0 -1 6010
box -12 -8 112 252
use AOI21X1  _2102_
timestamp 1728304211
transform 1 0 7810 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2103_
timestamp 1728305047
transform 1 0 7270 0 1 5530
box -12 -8 112 252
use OAI21X1  _2104_
timestamp 1728305162
transform -1 0 7690 0 -1 6010
box -12 -8 112 252
use AOI21X1  _2105_
timestamp 1728304211
transform 1 0 7810 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2106_
timestamp 1728305162
transform -1 0 7890 0 1 5050
box -12 -8 112 252
use NAND2X1  _2107_
timestamp 1728304996
transform -1 0 7610 0 -1 5050
box -12 -8 92 252
use NAND3X1  _2108_
timestamp 1728305047
transform -1 0 7810 0 -1 5530
box -12 -8 112 252
use INVX1  _2109_
timestamp 1728304789
transform -1 0 7770 0 1 5530
box -12 -8 72 252
use AOI21X1  _2110_
timestamp 1728304211
transform 1 0 7370 0 1 5530
box -12 -8 112 252
use OAI21X1  _2111_
timestamp 1728305162
transform 1 0 7610 0 1 5530
box -12 -8 112 252
use NAND3X1  _2112_
timestamp 1728305047
transform 1 0 7610 0 -1 5050
box -12 -8 112 252
use NAND2X1  _2113_
timestamp 1728304996
transform 1 0 7810 0 1 4570
box -12 -8 92 252
use INVX1  _2114_
timestamp 1728304789
transform 1 0 7850 0 -1 3610
box -12 -8 72 252
use NOR2X1  _2115_
timestamp 1728305106
transform -1 0 7750 0 -1 3610
box -12 -8 92 252
use INVX1  _2116_
timestamp 1728304789
transform 1 0 7830 0 -1 4570
box -12 -8 72 252
use NOR3X1  _2117_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728303224
transform 1 0 7610 0 1 3130
box -12 -8 192 252
use OAI21X1  _2118_
timestamp 1728305162
transform -1 0 7850 0 -1 3610
box -12 -8 112 252
use NAND2X1  _2119_
timestamp 1728304996
transform 1 0 7830 0 1 3130
box -12 -8 92 252
use OAI22X1  _2120_
timestamp 1728305200
transform 1 0 7630 0 1 2650
box -12 -8 132 252
use INVX1  _2121_
timestamp 1728304789
transform 1 0 7830 0 -1 2650
box -12 -8 72 252
use NAND2X1  _2122_
timestamp 1728304996
transform 1 0 6270 0 1 5530
box -12 -8 92 252
use AOI21X1  _2123_
timestamp 1728304211
transform 1 0 6990 0 1 6010
box -12 -8 112 252
use OAI21X1  _2124_
timestamp 1728305162
transform -1 0 7190 0 1 6010
box -12 -8 112 252
use AOI22X1  _2125_
timestamp 1728304278
transform -1 0 6150 0 1 6010
box -14 -8 132 252
use INVX1  _2126_
timestamp 1728304789
transform -1 0 5950 0 -1 6010
box -12 -8 72 252
use NAND2X1  _2127_
timestamp 1728304996
transform -1 0 5270 0 1 5530
box -12 -8 92 252
use NAND2X1  _2128_
timestamp 1728304996
transform -1 0 5130 0 1 5050
box -12 -8 92 252
use NAND2X1  _2129_
timestamp 1728304996
transform -1 0 4570 0 1 5050
box -12 -8 92 252
use OAI21X1  _2130_
timestamp 1728305162
transform 1 0 4830 0 1 5050
box -12 -8 112 252
use OAI21X1  _2131_
timestamp 1728305162
transform -1 0 5230 0 1 5050
box -12 -8 112 252
use OR2X2  _2132_
timestamp 1728305284
transform 1 0 5450 0 -1 6010
box -12 -8 112 252
use OAI21X1  _2133_
timestamp 1728305162
transform -1 0 5610 0 1 5530
box -12 -8 112 252
use NAND3X1  _2134_
timestamp 1728305047
transform 1 0 5990 0 -1 6010
box -12 -8 112 252
use NOR2X1  _2135_
timestamp 1728305106
transform -1 0 5210 0 -1 6010
box -12 -8 92 252
use AND2X2  _2136_
timestamp 1728304163
transform -1 0 5430 0 -1 6010
box -12 -8 112 252
use OAI21X1  _2137_
timestamp 1728305162
transform 1 0 5790 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2138_
timestamp 1728305047
transform 1 0 6490 0 -1 6010
box -12 -8 112 252
use OAI21X1  _2139_
timestamp 1728305162
transform 1 0 5690 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2140_
timestamp 1728305047
transform 1 0 6110 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2141_
timestamp 1728305047
transform 1 0 6210 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2142_
timestamp 1728305047
transform -1 0 7030 0 -1 6010
box -12 -8 112 252
use INVX1  _2143_
timestamp 1728304789
transform 1 0 7610 0 1 6010
box -12 -8 72 252
use AOI21X1  _2144_
timestamp 1728304211
transform -1 0 7610 0 1 6010
box -12 -8 112 252
use AOI21X1  _2145_
timestamp 1728304211
transform 1 0 6350 0 -1 6010
box -12 -8 112 252
use AOI21X1  _2146_
timestamp 1728304211
transform 1 0 6590 0 -1 6010
box -12 -8 112 252
use OAI21X1  _2147_
timestamp 1728305162
transform 1 0 7150 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2148_
timestamp 1728305047
transform 1 0 6970 0 1 5530
box -12 -8 112 252
use INVX1  _2149_
timestamp 1728304789
transform 1 0 6910 0 1 5530
box -12 -8 72 252
use OAI21X1  _2150_
timestamp 1728305162
transform -1 0 7130 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2151_
timestamp 1728305047
transform 1 0 7270 0 -1 6010
box -12 -8 112 252
use NAND3X1  _2152_
timestamp 1728305047
transform 1 0 7170 0 1 5530
box -12 -8 112 252
use AOI22X1  _2153_
timestamp 1728304278
transform -1 0 7410 0 -1 5530
box -14 -8 132 252
use OAI21X1  _2154_
timestamp 1728305162
transform -1 0 7570 0 1 5530
box -12 -8 112 252
use NAND3X1  _2155_
timestamp 1728305047
transform 1 0 7150 0 -1 5530
box -12 -8 112 252
use NAND3X1  _2156_
timestamp 1728305047
transform 1 0 7070 0 1 5530
box -12 -8 112 252
use AOI21X1  _2157_
timestamp 1728304211
transform 1 0 7370 0 1 5050
box -12 -8 112 252
use NOR2X1  _2158_
timestamp 1728305106
transform 1 0 7570 0 1 5050
box -12 -8 92 252
use AOI21X1  _2159_
timestamp 1728304211
transform 1 0 7590 0 1 4570
box -12 -8 112 252
use NAND2X1  _2160_
timestamp 1728304996
transform -1 0 7590 0 1 4570
box -12 -8 92 252
use NAND3X1  _2161_
timestamp 1728305047
transform 1 0 7470 0 1 5050
box -12 -8 112 252
use INVX1  _2162_
timestamp 1728304789
transform 1 0 7610 0 -1 5530
box -12 -8 72 252
use NAND3X1  _2163_
timestamp 1728305047
transform 1 0 7490 0 -1 5530
box -12 -8 112 252
use NAND2X1  _2164_
timestamp 1728304996
transform -1 0 7770 0 1 5050
box -12 -8 92 252
use NOR2X1  _2165_
timestamp 1728305106
transform -1 0 7830 0 -1 4570
box -12 -8 92 252
use OAI21X1  _2166_
timestamp 1728305162
transform 1 0 7770 0 1 250
box -12 -8 112 252
use OAI21X1  _2167_
timestamp 1728305162
transform -1 0 7910 0 -1 2170
box -12 -8 112 252
use INVX1  _2168_
timestamp 1728304789
transform -1 0 7910 0 1 1210
box -12 -8 72 252
use NAND3X1  _2169_
timestamp 1728305047
transform 1 0 7690 0 1 4570
box -12 -8 112 252
use AOI21X1  _2170_
timestamp 1728304211
transform 1 0 7610 0 1 3610
box -12 -8 112 252
use OAI21X1  _2171_
timestamp 1728305162
transform 1 0 7810 0 -1 5050
box -12 -8 112 252
use NOR2X1  _2172_
timestamp 1728305106
transform -1 0 7870 0 -1 4090
box -12 -8 92 252
use NOR2X1  _2173_
timestamp 1728305106
transform -1 0 5130 0 -1 6010
box -12 -8 92 252
use NAND2X1  _2174_
timestamp 1728304996
transform -1 0 4230 0 1 5530
box -12 -8 92 252
use NAND2X1  _2175_
timestamp 1728304996
transform -1 0 4430 0 -1 5530
box -12 -8 92 252
use OAI21X1  _2176_
timestamp 1728305162
transform 1 0 4390 0 1 5530
box -12 -8 112 252
use OAI21X1  _2177_
timestamp 1728305162
transform 1 0 4390 0 -1 6010
box -12 -8 112 252
use OAI21X1  _2178_
timestamp 1728305162
transform -1 0 4590 0 -1 6010
box -12 -8 112 252
use NOR2X1  _2179_
timestamp 1728305106
transform -1 0 4290 0 -1 6010
box -12 -8 92 252
use NOR2X1  _2180_
timestamp 1728305106
transform -1 0 4370 0 -1 6010
box -12 -8 92 252
use INVX1  _2181_
timestamp 1728304789
transform 1 0 4670 0 1 6010
box -12 -8 72 252
use NAND3X1  _2182_
timestamp 1728305047
transform 1 0 4730 0 1 6010
box -12 -8 112 252
use AND2X2  _2183_
timestamp 1728304163
transform 1 0 5170 0 1 6010
box -12 -8 112 252
use OAI21X1  _2184_
timestamp 1728305162
transform -1 0 5310 0 -1 6010
box -12 -8 112 252
use NOR2X1  _2185_
timestamp 1728305106
transform 1 0 5370 0 1 6010
box -12 -8 92 252
use NAND2X1  _2186_
timestamp 1728304996
transform 1 0 5270 0 1 6010
box -12 -8 92 252
use NAND2X1  _2187_
timestamp 1728304996
transform 1 0 5490 0 1 6010
box -12 -8 92 252
use NAND2X1  _2188_
timestamp 1728304996
transform 1 0 6690 0 -1 6010
box -12 -8 92 252
use NAND3X1  _2189_
timestamp 1728305047
transform 1 0 6790 0 -1 6010
box -12 -8 112 252
use NAND2X1  _2190_
timestamp 1728304996
transform 1 0 6490 0 1 5530
box -12 -8 92 252
use NAND3X1  _2191_
timestamp 1728305047
transform 1 0 6390 0 1 5530
box -12 -8 112 252
use NAND2X1  _2192_
timestamp 1728304996
transform -1 0 7010 0 1 5050
box -12 -8 92 252
use NAND3X1  _2193_
timestamp 1728305047
transform 1 0 7230 0 1 5050
box -12 -8 112 252
use NAND2X1  _2194_
timestamp 1728304996
transform 1 0 7150 0 1 5050
box -12 -8 92 252
use NAND3X1  _2195_
timestamp 1728305047
transform 1 0 7010 0 1 5050
box -12 -8 112 252
use NAND2X1  _2196_
timestamp 1728304996
transform 1 0 7390 0 1 4570
box -12 -8 92 252
use AND2X2  _2197_
timestamp 1728304163
transform 1 0 7710 0 -1 2650
box -12 -8 112 252
use OAI21X1  _2198_
timestamp 1728305162
transform -1 0 7850 0 -1 3130
box -12 -8 112 252
use OAI22X1  _2199_
timestamp 1728305200
transform -1 0 7870 0 1 2650
box -12 -8 132 252
use NAND2X1  _2200_
timestamp 1728304996
transform -1 0 7570 0 1 2170
box -12 -8 92 252
use INVX1  _2201_
timestamp 1728304789
transform 1 0 7630 0 1 4090
box -12 -8 72 252
use OAI21X1  _2202_
timestamp 1728305162
transform -1 0 7830 0 1 4090
box -12 -8 112 252
use AOI21X1  _2203_
timestamp 1728304211
transform 1 0 4550 0 1 6010
box -12 -8 112 252
use NOR2X1  _2204_
timestamp 1728305106
transform -1 0 4690 0 1 5530
box -12 -8 92 252
use INVX1  _2205_
timestamp 1728304789
transform -1 0 4750 0 1 5530
box -12 -8 72 252
use OAI21X1  _2206_
timestamp 1728305162
transform -1 0 4370 0 1 5530
box -12 -8 112 252
use OAI21X1  _2207_
timestamp 1728305162
transform -1 0 4590 0 1 5530
box -12 -8 112 252
use OR2X2  _2208_
timestamp 1728305284
transform -1 0 4950 0 1 6010
box -12 -8 112 252
use NAND2X1  _2209_
timestamp 1728304996
transform 1 0 4950 0 1 6010
box -12 -8 92 252
use NAND2X1  _2210_
timestamp 1728304996
transform 1 0 5050 0 1 6010
box -12 -8 92 252
use AND2X2  _2211_
timestamp 1728304163
transform 1 0 6670 0 1 5530
box -12 -8 112 252
use NOR2X1  _2212_
timestamp 1728305106
transform -1 0 6650 0 1 5530
box -12 -8 92 252
use OAI21X1  _2213_
timestamp 1728305162
transform 1 0 6770 0 -1 5530
box -12 -8 112 252
use INVX1  _2214_
timestamp 1728304789
transform -1 0 7010 0 -1 5530
box -12 -8 72 252
use NOR2X1  _2215_
timestamp 1728305106
transform 1 0 6790 0 1 5530
box -12 -8 92 252
use NAND2X1  _2216_
timestamp 1728304996
transform 1 0 6870 0 -1 5530
box -12 -8 92 252
use NAND2X1  _2217_
timestamp 1728304996
transform 1 0 7050 0 -1 5530
box -12 -8 92 252
use NAND3X1  _2218_
timestamp 1728305047
transform 1 0 7650 0 -1 4570
box -12 -8 112 252
use INVX1  _2219_
timestamp 1728304789
transform -1 0 7650 0 -1 4570
box -12 -8 72 252
use NOR2X1  _2220_
timestamp 1728305106
transform 1 0 7830 0 1 4090
box -12 -8 92 252
use OAI21X1  _2221_
timestamp 1728305162
transform -1 0 7850 0 1 3610
box -12 -8 112 252
use INVX1  _2222_
timestamp 1728304789
transform 1 0 7770 0 1 5530
box -12 -8 72 252
use AOI21X1  _2223_
timestamp 1728304211
transform -1 0 7750 0 -1 4090
box -12 -8 112 252
use INVX1  _2224_
timestamp 1728304789
transform 1 0 7230 0 1 4090
box -12 -8 72 252
use OAI21X1  _2225_
timestamp 1728305162
transform 1 0 7530 0 1 4090
box -12 -8 112 252
use NAND3X1  _2226_
timestamp 1728305047
transform -1 0 7590 0 1 3610
box -12 -8 112 252
use NAND2X1  _2227_
timestamp 1728304996
transform 1 0 7570 0 1 2170
box -12 -8 92 252
use NAND2X1  _2228_
timestamp 1728304996
transform -1 0 7070 0 1 730
box -12 -8 92 252
use OAI21X1  _2229_
timestamp 1728305162
transform -1 0 7370 0 1 4570
box -12 -8 112 252
use NOR2X1  _2230_
timestamp 1728305106
transform -1 0 7490 0 1 4090
box -12 -8 92 252
use AOI21X1  _2231_
timestamp 1728304211
transform -1 0 7390 0 1 4090
box -12 -8 112 252
use NAND3X1  _2232_
timestamp 1728305047
transform -1 0 7630 0 -1 4090
box -12 -8 112 252
use OAI21X1  _2233_
timestamp 1728305162
transform 1 0 4750 0 1 5530
box -12 -8 112 252
use OAI21X1  _2234_
timestamp 1728305162
transform 1 0 4610 0 -1 6010
box -12 -8 112 252
use OR2X2  _2235_
timestamp 1728305284
transform -1 0 4810 0 -1 6010
box -12 -8 112 252
use AND2X2  _2236_
timestamp 1728304163
transform 1 0 4850 0 -1 6010
box -12 -8 112 252
use OR2X2  _2237_
timestamp 1728305284
transform 1 0 6550 0 -1 5530
box -12 -8 112 252
use NAND2X1  _2238_
timestamp 1728304996
transform -1 0 6550 0 -1 5530
box -12 -8 92 252
use NAND2X1  _2239_
timestamp 1728304996
transform 1 0 6650 0 -1 5530
box -12 -8 92 252
use NAND3X1  _2240_
timestamp 1728305047
transform 1 0 7310 0 -1 4090
box -12 -8 112 252
use NAND2X1  _2241_
timestamp 1728304996
transform 1 0 7410 0 -1 4090
box -12 -8 92 252
use INVX1  _2242_
timestamp 1728304789
transform 1 0 7210 0 -1 4090
box -12 -8 72 252
use NAND2X1  _2243_
timestamp 1728304996
transform 1 0 7410 0 -1 5530
box -12 -8 92 252
use NAND3X1  _2244_
timestamp 1728305047
transform 1 0 7370 0 -1 2650
box -12 -8 112 252
use NAND2X1  _2245_
timestamp 1728304996
transform 1 0 7330 0 1 730
box -12 -8 92 252
use INVX1  _2246_
timestamp 1728304789
transform 1 0 7210 0 1 2170
box -12 -8 72 252
use INVX1  _2247_
timestamp 1728304789
transform 1 0 4990 0 -1 6010
box -12 -8 72 252
use OAI21X1  _2248_
timestamp 1728305162
transform 1 0 4850 0 1 5530
box -12 -8 112 252
use NOR2X1  _2249_
timestamp 1728305106
transform 1 0 4970 0 1 5530
box -12 -8 92 252
use AND2X2  _2250_
timestamp 1728304163
transform -1 0 6450 0 -1 5530
box -12 -8 112 252
use AOI22X1  _2251_
timestamp 1728304278
transform -1 0 7270 0 -1 2650
box -14 -8 132 252
use INVX1  _2252_
timestamp 1728304789
transform 1 0 4870 0 1 2650
box -12 -8 72 252
use NOR2X1  _2253_
timestamp 1728305106
transform 1 0 5070 0 1 2650
box -12 -8 92 252
use INVX1  _2254_
timestamp 1728304789
transform 1 0 5150 0 1 2650
box -12 -8 72 252
use NAND2X1  _2255_
timestamp 1728304996
transform -1 0 5050 0 1 2650
box -12 -8 92 252
use NAND2X1  _2256_
timestamp 1728304996
transform -1 0 5010 0 -1 2650
box -12 -8 92 252
use NAND2X1  _2257_
timestamp 1728304996
transform 1 0 4970 0 1 1690
box -12 -8 92 252
use OAI21X1  _2258_
timestamp 1728305162
transform -1 0 5010 0 1 2170
box -12 -8 112 252
use INVX1  _2259_
timestamp 1728304789
transform 1 0 4470 0 -1 2650
box -12 -8 72 252
use NOR2X1  _2260_
timestamp 1728305106
transform -1 0 4690 0 -1 2650
box -12 -8 92 252
use NOR2X1  _2261_
timestamp 1728305106
transform -1 0 4430 0 -1 2650
box -12 -8 92 252
use NOR2X1  _2262_
timestamp 1728305106
transform 1 0 4730 0 -1 2650
box -12 -8 92 252
use NAND2X1  _2263_
timestamp 1728304996
transform 1 0 5210 0 1 2650
box -12 -8 92 252
use OAI21X1  _2264_
timestamp 1728305162
transform 1 0 4830 0 -1 2650
box -12 -8 112 252
use NAND2X1  _2265_
timestamp 1728304996
transform 1 0 5230 0 1 2170
box -12 -8 92 252
use NAND2X1  _2266_
timestamp 1728304996
transform 1 0 5050 0 1 2170
box -12 -8 92 252
use OAI21X1  _2267_
timestamp 1728305162
transform -1 0 5230 0 1 2170
box -12 -8 112 252
use OAI21X1  _2268_
timestamp 1728305162
transform 1 0 5030 0 -1 2650
box -12 -8 112 252
use INVX1  _2269_
timestamp 1728304789
transform 1 0 6070 0 1 2650
box -12 -8 72 252
use NOR2X1  _2270_
timestamp 1728305106
transform 1 0 6170 0 1 2650
box -12 -8 92 252
use NOR2X1  _2271_
timestamp 1728305106
transform -1 0 6010 0 1 2650
box -12 -8 92 252
use NOR2X1  _2272_
timestamp 1728305106
transform -1 0 6010 0 -1 2650
box -12 -8 92 252
use NAND2X1  _2273_
timestamp 1728304996
transform -1 0 6090 0 -1 2650
box -12 -8 92 252
use OR2X2  _2274_
timestamp 1728305284
transform 1 0 6130 0 -1 2650
box -12 -8 112 252
use NAND2X1  _2275_
timestamp 1728304996
transform 1 0 6090 0 1 2170
box -12 -8 92 252
use NAND2X1  _2276_
timestamp 1728304996
transform 1 0 6310 0 1 2170
box -12 -8 92 252
use OAI21X1  _2277_
timestamp 1728305162
transform 1 0 6210 0 1 2170
box -12 -8 112 252
use AOI21X1  _2278_
timestamp 1728304211
transform -1 0 5910 0 -1 2650
box -12 -8 112 252
use INVX1  _2279_
timestamp 1728304789
transform -1 0 5370 0 -1 2650
box -12 -8 72 252
use INVX1  _2280_
timestamp 1728304789
transform 1 0 5290 0 1 2650
box -12 -8 72 252
use NOR2X1  _2281_
timestamp 1728305106
transform 1 0 5470 0 1 2650
box -12 -8 92 252
use NOR2X1  _2282_
timestamp 1728305106
transform 1 0 5350 0 1 2650
box -12 -8 92 252
use NOR2X1  _2283_
timestamp 1728305106
transform 1 0 5530 0 -1 2650
box -12 -8 92 252
use NAND2X1  _2284_
timestamp 1728304996
transform 1 0 5210 0 -1 2650
box -12 -8 92 252
use OAI21X1  _2285_
timestamp 1728305162
transform -1 0 5510 0 -1 2650
box -12 -8 112 252
use NAND2X1  _2286_
timestamp 1728304996
transform -1 0 5210 0 -1 2650
box -12 -8 92 252
use NAND2X1  _2287_
timestamp 1728304996
transform 1 0 5250 0 -1 2170
box -12 -8 92 252
use OAI21X1  _2288_
timestamp 1728305162
transform 1 0 5130 0 -1 2170
box -12 -8 112 252
use NAND2X1  _2289_
timestamp 1728304996
transform -1 0 6510 0 1 2170
box -12 -8 92 252
use INVX1  _2290_
timestamp 1728304789
transform 1 0 6730 0 -1 2650
box -12 -8 72 252
use NOR2X1  _2291_
timestamp 1728305106
transform -1 0 6730 0 -1 2650
box -12 -8 92 252
use NOR2X1  _2292_
timestamp 1728305106
transform 1 0 6790 0 -1 2650
box -12 -8 92 252
use INVX1  _2293_
timestamp 1728304789
transform 1 0 5750 0 -1 2650
box -12 -8 72 252
use OAI21X1  _2294_
timestamp 1728305162
transform 1 0 5630 0 -1 2650
box -12 -8 112 252
use INVX1  _2295_
timestamp 1728304789
transform 1 0 7270 0 1 2170
box -12 -8 72 252
use OAI21X1  _2296_
timestamp 1728305162
transform 1 0 7110 0 1 2170
box -12 -8 112 252
use NOR2X1  _2297_
timestamp 1728305106
transform -1 0 6810 0 -1 2170
box -12 -8 92 252
use NAND2X1  _2298_
timestamp 1728304996
transform 1 0 6910 0 1 2170
box -12 -8 92 252
use NAND2X1  _2299_
timestamp 1728304996
transform 1 0 6990 0 1 2170
box -12 -8 92 252
use OAI21X1  _2300_
timestamp 1728305162
transform -1 0 6890 0 1 2170
box -12 -8 112 252
use INVX1  _2301_
timestamp 1728304789
transform 1 0 5850 0 -1 2170
box -12 -8 72 252
use AOI21X1  _2302_
timestamp 1728304211
transform -1 0 6670 0 -1 2170
box -12 -8 112 252
use NAND2X1  _2303_
timestamp 1728304996
transform 1 0 6690 0 -1 1690
box -12 -8 92 252
use INVX1  _2304_
timestamp 1728304789
transform -1 0 6610 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2305_
timestamp 1728305106
transform 1 0 6610 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2306_
timestamp 1728305106
transform -1 0 6510 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2307_
timestamp 1728305106
transform 1 0 6370 0 -1 2170
box -12 -8 92 252
use AND2X2  _2308_
timestamp 1728304163
transform -1 0 6370 0 -1 2170
box -12 -8 112 252
use OAI21X1  _2309_
timestamp 1728305162
transform -1 0 6230 0 -1 2170
box -12 -8 112 252
use OAI21X1  _2310_
timestamp 1728305162
transform 1 0 5910 0 -1 2170
box -12 -8 112 252
use NAND2X1  _2311_
timestamp 1728304996
transform 1 0 4990 0 -1 1690
box -12 -8 92 252
use INVX1  _2312_
timestamp 1728304789
transform -1 0 6730 0 -1 2170
box -12 -8 72 252
use OAI21X1  _2313_
timestamp 1728305162
transform 1 0 6610 0 1 1690
box -12 -8 112 252
use AND2X2  _2314_
timestamp 1728304163
transform -1 0 6550 0 -1 2170
box -12 -8 112 252
use AOI21X1  _2315_
timestamp 1728304211
transform -1 0 6490 0 1 1690
box -12 -8 112 252
use NAND2X1  _2316_
timestamp 1728304996
transform 1 0 6010 0 1 1690
box -12 -8 92 252
use INVX1  _2317_
timestamp 1728304789
transform -1 0 5830 0 1 1690
box -12 -8 72 252
use NOR2X1  _2318_
timestamp 1728305106
transform 1 0 5930 0 1 1690
box -12 -8 92 252
use OR2X2  _2319_
timestamp 1728305284
transform -1 0 5750 0 1 1690
box -12 -8 112 252
use AND2X2  _2320_
timestamp 1728304163
transform -1 0 5610 0 1 1690
box -12 -8 112 252
use OAI21X1  _2321_
timestamp 1728305162
transform -1 0 5510 0 1 1690
box -12 -8 112 252
use OAI21X1  _2322_
timestamp 1728305162
transform -1 0 5390 0 1 1690
box -12 -8 112 252
use INVX1  _2323_
timestamp 1728304789
transform 1 0 5370 0 -1 1210
box -12 -8 72 252
use OAI21X1  _2324_
timestamp 1728305162
transform 1 0 5830 0 1 1690
box -12 -8 112 252
use NAND2X1  _2325_
timestamp 1728304996
transform 1 0 6210 0 -1 1690
box -12 -8 92 252
use INVX1  _2326_
timestamp 1728304789
transform -1 0 6090 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2327_
timestamp 1728305106
transform 1 0 6110 0 -1 1690
box -12 -8 92 252
use OAI21X1  _2328_
timestamp 1728305162
transform -1 0 5910 0 -1 1690
box -12 -8 112 252
use INVX1  _2329_
timestamp 1728304789
transform -1 0 5790 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2330_
timestamp 1728305106
transform 1 0 5950 0 -1 1690
box -12 -8 92 252
use AOI21X1  _2331_
timestamp 1728304211
transform -1 0 5730 0 -1 1690
box -12 -8 112 252
use AOI22X1  _2332_
timestamp 1728304278
transform 1 0 5550 0 1 1210
box -14 -8 132 252
use NAND2X1  _2333_
timestamp 1728304996
transform 1 0 7350 0 -1 1210
box -12 -8 92 252
use INVX1  _2334_
timestamp 1728304789
transform -1 0 7130 0 1 1690
box -12 -8 72 252
use NOR2X1  _2335_
timestamp 1728305106
transform 1 0 7230 0 1 1690
box -12 -8 92 252
use NOR2X1  _2336_
timestamp 1728305106
transform 1 0 7150 0 1 1690
box -12 -8 92 252
use NOR2X1  _2337_
timestamp 1728305106
transform -1 0 7390 0 1 1690
box -12 -8 92 252
use INVX1  _2338_
timestamp 1728304789
transform 1 0 7530 0 1 1210
box -12 -8 72 252
use OAI21X1  _2339_
timestamp 1728305162
transform 1 0 6090 0 1 1690
box -12 -8 112 252
use INVX1  _2340_
timestamp 1728304789
transform 1 0 6210 0 1 1690
box -12 -8 72 252
use NOR2X1  _2341_
timestamp 1728305106
transform 1 0 6270 0 1 1690
box -12 -8 92 252
use AOI21X1  _2342_
timestamp 1728304211
transform 1 0 6750 0 1 1690
box -12 -8 112 252
use NAND3X1  _2343_
timestamp 1728305047
transform 1 0 6490 0 1 1690
box -12 -8 112 252
use AND2X2  _2344_
timestamp 1728304163
transform 1 0 6850 0 1 1690
box -12 -8 112 252
use AND2X2  _2345_
timestamp 1728304163
transform -1 0 7810 0 1 1210
box -12 -8 112 252
use OAI21X1  _2346_
timestamp 1728305162
transform 1 0 7550 0 -1 1210
box -12 -8 112 252
use OAI21X1  _2347_
timestamp 1728305162
transform -1 0 7550 0 -1 1210
box -12 -8 112 252
use INVX1  _2348_
timestamp 1728304789
transform 1 0 7170 0 -1 1690
box -12 -8 72 252
use INVX1  _2349_
timestamp 1728304789
transform 1 0 7530 0 1 1690
box -12 -8 72 252
use OAI21X1  _2350_
timestamp 1728305162
transform 1 0 7390 0 1 1690
box -12 -8 112 252
use INVX1  _2351_
timestamp 1728304789
transform 1 0 7770 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2352_
timestamp 1728305106
transform 1 0 7830 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2353_
timestamp 1728305106
transform 1 0 7830 0 1 1690
box -12 -8 92 252
use NOR2X1  _2354_
timestamp 1728305106
transform 1 0 7670 0 -1 1690
box -12 -8 92 252
use INVX1  _2355_
timestamp 1728304789
transform -1 0 7670 0 -1 1690
box -12 -8 72 252
use OR2X2  _2356_
timestamp 1728305284
transform 1 0 7490 0 -1 1690
box -12 -8 112 252
use AOI21X1  _2357_
timestamp 1728304211
transform -1 0 7490 0 -1 1690
box -12 -8 112 252
use AOI22X1  _2358_
timestamp 1728304278
transform 1 0 7230 0 -1 1690
box -14 -8 132 252
use NAND2X1  _2359_
timestamp 1728304996
transform -1 0 7090 0 -1 730
box -12 -8 92 252
use NOR2X1  _2360_
timestamp 1728305106
transform -1 0 7670 0 1 1210
box -12 -8 92 252
use INVX1  _2361_
timestamp 1728304789
transform 1 0 7850 0 -1 1210
box -12 -8 72 252
use NOR2X1  _2362_
timestamp 1728305106
transform 1 0 7750 0 -1 1210
box -12 -8 92 252
use INVX1  _2363_
timestamp 1728304789
transform 1 0 7730 0 1 1690
box -12 -8 72 252
use OAI21X1  _2364_
timestamp 1728305162
transform 1 0 7630 0 1 1690
box -12 -8 112 252
use NOR2X1  _2365_
timestamp 1728305106
transform 1 0 7650 0 -1 1210
box -12 -8 92 252
use INVX1  _2366_
timestamp 1728304789
transform 1 0 7850 0 -1 730
box -12 -8 72 252
use NOR2X1  _2367_
timestamp 1728305106
transform -1 0 7830 0 -1 730
box -12 -8 92 252
use NOR2X1  _2368_
timestamp 1728305106
transform 1 0 7830 0 1 730
box -12 -8 92 252
use OAI21X1  _2369_
timestamp 1728305162
transform -1 0 7690 0 1 730
box -12 -8 112 252
use NOR2X1  _2370_
timestamp 1728305106
transform 1 0 7710 0 1 730
box -12 -8 92 252
use OAI21X1  _2371_
timestamp 1728305162
transform -1 0 7650 0 -1 730
box -12 -8 112 252
use NAND2X1  _2372_
timestamp 1728304996
transform -1 0 7550 0 -1 730
box -12 -8 92 252
use OAI21X1  _2373_
timestamp 1728305162
transform -1 0 7430 0 -1 730
box -12 -8 112 252
use INVX1  _2374_
timestamp 1728304789
transform 1 0 7390 0 -1 250
box -12 -8 72 252
use OAI21X1  _2375_
timestamp 1728305162
transform -1 0 7750 0 -1 730
box -12 -8 112 252
use AND2X2  _2376_
timestamp 1728304163
transform 1 0 6750 0 1 250
box -12 -8 112 252
use NOR2X1  _2377_
timestamp 1728305106
transform 1 0 6850 0 1 250
box -12 -8 92 252
use NOR2X1  _2378_
timestamp 1728305106
transform 1 0 6930 0 1 250
box -12 -8 92 252
use INVX1  _2379_
timestamp 1728304789
transform 1 0 7830 0 -1 250
box -12 -8 72 252
use OR2X2  _2380_
timestamp 1728305284
transform 1 0 7690 0 -1 250
box -12 -8 112 252
use AOI21X1  _2381_
timestamp 1728304211
transform -1 0 7690 0 -1 250
box -12 -8 112 252
use AOI22X1  _2382_
timestamp 1728304278
transform 1 0 7450 0 -1 250
box -14 -8 132 252
use NAND2X1  _2383_
timestamp 1728304996
transform -1 0 5390 0 1 250
box -12 -8 92 252
use AOI21X1  _2384_
timestamp 1728304211
transform 1 0 7010 0 1 250
box -12 -8 112 252
use AND2X2  _2385_
timestamp 1728304163
transform -1 0 7510 0 1 250
box -12 -8 112 252
use NAND2X1  _2386_
timestamp 1728304996
transform -1 0 7390 0 1 250
box -12 -8 92 252
use NAND2X1  _2387_
timestamp 1728304996
transform 1 0 7230 0 1 250
box -12 -8 92 252
use NAND2X1  _2388_
timestamp 1728304996
transform 1 0 7510 0 1 730
box -12 -8 92 252
use NOR2X1  _2389_
timestamp 1728305106
transform -1 0 7510 0 1 730
box -12 -8 92 252
use NOR2X1  _2390_
timestamp 1728305106
transform -1 0 7190 0 1 250
box -12 -8 92 252
use INVX1  _2391_
timestamp 1728304789
transform -1 0 5690 0 1 250
box -12 -8 72 252
use INVX1  _2392_
timestamp 1728304789
transform 1 0 6070 0 1 250
box -12 -8 72 252
use INVX1  _2393_
timestamp 1728304789
transform -1 0 6310 0 1 250
box -12 -8 72 252
use NOR2X1  _2394_
timestamp 1728305106
transform 1 0 6170 0 1 250
box -12 -8 92 252
use NOR2X1  _2395_
timestamp 1728305106
transform 1 0 6610 0 -1 250
box -12 -8 92 252
use NOR2X1  _2396_
timestamp 1728305106
transform -1 0 6610 0 -1 250
box -12 -8 92 252
use NOR2X1  _2397_
timestamp 1728305106
transform -1 0 5590 0 1 250
box -12 -8 92 252
use INVX1  _2398_
timestamp 1728304789
transform 1 0 5830 0 1 250
box -12 -8 72 252
use OAI21X1  _2399_
timestamp 1728305162
transform -1 0 5790 0 1 250
box -12 -8 112 252
use OAI21X1  _2400_
timestamp 1728305162
transform -1 0 5510 0 1 250
box -12 -8 112 252
use INVX1  _2401_
timestamp 1728304789
transform 1 0 6090 0 -1 250
box -12 -8 72 252
use INVX1  _2402_
timestamp 1728304789
transform 1 0 6830 0 -1 250
box -12 -8 72 252
use OAI21X1  _2403_
timestamp 1728305162
transform 1 0 6690 0 -1 250
box -12 -8 112 252
use AND2X2  _2404_
timestamp 1728304163
transform 1 0 6170 0 1 730
box -12 -8 112 252
use NOR2X1  _2405_
timestamp 1728305106
transform 1 0 6270 0 1 730
box -12 -8 92 252
use NOR2X1  _2406_
timestamp 1728305106
transform 1 0 6450 0 -1 730
box -12 -8 92 252
use INVX1  _2407_
timestamp 1728304789
transform 1 0 6530 0 -1 730
box -12 -8 72 252
use OR2X2  _2408_
timestamp 1728305284
transform -1 0 6510 0 -1 250
box -12 -8 112 252
use AOI21X1  _2409_
timestamp 1728304211
transform -1 0 6390 0 -1 250
box -12 -8 112 252
use AOI22X1  _2410_
timestamp 1728304278
transform 1 0 6170 0 -1 250
box -14 -8 132 252
use NAND2X1  _2411_
timestamp 1728304996
transform -1 0 6450 0 1 730
box -12 -8 92 252
use AOI21X1  _2412_
timestamp 1728304211
transform -1 0 6410 0 -1 730
box -12 -8 112 252
use NOR2X1  _2413_
timestamp 1728305106
transform -1 0 6010 0 1 250
box -12 -8 92 252
use INVX1  _2414_
timestamp 1728304789
transform 1 0 6010 0 1 250
box -12 -8 72 252
use OAI21X1  _2415_
timestamp 1728305162
transform 1 0 6210 0 -1 730
box -12 -8 112 252
use NOR2X1  _2416_
timestamp 1728305106
transform -1 0 6390 0 -1 1210
box -12 -8 92 252
use INVX1  _2417_
timestamp 1728304789
transform 1 0 6410 0 1 1210
box -12 -8 72 252
use INVX1  _2418_
timestamp 1728304789
transform 1 0 6130 0 -1 1210
box -12 -8 72 252
use OAI21X1  _2419_
timestamp 1728305162
transform 1 0 6210 0 -1 1210
box -12 -8 112 252
use OAI21X1  _2420_
timestamp 1728305162
transform 1 0 6390 0 -1 1210
box -12 -8 112 252
use NAND2X1  _2421_
timestamp 1728304996
transform 1 0 5910 0 -1 730
box -12 -8 92 252
use NAND3X1  _2422_
timestamp 1728305047
transform -1 0 6130 0 -1 1210
box -12 -8 112 252
use INVX1  _2423_
timestamp 1728304789
transform 1 0 5670 0 -1 1210
box -12 -8 72 252
use OAI21X1  _2424_
timestamp 1728305162
transform -1 0 5910 0 -1 1210
box -12 -8 112 252
use NAND2X1  _2425_
timestamp 1728304996
transform -1 0 6030 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2426_
timestamp 1728305162
transform -1 0 6070 0 1 730
box -12 -8 112 252
use DFFPOSX1  _2427_
timestamp 1728340458
transform 1 0 3590 0 1 4090
box -13 -8 253 252
use DFFPOSX1  _2428_
timestamp 1728340458
transform 1 0 4030 0 -1 5530
box -13 -8 253 252
use DFFPOSX1  _2429_
timestamp 1728340458
transform 1 0 4470 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _2430_
timestamp 1728340458
transform 1 0 4070 0 1 6010
box -13 -8 253 252
use DFFPOSX1  _2431_
timestamp 1728340458
transform 1 0 4390 0 1 4570
box -13 -8 253 252
use DFFPOSX1  _2432_
timestamp 1728340458
transform 1 0 3870 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _2433_
timestamp 1728340458
transform 1 0 4630 0 -1 3610
box -13 -8 253 252
use DFFPOSX1  _2434_
timestamp 1728340458
transform 1 0 4250 0 -1 3610
box -13 -8 253 252
use DFFPOSX1  _2435_
timestamp 1728340458
transform 1 0 4830 0 1 3130
box -13 -8 253 252
use DFFPOSX1  _2436_
timestamp 1728340458
transform 1 0 4650 0 -1 4090
box -13 -8 253 252
use DFFPOSX1  _2437_
timestamp 1728340458
transform 1 0 4330 0 1 3610
box -13 -8 253 252
use DFFPOSX1  _2438_
timestamp 1728340458
transform 1 0 3950 0 1 4090
box -13 -8 253 252
use DFFPOSX1  _2439_
timestamp 1728340458
transform 1 0 3130 0 -1 5530
box -13 -8 253 252
use DFFPOSX1  _2440_
timestamp 1728340458
transform 1 0 3790 0 1 5530
box -13 -8 253 252
use DFFPOSX1  _2441_
timestamp 1728340458
transform 1 0 4590 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _2442_
timestamp 1728340458
transform -1 0 4770 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _2443_
timestamp 1728340458
transform 1 0 5550 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _2444_
timestamp 1728340458
transform 1 0 5210 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _2445_
timestamp 1728340458
transform 1 0 6230 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _2446_
timestamp 1728340458
transform -1 0 7130 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _2447_
timestamp 1728340458
transform -1 0 7310 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _2448_
timestamp 1728340458
transform -1 0 7370 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _2449_
timestamp 1728340458
transform -1 0 7710 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _2450_
timestamp 1728340458
transform 1 0 7650 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _2451_
timestamp 1728340458
transform 1 0 7510 0 1 250
box -13 -8 253 252
use DFFPOSX1  _2452_
timestamp 1728340458
transform -1 0 7810 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _2453_
timestamp 1728340458
transform -1 0 7310 0 1 730
box -13 -8 253 252
use DFFPOSX1  _2454_
timestamp 1728340458
transform -1 0 7110 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _2455_
timestamp 1728340458
transform -1 0 5130 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _2456_
timestamp 1728340458
transform -1 0 4910 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _2457_
timestamp 1728340458
transform -1 0 6090 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _2458_
timestamp 1728340458
transform 1 0 5050 0 1 1690
box -13 -8 253 252
use DFFPOSX1  _2459_
timestamp 1728340458
transform -1 0 6750 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _2460_
timestamp 1728340458
transform -1 0 5850 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _2461_
timestamp 1728340458
transform -1 0 4950 0 1 1690
box -13 -8 253 252
use DFFPOSX1  _2462_
timestamp 1728340458
transform -1 0 5530 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _2463_
timestamp 1728340458
transform -1 0 7350 0 -1 1210
box -13 -8 253 252
use DFFPOSX1  _2464_
timestamp 1728340458
transform 1 0 6930 0 -1 1690
box -13 -8 253 252
use DFFPOSX1  _2465_
timestamp 1728340458
transform -1 0 7330 0 -1 730
box -13 -8 253 252
use DFFPOSX1  _2466_
timestamp 1728340458
transform -1 0 7370 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _2467_
timestamp 1728340458
transform -1 0 5850 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _2468_
timestamp 1728340458
transform 1 0 5850 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _2469_
timestamp 1728340458
transform -1 0 6830 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _2470_
timestamp 1728340458
transform -1 0 5970 0 1 730
box -13 -8 253 252
use NOR2X1  _2471_
timestamp 1728305106
transform 1 0 1690 0 -1 5530
box -12 -8 92 252
use INVX1  _2472_
timestamp 1728304789
transform 1 0 1750 0 1 5050
box -12 -8 72 252
use INVX1  _2473_
timestamp 1728304789
transform 1 0 2990 0 1 5530
box -12 -8 72 252
use INVX1  _2474_
timestamp 1728304789
transform 1 0 3070 0 -1 5530
box -12 -8 72 252
use NAND2X1  _2475_
timestamp 1728304996
transform -1 0 2570 0 -1 5530
box -12 -8 92 252
use INVX2  _2476_
timestamp 1728304826
transform 1 0 3390 0 -1 6010
box -12 -8 72 252
use AOI21X1  _2477_
timestamp 1728304211
transform -1 0 3150 0 1 5530
box -12 -8 112 252
use NAND2X1  _2478_
timestamp 1728304996
transform -1 0 3250 0 1 5530
box -12 -8 92 252
use INVX1  _2479_
timestamp 1728304789
transform -1 0 2970 0 1 5050
box -12 -8 72 252
use NAND2X1  _2480_
timestamp 1728304996
transform 1 0 3430 0 1 6010
box -12 -8 92 252
use INVX1  _2481_
timestamp 1728304789
transform 1 0 3510 0 1 6010
box -12 -8 72 252
use NOR2X1  _2482_
timestamp 1728305106
transform -1 0 2910 0 1 5530
box -12 -8 92 252
use INVX1  _2483_
timestamp 1728304789
transform -1 0 2490 0 -1 5530
box -12 -8 72 252
use NOR3X1  _2484_
timestamp 1728303224
transform 1 0 2310 0 1 5530
box -12 -8 192 252
use NAND2X1  _2485_
timestamp 1728304996
transform 1 0 2350 0 -1 5530
box -12 -8 92 252
use NOR2X1  _2486_
timestamp 1728305106
transform -1 0 3070 0 1 5050
box -12 -8 92 252
use INVX1  _2487_
timestamp 1728304789
transform 1 0 2350 0 1 5050
box -12 -8 72 252
use AOI21X1  _2488_
timestamp 1728304211
transform 1 0 2430 0 1 5050
box -12 -8 112 252
use INVX1  _2489_
timestamp 1728304789
transform 1 0 2130 0 1 5050
box -12 -8 72 252
use AOI21X1  _2490_
timestamp 1728304211
transform -1 0 2270 0 1 5530
box -12 -8 112 252
use AOI22X1  _2491_
timestamp 1728304278
transform 1 0 2230 0 1 5050
box -14 -8 132 252
use INVX1  _2492_
timestamp 1728304789
transform 1 0 1970 0 -1 5530
box -12 -8 72 252
use AOI22X1  _2493_
timestamp 1728304278
transform -1 0 2170 0 -1 5530
box -14 -8 132 252
use INVX1  _2494_
timestamp 1728304789
transform -1 0 2230 0 -1 5530
box -12 -8 72 252
use MUX2X1  _2495_
timestamp 1728304958
transform -1 0 2390 0 -1 5050
box -12 -8 131 252
use INVX1  _2496_
timestamp 1728304789
transform -1 0 2950 0 -1 5050
box -12 -8 72 252
use NOR2X1  _2497_
timestamp 1728305106
transform 1 0 2810 0 -1 5050
box -12 -8 92 252
use INVX1  _2498_
timestamp 1728304789
transform -1 0 3250 0 1 4570
box -12 -8 72 252
use NOR2X1  _2499_
timestamp 1728305106
transform 1 0 3110 0 1 4570
box -12 -8 92 252
use INVX1  _2500_
timestamp 1728304789
transform -1 0 3350 0 -1 6010
box -12 -8 72 252
use OAI21X1  _2501_
timestamp 1728305162
transform 1 0 3190 0 -1 6010
box -12 -8 112 252
use NAND2X1  _2502_
timestamp 1728304996
transform 1 0 2910 0 1 5530
box -12 -8 92 252
use OAI21X1  _2503_
timestamp 1728305162
transform -1 0 2710 0 -1 5530
box -12 -8 112 252
use NAND2X1  _2504_
timestamp 1728304996
transform -1 0 2810 0 1 5530
box -12 -8 92 252
use INVX1  _2505_
timestamp 1728304789
transform -1 0 1970 0 -1 5530
box -12 -8 72 252
use OAI21X1  _2506_
timestamp 1728305162
transform -1 0 1910 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2507_
timestamp 1728305162
transform -1 0 1690 0 -1 5530
box -12 -8 112 252
use AOI21X1  _2508_
timestamp 1728304211
transform -1 0 2350 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2509_
timestamp 1728305162
transform 1 0 2710 0 -1 5530
box -12 -8 112 252
use OAI21X1  _2510_
timestamp 1728305162
transform -1 0 2910 0 1 5050
box -12 -8 112 252
use OAI21X1  _2511_
timestamp 1728305162
transform 1 0 3250 0 1 5530
box -12 -8 112 252
use NOR2X1  _2512_
timestamp 1728305106
transform -1 0 3290 0 -1 5050
box -12 -8 92 252
use NOR2X1  _2513_
timestamp 1728305106
transform -1 0 3150 0 1 6010
box -12 -8 92 252
use AND2X2  _2514_
timestamp 1728304163
transform 1 0 2970 0 1 6010
box -12 -8 112 252
use DFFPOSX1  _2515_
timestamp 1728340458
transform 1 0 2530 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _2516_
timestamp 1728340458
transform 1 0 2390 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _2517_
timestamp 1728340458
transform 1 0 3070 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _2518_
timestamp 1728340458
transform 1 0 2950 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _2519_
timestamp 1728340458
transform -1 0 3530 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _2520_
timestamp 1728340458
transform 1 0 3150 0 1 6010
box -13 -8 253 252
use DFFPOSX1  _2521_
timestamp 1728340458
transform -1 0 2730 0 1 5530
box -13 -8 253 252
use DFFPOSX1  _2522_
timestamp 1728340458
transform 1 0 1350 0 -1 5530
box -13 -8 253 252
use DFFPOSX1  _2523_
timestamp 1728340458
transform 1 0 2810 0 -1 5530
box -13 -8 253 252
use DFFPOSX1  _2524_
timestamp 1728340458
transform -1 0 3590 0 1 5530
box -13 -8 253 252
use INVX1  _2525_
timestamp 1728304789
transform -1 0 2990 0 -1 6010
box -12 -8 72 252
use INVX1  _2526_
timestamp 1728304789
transform -1 0 3170 0 -1 6010
box -12 -8 72 252
use NAND2X1  _2527_
timestamp 1728304996
transform 1 0 2850 0 -1 6010
box -12 -8 92 252
use NAND2X1  _2528_
timestamp 1728304996
transform -1 0 2510 0 -1 6010
box -12 -8 92 252
use INVX1  _2529_
timestamp 1728304789
transform -1 0 3730 0 -1 6010
box -12 -8 72 252
use NOR2X1  _2530_
timestamp 1728305106
transform 1 0 3010 0 -1 6010
box -12 -8 92 252
use AOI21X1  _2531_
timestamp 1728304211
transform 1 0 2510 0 -1 6010
box -12 -8 112 252
use NOR2X1  _2532_
timestamp 1728305106
transform 1 0 3470 0 -1 6010
box -12 -8 92 252
use OAI21X1  _2533_
timestamp 1728305162
transform -1 0 3670 0 -1 6010
box -12 -8 112 252
use DFFPOSX1  _2534_
timestamp 1728340458
transform 1 0 2610 0 -1 6010
box -13 -8 253 252
use DFFPOSX1  _2535_
timestamp 1728340458
transform -1 0 3970 0 -1 6010
box -13 -8 253 252
use INVX1  _2536_
timestamp 1728304789
transform -1 0 70 0 -1 2170
box -12 -8 72 252
use INVX1  _2537_
timestamp 1728304789
transform -1 0 2650 0 -1 3610
box -12 -8 72 252
use INVX4  _2538_
timestamp 1728304878
transform 1 0 2410 0 1 3610
box -12 -8 92 252
use INVX1  _2539_
timestamp 1728304789
transform -1 0 2570 0 1 3610
box -12 -8 72 252
use NAND3X1  _2540_
timestamp 1728305047
transform -1 0 2550 0 -1 3610
box -12 -8 112 252
use NAND2X1  _2541_
timestamp 1728304996
transform 1 0 2810 0 1 3610
box -12 -8 92 252
use INVX4  _2542_
timestamp 1728304878
transform 1 0 3370 0 -1 4090
box -12 -8 92 252
use INVX4  _2543_
timestamp 1728304878
transform -1 0 3170 0 1 3610
box -12 -8 92 252
use NAND2X1  _2544_
timestamp 1728304996
transform 1 0 2210 0 -1 3610
box -12 -8 92 252
use INVX1  _2545_
timestamp 1728304789
transform -1 0 2610 0 1 4090
box -12 -8 72 252
use NAND3X1  _2546_
timestamp 1728305047
transform -1 0 2710 0 1 4090
box -12 -8 112 252
use OAI22X1  _2547_
timestamp 1728305200
transform -1 0 2110 0 -1 3610
box -12 -8 132 252
use NOR2X1  _2548_
timestamp 1728305106
transform 1 0 2850 0 1 4090
box -12 -8 92 252
use NAND2X1  _2549_
timestamp 1728304996
transform 1 0 3050 0 1 4090
box -12 -8 92 252
use NOR2X1  _2550_
timestamp 1728305106
transform -1 0 3010 0 1 4090
box -12 -8 92 252
use NAND2X1  _2551_
timestamp 1728304996
transform -1 0 2830 0 -1 4090
box -12 -8 92 252
use NOR2X1  _2552_
timestamp 1728305106
transform -1 0 630 0 -1 2170
box -12 -8 92 252
use NOR2X1  _2553_
timestamp 1728305106
transform 1 0 2290 0 -1 3610
box -12 -8 92 252
use OAI21X1  _2554_
timestamp 1728305162
transform -1 0 310 0 -1 2170
box -12 -8 112 252
use OAI22X1  _2555_
timestamp 1728305200
transform 1 0 70 0 -1 2170
box -12 -8 132 252
use INVX1  _2556_
timestamp 1728304789
transform 1 0 1810 0 -1 3130
box -12 -8 72 252
use NOR2X1  _2557_
timestamp 1728305106
transform -1 0 1410 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2558_
timestamp 1728305162
transform -1 0 1330 0 -1 3130
box -12 -8 112 252
use OAI22X1  _2559_
timestamp 1728305200
transform -1 0 1530 0 -1 3130
box -12 -8 132 252
use INVX1  _2560_
timestamp 1728304789
transform -1 0 2850 0 1 2170
box -12 -8 72 252
use NOR2X1  _2561_
timestamp 1728305106
transform -1 0 2650 0 -1 2170
box -12 -8 92 252
use OAI21X1  _2562_
timestamp 1728305162
transform 1 0 2530 0 1 2170
box -12 -8 112 252
use OAI22X1  _2563_
timestamp 1728305200
transform -1 0 2750 0 1 2170
box -12 -8 132 252
use INVX1  _2564_
timestamp 1728304789
transform 1 0 790 0 1 2650
box -12 -8 72 252
use NOR2X1  _2565_
timestamp 1728305106
transform 1 0 510 0 -1 2650
box -12 -8 92 252
use OAI21X1  _2566_
timestamp 1728305162
transform 1 0 250 0 1 2650
box -12 -8 112 252
use OAI22X1  _2567_
timestamp 1728305200
transform -1 0 510 0 1 2650
box -12 -8 132 252
use INVX1  _2568_
timestamp 1728304789
transform -1 0 1130 0 -1 2170
box -12 -8 72 252
use NOR2X1  _2569_
timestamp 1728305106
transform -1 0 910 0 -1 2170
box -12 -8 92 252
use OAI21X1  _2570_
timestamp 1728305162
transform 1 0 630 0 -1 2170
box -12 -8 112 252
use OAI22X1  _2571_
timestamp 1728305200
transform -1 0 1070 0 -1 2170
box -12 -8 132 252
use INVX1  _2572_
timestamp 1728304789
transform 1 0 3090 0 1 2650
box -12 -8 72 252
use NOR2X1  _2573_
timestamp 1728305106
transform -1 0 2910 0 -1 2650
box -12 -8 92 252
use OAI21X1  _2574_
timestamp 1728305162
transform 1 0 2830 0 1 2650
box -12 -8 112 252
use OAI22X1  _2575_
timestamp 1728305200
transform -1 0 3090 0 1 2650
box -12 -8 132 252
use INVX1  _2576_
timestamp 1728304789
transform 1 0 350 0 -1 3610
box -12 -8 72 252
use NOR2X1  _2577_
timestamp 1728305106
transform 1 0 590 0 -1 3610
box -12 -8 92 252
use OAI21X1  _2578_
timestamp 1728305162
transform -1 0 770 0 -1 3610
box -12 -8 112 252
use OAI22X1  _2579_
timestamp 1728305200
transform 1 0 450 0 -1 3610
box -12 -8 132 252
use INVX1  _2580_
timestamp 1728304789
transform -1 0 1530 0 1 3610
box -12 -8 72 252
use NOR2X1  _2581_
timestamp 1728305106
transform -1 0 1310 0 -1 3610
box -12 -8 92 252
use OAI21X1  _2582_
timestamp 1728305162
transform 1 0 1110 0 -1 3610
box -12 -8 112 252
use OAI22X1  _2583_
timestamp 1728305200
transform -1 0 1450 0 -1 3610
box -12 -8 132 252
use INVX4  _2584_
timestamp 1728304878
transform -1 0 2770 0 -1 4570
box -12 -8 92 252
use NAND2X1  _2585_
timestamp 1728304996
transform -1 0 1390 0 -1 1690
box -12 -8 92 252
use MUX2X1  _2586_
timestamp 1728304958
transform 1 0 1850 0 1 1690
box -12 -8 131 252
use MUX2X1  _2587_
timestamp 1728304958
transform 1 0 1550 0 1 1690
box -12 -8 131 252
use MUX2X1  _2588_
timestamp 1728304958
transform -1 0 1810 0 1 1690
box -12 -8 131 252
use MUX2X1  _2589_
timestamp 1728304958
transform -1 0 2710 0 -1 1210
box -12 -8 131 252
use MUX2X1  _2590_
timestamp 1728304958
transform 1 0 1890 0 1 730
box -12 -8 131 252
use MUX2X1  _2591_
timestamp 1728304958
transform -1 0 2250 0 1 1210
box -12 -8 131 252
use MUX2X1  _2592_
timestamp 1728304958
transform -1 0 1630 0 -1 1690
box -12 -8 131 252
use OAI21X1  _2593_
timestamp 1728305162
transform -1 0 1490 0 -1 1690
box -12 -8 112 252
use INVX1  _2594_
timestamp 1728304789
transform -1 0 2990 0 -1 3130
box -12 -8 72 252
use INVX2  _2595_
timestamp 1728304826
transform 1 0 1950 0 1 2650
box -12 -8 72 252
use MUX2X1  _2596_
timestamp 1728304958
transform -1 0 2630 0 1 3130
box -12 -8 131 252
use MUX2X1  _2597_
timestamp 1728304958
transform -1 0 3210 0 1 3130
box -12 -8 131 252
use MUX2X1  _2598_
timestamp 1728304958
transform 1 0 2770 0 1 3130
box -12 -8 131 252
use AOI22X1  _2599_
timestamp 1728304278
transform 1 0 2650 0 -1 3130
box -14 -8 132 252
use INVX1  _2600_
timestamp 1728304789
transform 1 0 3030 0 1 3130
box -12 -8 72 252
use NAND3X1  _2601_
timestamp 1728305047
transform -1 0 2790 0 -1 3610
box -12 -8 112 252
use NAND2X1  _2602_
timestamp 1728304996
transform 1 0 2370 0 -1 3610
box -12 -8 92 252
use MUX2X1  _2603_
timestamp 1728304958
transform 1 0 3330 0 1 3130
box -12 -8 131 252
use OAI22X1  _2604_
timestamp 1728305200
transform 1 0 3190 0 -1 3130
box -12 -8 132 252
use NOR2X1  _2605_
timestamp 1728305106
transform 1 0 3110 0 -1 3130
box -12 -8 92 252
use AOI22X1  _2606_
timestamp 1728304278
transform -1 0 2890 0 -1 3130
box -14 -8 132 252
use INVX1  _2607_
timestamp 1728304789
transform -1 0 2790 0 1 1690
box -12 -8 72 252
use MUX2X1  _2608_
timestamp 1728304958
transform -1 0 790 0 1 1210
box -12 -8 131 252
use MUX2X1  _2609_
timestamp 1728304958
transform -1 0 3250 0 1 1210
box -12 -8 131 252
use MUX2X1  _2610_
timestamp 1728304958
transform 1 0 2250 0 1 1210
box -12 -8 131 252
use AOI22X1  _2611_
timestamp 1728304278
transform -1 0 2450 0 -1 1690
box -14 -8 132 252
use INVX1  _2612_
timestamp 1728304789
transform -1 0 2370 0 1 1690
box -12 -8 72 252
use MUX2X1  _2613_
timestamp 1728304958
transform 1 0 3350 0 1 1690
box -12 -8 131 252
use OAI22X1  _2614_
timestamp 1728305200
transform 1 0 2790 0 1 1690
box -12 -8 132 252
use NOR2X1  _2615_
timestamp 1728305106
transform -1 0 2590 0 1 1690
box -12 -8 92 252
use AOI22X1  _2616_
timestamp 1728304278
transform -1 0 2710 0 1 1690
box -14 -8 132 252
use INVX1  _2617_
timestamp 1728304789
transform 1 0 1250 0 1 2650
box -12 -8 72 252
use MUX2X1  _2618_
timestamp 1728304958
transform -1 0 1030 0 -1 730
box -12 -8 131 252
use MUX2X1  _2619_
timestamp 1728304958
transform -1 0 1390 0 1 730
box -12 -8 131 252
use MUX2X1  _2620_
timestamp 1728304958
transform 1 0 1070 0 1 730
box -12 -8 131 252
use MUX2X1  _2621_
timestamp 1728304958
transform -1 0 1030 0 1 2170
box -12 -8 131 252
use OAI22X1  _2622_
timestamp 1728305200
transform -1 0 990 0 1 2650
box -12 -8 132 252
use AOI21X1  _2623_
timestamp 1728304211
transform 1 0 990 0 1 2650
box -12 -8 112 252
use INVX1  _2624_
timestamp 1728304789
transform 1 0 1450 0 1 2650
box -12 -8 72 252
use AOI21X1  _2625_
timestamp 1728304211
transform -1 0 1410 0 1 2650
box -12 -8 112 252
use AOI22X1  _2626_
timestamp 1728304278
transform -1 0 1230 0 1 2650
box -14 -8 132 252
use INVX1  _2627_
timestamp 1728304789
transform 1 0 850 0 1 1210
box -12 -8 72 252
use MUX2X1  _2628_
timestamp 1728304958
transform -1 0 1190 0 -1 730
box -12 -8 131 252
use MUX2X1  _2629_
timestamp 1728304958
transform -1 0 1390 0 1 1210
box -12 -8 131 252
use MUX2X1  _2630_
timestamp 1728304958
transform -1 0 1110 0 -1 1210
box -12 -8 131 252
use AOI22X1  _2631_
timestamp 1728304278
transform -1 0 1070 0 -1 1690
box -14 -8 132 252
use INVX1  _2632_
timestamp 1728304789
transform 1 0 1210 0 1 1690
box -12 -8 72 252
use MUX2X1  _2633_
timestamp 1728304958
transform 1 0 930 0 1 1690
box -12 -8 131 252
use OAI22X1  _2634_
timestamp 1728305200
transform -1 0 1170 0 1 1690
box -12 -8 132 252
use NOR2X1  _2635_
timestamp 1728305106
transform 1 0 1070 0 1 1210
box -12 -8 92 252
use AOI22X1  _2636_
timestamp 1728304278
transform 1 0 910 0 1 1210
box -14 -8 132 252
use INVX1  _2637_
timestamp 1728304789
transform -1 0 2870 0 -1 2170
box -12 -8 72 252
use MUX2X1  _2638_
timestamp 1728304958
transform 1 0 2030 0 1 250
box -12 -8 131 252
use MUX2X1  _2639_
timestamp 1728304958
transform 1 0 2830 0 1 730
box -12 -8 131 252
use MUX2X1  _2640_
timestamp 1728304958
transform 1 0 2470 0 1 730
box -12 -8 131 252
use AOI22X1  _2641_
timestamp 1728304278
transform -1 0 2790 0 -1 2170
box -14 -8 132 252
use INVX1  _2642_
timestamp 1728304789
transform 1 0 3150 0 -1 2650
box -12 -8 72 252
use MUX2X1  _2643_
timestamp 1728304958
transform -1 0 3310 0 1 1690
box -12 -8 131 252
use OAI22X1  _2644_
timestamp 1728305200
transform 1 0 3230 0 -1 2170
box -12 -8 132 252
use NOR2X1  _2645_
timestamp 1728305106
transform 1 0 3370 0 -1 2170
box -12 -8 92 252
use AOI22X1  _2646_
timestamp 1728304278
transform 1 0 2870 0 -1 2170
box -14 -8 132 252
use INVX1  _2647_
timestamp 1728304789
transform 1 0 890 0 1 3610
box -12 -8 72 252
use MUX2X1  _2648_
timestamp 1728304958
transform 1 0 970 0 -1 4570
box -12 -8 131 252
use MUX2X1  _2649_
timestamp 1728304958
transform -1 0 1670 0 -1 5050
box -12 -8 131 252
use MUX2X1  _2650_
timestamp 1728304958
transform 1 0 1090 0 -1 4570
box -12 -8 131 252
use AOI22X1  _2651_
timestamp 1728304278
transform 1 0 1110 0 1 3610
box -14 -8 132 252
use INVX1  _2652_
timestamp 1728304789
transform -1 0 1410 0 -1 4090
box -12 -8 72 252
use MUX2X1  _2653_
timestamp 1728304958
transform -1 0 830 0 -1 4090
box -12 -8 131 252
use OAI22X1  _2654_
timestamp 1728305200
transform -1 0 1470 0 1 3610
box -12 -8 132 252
use NOR2X1  _2655_
timestamp 1728305106
transform 1 0 1230 0 1 3610
box -12 -8 92 252
use AOI22X1  _2656_
timestamp 1728304278
transform 1 0 970 0 1 3610
box -14 -8 132 252
use INVX1  _2657_
timestamp 1728304789
transform 1 0 1430 0 -1 4570
box -12 -8 72 252
use MUX2X1  _2658_
timestamp 1728304958
transform 1 0 930 0 -1 5050
box -12 -8 131 252
use MUX2X1  _2659_
timestamp 1728304958
transform -1 0 1790 0 1 4570
box -12 -8 131 252
use MUX2X1  _2660_
timestamp 1728304958
transform 1 0 1230 0 1 4570
box -12 -8 131 252
use MUX2X1  _2661_
timestamp 1728304958
transform 1 0 830 0 -1 4090
box -12 -8 131 252
use OAI22X1  _2662_
timestamp 1728305200
transform 1 0 1130 0 -1 4090
box -12 -8 132 252
use AOI21X1  _2663_
timestamp 1728304211
transform -1 0 1310 0 -1 4570
box -12 -8 112 252
use AOI21X1  _2664_
timestamp 1728304211
transform -1 0 1470 0 1 3130
box -12 -8 112 252
use AOI22X1  _2665_
timestamp 1728304278
transform -1 0 1430 0 -1 4570
box -14 -8 132 252
use INVX1  _2666_
timestamp 1728304789
transform 1 0 2750 0 -1 1210
box -12 -8 72 252
use NAND2X1  _2667_
timestamp 1728304996
transform -1 0 2150 0 1 4090
box -12 -8 92 252
use NAND3X1  _2668_
timestamp 1728305047
transform -1 0 2670 0 1 3610
box -12 -8 112 252
use NAND2X1  _2669_
timestamp 1728304996
transform -1 0 2630 0 -1 4090
box -12 -8 92 252
use OAI22X1  _2670_
timestamp 1728305200
transform 1 0 2130 0 -1 4090
box -12 -8 132 252
use NOR2X1  _2671_
timestamp 1728305106
transform 1 0 3190 0 1 3610
box -12 -8 92 252
use NAND2X1  _2672_
timestamp 1728304996
transform -1 0 2510 0 1 4090
box -12 -8 92 252
use NOR2X1  _2673_
timestamp 1728305106
transform 1 0 2110 0 -1 1210
box -12 -8 92 252
use NOR2X1  _2674_
timestamp 1728305106
transform -1 0 2430 0 1 4090
box -12 -8 92 252
use OAI21X1  _2675_
timestamp 1728305162
transform 1 0 2210 0 -1 1210
box -12 -8 112 252
use OAI22X1  _2676_
timestamp 1728305200
transform -1 0 2430 0 -1 1210
box -12 -8 132 252
use INVX1  _2677_
timestamp 1728304789
transform 1 0 3310 0 -1 3610
box -12 -8 72 252
use NOR2X1  _2678_
timestamp 1728305106
transform 1 0 2990 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2679_
timestamp 1728305162
transform -1 0 2910 0 -1 3610
box -12 -8 112 252
use OAI22X1  _2680_
timestamp 1728305200
transform -1 0 3030 0 -1 3610
box -12 -8 132 252
use INVX1  _2681_
timestamp 1728304789
transform 1 0 3290 0 1 1210
box -12 -8 72 252
use NOR2X1  _2682_
timestamp 1728305106
transform -1 0 2450 0 1 1210
box -12 -8 92 252
use OAI21X1  _2683_
timestamp 1728305162
transform -1 0 2690 0 1 1210
box -12 -8 112 252
use OAI22X1  _2684_
timestamp 1728305200
transform -1 0 2850 0 1 1210
box -12 -8 132 252
use INVX1  _2685_
timestamp 1728304789
transform 1 0 1350 0 -1 1210
box -12 -8 72 252
use NOR2X1  _2686_
timestamp 1728305106
transform 1 0 1890 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2687_
timestamp 1728305162
transform -1 0 1670 0 -1 1210
box -12 -8 112 252
use OAI22X1  _2688_
timestamp 1728305200
transform 1 0 1450 0 -1 1210
box -12 -8 132 252
use INVX1  _2689_
timestamp 1728304789
transform 1 0 1890 0 1 1210
box -12 -8 72 252
use NOR2X1  _2690_
timestamp 1728305106
transform 1 0 1790 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2691_
timestamp 1728305162
transform 1 0 1630 0 1 1210
box -12 -8 112 252
use OAI22X1  _2692_
timestamp 1728305200
transform -1 0 1890 0 1 1210
box -12 -8 132 252
use INVX1  _2693_
timestamp 1728304789
transform 1 0 3170 0 -1 1210
box -12 -8 72 252
use NOR2X1  _2694_
timestamp 1728305106
transform -1 0 3170 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2695_
timestamp 1728305162
transform 1 0 2810 0 -1 1210
box -12 -8 112 252
use OAI22X1  _2696_
timestamp 1728305200
transform -1 0 3070 0 -1 1210
box -12 -8 132 252
use INVX1  _2697_
timestamp 1728304789
transform 1 0 1910 0 -1 5050
box -12 -8 72 252
use NOR2X1  _2698_
timestamp 1728305106
transform -1 0 1630 0 1 4090
box -12 -8 92 252
use OAI21X1  _2699_
timestamp 1728305162
transform 1 0 1970 0 1 4090
box -12 -8 112 252
use OAI22X1  _2700_
timestamp 1728305200
transform -1 0 1850 0 1 4090
box -12 -8 132 252
use INVX1  _2701_
timestamp 1728304789
transform 1 0 1850 0 -1 4570
box -12 -8 72 252
use NOR2X1  _2702_
timestamp 1728305106
transform -1 0 1710 0 1 4090
box -12 -8 92 252
use OAI21X1  _2703_
timestamp 1728305162
transform 1 0 1850 0 -1 4090
box -12 -8 112 252
use OAI22X1  _2704_
timestamp 1728305200
transform -1 0 1970 0 1 4090
box -12 -8 132 252
use INVX1  _2705_
timestamp 1728304789
transform -1 0 2350 0 -1 730
box -12 -8 72 252
use NAND3X1  _2706_
timestamp 1728305047
transform -1 0 2770 0 1 3610
box -12 -8 112 252
use NAND3X1  _2707_
timestamp 1728305047
transform 1 0 2750 0 1 4090
box -12 -8 112 252
use OAI22X1  _2708_
timestamp 1728305200
transform 1 0 2150 0 1 4090
box -12 -8 132 252
use INVX1  _2709_
timestamp 1728304789
transform -1 0 3010 0 -1 4090
box -12 -8 72 252
use NAND2X1  _2710_
timestamp 1728304996
transform 1 0 3010 0 -1 4090
box -12 -8 92 252
use NOR2X1  _2711_
timestamp 1728305106
transform 1 0 2150 0 1 730
box -12 -8 92 252
use NOR2X1  _2712_
timestamp 1728305106
transform 1 0 2270 0 1 4090
box -12 -8 92 252
use OAI21X1  _2713_
timestamp 1728305162
transform 1 0 2050 0 -1 730
box -12 -8 112 252
use OAI22X1  _2714_
timestamp 1728305200
transform -1 0 2270 0 -1 730
box -12 -8 132 252
use INVX1  _2715_
timestamp 1728304789
transform 1 0 3990 0 1 2650
box -12 -8 72 252
use NOR2X1  _2716_
timestamp 1728305106
transform 1 0 3610 0 1 2650
box -12 -8 92 252
use OAI21X1  _2717_
timestamp 1728305162
transform 1 0 3390 0 1 2650
box -12 -8 112 252
use OAI22X1  _2718_
timestamp 1728305200
transform -1 0 3850 0 1 2650
box -12 -8 132 252
use INVX1  _2719_
timestamp 1728304789
transform -1 0 2910 0 -1 730
box -12 -8 72 252
use NOR2X1  _2720_
timestamp 1728305106
transform -1 0 2790 0 1 730
box -12 -8 92 252
use OAI21X1  _2721_
timestamp 1728305162
transform -1 0 2690 0 -1 730
box -12 -8 112 252
use OAI22X1  _2722_
timestamp 1728305200
transform -1 0 2850 0 -1 730
box -12 -8 132 252
use INVX1  _2723_
timestamp 1728304789
transform 1 0 1310 0 -1 250
box -12 -8 72 252
use NOR2X1  _2724_
timestamp 1728305106
transform -1 0 1430 0 1 250
box -12 -8 92 252
use OAI21X1  _2725_
timestamp 1728305162
transform -1 0 1570 0 -1 730
box -12 -8 112 252
use OAI22X1  _2726_
timestamp 1728305200
transform 1 0 1410 0 -1 250
box -12 -8 132 252
use INVX1  _2727_
timestamp 1728304789
transform -1 0 1830 0 -1 250
box -12 -8 72 252
use NOR2X1  _2728_
timestamp 1728305106
transform -1 0 1330 0 1 250
box -12 -8 92 252
use OAI21X1  _2729_
timestamp 1728305162
transform -1 0 1530 0 1 250
box -12 -8 112 252
use OAI22X1  _2730_
timestamp 1728305200
transform -1 0 1690 0 1 250
box -12 -8 132 252
use INVX1  _2731_
timestamp 1728304789
transform -1 0 2610 0 -1 250
box -12 -8 72 252
use NOR2X1  _2732_
timestamp 1728305106
transform -1 0 2350 0 1 250
box -12 -8 92 252
use OAI21X1  _2733_
timestamp 1728305162
transform -1 0 2450 0 1 250
box -12 -8 112 252
use OAI22X1  _2734_
timestamp 1728305200
transform -1 0 2550 0 -1 250
box -12 -8 132 252
use INVX1  _2735_
timestamp 1728304789
transform -1 0 1430 0 1 4570
box -12 -8 72 252
use NOR2X1  _2736_
timestamp 1728305106
transform -1 0 1330 0 -1 4090
box -12 -8 92 252
use OAI21X1  _2737_
timestamp 1728305162
transform -1 0 1530 0 1 4090
box -12 -8 112 252
use OAI22X1  _2738_
timestamp 1728305200
transform -1 0 1390 0 1 4090
box -12 -8 132 252
use INVX1  _2739_
timestamp 1728304789
transform -1 0 1830 0 -1 4570
box -12 -8 72 252
use NOR2X1  _2740_
timestamp 1728305106
transform 1 0 1650 0 -1 4090
box -12 -8 92 252
use OAI21X1  _2741_
timestamp 1728305162
transform 1 0 1530 0 -1 4570
box -12 -8 112 252
use OAI22X1  _2742_
timestamp 1728305200
transform -1 0 1750 0 -1 4570
box -12 -8 132 252
use NAND2X1  _2743_
timestamp 1728304996
transform 1 0 2330 0 1 3610
box -12 -8 92 252
use OR2X2  _2744_
timestamp 1728305284
transform 1 0 2210 0 1 3610
box -12 -8 112 252
use NAND2X1  _2745_
timestamp 1728304996
transform 1 0 2990 0 1 3610
box -12 -8 92 252
use INVX2  _2746_
timestamp 1728304826
transform -1 0 2950 0 1 3610
box -12 -8 72 252
use NAND2X1  _2747_
timestamp 1728304996
transform 1 0 2410 0 -1 4570
box -12 -8 92 252
use NAND3X1  _2748_
timestamp 1728305047
transform -1 0 1790 0 -1 730
box -12 -8 112 252
use NOR2X1  _2749_
timestamp 1728305106
transform 1 0 1770 0 1 730
box -12 -8 92 252
use NOR2X1  _2750_
timestamp 1728305106
transform 1 0 2130 0 1 3610
box -12 -8 92 252
use NOR2X1  _2751_
timestamp 1728305106
transform 1 0 1890 0 -1 3610
box -12 -8 92 252
use AOI21X1  _2752_
timestamp 1728304211
transform 1 0 1530 0 1 730
box -12 -8 112 252
use OAI21X1  _2753_
timestamp 1728305162
transform -1 0 1730 0 1 730
box -12 -8 112 252
use NAND3X1  _2754_
timestamp 1728305047
transform -1 0 2170 0 -1 3130
box -12 -8 112 252
use NOR2X1  _2755_
timestamp 1728305106
transform -1 0 1950 0 -1 3130
box -12 -8 92 252
use AOI21X1  _2756_
timestamp 1728304211
transform 1 0 1930 0 1 3130
box -12 -8 112 252
use OAI21X1  _2757_
timestamp 1728305162
transform 1 0 1950 0 -1 3130
box -12 -8 112 252
use NAND3X1  _2758_
timestamp 1728305047
transform 1 0 230 0 -1 1210
box -12 -8 112 252
use NOR2X1  _2759_
timestamp 1728305106
transform -1 0 430 0 1 730
box -12 -8 92 252
use AOI21X1  _2760_
timestamp 1728304211
transform -1 0 570 0 1 730
box -12 -8 112 252
use OAI21X1  _2761_
timestamp 1728305162
transform -1 0 350 0 1 730
box -12 -8 112 252
use NAND3X1  _2762_
timestamp 1728305047
transform -1 0 590 0 -1 250
box -12 -8 112 252
use NOR2X1  _2763_
timestamp 1728305106
transform 1 0 470 0 1 250
box -12 -8 92 252
use AOI21X1  _2764_
timestamp 1728304211
transform 1 0 370 0 1 250
box -12 -8 112 252
use OAI21X1  _2765_
timestamp 1728305162
transform -1 0 470 0 -1 250
box -12 -8 112 252
use NAND3X1  _2766_
timestamp 1728305047
transform -1 0 370 0 -1 250
box -12 -8 112 252
use NOR2X1  _2767_
timestamp 1728305106
transform 1 0 130 0 1 250
box -12 -8 92 252
use AOI21X1  _2768_
timestamp 1728304211
transform -1 0 330 0 1 250
box -12 -8 112 252
use OAI21X1  _2769_
timestamp 1728305162
transform -1 0 130 0 1 250
box -12 -8 112 252
use NAND3X1  _2770_
timestamp 1728305047
transform -1 0 2170 0 -1 250
box -12 -8 112 252
use NOR2X1  _2771_
timestamp 1728305106
transform -1 0 1810 0 1 250
box -12 -8 92 252
use AOI21X1  _2772_
timestamp 1728304211
transform 1 0 1810 0 1 250
box -12 -8 112 252
use OAI21X1  _2773_
timestamp 1728305162
transform 1 0 1930 0 1 250
box -12 -8 112 252
use NAND3X1  _2774_
timestamp 1728305047
transform -1 0 550 0 -1 4570
box -12 -8 112 252
use NOR2X1  _2775_
timestamp 1728305106
transform -1 0 330 0 -1 4570
box -12 -8 92 252
use AOI21X1  _2776_
timestamp 1728304211
transform -1 0 350 0 -1 3610
box -12 -8 112 252
use OAI21X1  _2777_
timestamp 1728305162
transform 1 0 350 0 -1 4570
box -12 -8 112 252
use NAND3X1  _2778_
timestamp 1728305047
transform -1 0 890 0 -1 4570
box -12 -8 112 252
use NOR2X1  _2779_
timestamp 1728305106
transform -1 0 670 0 -1 4570
box -12 -8 92 252
use AOI21X1  _2780_
timestamp 1728304211
transform -1 0 870 0 -1 3610
box -12 -8 112 252
use OAI21X1  _2781_
timestamp 1728305162
transform 1 0 690 0 -1 4570
box -12 -8 112 252
use INVX1  _2782_
timestamp 1728304789
transform -1 0 1930 0 -1 1690
box -12 -8 72 252
use NAND2X1  _2783_
timestamp 1728304996
transform 1 0 2670 0 -1 4090
box -12 -8 92 252
use OAI22X1  _2784_
timestamp 1728305200
transform -1 0 2370 0 -1 4090
box -12 -8 132 252
use NOR2X1  _2785_
timestamp 1728305106
transform 1 0 3290 0 -1 4090
box -12 -8 92 252
use NAND2X1  _2786_
timestamp 1728304996
transform 1 0 3210 0 -1 4090
box -12 -8 92 252
use NOR2X1  _2787_
timestamp 1728305106
transform -1 0 1710 0 -1 1690
box -12 -8 92 252
use NOR2X1  _2788_
timestamp 1728305106
transform 1 0 2050 0 -1 4090
box -12 -8 92 252
use OAI21X1  _2789_
timestamp 1728305162
transform 1 0 1970 0 1 1690
box -12 -8 112 252
use OAI22X1  _2790_
timestamp 1728305200
transform -1 0 1870 0 -1 1690
box -12 -8 132 252
use INVX1  _2791_
timestamp 1728304789
transform 1 0 3610 0 1 3130
box -12 -8 72 252
use NOR2X1  _2792_
timestamp 1728305106
transform -1 0 3530 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2793_
timestamp 1728305162
transform 1 0 3210 0 1 3130
box -12 -8 112 252
use OAI22X1  _2794_
timestamp 1728305200
transform -1 0 3610 0 1 3130
box -12 -8 132 252
use INVX1  _2795_
timestamp 1728304789
transform -1 0 3390 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2796_
timestamp 1728305106
transform -1 0 3170 0 -1 1690
box -12 -8 92 252
use OAI21X1  _2797_
timestamp 1728305162
transform -1 0 3070 0 -1 1690
box -12 -8 112 252
use OAI22X1  _2798_
timestamp 1728305200
transform -1 0 3330 0 -1 1690
box -12 -8 132 252
use INVX1  _2799_
timestamp 1728304789
transform 1 0 850 0 1 2170
box -12 -8 72 252
use NOR2X1  _2800_
timestamp 1728305106
transform -1 0 810 0 -1 2170
box -12 -8 92 252
use OAI21X1  _2801_
timestamp 1728305162
transform -1 0 730 0 1 2170
box -12 -8 112 252
use OAI22X1  _2802_
timestamp 1728305200
transform -1 0 850 0 1 2170
box -12 -8 132 252
use INVX1  _2803_
timestamp 1728304789
transform -1 0 170 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2804_
timestamp 1728305106
transform -1 0 90 0 -1 1690
box -12 -8 92 252
use OAI21X1  _2805_
timestamp 1728305162
transform 1 0 330 0 -1 1690
box -12 -8 112 252
use OAI22X1  _2806_
timestamp 1728305200
transform 1 0 170 0 -1 1690
box -12 -8 132 252
use INVX1  _2807_
timestamp 1728304789
transform -1 0 2730 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2808_
timestamp 1728305106
transform -1 0 2530 0 -1 1690
box -12 -8 92 252
use OAI21X1  _2809_
timestamp 1728305162
transform 1 0 2210 0 -1 1690
box -12 -8 112 252
use OAI22X1  _2810_
timestamp 1728305200
transform -1 0 2650 0 -1 1690
box -12 -8 132 252
use INVX1  _2811_
timestamp 1728304789
transform -1 0 210 0 -1 4570
box -12 -8 72 252
use NOR2X1  _2812_
timestamp 1728305106
transform -1 0 90 0 1 4090
box -12 -8 92 252
use OAI21X1  _2813_
timestamp 1728305162
transform -1 0 230 0 1 4090
box -12 -8 112 252
use OAI22X1  _2814_
timestamp 1728305200
transform -1 0 130 0 -1 4570
box -12 -8 132 252
use INVX1  _2815_
timestamp 1728304789
transform -1 0 650 0 1 4090
box -12 -8 72 252
use NOR2X1  _2816_
timestamp 1728305106
transform -1 0 570 0 1 4090
box -12 -8 92 252
use OAI21X1  _2817_
timestamp 1728305162
transform -1 0 350 0 1 4090
box -12 -8 112 252
use OAI22X1  _2818_
timestamp 1728305200
transform -1 0 490 0 1 4090
box -12 -8 132 252
use OAI22X1  _2819_
timestamp 1728305200
transform -1 0 2130 0 1 3610
box -12 -8 132 252
use INVX2  _2820_
timestamp 1728304826
transform 1 0 610 0 1 730
box -12 -8 72 252
use NAND2X1  _2821_
timestamp 1728304996
transform -1 0 750 0 -1 1210
box -12 -8 92 252
use NOR2X1  _2822_
timestamp 1728305106
transform 1 0 1810 0 -1 3610
box -12 -8 92 252
use INVX2  _2823_
timestamp 1728304826
transform 1 0 890 0 -1 1690
box -12 -8 72 252
use NOR2X1  _2824_
timestamp 1728305106
transform -1 0 670 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2825_
timestamp 1728305162
transform 1 0 870 0 -1 1210
box -12 -8 112 252
use OAI21X1  _2826_
timestamp 1728305162
transform -1 0 870 0 -1 1210
box -12 -8 112 252
use NAND2X1  _2827_
timestamp 1728304996
transform 1 0 1010 0 -1 3130
box -12 -8 92 252
use NOR2X1  _2828_
timestamp 1728305106
transform -1 0 1210 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2829_
timestamp 1728305162
transform -1 0 890 0 -1 3130
box -12 -8 112 252
use OAI21X1  _2830_
timestamp 1728305162
transform 1 0 910 0 -1 3130
box -12 -8 112 252
use NAND2X1  _2831_
timestamp 1728304996
transform 1 0 590 0 1 1210
box -12 -8 92 252
use NOR2X1  _2832_
timestamp 1728305106
transform -1 0 450 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2833_
timestamp 1728305162
transform -1 0 550 0 -1 1210
box -12 -8 112 252
use OAI21X1  _2834_
timestamp 1728305162
transform 1 0 490 0 1 1210
box -12 -8 112 252
use NAND2X1  _2835_
timestamp 1728304996
transform -1 0 370 0 -1 730
box -12 -8 92 252
use NOR2X1  _2836_
timestamp 1728305106
transform 1 0 470 0 -1 730
box -12 -8 92 252
use OAI21X1  _2837_
timestamp 1728305162
transform 1 0 570 0 -1 730
box -12 -8 112 252
use OAI21X1  _2838_
timestamp 1728305162
transform -1 0 470 0 -1 730
box -12 -8 112 252
use NAND2X1  _2839_
timestamp 1728304996
transform -1 0 930 0 1 250
box -12 -8 92 252
use NOR2X1  _2840_
timestamp 1728305106
transform -1 0 630 0 1 250
box -12 -8 92 252
use OAI21X1  _2841_
timestamp 1728305162
transform 1 0 690 0 1 730
box -12 -8 112 252
use OAI21X1  _2842_
timestamp 1728305162
transform 1 0 710 0 1 250
box -12 -8 112 252
use NAND2X1  _2843_
timestamp 1728304996
transform -1 0 1050 0 1 250
box -12 -8 92 252
use NOR2X1  _2844_
timestamp 1728305106
transform -1 0 1130 0 1 250
box -12 -8 92 252
use OAI21X1  _2845_
timestamp 1728305162
transform 1 0 1590 0 -1 730
box -12 -8 112 252
use OAI21X1  _2846_
timestamp 1728305162
transform -1 0 1230 0 1 250
box -12 -8 112 252
use NAND2X1  _2847_
timestamp 1728304996
transform 1 0 290 0 1 3130
box -12 -8 92 252
use NOR2X1  _2848_
timestamp 1728305106
transform -1 0 550 0 1 3130
box -12 -8 92 252
use OAI21X1  _2849_
timestamp 1728305162
transform 1 0 570 0 1 3130
box -12 -8 112 252
use OAI21X1  _2850_
timestamp 1728305162
transform -1 0 470 0 1 3130
box -12 -8 112 252
use NAND2X1  _2851_
timestamp 1728304996
transform 1 0 1030 0 1 3130
box -12 -8 92 252
use NOR2X1  _2852_
timestamp 1728305106
transform -1 0 870 0 1 3130
box -12 -8 92 252
use OAI21X1  _2853_
timestamp 1728305162
transform -1 0 770 0 1 3130
box -12 -8 112 252
use OAI21X1  _2854_
timestamp 1728305162
transform 1 0 910 0 1 3130
box -12 -8 112 252
use NOR2X1  _2855_
timestamp 1728305106
transform 1 0 2150 0 1 3130
box -12 -8 92 252
use NAND2X1  _2856_
timestamp 1728304996
transform 1 0 2850 0 -1 4090
box -12 -8 92 252
use NAND3X1  _2857_
timestamp 1728305047
transform 1 0 2210 0 -1 2650
box -12 -8 112 252
use OR2X2  _2858_
timestamp 1728305284
transform 1 0 2050 0 1 2650
box -12 -8 112 252
use NAND3X1  _2859_
timestamp 1728305047
transform 1 0 1890 0 -1 2650
box -12 -8 112 252
use NOR2X1  _2860_
timestamp 1728305106
transform -1 0 2210 0 -1 3610
box -12 -8 92 252
use NAND2X1  _2861_
timestamp 1728304996
transform 1 0 2130 0 -1 2650
box -12 -8 92 252
use NAND3X1  _2862_
timestamp 1728305047
transform -1 0 2130 0 -1 2650
box -12 -8 112 252
use NAND3X1  _2863_
timestamp 1728305047
transform 1 0 2150 0 1 2650
box -12 -8 112 252
use NAND3X1  _2864_
timestamp 1728305047
transform -1 0 2590 0 1 2650
box -12 -8 112 252
use NAND2X1  _2865_
timestamp 1728304996
transform -1 0 2330 0 1 2650
box -12 -8 92 252
use NAND3X1  _2866_
timestamp 1728305047
transform 1 0 2370 0 1 2650
box -12 -8 112 252
use NAND3X1  _2867_
timestamp 1728305047
transform 1 0 1970 0 1 2170
box -12 -8 112 252
use NAND3X1  _2868_
timestamp 1728305047
transform -1 0 2270 0 1 2170
box -12 -8 112 252
use NAND2X1  _2869_
timestamp 1728304996
transform -1 0 1970 0 1 2170
box -12 -8 92 252
use NAND3X1  _2870_
timestamp 1728305047
transform 1 0 2070 0 1 2170
box -12 -8 112 252
use NAND3X1  _2871_
timestamp 1728305047
transform 1 0 1730 0 1 2650
box -12 -8 112 252
use NAND3X1  _2872_
timestamp 1728305047
transform 1 0 1510 0 1 2650
box -12 -8 112 252
use NAND2X1  _2873_
timestamp 1728304996
transform 1 0 1870 0 1 2650
box -12 -8 92 252
use NAND3X1  _2874_
timestamp 1728305047
transform -1 0 1710 0 1 2650
box -12 -8 112 252
use NAND3X1  _2875_
timestamp 1728305047
transform 1 0 1630 0 1 2170
box -12 -8 112 252
use NAND3X1  _2876_
timestamp 1728305047
transform 1 0 1410 0 1 2170
box -12 -8 112 252
use NAND2X1  _2877_
timestamp 1728304996
transform 1 0 1770 0 1 2170
box -12 -8 92 252
use NAND3X1  _2878_
timestamp 1728305047
transform -1 0 1610 0 1 2170
box -12 -8 112 252
use OAI21X1  _2879_
timestamp 1728305162
transform 1 0 2050 0 1 3130
box -12 -8 112 252
use NOR2X1  _2880_
timestamp 1728305106
transform -1 0 2690 0 -1 2650
box -12 -8 92 252
use AOI21X1  _2881_
timestamp 1728304211
transform 1 0 2350 0 -1 2650
box -12 -8 112 252
use OAI22X1  _2882_
timestamp 1728305200
transform -1 0 2810 0 -1 2650
box -12 -8 132 252
use NOR2X1  _2883_
timestamp 1728305106
transform 1 0 1830 0 1 3610
box -12 -8 92 252
use AOI21X1  _2884_
timestamp 1728304211
transform 1 0 1690 0 -1 3610
box -12 -8 112 252
use OAI22X1  _2885_
timestamp 1728305200
transform 1 0 1690 0 1 3610
box -12 -8 132 252
use INVX1  _2886_
timestamp 1728304789
transform -1 0 1550 0 1 3130
box -12 -8 72 252
use NOR2X1  _2887_
timestamp 1728305106
transform 1 0 1670 0 1 3130
box -12 -8 92 252
use AOI21X1  _2888_
timestamp 1728304211
transform -1 0 1890 0 1 3130
box -12 -8 112 252
use OAI22X1  _2889_
timestamp 1728305200
transform 1 0 1550 0 1 3130
box -12 -8 132 252
use INVX4  _2890_
timestamp 1728304878
transform 1 0 3150 0 1 4090
box -12 -8 92 252
use INVX1  _2891_
timestamp 1728304789
transform 1 0 4210 0 -1 2170
box -12 -8 72 252
use INVX1  _2892_
timestamp 1728304789
transform 1 0 2050 0 1 730
box -12 -8 72 252
use NAND2X1  _2893_
timestamp 1728304996
transform -1 0 2510 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2894_
timestamp 1728305162
transform -1 0 3350 0 -1 1210
box -12 -8 112 252
use AOI21X1  _2895_
timestamp 1728304211
transform 1 0 3710 0 1 1690
box -12 -8 112 252
use MUX2X1  _2896_
timestamp 1728304958
transform -1 0 2230 0 1 1690
box -12 -8 131 252
use MUX2X1  _2897_
timestamp 1728304958
transform 1 0 1490 0 -1 2170
box -12 -8 131 252
use MUX2X1  _2898_
timestamp 1728304958
transform 1 0 2170 0 -1 2170
box -12 -8 131 252
use NAND2X1  _2899_
timestamp 1728304996
transform 1 0 2510 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2900_
timestamp 1728305162
transform 1 0 2490 0 1 1210
box -12 -8 112 252
use AOI22X1  _2901_
timestamp 1728304278
transform -1 0 2570 0 -1 2170
box -14 -8 132 252
use AOI22X1  _2902_
timestamp 1728304278
transform -1 0 4210 0 -1 2170
box -14 -8 132 252
use INVX1  _2903_
timestamp 1728304789
transform 1 0 3990 0 -1 3610
box -12 -8 72 252
use INVX1  _2904_
timestamp 1728304789
transform -1 0 2490 0 1 3130
box -12 -8 72 252
use NAND2X1  _2905_
timestamp 1728304996
transform -1 0 2330 0 1 3130
box -12 -8 92 252
use OAI21X1  _2906_
timestamp 1728305162
transform -1 0 2430 0 1 3130
box -12 -8 112 252
use AOI21X1  _2907_
timestamp 1728304211
transform 1 0 3310 0 1 3610
box -12 -8 112 252
use MUX2X1  _2908_
timestamp 1728304958
transform 1 0 3790 0 1 3130
box -12 -8 131 252
use MUX2X1  _2909_
timestamp 1728304958
transform 1 0 2910 0 1 3130
box -12 -8 131 252
use MUX2X1  _2910_
timestamp 1728304958
transform -1 0 3790 0 1 3130
box -12 -8 131 252
use NAND2X1  _2911_
timestamp 1728304996
transform 1 0 3510 0 -1 3610
box -12 -8 92 252
use OAI21X1  _2912_
timestamp 1728305162
transform 1 0 3370 0 -1 3610
box -12 -8 112 252
use AOI22X1  _2913_
timestamp 1728304278
transform 1 0 3610 0 -1 3610
box -14 -8 132 252
use AOI22X1  _2914_
timestamp 1728304278
transform -1 0 3850 0 -1 3610
box -14 -8 132 252
use INVX1  _2915_
timestamp 1728304789
transform -1 0 4530 0 -1 2170
box -12 -8 72 252
use INVX1  _2916_
timestamp 1728304789
transform 1 0 790 0 1 1210
box -12 -8 72 252
use NAND2X1  _2917_
timestamp 1728304996
transform -1 0 750 0 -1 1690
box -12 -8 92 252
use OAI21X1  _2918_
timestamp 1728305162
transform -1 0 890 0 -1 1690
box -12 -8 112 252
use AOI21X1  _2919_
timestamp 1728304211
transform 1 0 3910 0 1 1690
box -12 -8 112 252
use MUX2X1  _2920_
timestamp 1728304958
transform 1 0 3410 0 -1 1690
box -12 -8 131 252
use MUX2X1  _2921_
timestamp 1728304958
transform -1 0 2490 0 1 1690
box -12 -8 131 252
use MUX2X1  _2922_
timestamp 1728304958
transform 1 0 3590 0 1 1690
box -12 -8 131 252
use NAND2X1  _2923_
timestamp 1728304996
transform -1 0 3430 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2924_
timestamp 1728305162
transform 1 0 3370 0 1 1210
box -12 -8 112 252
use AOI22X1  _2925_
timestamp 1728304278
transform 1 0 3870 0 -1 2170
box -14 -8 132 252
use AOI22X1  _2926_
timestamp 1728304278
transform -1 0 4430 0 -1 2170
box -14 -8 132 252
use INVX1  _2927_
timestamp 1728304789
transform -1 0 4350 0 -1 3130
box -12 -8 72 252
use INVX1  _2928_
timestamp 1728304789
transform -1 0 710 0 1 250
box -12 -8 72 252
use NAND2X1  _2929_
timestamp 1728304996
transform -1 0 750 0 -1 730
box -12 -8 92 252
use OAI21X1  _2930_
timestamp 1728305162
transform 1 0 790 0 -1 730
box -12 -8 112 252
use AOI21X1  _2931_
timestamp 1728304211
transform 1 0 3810 0 1 1690
box -12 -8 112 252
use MUX2X1  _2932_
timestamp 1728304958
transform 1 0 1050 0 1 2170
box -12 -8 131 252
use MUX2X1  _2933_
timestamp 1728304958
transform 1 0 1070 0 -1 2650
box -12 -8 131 252
use MUX2X1  _2934_
timestamp 1728304958
transform 1 0 1210 0 -1 2650
box -12 -8 131 252
use NAND2X1  _2935_
timestamp 1728304996
transform -1 0 1490 0 1 730
box -12 -8 92 252
use OAI21X1  _2936_
timestamp 1728305162
transform 1 0 1670 0 -1 1210
box -12 -8 112 252
use AOI22X1  _2937_
timestamp 1728304278
transform -1 0 2610 0 -1 2650
box -14 -8 132 252
use AOI22X1  _2938_
timestamp 1728304278
transform -1 0 4190 0 -1 3130
box -14 -8 132 252
use INVX1  _2939_
timestamp 1728304789
transform -1 0 3650 0 -1 2650
box -12 -8 72 252
use INVX1  _2940_
timestamp 1728304789
transform 1 0 1310 0 -1 730
box -12 -8 72 252
use NAND2X1  _2941_
timestamp 1728304996
transform -1 0 1310 0 -1 730
box -12 -8 92 252
use OAI21X1  _2942_
timestamp 1728305162
transform 1 0 1370 0 -1 730
box -12 -8 112 252
use AOI21X1  _2943_
timestamp 1728304211
transform 1 0 3350 0 -1 2650
box -12 -8 112 252
use MUX2X1  _2944_
timestamp 1728304958
transform 1 0 810 0 1 1690
box -12 -8 131 252
use MUX2X1  _2945_
timestamp 1728304958
transform 1 0 1310 0 1 1690
box -12 -8 131 252
use MUX2X1  _2946_
timestamp 1728304958
transform 1 0 1430 0 1 1690
box -12 -8 131 252
use NAND2X1  _2947_
timestamp 1728304996
transform 1 0 1990 0 -1 1210
box -12 -8 92 252
use OAI21X1  _2948_
timestamp 1728305162
transform 1 0 1950 0 1 1210
box -12 -8 112 252
use AOI22X1  _2949_
timestamp 1728304278
transform -1 0 2450 0 -1 2170
box -14 -8 132 252
use AOI22X1  _2950_
timestamp 1728304278
transform -1 0 3570 0 -1 2650
box -14 -8 132 252
use INVX1  _2951_
timestamp 1728304789
transform -1 0 4190 0 -1 2650
box -12 -8 72 252
use INVX1  _2952_
timestamp 1728304789
transform 1 0 2190 0 1 250
box -12 -8 72 252
use NAND2X1  _2953_
timestamp 1728304996
transform -1 0 2530 0 1 250
box -12 -8 92 252
use OAI21X1  _2954_
timestamp 1728305162
transform 1 0 2550 0 1 250
box -12 -8 112 252
use AOI21X1  _2955_
timestamp 1728304211
transform 1 0 3990 0 -1 2170
box -12 -8 112 252
use MUX2X1  _2956_
timestamp 1728304958
transform 1 0 3490 0 -1 2170
box -12 -8 131 252
use MUX2X1  _2957_
timestamp 1728304958
transform 1 0 3490 0 1 2650
box -12 -8 131 252
use MUX2X1  _2958_
timestamp 1728304958
transform 1 0 3630 0 -1 2170
box -12 -8 131 252
use NAND2X1  _2959_
timestamp 1728304996
transform -1 0 3030 0 1 730
box -12 -8 92 252
use OAI21X1  _2960_
timestamp 1728305162
transform 1 0 3470 0 -1 1210
box -12 -8 112 252
use AOI22X1  _2961_
timestamp 1728304278
transform -1 0 3870 0 -1 2170
box -14 -8 132 252
use AOI22X1  _2962_
timestamp 1728304278
transform -1 0 4190 0 1 2170
box -14 -8 132 252
use INVX1  _2963_
timestamp 1728304789
transform -1 0 2670 0 -1 4570
box -12 -8 72 252
use INVX1  _2964_
timestamp 1728304789
transform 1 0 770 0 1 4570
box -12 -8 72 252
use NAND2X1  _2965_
timestamp 1728304996
transform 1 0 890 0 -1 4570
box -12 -8 92 252
use OAI21X1  _2966_
timestamp 1728305162
transform 1 0 850 0 1 4570
box -12 -8 112 252
use AOI21X1  _2967_
timestamp 1728304211
transform 1 0 2390 0 1 4570
box -12 -8 112 252
use MUX2X1  _2968_
timestamp 1728304958
transform -1 0 790 0 1 4090
box -12 -8 131 252
use MUX2X1  _2969_
timestamp 1728304958
transform 1 0 970 0 -1 4090
box -12 -8 131 252
use MUX2X1  _2970_
timestamp 1728304958
transform -1 0 1150 0 1 4090
box -12 -8 131 252
use NAND2X1  _2971_
timestamp 1728304996
transform -1 0 2150 0 1 4570
box -12 -8 92 252
use OAI21X1  _2972_
timestamp 1728305162
transform 1 0 2150 0 1 4570
box -12 -8 112 252
use AOI22X1  _2973_
timestamp 1728304278
transform -1 0 2390 0 -1 4570
box -14 -8 132 252
use AOI22X1  _2974_
timestamp 1728304278
transform -1 0 2610 0 -1 4570
box -14 -8 132 252
use INVX1  _2975_
timestamp 1728304789
transform -1 0 2070 0 -1 5050
box -12 -8 72 252
use INVX1  _2976_
timestamp 1728304789
transform 1 0 950 0 1 4570
box -12 -8 72 252
use NAND2X1  _2977_
timestamp 1728304996
transform -1 0 1110 0 1 4570
box -12 -8 92 252
use OAI21X1  _2978_
timestamp 1728305162
transform 1 0 1110 0 1 4570
box -12 -8 112 252
use AOI21X1  _2979_
timestamp 1728304211
transform 1 0 2290 0 1 4570
box -12 -8 112 252
use MUX2X1  _2980_
timestamp 1728304958
transform 1 0 790 0 1 4090
box -12 -8 131 252
use MUX2X1  _2981_
timestamp 1728304958
transform -1 0 1670 0 1 3610
box -12 -8 131 252
use MUX2X1  _2982_
timestamp 1728304958
transform 1 0 1150 0 1 4090
box -12 -8 131 252
use NAND2X1  _2983_
timestamp 1728304996
transform -1 0 2030 0 -1 4570
box -12 -8 92 252
use OAI21X1  _2984_
timestamp 1728305162
transform 1 0 2030 0 -1 4570
box -12 -8 112 252
use AOI22X1  _2985_
timestamp 1728304278
transform -1 0 2250 0 -1 4570
box -14 -8 132 252
use AOI22X1  _2986_
timestamp 1728304278
transform 1 0 2110 0 -1 5050
box -14 -8 132 252
use INVX1  _2987_
timestamp 1728304789
transform 1 0 1850 0 -1 2170
box -12 -8 72 252
use OAI22X1  _2988_
timestamp 1728305200
transform 1 0 2390 0 -1 4090
box -12 -8 132 252
use NAND2X1  _2989_
timestamp 1728304996
transform -1 0 3170 0 -1 4090
box -12 -8 92 252
use NOR2X1  _2990_
timestamp 1728305106
transform -1 0 1730 0 -1 2170
box -12 -8 92 252
use NOR2X1  _2991_
timestamp 1728305106
transform -1 0 2030 0 -1 4090
box -12 -8 92 252
use OAI21X1  _2992_
timestamp 1728305162
transform 1 0 1390 0 -1 2170
box -12 -8 112 252
use OAI22X1  _2993_
timestamp 1728305200
transform -1 0 1850 0 -1 2170
box -12 -8 132 252
use INVX1  _2994_
timestamp 1728304789
transform 1 0 3770 0 -1 3130
box -12 -8 72 252
use NOR2X1  _2995_
timestamp 1728305106
transform -1 0 3610 0 -1 3130
box -12 -8 92 252
use OAI21X1  _2996_
timestamp 1728305162
transform 1 0 3330 0 -1 3130
box -12 -8 112 252
use OAI22X1  _2997_
timestamp 1728305200
transform -1 0 3730 0 -1 3130
box -12 -8 132 252
use INVX1  _2998_
timestamp 1728304789
transform 1 0 3990 0 1 2170
box -12 -8 72 252
use NOR2X1  _2999_
timestamp 1728305106
transform 1 0 3510 0 1 2170
box -12 -8 92 252
use OAI21X1  _3000_
timestamp 1728305162
transform 1 0 3230 0 -1 2650
box -12 -8 112 252
use OAI22X1  _3001_
timestamp 1728305200
transform -1 0 3950 0 1 2170
box -12 -8 132 252
use INVX1  _3002_
timestamp 1728304789
transform 1 0 270 0 1 2170
box -12 -8 72 252
use NOR2X1  _3003_
timestamp 1728305106
transform 1 0 430 0 -1 2170
box -12 -8 92 252
use OAI21X1  _3004_
timestamp 1728305162
transform -1 0 590 0 1 2170
box -12 -8 112 252
use OAI22X1  _3005_
timestamp 1728305200
transform 1 0 370 0 1 2170
box -12 -8 132 252
use INVX1  _3006_
timestamp 1728304789
transform -1 0 710 0 1 1690
box -12 -8 72 252
use NOR2X1  _3007_
timestamp 1728305106
transform 1 0 730 0 1 1690
box -12 -8 92 252
use OAI21X1  _3008_
timestamp 1728305162
transform -1 0 410 0 -1 2170
box -12 -8 112 252
use OAI22X1  _3009_
timestamp 1728305200
transform -1 0 650 0 1 1690
box -12 -8 132 252
use INVX1  _3010_
timestamp 1728304789
transform 1 0 3450 0 1 2170
box -12 -8 72 252
use NOR2X1  _3011_
timestamp 1728305106
transform 1 0 3210 0 1 2170
box -12 -8 92 252
use OAI21X1  _3012_
timestamp 1728305162
transform 1 0 3090 0 1 2170
box -12 -8 112 252
use OAI22X1  _3013_
timestamp 1728305200
transform -1 0 3450 0 1 2170
box -12 -8 132 252
use INVX1  _3014_
timestamp 1728304789
transform 1 0 650 0 -1 4090
box -12 -8 72 252
use NOR2X1  _3015_
timestamp 1728305106
transform 1 0 770 0 1 3610
box -12 -8 92 252
use OAI21X1  _3016_
timestamp 1728305162
transform 1 0 490 0 1 3610
box -12 -8 112 252
use OAI22X1  _3017_
timestamp 1728305200
transform 1 0 630 0 1 3610
box -12 -8 132 252
use INVX1  _3018_
timestamp 1728304789
transform 1 0 250 0 -1 4090
box -12 -8 72 252
use NOR2X1  _3019_
timestamp 1728305106
transform 1 0 570 0 -1 4090
box -12 -8 92 252
use OAI21X1  _3020_
timestamp 1728305162
transform 1 0 470 0 -1 4090
box -12 -8 112 252
use OAI22X1  _3021_
timestamp 1728305200
transform 1 0 310 0 -1 4090
box -12 -8 132 252
use DFFPOSX1  _3022_
timestamp 1728340458
transform 1 0 10 0 1 1690
box -13 -8 253 252
use DFFPOSX1  _3023_
timestamp 1728340458
transform 1 0 1530 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _3024_
timestamp 1728340458
transform -1 0 3090 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _3025_
timestamp 1728340458
transform 1 0 510 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _3026_
timestamp 1728340458
transform 1 0 1130 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _3027_
timestamp 1728340458
transform 1 0 3150 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _3028_
timestamp 1728340458
transform 1 0 10 0 -1 3610
box -13 -8 253 252
use DFFPOSX1  _3029_
timestamp 1728340458
transform 1 0 1450 0 -1 3610
box -13 -8 253 252
use DFFPOSX1  _3030_
timestamp 1728340458
transform -1 0 1310 0 -1 1690
box -13 -8 253 252
use DFFPOSX1  _3031_
timestamp 1728340458
transform -1 0 2650 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _3032_
timestamp 1728340458
transform 1 0 2910 0 1 1690
box -13 -8 253 252
use DFFPOSX1  _3033_
timestamp 1728340458
transform -1 0 1070 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _3034_
timestamp 1728340458
transform 1 0 10 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _3035_
timestamp 1728340458
transform 1 0 2990 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _3036_
timestamp 1728340458
transform 1 0 10 0 1 3610
box -13 -8 253 252
use DFFPOSX1  _3037_
timestamp 1728340458
transform -1 0 1290 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _3038_
timestamp 1728340458
transform 1 0 2230 0 1 730
box -13 -8 253 252
use DFFPOSX1  _3039_
timestamp 1728340458
transform 1 0 3030 0 -1 3610
box -13 -8 253 252
use DFFPOSX1  _3040_
timestamp 1728340458
transform -1 0 3790 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _3041_
timestamp 1728340458
transform 1 0 1110 0 -1 1210
box -13 -8 253 252
use DFFPOSX1  _3042_
timestamp 1728340458
transform -1 0 1630 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _3043_
timestamp 1728340458
transform -1 0 3090 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _3044_
timestamp 1728340458
transform 1 0 1670 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _3045_
timestamp 1728340458
transform -1 0 2030 0 1 4570
box -13 -8 253 252
use DFFPOSX1  _3046_
timestamp 1728340458
transform 1 0 2350 0 -1 730
box -13 -8 253 252
use DFFPOSX1  _3047_
timestamp 1728340458
transform -1 0 4290 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _3048_
timestamp 1728340458
transform 1 0 3050 0 -1 730
box -13 -8 253 252
use DFFPOSX1  _3049_
timestamp 1728340458
transform 1 0 1070 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3050_
timestamp 1728340458
transform 1 0 1830 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3051_
timestamp 1728340458
transform 1 0 2610 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3052_
timestamp 1728340458
transform 1 0 1290 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _3053_
timestamp 1728340458
transform 1 0 1430 0 1 4570
box -13 -8 253 252
use DFFPOSX1  _3054_
timestamp 1728340458
transform 1 0 1790 0 -1 730
box -13 -8 253 252
use DFFPOSX1  _3055_
timestamp 1728340458
transform 1 0 2170 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _3056_
timestamp 1728340458
transform 1 0 10 0 1 730
box -13 -8 253 252
use DFFPOSX1  _3057_
timestamp 1728340458
transform 1 0 590 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3058_
timestamp 1728340458
transform 1 0 10 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3059_
timestamp 1728340458
transform -1 0 2410 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3060_
timestamp 1728340458
transform 1 0 250 0 1 4570
box -13 -8 253 252
use DFFPOSX1  _3061_
timestamp 1728340458
transform 1 0 650 0 -1 5050
box -13 -8 253 252
use DFFPOSX1  _3062_
timestamp 1728340458
transform 1 0 1930 0 -1 1690
box -13 -8 253 252
use DFFPOSX1  _3063_
timestamp 1728340458
transform -1 0 4150 0 1 3130
box -13 -8 253 252
use DFFPOSX1  _3064_
timestamp 1728340458
transform -1 0 3770 0 -1 1690
box -13 -8 253 252
use DFFPOSX1  _3065_
timestamp 1728340458
transform 1 0 590 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _3066_
timestamp 1728340458
transform 1 0 250 0 1 1690
box -13 -8 253 252
use DFFPOSX1  _3067_
timestamp 1728340458
transform 1 0 2730 0 -1 1690
box -13 -8 253 252
use DFFPOSX1  _3068_
timestamp 1728340458
transform 1 0 10 0 1 4570
box -13 -8 253 252
use DFFPOSX1  _3069_
timestamp 1728340458
transform 1 0 490 0 1 4570
box -13 -8 253 252
use DFFPOSX1  _3070_
timestamp 1728340458
transform 1 0 790 0 1 730
box -13 -8 253 252
use DFFPOSX1  _3071_
timestamp 1728340458
transform 1 0 550 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _3072_
timestamp 1728340458
transform 1 0 250 0 1 1210
box -13 -8 253 252
use DFFPOSX1  _3073_
timestamp 1728340458
transform 1 0 10 0 -1 730
box -13 -8 253 252
use DFFPOSX1  _3074_
timestamp 1728340458
transform 1 0 830 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3075_
timestamp 1728340458
transform 1 0 1530 0 -1 250
box -13 -8 253 252
use DFFPOSX1  _3076_
timestamp 1728340458
transform 1 0 10 0 1 3130
box -13 -8 253 252
use DFFPOSX1  _3077_
timestamp 1728340458
transform 1 0 870 0 -1 3610
box -13 -8 253 252
use DFFPOSX1  _3078_
timestamp 1728340458
transform -1 0 1890 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _3079_
timestamp 1728340458
transform 1 0 2590 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _3080_
timestamp 1728340458
transform -1 0 2510 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _3081_
timestamp 1728340458
transform -1 0 1650 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _3082_
timestamp 1728340458
transform -1 0 1410 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _3083_
timestamp 1728340458
transform 1 0 2910 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _3084_
timestamp 1728340458
transform -1 0 1650 0 -1 4090
box -13 -8 253 252
use DFFPOSX1  _3085_
timestamp 1728340458
transform 1 0 1110 0 1 3130
box -13 -8 253 252
use DFFPOSX1  _3086_
timestamp 1728340458
transform 1 0 3890 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _3087_
timestamp 1728340458
transform 1 0 3410 0 1 3610
box -13 -8 253 252
use DFFPOSX1  _3088_
timestamp 1728340458
transform 1 0 4430 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _3089_
timestamp 1728340458
transform 1 0 4350 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _3090_
timestamp 1728340458
transform 1 0 3650 0 -1 2650
box -13 -8 253 252
use DFFPOSX1  _3091_
timestamp 1728340458
transform -1 0 4530 0 1 2650
box -13 -8 253 252
use DFFPOSX1  _3092_
timestamp 1728340458
transform 1 0 2490 0 1 4570
box -13 -8 253 252
use DFFPOSX1  _3093_
timestamp 1728340458
transform 1 0 1870 0 1 5050
box -13 -8 253 252
use DFFPOSX1  _3094_
timestamp 1728340458
transform 1 0 1910 0 -1 2170
box -13 -8 253 252
use DFFPOSX1  _3095_
timestamp 1728340458
transform -1 0 4070 0 -1 3130
box -13 -8 253 252
use DFFPOSX1  _3096_
timestamp 1728340458
transform -1 0 4430 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _3097_
timestamp 1728340458
transform 1 0 10 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _3098_
timestamp 1728340458
transform 1 0 430 0 -1 1690
box -13 -8 253 252
use DFFPOSX1  _3099_
timestamp 1728340458
transform -1 0 3830 0 1 2170
box -13 -8 253 252
use DFFPOSX1  _3100_
timestamp 1728340458
transform 1 0 250 0 1 3610
box -13 -8 253 252
use DFFPOSX1  _3101_
timestamp 1728340458
transform 1 0 10 0 -1 4090
box -13 -8 253 252
use BUFX2  _3102_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304320
transform -1 0 110 0 1 6010
box -12 -8 92 252
use BUFX2  _3103_
timestamp 1728304320
transform 1 0 3910 0 -1 730
box -12 -8 92 252
use BUFX2  _3104_
timestamp 1728304320
transform -1 0 3530 0 1 250
box -12 -8 92 252
use BUFX2  _3105_
timestamp 1728304320
transform -1 0 3610 0 1 250
box -12 -8 92 252
use BUFX2  _3106_
timestamp 1728304320
transform -1 0 3870 0 -1 250
box -12 -8 92 252
use BUFX2  _3107_
timestamp 1728304320
transform -1 0 4430 0 -1 250
box -12 -8 92 252
use BUFX2  _3108_
timestamp 1728304320
transform -1 0 3710 0 -1 250
box -12 -8 92 252
use BUFX2  _3109_
timestamp 1728304320
transform -1 0 4730 0 -1 250
box -12 -8 92 252
use BUFX2  _3110_
timestamp 1728304320
transform 1 0 4990 0 -1 250
box -12 -8 92 252
use BUFX2  BUFX2_insert13
timestamp 1728304320
transform 1 0 6850 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert14
timestamp 1728304320
transform -1 0 5950 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert15
timestamp 1728304320
transform 1 0 5470 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert16
timestamp 1728304320
transform 1 0 6870 0 1 730
box -12 -8 92 252
use BUFX2  BUFX2_insert17
timestamp 1728304320
transform -1 0 6150 0 1 730
box -12 -8 92 252
use BUFX2  BUFX2_insert18
timestamp 1728304320
transform 1 0 5770 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert19
timestamp 1728304320
transform -1 0 4850 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert20
timestamp 1728304320
transform -1 0 4130 0 1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert21
timestamp 1728304320
transform 1 0 5670 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert22
timestamp 1728304320
transform 1 0 1930 0 1 3610
box -12 -8 92 252
use BUFX2  BUFX2_insert23
timestamp 1728304320
transform -1 0 2130 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert24
timestamp 1728304320
transform -1 0 1030 0 1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert25
timestamp 1728304320
transform 1 0 3470 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert26
timestamp 1728304320
transform 1 0 1330 0 -1 2650
box -12 -8 92 252
use BUFX2  BUFX2_insert27
timestamp 1728304320
transform 1 0 3490 0 -1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert28
timestamp 1728304320
transform 1 0 2230 0 1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert29
timestamp 1728304320
transform 1 0 110 0 -1 6010
box -12 -8 92 252
use BUFX2  BUFX2_insert30
timestamp 1728304320
transform -1 0 530 0 -1 5530
box -12 -8 92 252
use BUFX2  BUFX2_insert31
timestamp 1728304320
transform -1 0 130 0 1 5050
box -12 -8 92 252
use BUFX2  BUFX2_insert32
timestamp 1728304320
transform -1 0 90 0 -1 6010
box -12 -8 92 252
use BUFX2  BUFX2_insert33
timestamp 1728304320
transform 1 0 5350 0 -1 2170
box -12 -8 92 252
use BUFX2  BUFX2_insert34
timestamp 1728304320
transform 1 0 6770 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert35
timestamp 1728304320
transform -1 0 6410 0 -1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert36
timestamp 1728304320
transform -1 0 4390 0 1 1690
box -12 -8 92 252
use BUFX2  BUFX2_insert37
timestamp 1728304320
transform 1 0 2650 0 1 3130
box -12 -8 92 252
use BUFX2  BUFX2_insert38
timestamp 1728304320
transform -1 0 1810 0 -1 4090
box -12 -8 92 252
use BUFX2  BUFX2_insert39
timestamp 1728304320
transform -1 0 1270 0 1 1210
box -12 -8 92 252
use BUFX2  BUFX2_insert40
timestamp 1728304320
transform 1 0 1190 0 1 730
box -12 -8 92 252
use BUFX2  BUFX2_insert41
timestamp 1728304320
transform 1 0 2610 0 1 730
box -12 -8 92 252
use CLKBUF1  CLKBUF1_insert0 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728304421
transform 1 0 10 0 -1 1210
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert1
timestamp 1728304421
transform -1 0 4230 0 1 1210
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert2
timestamp 1728304421
transform -1 0 4090 0 -1 1690
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert3
timestamp 1728304421
transform 1 0 6350 0 1 2650
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert4
timestamp 1728304421
transform -1 0 2930 0 1 6010
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert5
timestamp 1728304421
transform -1 0 4550 0 1 6010
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert6
timestamp 1728304421
transform 1 0 4390 0 1 3130
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert7
timestamp 1728304421
transform -1 0 650 0 1 5050
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert8
timestamp 1728304421
transform -1 0 4850 0 1 730
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert9
timestamp 1728304421
transform 1 0 4850 0 1 730
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert10
timestamp 1728304421
transform -1 0 510 0 -1 2650
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert11
timestamp 1728304421
transform -1 0 4490 0 -1 4090
box -12 -8 212 252
use CLKBUF1  CLKBUF1_insert12
timestamp 1728304421
transform 1 0 450 0 -1 5050
box -12 -8 212 252
use FILL  FILL117750x43350 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1728341909
transform -1 0 7870 0 -1 3130
box -12 -8 32 252
use FILL  FILL117750x54150
timestamp 1728341909
transform 1 0 7850 0 1 3610
box -12 -8 32 252
use FILL  FILL118050x3750
timestamp 1728341909
transform 1 0 7870 0 1 250
box -12 -8 32 252
use FILL  FILL118050x39750
timestamp 1728341909
transform 1 0 7870 0 1 2650
box -12 -8 32 252
use FILL  FILL118050x43350
timestamp 1728341909
transform -1 0 7890 0 -1 3130
box -12 -8 32 252
use FILL  FILL118050x54150
timestamp 1728341909
transform 1 0 7870 0 1 3610
box -12 -8 32 252
use FILL  FILL118050x57750
timestamp 1728341909
transform -1 0 7890 0 -1 4090
box -12 -8 32 252
use FILL  FILL118350x150
timestamp 1728341909
transform -1 0 7910 0 -1 250
box -12 -8 32 252
use FILL  FILL118350x3750
timestamp 1728341909
transform 1 0 7890 0 1 250
box -12 -8 32 252
use FILL  FILL118350x32550
timestamp 1728341909
transform 1 0 7890 0 1 2170
box -12 -8 32 252
use FILL  FILL118350x36150
timestamp 1728341909
transform -1 0 7910 0 -1 2650
box -12 -8 32 252
use FILL  FILL118350x39750
timestamp 1728341909
transform 1 0 7890 0 1 2650
box -12 -8 32 252
use FILL  FILL118350x43350
timestamp 1728341909
transform -1 0 7910 0 -1 3130
box -12 -8 32 252
use FILL  FILL118350x54150
timestamp 1728341909
transform 1 0 7890 0 1 3610
box -12 -8 32 252
use FILL  FILL118350x57750
timestamp 1728341909
transform -1 0 7910 0 -1 4090
box -12 -8 32 252
use FILL  FILL118350x64950
timestamp 1728341909
transform -1 0 7910 0 -1 4570
box -12 -8 32 252
use FILL  FILL118350x68550
timestamp 1728341909
transform 1 0 7890 0 1 4570
box -12 -8 32 252
use FILL  FILL118350x75750
timestamp 1728341909
transform 1 0 7890 0 1 5050
box -12 -8 32 252
use FILL  FILL118350x82950
timestamp 1728341909
transform 1 0 7890 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1434_
timestamp 1728341909
transform -1 0 4550 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1436_
timestamp 1728341909
transform -1 0 4270 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1438_
timestamp 1728341909
transform 1 0 4090 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1440_
timestamp 1728341909
transform -1 0 4490 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1443_
timestamp 1728341909
transform 1 0 4250 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1445_
timestamp 1728341909
transform 1 0 5070 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1447_
timestamp 1728341909
transform -1 0 5170 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1449_
timestamp 1728341909
transform -1 0 4890 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1451_
timestamp 1728341909
transform -1 0 4750 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1453_
timestamp 1728341909
transform -1 0 3870 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1455_
timestamp 1728341909
transform -1 0 3990 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1457_
timestamp 1728341909
transform 1 0 4150 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1459_
timestamp 1728341909
transform -1 0 4450 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1460_
timestamp 1728341909
transform 1 0 4490 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1462_
timestamp 1728341909
transform 1 0 3970 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1464_
timestamp 1728341909
transform -1 0 4670 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1466_
timestamp 1728341909
transform -1 0 3870 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1468_
timestamp 1728341909
transform -1 0 3630 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1470_
timestamp 1728341909
transform -1 0 3890 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1472_
timestamp 1728341909
transform 1 0 4430 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1474_
timestamp 1728341909
transform -1 0 4230 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1477_
timestamp 1728341909
transform 1 0 5170 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1479_
timestamp 1728341909
transform 1 0 4190 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1481_
timestamp 1728341909
transform 1 0 4730 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1483_
timestamp 1728341909
transform -1 0 4530 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1485_
timestamp 1728341909
transform -1 0 2850 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1487_
timestamp 1728341909
transform 1 0 2850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1489_
timestamp 1728341909
transform 1 0 3350 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1491_
timestamp 1728341909
transform 1 0 2770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1493_
timestamp 1728341909
transform 1 0 3050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1494_
timestamp 1728341909
transform 1 0 3250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1496_
timestamp 1728341909
transform 1 0 3330 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1498_
timestamp 1728341909
transform 1 0 2950 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1500_
timestamp 1728341909
transform -1 0 30 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1502_
timestamp 1728341909
transform 1 0 130 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1504_
timestamp 1728341909
transform -1 0 30 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1506_
timestamp 1728341909
transform -1 0 210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1508_
timestamp 1728341909
transform 1 0 270 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1511_
timestamp 1728341909
transform -1 0 110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1513_
timestamp 1728341909
transform -1 0 330 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1515_
timestamp 1728341909
transform -1 0 230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1517_
timestamp 1728341909
transform -1 0 110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1519_
timestamp 1728341909
transform -1 0 130 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1521_
timestamp 1728341909
transform -1 0 270 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1523_
timestamp 1728341909
transform 1 0 330 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1526_
timestamp 1728341909
transform 1 0 1430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1528_
timestamp 1728341909
transform -1 0 970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1530_
timestamp 1728341909
transform 1 0 530 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1532_
timestamp 1728341909
transform -1 0 830 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1534_
timestamp 1728341909
transform 1 0 1350 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1536_
timestamp 1728341909
transform -1 0 1070 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1538_
timestamp 1728341909
transform -1 0 1130 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1540_
timestamp 1728341909
transform 1 0 2050 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1542_
timestamp 1728341909
transform -1 0 1950 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1543_
timestamp 1728341909
transform -1 0 1810 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1545_
timestamp 1728341909
transform -1 0 1170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1547_
timestamp 1728341909
transform -1 0 1490 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1549_
timestamp 1728341909
transform 1 0 1570 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1551_
timestamp 1728341909
transform -1 0 3650 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1553_
timestamp 1728341909
transform -1 0 1150 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1555_
timestamp 1728341909
transform 1 0 1230 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1572_
timestamp 1728341909
transform -1 0 3790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1575_
timestamp 1728341909
transform 1 0 3850 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1577_
timestamp 1728341909
transform -1 0 3490 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1579_
timestamp 1728341909
transform -1 0 3330 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1581_
timestamp 1728341909
transform -1 0 3310 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1583_
timestamp 1728341909
transform -1 0 3290 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1585_
timestamp 1728341909
transform 1 0 4530 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1587_
timestamp 1728341909
transform 1 0 4770 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1589_
timestamp 1728341909
transform -1 0 4230 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1591_
timestamp 1728341909
transform 1 0 5510 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1592_
timestamp 1728341909
transform 1 0 5750 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1594_
timestamp 1728341909
transform 1 0 4650 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1596_
timestamp 1728341909
transform -1 0 4870 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1598_
timestamp 1728341909
transform 1 0 6010 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__1600_
timestamp 1728341909
transform 1 0 5070 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1602_
timestamp 1728341909
transform -1 0 5370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1604_
timestamp 1728341909
transform 1 0 4670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__1606_
timestamp 1728341909
transform -1 0 4890 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1609_
timestamp 1728341909
transform -1 0 6510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1611_
timestamp 1728341909
transform 1 0 7070 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1613_
timestamp 1728341909
transform 1 0 7290 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1615_
timestamp 1728341909
transform -1 0 6610 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1617_
timestamp 1728341909
transform -1 0 6810 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1619_
timestamp 1728341909
transform -1 0 6630 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1621_
timestamp 1728341909
transform -1 0 4790 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1623_
timestamp 1728341909
transform -1 0 5010 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1625_
timestamp 1728341909
transform 1 0 6090 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1626_
timestamp 1728341909
transform -1 0 6010 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1628_
timestamp 1728341909
transform 1 0 6470 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1630_
timestamp 1728341909
transform 1 0 5290 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1632_
timestamp 1728341909
transform -1 0 5550 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1634_
timestamp 1728341909
transform 1 0 3810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1636_
timestamp 1728341909
transform 1 0 1210 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1638_
timestamp 1728341909
transform 1 0 3790 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1640_
timestamp 1728341909
transform 1 0 3630 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1643_
timestamp 1728341909
transform -1 0 3510 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1645_
timestamp 1728341909
transform -1 0 2930 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1647_
timestamp 1728341909
transform -1 0 3190 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1649_
timestamp 1728341909
transform -1 0 2910 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1651_
timestamp 1728341909
transform -1 0 4410 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__1653_
timestamp 1728341909
transform -1 0 5570 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1655_
timestamp 1728341909
transform -1 0 5530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__1658_
timestamp 1728341909
transform -1 0 5010 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1660_
timestamp 1728341909
transform -1 0 7190 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__1662_
timestamp 1728341909
transform 1 0 6470 0 1 250
box -12 -8 32 252
use FILL  FILL_0__1664_
timestamp 1728341909
transform -1 0 5690 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__1666_
timestamp 1728341909
transform -1 0 5410 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1668_
timestamp 1728341909
transform -1 0 3910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1670_
timestamp 1728341909
transform 1 0 3450 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__1672_
timestamp 1728341909
transform -1 0 3870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1674_
timestamp 1728341909
transform 1 0 1470 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1675_
timestamp 1728341909
transform -1 0 1370 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1705_
timestamp 1728341909
transform 1 0 4050 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1707_
timestamp 1728341909
transform -1 0 3470 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1709_
timestamp 1728341909
transform -1 0 3490 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1711_
timestamp 1728341909
transform -1 0 3250 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1713_
timestamp 1728341909
transform 1 0 3930 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1715_
timestamp 1728341909
transform 1 0 3570 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1717_
timestamp 1728341909
transform 1 0 3690 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1720_
timestamp 1728341909
transform 1 0 3830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1722_
timestamp 1728341909
transform -1 0 3630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1724_
timestamp 1728341909
transform 1 0 3590 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1730_
timestamp 1728341909
transform 1 0 2210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1732_
timestamp 1728341909
transform 1 0 2090 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1734_
timestamp 1728341909
transform 1 0 2290 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1736_
timestamp 1728341909
transform 1 0 2210 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__1740_
timestamp 1728341909
transform -1 0 4910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1742_
timestamp 1728341909
transform 1 0 3830 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1743_
timestamp 1728341909
transform -1 0 4650 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1745_
timestamp 1728341909
transform -1 0 4210 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1747_
timestamp 1728341909
transform -1 0 4290 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1749_
timestamp 1728341909
transform -1 0 4350 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1751_
timestamp 1728341909
transform -1 0 4070 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__1753_
timestamp 1728341909
transform -1 0 4190 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1755_
timestamp 1728341909
transform -1 0 3890 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1757_
timestamp 1728341909
transform -1 0 3750 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1760_
timestamp 1728341909
transform -1 0 4510 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1762_
timestamp 1728341909
transform -1 0 4070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1764_
timestamp 1728341909
transform -1 0 4730 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1766_
timestamp 1728341909
transform -1 0 4730 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1768_
timestamp 1728341909
transform 1 0 4590 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1770_
timestamp 1728341909
transform -1 0 4730 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1772_
timestamp 1728341909
transform -1 0 4210 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1774_
timestamp 1728341909
transform 1 0 4190 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1776_
timestamp 1728341909
transform -1 0 3810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__1777_
timestamp 1728341909
transform -1 0 3330 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__1779_
timestamp 1728341909
transform 1 0 4030 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1781_
timestamp 1728341909
transform -1 0 3690 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__1783_
timestamp 1728341909
transform -1 0 4890 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1785_
timestamp 1728341909
transform -1 0 4290 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__1787_
timestamp 1728341909
transform -1 0 4650 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1789_
timestamp 1728341909
transform -1 0 5150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1791_
timestamp 1728341909
transform 1 0 4990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1794_
timestamp 1728341909
transform 1 0 5230 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1796_
timestamp 1728341909
transform -1 0 5610 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1798_
timestamp 1728341909
transform 1 0 5270 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1800_
timestamp 1728341909
transform 1 0 5070 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1802_
timestamp 1728341909
transform 1 0 6030 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1804_
timestamp 1728341909
transform 1 0 6270 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1806_
timestamp 1728341909
transform -1 0 5810 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1809_
timestamp 1728341909
transform -1 0 4770 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1811_
timestamp 1728341909
transform 1 0 5010 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1813_
timestamp 1728341909
transform 1 0 5470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1815_
timestamp 1728341909
transform 1 0 5650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1817_
timestamp 1728341909
transform -1 0 5250 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1819_
timestamp 1728341909
transform 1 0 5870 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1821_
timestamp 1728341909
transform 1 0 5890 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1823_
timestamp 1728341909
transform -1 0 5790 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1825_
timestamp 1728341909
transform -1 0 5470 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1826_
timestamp 1728341909
transform 1 0 5870 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1828_
timestamp 1728341909
transform 1 0 6130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1830_
timestamp 1728341909
transform 1 0 5510 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1832_
timestamp 1728341909
transform 1 0 6450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1834_
timestamp 1728341909
transform 1 0 6070 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1836_
timestamp 1728341909
transform -1 0 5170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1838_
timestamp 1728341909
transform 1 0 4590 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1840_
timestamp 1728341909
transform 1 0 5270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1843_
timestamp 1728341909
transform 1 0 5690 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1845_
timestamp 1728341909
transform 1 0 5770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1847_
timestamp 1728341909
transform -1 0 5370 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1849_
timestamp 1728341909
transform 1 0 6110 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1851_
timestamp 1728341909
transform 1 0 6030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1853_
timestamp 1728341909
transform 1 0 6310 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1855_
timestamp 1728341909
transform 1 0 6450 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1857_
timestamp 1728341909
transform -1 0 6010 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1859_
timestamp 1728341909
transform 1 0 6370 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1860_
timestamp 1728341909
transform 1 0 6110 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1862_
timestamp 1728341909
transform -1 0 6350 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1864_
timestamp 1728341909
transform 1 0 6650 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1866_
timestamp 1728341909
transform 1 0 6930 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1868_
timestamp 1728341909
transform 1 0 6830 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1870_
timestamp 1728341909
transform -1 0 6570 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1872_
timestamp 1728341909
transform 1 0 6450 0 1 730
box -12 -8 32 252
use FILL  FILL_0__1874_
timestamp 1728341909
transform -1 0 6850 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1877_
timestamp 1728341909
transform -1 0 4650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1879_
timestamp 1728341909
transform 1 0 4890 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1881_
timestamp 1728341909
transform -1 0 4370 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1883_
timestamp 1728341909
transform 1 0 4770 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1885_
timestamp 1728341909
transform 1 0 5230 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1887_
timestamp 1728341909
transform 1 0 4750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1889_
timestamp 1728341909
transform -1 0 4970 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1891_
timestamp 1728341909
transform 1 0 5530 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1893_
timestamp 1728341909
transform 1 0 5810 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1894_
timestamp 1728341909
transform -1 0 5090 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1896_
timestamp 1728341909
transform 1 0 6030 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1898_
timestamp 1728341909
transform 1 0 4370 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1900_
timestamp 1728341909
transform 1 0 5090 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1902_
timestamp 1728341909
transform 1 0 5230 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1904_
timestamp 1728341909
transform 1 0 5850 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1906_
timestamp 1728341909
transform -1 0 6110 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1908_
timestamp 1728341909
transform 1 0 6210 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1911_
timestamp 1728341909
transform -1 0 6450 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1913_
timestamp 1728341909
transform 1 0 7090 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1915_
timestamp 1728341909
transform -1 0 6650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1917_
timestamp 1728341909
transform 1 0 6970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1919_
timestamp 1728341909
transform 1 0 6470 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1921_
timestamp 1728341909
transform -1 0 6770 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__1923_
timestamp 1728341909
transform -1 0 6990 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1926_
timestamp 1728341909
transform -1 0 7350 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__1928_
timestamp 1728341909
transform 1 0 7210 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1930_
timestamp 1728341909
transform 1 0 7050 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1932_
timestamp 1728341909
transform 1 0 6390 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1934_
timestamp 1728341909
transform 1 0 5130 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1936_
timestamp 1728341909
transform -1 0 5010 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1938_
timestamp 1728341909
transform -1 0 5350 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1940_
timestamp 1728341909
transform -1 0 5130 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1942_
timestamp 1728341909
transform -1 0 4910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1943_
timestamp 1728341909
transform 1 0 5010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1945_
timestamp 1728341909
transform -1 0 5390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1947_
timestamp 1728341909
transform -1 0 5890 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1949_
timestamp 1728341909
transform 1 0 5530 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1951_
timestamp 1728341909
transform 1 0 6110 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1953_
timestamp 1728341909
transform 1 0 5650 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1955_
timestamp 1728341909
transform 1 0 5790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__1957_
timestamp 1728341909
transform 1 0 6270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1960_
timestamp 1728341909
transform 1 0 5970 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1962_
timestamp 1728341909
transform 1 0 6510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1964_
timestamp 1728341909
transform 1 0 6430 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__1966_
timestamp 1728341909
transform -1 0 6650 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1968_
timestamp 1728341909
transform 1 0 6750 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1970_
timestamp 1728341909
transform 1 0 6750 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1972_
timestamp 1728341909
transform 1 0 6870 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__1974_
timestamp 1728341909
transform -1 0 5630 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1976_
timestamp 1728341909
transform -1 0 6530 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1977_
timestamp 1728341909
transform 1 0 6970 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1979_
timestamp 1728341909
transform 1 0 6750 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1981_
timestamp 1728341909
transform 1 0 6850 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__1983_
timestamp 1728341909
transform 1 0 7090 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1985_
timestamp 1728341909
transform 1 0 7290 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__1987_
timestamp 1728341909
transform 1 0 7310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__1989_
timestamp 1728341909
transform 1 0 6910 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1991_
timestamp 1728341909
transform 1 0 7310 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__1994_
timestamp 1728341909
transform 1 0 7370 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__1996_
timestamp 1728341909
transform 1 0 6910 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__1998_
timestamp 1728341909
transform -1 0 4950 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2000_
timestamp 1728341909
transform 1 0 7250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2002_
timestamp 1728341909
transform 1 0 6670 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2004_
timestamp 1728341909
transform -1 0 4450 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2006_
timestamp 1728341909
transform 1 0 4950 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2008_
timestamp 1728341909
transform 1 0 5050 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2010_
timestamp 1728341909
transform 1 0 4730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2011_
timestamp 1728341909
transform 1 0 4510 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2013_
timestamp 1728341909
transform -1 0 6150 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2015_
timestamp 1728341909
transform 1 0 5530 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2017_
timestamp 1728341909
transform -1 0 5710 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2019_
timestamp 1728341909
transform 1 0 5530 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2021_
timestamp 1728341909
transform 1 0 5870 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2023_
timestamp 1728341909
transform -1 0 5750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2025_
timestamp 1728341909
transform 1 0 5470 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2028_
timestamp 1728341909
transform 1 0 6090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2030_
timestamp 1728341909
transform 1 0 5750 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2032_
timestamp 1728341909
transform 1 0 6690 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2034_
timestamp 1728341909
transform 1 0 6430 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2036_
timestamp 1728341909
transform 1 0 6650 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2038_
timestamp 1728341909
transform 1 0 6810 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2040_
timestamp 1728341909
transform 1 0 6790 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2043_
timestamp 1728341909
transform 1 0 7130 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2045_
timestamp 1728341909
transform 1 0 7130 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2047_
timestamp 1728341909
transform 1 0 7430 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2049_
timestamp 1728341909
transform 1 0 7210 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2051_
timestamp 1728341909
transform -1 0 7010 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2053_
timestamp 1728341909
transform 1 0 7390 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2055_
timestamp 1728341909
transform 1 0 7610 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2057_
timestamp 1728341909
transform 1 0 7530 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2059_
timestamp 1728341909
transform -1 0 7390 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2060_
timestamp 1728341909
transform 1 0 7490 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2062_
timestamp 1728341909
transform 1 0 7390 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2064_
timestamp 1728341909
transform -1 0 7550 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2066_
timestamp 1728341909
transform -1 0 5270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2068_
timestamp 1728341909
transform 1 0 6310 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2070_
timestamp 1728341909
transform 1 0 5350 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2072_
timestamp 1728341909
transform -1 0 5990 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2074_
timestamp 1728341909
transform -1 0 5630 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2077_
timestamp 1728341909
transform 1 0 5910 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2079_
timestamp 1728341909
transform -1 0 5250 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2081_
timestamp 1728341909
transform 1 0 5550 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2083_
timestamp 1728341909
transform -1 0 5590 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2085_
timestamp 1728341909
transform 1 0 6230 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2087_
timestamp 1728341909
transform 1 0 6150 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2089_
timestamp 1728341909
transform 1 0 6370 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2091_
timestamp 1728341909
transform 1 0 6710 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2093_
timestamp 1728341909
transform 1 0 7430 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2094_
timestamp 1728341909
transform 1 0 6830 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2096_
timestamp 1728341909
transform 1 0 7770 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2098_
timestamp 1728341909
transform -1 0 7490 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2100_
timestamp 1728341909
transform 1 0 7190 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2102_
timestamp 1728341909
transform 1 0 7790 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2104_
timestamp 1728341909
transform -1 0 7570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2106_
timestamp 1728341909
transform -1 0 7790 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2108_
timestamp 1728341909
transform -1 0 7690 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2111_
timestamp 1728341909
transform 1 0 7570 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2113_
timestamp 1728341909
transform 1 0 7790 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2115_
timestamp 1728341909
transform -1 0 7650 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2117_
timestamp 1728341909
transform 1 0 7590 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2119_
timestamp 1728341909
transform 1 0 7790 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2121_
timestamp 1728341909
transform 1 0 7810 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2123_
timestamp 1728341909
transform 1 0 6950 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2125_
timestamp 1728341909
transform -1 0 6030 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2127_
timestamp 1728341909
transform -1 0 5190 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2128_
timestamp 1728341909
transform -1 0 5050 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2130_
timestamp 1728341909
transform 1 0 4790 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2132_
timestamp 1728341909
transform 1 0 5430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2134_
timestamp 1728341909
transform 1 0 5950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2136_
timestamp 1728341909
transform -1 0 5330 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2138_
timestamp 1728341909
transform 1 0 6450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2140_
timestamp 1728341909
transform 1 0 6090 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2142_
timestamp 1728341909
transform -1 0 6910 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2145_
timestamp 1728341909
transform 1 0 6310 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2147_
timestamp 1728341909
transform 1 0 7130 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2149_
timestamp 1728341909
transform 1 0 6870 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2151_
timestamp 1728341909
transform 1 0 7250 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2153_
timestamp 1728341909
transform -1 0 7270 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2155_
timestamp 1728341909
transform 1 0 7130 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2157_
timestamp 1728341909
transform 1 0 7330 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2160_
timestamp 1728341909
transform -1 0 7490 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2162_
timestamp 1728341909
transform 1 0 7590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2164_
timestamp 1728341909
transform -1 0 7670 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2166_
timestamp 1728341909
transform 1 0 7750 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2168_
timestamp 1728341909
transform -1 0 7830 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2170_
timestamp 1728341909
transform 1 0 7590 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2172_
timestamp 1728341909
transform -1 0 7770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2174_
timestamp 1728341909
transform -1 0 4150 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2176_
timestamp 1728341909
transform 1 0 4370 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2177_
timestamp 1728341909
transform 1 0 4370 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2179_
timestamp 1728341909
transform -1 0 4190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2181_
timestamp 1728341909
transform 1 0 4650 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2183_
timestamp 1728341909
transform 1 0 5130 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2185_
timestamp 1728341909
transform 1 0 5350 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2187_
timestamp 1728341909
transform 1 0 5450 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2189_
timestamp 1728341909
transform 1 0 6770 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2191_
timestamp 1728341909
transform 1 0 6350 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2194_
timestamp 1728341909
transform 1 0 7110 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2196_
timestamp 1728341909
transform 1 0 7370 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2198_
timestamp 1728341909
transform -1 0 7730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2200_
timestamp 1728341909
transform -1 0 7490 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2202_
timestamp 1728341909
transform -1 0 7710 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2204_
timestamp 1728341909
transform -1 0 4610 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2206_
timestamp 1728341909
transform -1 0 4250 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2208_
timestamp 1728341909
transform -1 0 4850 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2210_
timestamp 1728341909
transform 1 0 5030 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2211_
timestamp 1728341909
transform 1 0 6650 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2213_
timestamp 1728341909
transform 1 0 6730 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2215_
timestamp 1728341909
transform 1 0 6770 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2217_
timestamp 1728341909
transform 1 0 7010 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2219_
timestamp 1728341909
transform -1 0 7590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2221_
timestamp 1728341909
transform -1 0 7730 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2223_
timestamp 1728341909
transform -1 0 7650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2225_
timestamp 1728341909
transform 1 0 7490 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2228_
timestamp 1728341909
transform -1 0 6970 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2230_
timestamp 1728341909
transform -1 0 7410 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2232_
timestamp 1728341909
transform -1 0 7510 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2234_
timestamp 1728341909
transform 1 0 4590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2236_
timestamp 1728341909
transform 1 0 4810 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2238_
timestamp 1728341909
transform -1 0 6470 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2240_
timestamp 1728341909
transform 1 0 7270 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2242_
timestamp 1728341909
transform 1 0 7190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2244_
timestamp 1728341909
transform 1 0 7350 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2245_
timestamp 1728341909
transform 1 0 7310 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2247_
timestamp 1728341909
transform 1 0 4950 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2249_
timestamp 1728341909
transform 1 0 4950 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2251_
timestamp 1728341909
transform -1 0 7130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2253_
timestamp 1728341909
transform 1 0 5050 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2255_
timestamp 1728341909
transform -1 0 4950 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2257_
timestamp 1728341909
transform 1 0 4950 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2259_
timestamp 1728341909
transform 1 0 4430 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2262_
timestamp 1728341909
transform 1 0 4690 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2264_
timestamp 1728341909
transform 1 0 4810 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2266_
timestamp 1728341909
transform 1 0 5010 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2268_
timestamp 1728341909
transform 1 0 5010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2270_
timestamp 1728341909
transform 1 0 6130 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2272_
timestamp 1728341909
transform -1 0 5930 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2274_
timestamp 1728341909
transform 1 0 6090 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2277_
timestamp 1728341909
transform 1 0 6170 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2279_
timestamp 1728341909
transform -1 0 5310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2281_
timestamp 1728341909
transform 1 0 5430 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2283_
timestamp 1728341909
transform 1 0 5510 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2285_
timestamp 1728341909
transform -1 0 5390 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2287_
timestamp 1728341909
transform 1 0 5230 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2289_
timestamp 1728341909
transform -1 0 6410 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2291_
timestamp 1728341909
transform -1 0 6650 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2293_
timestamp 1728341909
transform 1 0 5730 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2294_
timestamp 1728341909
transform 1 0 5610 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2296_
timestamp 1728341909
transform 1 0 7070 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2298_
timestamp 1728341909
transform 1 0 6890 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2300_
timestamp 1728341909
transform -1 0 6770 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2302_
timestamp 1728341909
transform -1 0 6570 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2304_
timestamp 1728341909
transform -1 0 6530 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2306_
timestamp 1728341909
transform -1 0 6430 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2308_
timestamp 1728341909
transform -1 0 6250 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2311_
timestamp 1728341909
transform 1 0 4950 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2313_
timestamp 1728341909
transform 1 0 6590 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2315_
timestamp 1728341909
transform -1 0 6370 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2317_
timestamp 1728341909
transform -1 0 5770 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2319_
timestamp 1728341909
transform -1 0 5630 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2321_
timestamp 1728341909
transform -1 0 5410 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2323_
timestamp 1728341909
transform 1 0 5330 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2325_
timestamp 1728341909
transform 1 0 6190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2327_
timestamp 1728341909
transform 1 0 6090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2328_
timestamp 1728341909
transform -1 0 5810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2330_
timestamp 1728341909
transform 1 0 5910 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2332_
timestamp 1728341909
transform 1 0 5530 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2334_
timestamp 1728341909
transform -1 0 7050 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2336_
timestamp 1728341909
transform 1 0 7130 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2338_
timestamp 1728341909
transform 1 0 7490 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2340_
timestamp 1728341909
transform 1 0 6190 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2342_
timestamp 1728341909
transform 1 0 6710 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2345_
timestamp 1728341909
transform -1 0 7690 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2347_
timestamp 1728341909
transform -1 0 7450 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2349_
timestamp 1728341909
transform 1 0 7490 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2351_
timestamp 1728341909
transform 1 0 7750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2353_
timestamp 1728341909
transform 1 0 7790 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2355_
timestamp 1728341909
transform -1 0 7610 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2357_
timestamp 1728341909
transform -1 0 7370 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2359_
timestamp 1728341909
transform -1 0 7010 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2361_
timestamp 1728341909
transform 1 0 7830 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2362_
timestamp 1728341909
transform 1 0 7730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2364_
timestamp 1728341909
transform 1 0 7590 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2366_
timestamp 1728341909
transform 1 0 7830 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2368_
timestamp 1728341909
transform 1 0 7790 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2370_
timestamp 1728341909
transform 1 0 7690 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2372_
timestamp 1728341909
transform -1 0 7450 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2374_
timestamp 1728341909
transform 1 0 7370 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2376_
timestamp 1728341909
transform 1 0 6710 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2379_
timestamp 1728341909
transform 1 0 7790 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2381_
timestamp 1728341909
transform -1 0 7590 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2383_
timestamp 1728341909
transform -1 0 5290 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2385_
timestamp 1728341909
transform -1 0 7410 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2387_
timestamp 1728341909
transform 1 0 7190 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2389_
timestamp 1728341909
transform -1 0 7430 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2391_
timestamp 1728341909
transform -1 0 5610 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2394_
timestamp 1728341909
transform 1 0 6130 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2396_
timestamp 1728341909
transform -1 0 6530 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2398_
timestamp 1728341909
transform 1 0 5790 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2400_
timestamp 1728341909
transform -1 0 5410 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2402_
timestamp 1728341909
transform 1 0 6790 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2404_
timestamp 1728341909
transform 1 0 6150 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2406_
timestamp 1728341909
transform 1 0 6410 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2408_
timestamp 1728341909
transform -1 0 6410 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2410_
timestamp 1728341909
transform 1 0 6150 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2411_
timestamp 1728341909
transform -1 0 6370 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2413_
timestamp 1728341909
transform -1 0 5910 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2415_
timestamp 1728341909
transform 1 0 6190 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2417_
timestamp 1728341909
transform 1 0 6370 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2419_
timestamp 1728341909
transform 1 0 6190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2421_
timestamp 1728341909
transform 1 0 5870 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2423_
timestamp 1728341909
transform 1 0 5650 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2425_
timestamp 1728341909
transform -1 0 5930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2472_
timestamp 1728341909
transform 1 0 1710 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2474_
timestamp 1728341909
transform 1 0 3050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2476_
timestamp 1728341909
transform 1 0 3350 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2478_
timestamp 1728341909
transform -1 0 3170 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2480_
timestamp 1728341909
transform 1 0 3390 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2482_
timestamp 1728341909
transform -1 0 2830 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2484_
timestamp 1728341909
transform 1 0 2270 0 1 5530
box -12 -8 32 252
use FILL  FILL_0__2486_
timestamp 1728341909
transform -1 0 2990 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2488_
timestamp 1728341909
transform 1 0 2410 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2489_
timestamp 1728341909
transform 1 0 2110 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2491_
timestamp 1728341909
transform 1 0 2190 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2493_
timestamp 1728341909
transform -1 0 2050 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2495_
timestamp 1728341909
transform -1 0 2250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2497_
timestamp 1728341909
transform 1 0 2790 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2499_
timestamp 1728341909
transform 1 0 3070 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2501_
timestamp 1728341909
transform 1 0 3170 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2503_
timestamp 1728341909
transform -1 0 2590 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2506_
timestamp 1728341909
transform -1 0 1790 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2508_
timestamp 1728341909
transform -1 0 2250 0 -1 5530
box -12 -8 32 252
use FILL  FILL_0__2510_
timestamp 1728341909
transform -1 0 2790 0 1 5050
box -12 -8 32 252
use FILL  FILL_0__2512_
timestamp 1728341909
transform -1 0 3210 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2514_
timestamp 1728341909
transform 1 0 2930 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__2526_
timestamp 1728341909
transform -1 0 3110 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2528_
timestamp 1728341909
transform -1 0 2410 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2530_
timestamp 1728341909
transform 1 0 2990 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2532_
timestamp 1728341909
transform 1 0 3450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2533_
timestamp 1728341909
transform -1 0 3570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0__2537_
timestamp 1728341909
transform -1 0 2570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2539_
timestamp 1728341909
transform -1 0 2510 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2541_
timestamp 1728341909
transform 1 0 2770 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2543_
timestamp 1728341909
transform -1 0 3090 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2545_
timestamp 1728341909
transform -1 0 2530 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2547_
timestamp 1728341909
transform -1 0 1990 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2549_
timestamp 1728341909
transform 1 0 3010 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2552_
timestamp 1728341909
transform -1 0 530 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2554_
timestamp 1728341909
transform -1 0 210 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2556_
timestamp 1728341909
transform 1 0 1770 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2558_
timestamp 1728341909
transform -1 0 1230 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2560_
timestamp 1728341909
transform -1 0 2770 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2562_
timestamp 1728341909
transform 1 0 2510 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2564_
timestamp 1728341909
transform 1 0 750 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2567_
timestamp 1728341909
transform -1 0 370 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2569_
timestamp 1728341909
transform -1 0 830 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2571_
timestamp 1728341909
transform -1 0 930 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2573_
timestamp 1728341909
transform -1 0 2830 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2575_
timestamp 1728341909
transform -1 0 2950 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2577_
timestamp 1728341909
transform 1 0 570 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2579_
timestamp 1728341909
transform 1 0 410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2581_
timestamp 1728341909
transform -1 0 1230 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2583_
timestamp 1728341909
transform -1 0 1330 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2584_
timestamp 1728341909
transform -1 0 2690 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2586_
timestamp 1728341909
transform 1 0 1810 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2588_
timestamp 1728341909
transform -1 0 1690 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2590_
timestamp 1728341909
transform 1 0 1850 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2592_
timestamp 1728341909
transform -1 0 1510 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2594_
timestamp 1728341909
transform -1 0 2910 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2596_
timestamp 1728341909
transform -1 0 2510 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2598_
timestamp 1728341909
transform 1 0 2730 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2601_
timestamp 1728341909
transform -1 0 2670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2603_
timestamp 1728341909
transform 1 0 3310 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2605_
timestamp 1728341909
transform 1 0 3070 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2607_
timestamp 1728341909
transform -1 0 2730 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2609_
timestamp 1728341909
transform -1 0 3110 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2611_
timestamp 1728341909
transform -1 0 2330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2613_
timestamp 1728341909
transform 1 0 3310 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2615_
timestamp 1728341909
transform -1 0 2510 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2617_
timestamp 1728341909
transform 1 0 1230 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2618_
timestamp 1728341909
transform -1 0 910 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2620_
timestamp 1728341909
transform 1 0 1030 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2622_
timestamp 1728341909
transform -1 0 870 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2624_
timestamp 1728341909
transform 1 0 1410 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2626_
timestamp 1728341909
transform -1 0 1110 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2628_
timestamp 1728341909
transform -1 0 1050 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2630_
timestamp 1728341909
transform -1 0 990 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2632_
timestamp 1728341909
transform 1 0 1170 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2635_
timestamp 1728341909
transform 1 0 1030 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2637_
timestamp 1728341909
transform -1 0 2810 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2639_
timestamp 1728341909
transform 1 0 2790 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2641_
timestamp 1728341909
transform -1 0 2670 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2643_
timestamp 1728341909
transform -1 0 3170 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2645_
timestamp 1728341909
transform 1 0 3350 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2647_
timestamp 1728341909
transform 1 0 850 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2649_
timestamp 1728341909
transform -1 0 1550 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2651_
timestamp 1728341909
transform 1 0 1090 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2652_
timestamp 1728341909
transform -1 0 1350 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2654_
timestamp 1728341909
transform -1 0 1330 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2656_
timestamp 1728341909
transform 1 0 950 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2658_
timestamp 1728341909
transform 1 0 890 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2660_
timestamp 1728341909
transform 1 0 1210 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2662_
timestamp 1728341909
transform 1 0 1090 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2664_
timestamp 1728341909
transform -1 0 1370 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2666_
timestamp 1728341909
transform 1 0 2710 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2669_
timestamp 1728341909
transform -1 0 2530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2671_
timestamp 1728341909
transform 1 0 3170 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2673_
timestamp 1728341909
transform 1 0 2070 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2675_
timestamp 1728341909
transform 1 0 2190 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2677_
timestamp 1728341909
transform 1 0 3270 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2679_
timestamp 1728341909
transform -1 0 2810 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2681_
timestamp 1728341909
transform 1 0 3250 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2684_
timestamp 1728341909
transform -1 0 2710 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2686_
timestamp 1728341909
transform 1 0 1870 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2688_
timestamp 1728341909
transform 1 0 1410 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2690_
timestamp 1728341909
transform 1 0 1770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2692_
timestamp 1728341909
transform -1 0 1750 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2694_
timestamp 1728341909
transform -1 0 3090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2696_
timestamp 1728341909
transform -1 0 2930 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2698_
timestamp 1728341909
transform -1 0 1550 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2700_
timestamp 1728341909
transform -1 0 1730 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2701_
timestamp 1728341909
transform 1 0 1830 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2703_
timestamp 1728341909
transform 1 0 1810 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2705_
timestamp 1728341909
transform -1 0 2290 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2707_
timestamp 1728341909
transform 1 0 2710 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2709_
timestamp 1728341909
transform -1 0 2950 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2711_
timestamp 1728341909
transform 1 0 2110 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2713_
timestamp 1728341909
transform 1 0 2030 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2715_
timestamp 1728341909
transform 1 0 3950 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2718_
timestamp 1728341909
transform -1 0 3710 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2720_
timestamp 1728341909
transform -1 0 2710 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2722_
timestamp 1728341909
transform -1 0 2710 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2724_
timestamp 1728341909
transform -1 0 1350 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2726_
timestamp 1728341909
transform 1 0 1370 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2728_
timestamp 1728341909
transform -1 0 1250 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2730_
timestamp 1728341909
transform -1 0 1550 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2732_
timestamp 1728341909
transform -1 0 2270 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2734_
timestamp 1728341909
transform -1 0 2430 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2735_
timestamp 1728341909
transform -1 0 1370 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2737_
timestamp 1728341909
transform -1 0 1410 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2739_
timestamp 1728341909
transform -1 0 1770 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2741_
timestamp 1728341909
transform 1 0 1490 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2743_
timestamp 1728341909
transform 1 0 2310 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2745_
timestamp 1728341909
transform 1 0 2950 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2747_
timestamp 1728341909
transform 1 0 2390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2749_
timestamp 1728341909
transform 1 0 1730 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2752_
timestamp 1728341909
transform 1 0 1490 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2754_
timestamp 1728341909
transform -1 0 2070 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2756_
timestamp 1728341909
transform 1 0 1890 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2758_
timestamp 1728341909
transform 1 0 210 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2760_
timestamp 1728341909
transform -1 0 450 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2762_
timestamp 1728341909
transform -1 0 490 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2764_
timestamp 1728341909
transform 1 0 330 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2766_
timestamp 1728341909
transform -1 0 270 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__2768_
timestamp 1728341909
transform -1 0 230 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2769_
timestamp 1728341909
transform -1 0 30 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2771_
timestamp 1728341909
transform -1 0 1710 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2773_
timestamp 1728341909
transform 1 0 1910 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2775_
timestamp 1728341909
transform -1 0 230 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2777_
timestamp 1728341909
transform 1 0 330 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2779_
timestamp 1728341909
transform -1 0 570 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2781_
timestamp 1728341909
transform 1 0 670 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2783_
timestamp 1728341909
transform 1 0 2630 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2786_
timestamp 1728341909
transform 1 0 3170 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2788_
timestamp 1728341909
transform 1 0 2030 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2790_
timestamp 1728341909
transform -1 0 1730 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2792_
timestamp 1728341909
transform -1 0 3450 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2794_
timestamp 1728341909
transform -1 0 3470 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2796_
timestamp 1728341909
transform -1 0 3090 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2798_
timestamp 1728341909
transform -1 0 3190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2801_
timestamp 1728341909
transform -1 0 610 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2803_
timestamp 1728341909
transform -1 0 110 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2805_
timestamp 1728341909
transform 1 0 290 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2807_
timestamp 1728341909
transform -1 0 2670 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2809_
timestamp 1728341909
transform 1 0 2170 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2811_
timestamp 1728341909
transform -1 0 150 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2813_
timestamp 1728341909
transform -1 0 110 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2815_
timestamp 1728341909
transform -1 0 590 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2817_
timestamp 1728341909
transform -1 0 250 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2818_
timestamp 1728341909
transform -1 0 370 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2820_
timestamp 1728341909
transform 1 0 570 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2822_
timestamp 1728341909
transform 1 0 1790 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2824_
timestamp 1728341909
transform -1 0 570 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2826_
timestamp 1728341909
transform -1 0 770 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2828_
timestamp 1728341909
transform -1 0 1110 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2830_
timestamp 1728341909
transform 1 0 890 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2832_
timestamp 1728341909
transform -1 0 350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2835_
timestamp 1728341909
transform -1 0 270 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2837_
timestamp 1728341909
transform 1 0 550 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2839_
timestamp 1728341909
transform -1 0 830 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2841_
timestamp 1728341909
transform 1 0 670 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2843_
timestamp 1728341909
transform -1 0 950 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2845_
timestamp 1728341909
transform 1 0 1570 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2847_
timestamp 1728341909
transform 1 0 250 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2849_
timestamp 1728341909
transform 1 0 550 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2851_
timestamp 1728341909
transform 1 0 1010 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2852_
timestamp 1728341909
transform -1 0 790 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2854_
timestamp 1728341909
transform 1 0 870 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2856_
timestamp 1728341909
transform 1 0 2830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2858_
timestamp 1728341909
transform 1 0 2010 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2860_
timestamp 1728341909
transform -1 0 2130 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2862_
timestamp 1728341909
transform -1 0 2010 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2864_
timestamp 1728341909
transform -1 0 2490 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2866_
timestamp 1728341909
transform 1 0 2330 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2869_
timestamp 1728341909
transform -1 0 1870 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2871_
timestamp 1728341909
transform 1 0 1710 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2873_
timestamp 1728341909
transform 1 0 1830 0 1 2650
box -12 -8 32 252
use FILL  FILL_0__2875_
timestamp 1728341909
transform 1 0 1610 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2877_
timestamp 1728341909
transform 1 0 1730 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2879_
timestamp 1728341909
transform 1 0 2030 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2881_
timestamp 1728341909
transform 1 0 2310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2883_
timestamp 1728341909
transform 1 0 1810 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2885_
timestamp 1728341909
transform 1 0 1670 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2886_
timestamp 1728341909
transform -1 0 1490 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2888_
timestamp 1728341909
transform -1 0 1770 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2890_
timestamp 1728341909
transform 1 0 3130 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2892_
timestamp 1728341909
transform 1 0 2010 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2894_
timestamp 1728341909
transform -1 0 3250 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2896_
timestamp 1728341909
transform -1 0 2090 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2898_
timestamp 1728341909
transform 1 0 2150 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2900_
timestamp 1728341909
transform 1 0 2450 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2903_
timestamp 1728341909
transform 1 0 3950 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2905_
timestamp 1728341909
transform -1 0 2250 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2907_
timestamp 1728341909
transform 1 0 3270 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2909_
timestamp 1728341909
transform 1 0 2890 0 1 3130
box -12 -8 32 252
use FILL  FILL_0__2911_
timestamp 1728341909
transform 1 0 3470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2913_
timestamp 1728341909
transform 1 0 3590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_0__2915_
timestamp 1728341909
transform -1 0 4450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2918_
timestamp 1728341909
transform -1 0 770 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2920_
timestamp 1728341909
transform 1 0 3390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0__2922_
timestamp 1728341909
transform 1 0 3550 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2924_
timestamp 1728341909
transform 1 0 3350 0 1 1210
box -12 -8 32 252
use FILL  FILL_0__2926_
timestamp 1728341909
transform -1 0 4290 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2928_
timestamp 1728341909
transform -1 0 650 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2930_
timestamp 1728341909
transform 1 0 750 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2932_
timestamp 1728341909
transform 1 0 1030 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2934_
timestamp 1728341909
transform 1 0 1190 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2935_
timestamp 1728341909
transform -1 0 1410 0 1 730
box -12 -8 32 252
use FILL  FILL_0__2937_
timestamp 1728341909
transform -1 0 2470 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2939_
timestamp 1728341909
transform -1 0 3590 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2941_
timestamp 1728341909
transform -1 0 1210 0 -1 730
box -12 -8 32 252
use FILL  FILL_0__2943_
timestamp 1728341909
transform 1 0 3330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__2945_
timestamp 1728341909
transform 1 0 1270 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__2947_
timestamp 1728341909
transform 1 0 1970 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2949_
timestamp 1728341909
transform -1 0 2310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2952_
timestamp 1728341909
transform 1 0 2150 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2954_
timestamp 1728341909
transform 1 0 2530 0 1 250
box -12 -8 32 252
use FILL  FILL_0__2956_
timestamp 1728341909
transform 1 0 3450 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2958_
timestamp 1728341909
transform 1 0 3610 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2960_
timestamp 1728341909
transform 1 0 3430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_0__2962_
timestamp 1728341909
transform -1 0 4070 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__2964_
timestamp 1728341909
transform 1 0 730 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2966_
timestamp 1728341909
transform 1 0 830 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2968_
timestamp 1728341909
transform -1 0 670 0 1 4090
box -12 -8 32 252
use FILL  FILL_0__2969_
timestamp 1728341909
transform 1 0 950 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2971_
timestamp 1728341909
transform -1 0 2050 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2973_
timestamp 1728341909
transform -1 0 2270 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2975_
timestamp 1728341909
transform -1 0 1990 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2977_
timestamp 1728341909
transform -1 0 1030 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2979_
timestamp 1728341909
transform 1 0 2250 0 1 4570
box -12 -8 32 252
use FILL  FILL_0__2981_
timestamp 1728341909
transform -1 0 1550 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__2983_
timestamp 1728341909
transform -1 0 1930 0 -1 4570
box -12 -8 32 252
use FILL  FILL_0__2986_
timestamp 1728341909
transform 1 0 2070 0 -1 5050
box -12 -8 32 252
use FILL  FILL_0__2988_
timestamp 1728341909
transform 1 0 2370 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__2990_
timestamp 1728341909
transform -1 0 1630 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2992_
timestamp 1728341909
transform 1 0 1370 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__2994_
timestamp 1728341909
transform 1 0 3730 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2996_
timestamp 1728341909
transform 1 0 3310 0 -1 3130
box -12 -8 32 252
use FILL  FILL_0__2998_
timestamp 1728341909
transform 1 0 3950 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__3000_
timestamp 1728341909
transform 1 0 3210 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0__3002_
timestamp 1728341909
transform 1 0 250 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__3003_
timestamp 1728341909
transform 1 0 410 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0__3005_
timestamp 1728341909
transform 1 0 330 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__3007_
timestamp 1728341909
transform 1 0 710 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__3009_
timestamp 1728341909
transform -1 0 510 0 1 1690
box -12 -8 32 252
use FILL  FILL_0__3011_
timestamp 1728341909
transform 1 0 3190 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__3013_
timestamp 1728341909
transform -1 0 3310 0 1 2170
box -12 -8 32 252
use FILL  FILL_0__3015_
timestamp 1728341909
transform 1 0 750 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3017_
timestamp 1728341909
transform 1 0 590 0 1 3610
box -12 -8 32 252
use FILL  FILL_0__3020_
timestamp 1728341909
transform 1 0 430 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0__3102_
timestamp 1728341909
transform -1 0 30 0 1 6010
box -12 -8 32 252
use FILL  FILL_0__3104_
timestamp 1728341909
transform -1 0 3430 0 1 250
box -12 -8 32 252
use FILL  FILL_0__3106_
timestamp 1728341909
transform -1 0 3790 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3108_
timestamp 1728341909
transform -1 0 3610 0 -1 250
box -12 -8 32 252
use FILL  FILL_0__3110_
timestamp 1728341909
transform 1 0 4970 0 -1 250
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert14
timestamp 1728341909
transform -1 0 5870 0 1 1210
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert16
timestamp 1728341909
transform 1 0 6830 0 1 730
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert18
timestamp 1728341909
transform 1 0 5750 0 1 1210
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert20
timestamp 1728341909
transform -1 0 4030 0 1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert22
timestamp 1728341909
transform 1 0 1910 0 1 3610
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert24
timestamp 1728341909
transform -1 0 930 0 1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert27
timestamp 1728341909
transform 1 0 3450 0 -1 4090
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert29
timestamp 1728341909
transform 1 0 90 0 -1 6010
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert31
timestamp 1728341909
transform -1 0 30 0 1 5050
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert33
timestamp 1728341909
transform 1 0 5330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert35
timestamp 1728341909
transform -1 0 6310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert37
timestamp 1728341909
transform 1 0 2630 0 1 3130
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert39
timestamp 1728341909
transform -1 0 1170 0 1 1210
box -12 -8 32 252
use FILL  FILL_0_BUFX2_insert41
timestamp 1728341909
transform 1 0 2590 0 1 730
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert1
timestamp 1728341909
transform -1 0 4010 0 1 1210
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert3
timestamp 1728341909
transform 1 0 6330 0 1 2650
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert5
timestamp 1728341909
transform -1 0 4330 0 1 6010
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert7
timestamp 1728341909
transform -1 0 450 0 1 5050
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1728341909
transform -1 0 4650 0 1 730
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1728341909
transform -1 0 310 0 -1 2650
box -12 -8 32 252
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1728341909
transform 1 0 410 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1436_
timestamp 1728341909
transform -1 0 4290 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1440_
timestamp 1728341909
transform -1 0 4510 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1443_
timestamp 1728341909
transform 1 0 4270 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1447_
timestamp 1728341909
transform -1 0 5190 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1451_
timestamp 1728341909
transform -1 0 4770 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1455_
timestamp 1728341909
transform -1 0 4010 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1462_
timestamp 1728341909
transform 1 0 3990 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1466_
timestamp 1728341909
transform -1 0 3890 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1470_
timestamp 1728341909
transform -1 0 3910 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1474_
timestamp 1728341909
transform -1 0 4250 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1477_
timestamp 1728341909
transform 1 0 5190 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1481_
timestamp 1728341909
transform 1 0 4750 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1485_
timestamp 1728341909
transform -1 0 2870 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1489_
timestamp 1728341909
transform 1 0 3370 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1496_
timestamp 1728341909
transform 1 0 3350 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1500_
timestamp 1728341909
transform -1 0 50 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1504_
timestamp 1728341909
transform -1 0 50 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1508_
timestamp 1728341909
transform 1 0 290 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__1511_
timestamp 1728341909
transform -1 0 130 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__1515_
timestamp 1728341909
transform -1 0 250 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1519_
timestamp 1728341909
transform -1 0 150 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1523_
timestamp 1728341909
transform 1 0 350 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1526_
timestamp 1728341909
transform 1 0 1450 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__1530_
timestamp 1728341909
transform 1 0 550 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__1534_
timestamp 1728341909
transform 1 0 1370 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1538_
timestamp 1728341909
transform -1 0 1150 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1545_
timestamp 1728341909
transform -1 0 1190 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__1549_
timestamp 1728341909
transform 1 0 1590 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1553_
timestamp 1728341909
transform -1 0 1170 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1572_
timestamp 1728341909
transform -1 0 3810 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1575_
timestamp 1728341909
transform 1 0 3870 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1579_
timestamp 1728341909
transform -1 0 3350 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1583_
timestamp 1728341909
transform -1 0 3310 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1587_
timestamp 1728341909
transform 1 0 4790 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1594_
timestamp 1728341909
transform 1 0 4670 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1598_
timestamp 1728341909
transform 1 0 6030 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__1602_
timestamp 1728341909
transform -1 0 5390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__1606_
timestamp 1728341909
transform -1 0 4910 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1609_
timestamp 1728341909
transform -1 0 6530 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1613_
timestamp 1728341909
transform 1 0 7310 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1617_
timestamp 1728341909
transform -1 0 6830 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__1621_
timestamp 1728341909
transform -1 0 4810 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1628_
timestamp 1728341909
transform 1 0 6490 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1632_
timestamp 1728341909
transform -1 0 5570 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1636_
timestamp 1728341909
transform 1 0 1230 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1640_
timestamp 1728341909
transform 1 0 3650 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1643_
timestamp 1728341909
transform -1 0 3530 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1647_
timestamp 1728341909
transform -1 0 3210 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1651_
timestamp 1728341909
transform -1 0 4430 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__1655_
timestamp 1728341909
transform -1 0 5550 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__1658_
timestamp 1728341909
transform -1 0 5030 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__1662_
timestamp 1728341909
transform 1 0 6490 0 1 250
box -12 -8 32 252
use FILL  FILL_1__1666_
timestamp 1728341909
transform -1 0 5430 0 1 730
box -12 -8 32 252
use FILL  FILL_1__1670_
timestamp 1728341909
transform 1 0 3470 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__1705_
timestamp 1728341909
transform 1 0 4070 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1709_
timestamp 1728341909
transform -1 0 3510 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1713_
timestamp 1728341909
transform 1 0 3950 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1717_
timestamp 1728341909
transform 1 0 3710 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1720_
timestamp 1728341909
transform 1 0 3850 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1724_
timestamp 1728341909
transform 1 0 3610 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1732_
timestamp 1728341909
transform 1 0 2110 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1736_
timestamp 1728341909
transform 1 0 2230 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__1745_
timestamp 1728341909
transform -1 0 4230 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1749_
timestamp 1728341909
transform -1 0 4370 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1753_
timestamp 1728341909
transform -1 0 4210 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1757_
timestamp 1728341909
transform -1 0 3770 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__1760_
timestamp 1728341909
transform -1 0 4530 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1764_
timestamp 1728341909
transform -1 0 4750 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1768_
timestamp 1728341909
transform 1 0 4610 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1772_
timestamp 1728341909
transform -1 0 4230 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1779_
timestamp 1728341909
transform 1 0 4050 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__1783_
timestamp 1728341909
transform -1 0 4910 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1787_
timestamp 1728341909
transform -1 0 4670 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1791_
timestamp 1728341909
transform 1 0 5010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1794_
timestamp 1728341909
transform 1 0 5250 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1798_
timestamp 1728341909
transform 1 0 5290 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1802_
timestamp 1728341909
transform 1 0 6050 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1806_
timestamp 1728341909
transform -1 0 5830 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1809_
timestamp 1728341909
transform -1 0 4790 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1813_
timestamp 1728341909
transform 1 0 5490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1817_
timestamp 1728341909
transform -1 0 5270 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1821_
timestamp 1728341909
transform 1 0 5910 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1828_
timestamp 1728341909
transform 1 0 6150 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1832_
timestamp 1728341909
transform 1 0 6470 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1836_
timestamp 1728341909
transform -1 0 5190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1840_
timestamp 1728341909
transform 1 0 5290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1843_
timestamp 1728341909
transform 1 0 5710 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1847_
timestamp 1728341909
transform -1 0 5390 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1851_
timestamp 1728341909
transform 1 0 6050 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1855_
timestamp 1728341909
transform 1 0 6470 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1862_
timestamp 1728341909
transform -1 0 6370 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1866_
timestamp 1728341909
transform 1 0 6950 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1870_
timestamp 1728341909
transform -1 0 6590 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1874_
timestamp 1728341909
transform -1 0 6870 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1877_
timestamp 1728341909
transform -1 0 4670 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1881_
timestamp 1728341909
transform -1 0 4390 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1885_
timestamp 1728341909
transform 1 0 5250 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1889_
timestamp 1728341909
transform -1 0 4990 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1896_
timestamp 1728341909
transform 1 0 6050 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1900_
timestamp 1728341909
transform 1 0 5110 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1904_
timestamp 1728341909
transform 1 0 5870 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1908_
timestamp 1728341909
transform 1 0 6230 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1911_
timestamp 1728341909
transform -1 0 6470 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1915_
timestamp 1728341909
transform -1 0 6670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__1919_
timestamp 1728341909
transform 1 0 6490 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1923_
timestamp 1728341909
transform -1 0 7010 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1926_
timestamp 1728341909
transform -1 0 7370 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__1930_
timestamp 1728341909
transform 1 0 7070 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1934_
timestamp 1728341909
transform 1 0 5150 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1938_
timestamp 1728341909
transform -1 0 5370 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1945_
timestamp 1728341909
transform -1 0 5410 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1949_
timestamp 1728341909
transform 1 0 5550 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1953_
timestamp 1728341909
transform 1 0 5670 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__1957_
timestamp 1728341909
transform 1 0 6290 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1960_
timestamp 1728341909
transform 1 0 5990 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1964_
timestamp 1728341909
transform 1 0 6450 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__1968_
timestamp 1728341909
transform 1 0 6770 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__1972_
timestamp 1728341909
transform 1 0 6890 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__1979_
timestamp 1728341909
transform 1 0 6770 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__1983_
timestamp 1728341909
transform 1 0 7110 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__1987_
timestamp 1728341909
transform 1 0 7330 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__1991_
timestamp 1728341909
transform 1 0 7330 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__1994_
timestamp 1728341909
transform 1 0 7390 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__1998_
timestamp 1728341909
transform -1 0 4970 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2002_
timestamp 1728341909
transform 1 0 6690 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2006_
timestamp 1728341909
transform 1 0 4970 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2013_
timestamp 1728341909
transform -1 0 6170 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2017_
timestamp 1728341909
transform -1 0 5730 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2021_
timestamp 1728341909
transform 1 0 5890 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2025_
timestamp 1728341909
transform 1 0 5490 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2028_
timestamp 1728341909
transform 1 0 6110 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2032_
timestamp 1728341909
transform 1 0 6710 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2036_
timestamp 1728341909
transform 1 0 6670 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2040_
timestamp 1728341909
transform 1 0 6810 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2043_
timestamp 1728341909
transform 1 0 7150 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2047_
timestamp 1728341909
transform 1 0 7450 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2051_
timestamp 1728341909
transform -1 0 7030 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2055_
timestamp 1728341909
transform 1 0 7630 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2062_
timestamp 1728341909
transform 1 0 7410 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2066_
timestamp 1728341909
transform -1 0 5290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2070_
timestamp 1728341909
transform 1 0 5370 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2074_
timestamp 1728341909
transform -1 0 5650 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2077_
timestamp 1728341909
transform 1 0 5930 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2081_
timestamp 1728341909
transform 1 0 5570 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2085_
timestamp 1728341909
transform 1 0 6250 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2089_
timestamp 1728341909
transform 1 0 6390 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2096_
timestamp 1728341909
transform 1 0 7790 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2100_
timestamp 1728341909
transform 1 0 7210 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2104_
timestamp 1728341909
transform -1 0 7590 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2108_
timestamp 1728341909
transform -1 0 7710 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2111_
timestamp 1728341909
transform 1 0 7590 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2115_
timestamp 1728341909
transform -1 0 7670 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2119_
timestamp 1728341909
transform 1 0 7810 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2123_
timestamp 1728341909
transform 1 0 6970 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2130_
timestamp 1728341909
transform 1 0 4810 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2134_
timestamp 1728341909
transform 1 0 5970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2138_
timestamp 1728341909
transform 1 0 6470 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2142_
timestamp 1728341909
transform -1 0 6930 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2145_
timestamp 1728341909
transform 1 0 6330 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2149_
timestamp 1728341909
transform 1 0 6890 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2153_
timestamp 1728341909
transform -1 0 7290 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2157_
timestamp 1728341909
transform 1 0 7350 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2160_
timestamp 1728341909
transform -1 0 7510 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2164_
timestamp 1728341909
transform -1 0 7690 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2168_
timestamp 1728341909
transform -1 0 7850 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2172_
timestamp 1728341909
transform -1 0 7790 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2179_
timestamp 1728341909
transform -1 0 4210 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2183_
timestamp 1728341909
transform 1 0 5150 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2187_
timestamp 1728341909
transform 1 0 5470 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2191_
timestamp 1728341909
transform 1 0 6370 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2194_
timestamp 1728341909
transform 1 0 7130 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2198_
timestamp 1728341909
transform -1 0 7750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2202_
timestamp 1728341909
transform -1 0 7730 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2206_
timestamp 1728341909
transform -1 0 4270 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2213_
timestamp 1728341909
transform 1 0 6750 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2217_
timestamp 1728341909
transform 1 0 7030 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2221_
timestamp 1728341909
transform -1 0 7750 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2225_
timestamp 1728341909
transform 1 0 7510 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2228_
timestamp 1728341909
transform -1 0 6990 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2232_
timestamp 1728341909
transform -1 0 7530 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2236_
timestamp 1728341909
transform 1 0 4830 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2240_
timestamp 1728341909
transform 1 0 7290 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2247_
timestamp 1728341909
transform 1 0 4970 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2251_
timestamp 1728341909
transform -1 0 7150 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2255_
timestamp 1728341909
transform -1 0 4970 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2259_
timestamp 1728341909
transform 1 0 4450 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2262_
timestamp 1728341909
transform 1 0 4710 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2266_
timestamp 1728341909
transform 1 0 5030 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2270_
timestamp 1728341909
transform 1 0 6150 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2274_
timestamp 1728341909
transform 1 0 6110 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2277_
timestamp 1728341909
transform 1 0 6190 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2281_
timestamp 1728341909
transform 1 0 5450 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2285_
timestamp 1728341909
transform -1 0 5410 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2289_
timestamp 1728341909
transform -1 0 6430 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2296_
timestamp 1728341909
transform 1 0 7090 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2300_
timestamp 1728341909
transform -1 0 6790 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2304_
timestamp 1728341909
transform -1 0 6550 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2308_
timestamp 1728341909
transform -1 0 6270 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2311_
timestamp 1728341909
transform 1 0 4970 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2315_
timestamp 1728341909
transform -1 0 6390 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2319_
timestamp 1728341909
transform -1 0 5650 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2323_
timestamp 1728341909
transform 1 0 5350 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2330_
timestamp 1728341909
transform 1 0 5930 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2334_
timestamp 1728341909
transform -1 0 7070 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2338_
timestamp 1728341909
transform 1 0 7510 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2342_
timestamp 1728341909
transform 1 0 6730 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2345_
timestamp 1728341909
transform -1 0 7710 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2349_
timestamp 1728341909
transform 1 0 7510 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2353_
timestamp 1728341909
transform 1 0 7810 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2357_
timestamp 1728341909
transform -1 0 7390 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2364_
timestamp 1728341909
transform 1 0 7610 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2368_
timestamp 1728341909
transform 1 0 7810 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2372_
timestamp 1728341909
transform -1 0 7470 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2376_
timestamp 1728341909
transform 1 0 6730 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2379_
timestamp 1728341909
transform 1 0 7810 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2383_
timestamp 1728341909
transform -1 0 5310 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2387_
timestamp 1728341909
transform 1 0 7210 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2391_
timestamp 1728341909
transform -1 0 5630 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2394_
timestamp 1728341909
transform 1 0 6150 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2398_
timestamp 1728341909
transform 1 0 5810 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2402_
timestamp 1728341909
transform 1 0 6810 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2406_
timestamp 1728341909
transform 1 0 6430 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2413_
timestamp 1728341909
transform -1 0 5930 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2417_
timestamp 1728341909
transform 1 0 6390 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2421_
timestamp 1728341909
transform 1 0 5890 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2425_
timestamp 1728341909
transform -1 0 5950 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2472_
timestamp 1728341909
transform 1 0 1730 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2476_
timestamp 1728341909
transform 1 0 3370 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2480_
timestamp 1728341909
transform 1 0 3410 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2484_
timestamp 1728341909
transform 1 0 2290 0 1 5530
box -12 -8 32 252
use FILL  FILL_1__2491_
timestamp 1728341909
transform 1 0 2210 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2495_
timestamp 1728341909
transform -1 0 2270 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2499_
timestamp 1728341909
transform 1 0 3090 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2503_
timestamp 1728341909
transform -1 0 2610 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2506_
timestamp 1728341909
transform -1 0 1810 0 -1 5530
box -12 -8 32 252
use FILL  FILL_1__2510_
timestamp 1728341909
transform -1 0 2810 0 1 5050
box -12 -8 32 252
use FILL  FILL_1__2514_
timestamp 1728341909
transform 1 0 2950 0 1 6010
box -12 -8 32 252
use FILL  FILL_1__2528_
timestamp 1728341909
transform -1 0 2430 0 -1 6010
box -12 -8 32 252
use FILL  FILL_1__2537_
timestamp 1728341909
transform -1 0 2590 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2541_
timestamp 1728341909
transform 1 0 2790 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2545_
timestamp 1728341909
transform -1 0 2550 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2549_
timestamp 1728341909
transform 1 0 3030 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2552_
timestamp 1728341909
transform -1 0 550 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2556_
timestamp 1728341909
transform 1 0 1790 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2560_
timestamp 1728341909
transform -1 0 2790 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2564_
timestamp 1728341909
transform 1 0 770 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2567_
timestamp 1728341909
transform -1 0 390 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2571_
timestamp 1728341909
transform -1 0 950 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2575_
timestamp 1728341909
transform -1 0 2970 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2579_
timestamp 1728341909
transform 1 0 430 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2586_
timestamp 1728341909
transform 1 0 1830 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2590_
timestamp 1728341909
transform 1 0 1870 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2594_
timestamp 1728341909
transform -1 0 2930 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2598_
timestamp 1728341909
transform 1 0 2750 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2601_
timestamp 1728341909
transform -1 0 2690 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2605_
timestamp 1728341909
transform 1 0 3090 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2609_
timestamp 1728341909
transform -1 0 3130 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2613_
timestamp 1728341909
transform 1 0 3330 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2620_
timestamp 1728341909
transform 1 0 1050 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2624_
timestamp 1728341909
transform 1 0 1430 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2628_
timestamp 1728341909
transform -1 0 1070 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2632_
timestamp 1728341909
transform 1 0 1190 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2635_
timestamp 1728341909
transform 1 0 1050 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2639_
timestamp 1728341909
transform 1 0 2810 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2643_
timestamp 1728341909
transform -1 0 3190 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2647_
timestamp 1728341909
transform 1 0 870 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2654_
timestamp 1728341909
transform -1 0 1350 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2658_
timestamp 1728341909
transform 1 0 910 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2662_
timestamp 1728341909
transform 1 0 1110 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2666_
timestamp 1728341909
transform 1 0 2730 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2669_
timestamp 1728341909
transform -1 0 2550 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2673_
timestamp 1728341909
transform 1 0 2090 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2677_
timestamp 1728341909
transform 1 0 3290 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2681_
timestamp 1728341909
transform 1 0 3270 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2684_
timestamp 1728341909
transform -1 0 2730 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2688_
timestamp 1728341909
transform 1 0 1430 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2692_
timestamp 1728341909
transform -1 0 1770 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2696_
timestamp 1728341909
transform -1 0 2950 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2703_
timestamp 1728341909
transform 1 0 1830 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2707_
timestamp 1728341909
transform 1 0 2730 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2711_
timestamp 1728341909
transform 1 0 2130 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2715_
timestamp 1728341909
transform 1 0 3970 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2718_
timestamp 1728341909
transform -1 0 3730 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2722_
timestamp 1728341909
transform -1 0 2730 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2726_
timestamp 1728341909
transform 1 0 1390 0 -1 250
box -12 -8 32 252
use FILL  FILL_1__2730_
timestamp 1728341909
transform -1 0 1570 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2737_
timestamp 1728341909
transform -1 0 1430 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2741_
timestamp 1728341909
transform 1 0 1510 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2745_
timestamp 1728341909
transform 1 0 2970 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2749_
timestamp 1728341909
transform 1 0 1750 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2752_
timestamp 1728341909
transform 1 0 1510 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2756_
timestamp 1728341909
transform 1 0 1910 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2760_
timestamp 1728341909
transform -1 0 470 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2764_
timestamp 1728341909
transform 1 0 350 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2771_
timestamp 1728341909
transform -1 0 1730 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2775_
timestamp 1728341909
transform -1 0 250 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2779_
timestamp 1728341909
transform -1 0 590 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2783_
timestamp 1728341909
transform 1 0 2650 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2786_
timestamp 1728341909
transform 1 0 3190 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__2790_
timestamp 1728341909
transform -1 0 1750 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2794_
timestamp 1728341909
transform -1 0 3490 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2798_
timestamp 1728341909
transform -1 0 3210 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2801_
timestamp 1728341909
transform -1 0 630 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2805_
timestamp 1728341909
transform 1 0 310 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2809_
timestamp 1728341909
transform 1 0 2190 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2813_
timestamp 1728341909
transform -1 0 130 0 1 4090
box -12 -8 32 252
use FILL  FILL_1__2820_
timestamp 1728341909
transform 1 0 590 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2824_
timestamp 1728341909
transform -1 0 590 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2828_
timestamp 1728341909
transform -1 0 1130 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2832_
timestamp 1728341909
transform -1 0 370 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2835_
timestamp 1728341909
transform -1 0 290 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2839_
timestamp 1728341909
transform -1 0 850 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2843_
timestamp 1728341909
transform -1 0 970 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2847_
timestamp 1728341909
transform 1 0 270 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2854_
timestamp 1728341909
transform 1 0 890 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2858_
timestamp 1728341909
transform 1 0 2030 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2862_
timestamp 1728341909
transform -1 0 2030 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2866_
timestamp 1728341909
transform 1 0 2350 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2869_
timestamp 1728341909
transform -1 0 1890 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2873_
timestamp 1728341909
transform 1 0 1850 0 1 2650
box -12 -8 32 252
use FILL  FILL_1__2877_
timestamp 1728341909
transform 1 0 1750 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__2881_
timestamp 1728341909
transform 1 0 2330 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2888_
timestamp 1728341909
transform -1 0 1790 0 1 3130
box -12 -8 32 252
use FILL  FILL_1__2892_
timestamp 1728341909
transform 1 0 2030 0 1 730
box -12 -8 32 252
use FILL  FILL_1__2896_
timestamp 1728341909
transform -1 0 2110 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2900_
timestamp 1728341909
transform 1 0 2470 0 1 1210
box -12 -8 32 252
use FILL  FILL_1__2903_
timestamp 1728341909
transform 1 0 3970 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2907_
timestamp 1728341909
transform 1 0 3290 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__2911_
timestamp 1728341909
transform 1 0 3490 0 -1 3610
box -12 -8 32 252
use FILL  FILL_1__2915_
timestamp 1728341909
transform -1 0 4470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2918_
timestamp 1728341909
transform -1 0 790 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1__2922_
timestamp 1728341909
transform 1 0 3570 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2926_
timestamp 1728341909
transform -1 0 4310 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2930_
timestamp 1728341909
transform 1 0 770 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2937_
timestamp 1728341909
transform -1 0 2490 0 -1 2650
box -12 -8 32 252
use FILL  FILL_1__2941_
timestamp 1728341909
transform -1 0 1230 0 -1 730
box -12 -8 32 252
use FILL  FILL_1__2945_
timestamp 1728341909
transform 1 0 1290 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__2949_
timestamp 1728341909
transform -1 0 2330 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2952_
timestamp 1728341909
transform 1 0 2170 0 1 250
box -12 -8 32 252
use FILL  FILL_1__2956_
timestamp 1728341909
transform 1 0 3470 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2960_
timestamp 1728341909
transform 1 0 3450 0 -1 1210
box -12 -8 32 252
use FILL  FILL_1__2964_
timestamp 1728341909
transform 1 0 750 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2971_
timestamp 1728341909
transform -1 0 2070 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2975_
timestamp 1728341909
transform -1 0 2010 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2979_
timestamp 1728341909
transform 1 0 2270 0 1 4570
box -12 -8 32 252
use FILL  FILL_1__2983_
timestamp 1728341909
transform -1 0 1950 0 -1 4570
box -12 -8 32 252
use FILL  FILL_1__2986_
timestamp 1728341909
transform 1 0 2090 0 -1 5050
box -12 -8 32 252
use FILL  FILL_1__2990_
timestamp 1728341909
transform -1 0 1650 0 -1 2170
box -12 -8 32 252
use FILL  FILL_1__2994_
timestamp 1728341909
transform 1 0 3750 0 -1 3130
box -12 -8 32 252
use FILL  FILL_1__2998_
timestamp 1728341909
transform 1 0 3970 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__3005_
timestamp 1728341909
transform 1 0 350 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__3009_
timestamp 1728341909
transform -1 0 530 0 1 1690
box -12 -8 32 252
use FILL  FILL_1__3013_
timestamp 1728341909
transform -1 0 3330 0 1 2170
box -12 -8 32 252
use FILL  FILL_1__3017_
timestamp 1728341909
transform 1 0 610 0 1 3610
box -12 -8 32 252
use FILL  FILL_1__3020_
timestamp 1728341909
transform 1 0 450 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1__3104_
timestamp 1728341909
transform -1 0 3450 0 1 250
box -12 -8 32 252
use FILL  FILL_1__3108_
timestamp 1728341909
transform -1 0 3630 0 -1 250
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert16
timestamp 1728341909
transform 1 0 6850 0 1 730
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert20
timestamp 1728341909
transform -1 0 4050 0 1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert24
timestamp 1728341909
transform -1 0 950 0 1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert27
timestamp 1728341909
transform 1 0 3470 0 -1 4090
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert31
timestamp 1728341909
transform -1 0 50 0 1 5050
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert35
timestamp 1728341909
transform -1 0 6330 0 -1 1690
box -12 -8 32 252
use FILL  FILL_1_BUFX2_insert39
timestamp 1728341909
transform -1 0 1190 0 1 1210
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert1
timestamp 1728341909
transform -1 0 4030 0 1 1210
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert5
timestamp 1728341909
transform -1 0 4350 0 1 6010
box -12 -8 32 252
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1728341909
transform 1 0 430 0 -1 5050
box -12 -8 32 252
<< labels >>
flabel metal1 s 7922 2 7982 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s -24 3056 -16 3064 7 FreeSans 16 0 0 0 clk
port 2 nsew
flabel metal3 s -24 5416 -16 5424 7 FreeSans 16 0 0 0 rst
port 4 nsew
flabel metal2 s 177 6297 183 6303 3 FreeSans 16 90 0 0 x[6]
port 6 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 x[5]
port 7 nsew
flabel metal2 s 357 6297 363 6303 3 FreeSans 16 90 0 0 x[4]
port 8 nsew
flabel metal3 s -24 2516 -16 2524 7 FreeSans 16 0 0 0 x[3]
port 9 nsew
flabel metal3 s -24 6156 -16 6164 7 FreeSans 16 0 0 0 x[1]
port 11 nsew
flabel metal2 s 5017 -23 5023 -17 7 FreeSans 16 270 0 0 y[7]
port 13 nsew
flabel metal2 s 4657 -23 4663 -17 7 FreeSans 16 270 0 0 y[6]
port 14 nsew
flabel metal2 s 4397 -23 4403 -17 7 FreeSans 16 270 0 0 y[4]
port 16 nsew
flabel metal2 s 3837 -23 3843 -17 7 FreeSans 16 270 0 0 y[3]
port 17 nsew
flabel metal2 s 3917 -23 3923 -17 7 FreeSans 16 270 0 0 y[0]
port 20 nsew
flabel metal2 s 3637 -23 3643 -17 7 FreeSans 16 270 0 0 y[5]
port 15 nsew
flabel metal2 s 3577 -23 3583 -17 7 FreeSans 16 270 0 0 y[2]
port 18 nsew
flabel metal2 s 3457 -23 3463 -17 7 FreeSans 16 270 0 0 y[1]
port 19 nsew
flabel metal3 s -24 6096 -16 6104 7 FreeSans 16 0 0 0 ready
port 3 nsew
flabel metal2 s 277 6297 283 6303 3 FreeSans 16 90 0 0 x[0]
port 12 nsew
flabel metal2 s 457 6297 463 6303 3 FreeSans 16 90 0 0 x[7]
port 5 nsew
flabel metal2 s 537 6297 543 6303 3 FreeSans 16 90 0 0 x[2]
port 10 nsew
<< properties >>
string FIXED_BBOX -40 -40 7920 6300
<< end >>
