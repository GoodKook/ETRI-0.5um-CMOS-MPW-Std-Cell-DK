magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -56 -56 114 114
<< genericcontact >>
rect 12 40 18 46
rect 40 40 46 46
rect 12 12 18 18
rect 40 12 46 18
<< metal1 >>
rect 4 4 54 54
<< end >>
