magic
tech scmos
magscale 1 30
timestamp 1727158408
<< checkpaint >>
rect 87840 95160 90705 95248
rect -1545 81690 93660 95160
rect -1545 80760 93930 81690
rect -1545 77025 94305 80760
rect -1545 76965 94125 77025
rect -1545 22260 93660 76965
rect -1545 22080 93810 22260
rect -1545 20205 94350 22080
rect -1545 19665 94095 20205
rect -1545 -960 93660 19665
rect 69545 -980 71175 -960
<< error_p >>
rect 42495 88995 42705 89205
rect 51495 82995 51705 83205
rect 25695 45195 25905 45405
rect 29295 37395 29505 37605
rect 63495 29595 63705 29805
rect 79395 17295 79605 17505
rect 62295 13995 62505 14205
rect 8595 1695 8805 1905
<< nwell >>
rect 88955 93240 90005 93360
rect 33000 56265 33225 56340
<< metal1 >>
rect -945 93630 450 93870
rect -945 86070 -45 93630
rect 34305 92055 34995 92145
rect 38205 92055 39795 92145
rect 84105 92055 85395 92145
rect 58695 91845 58905 91995
rect 58455 91800 58905 91845
rect 58455 91755 58845 91800
rect 58455 91305 58545 91755
rect 60405 91845 60600 91905
rect 88500 91845 88695 91905
rect 60405 91695 60645 91845
rect 60555 91305 60645 91695
rect 88455 91695 88695 91845
rect 68805 91545 69000 91605
rect 68805 91455 69210 91545
rect 68805 91395 69000 91455
rect 88455 91305 88545 91695
rect 58455 91155 58695 91305
rect 58500 91095 58695 91155
rect 60555 91155 60795 91305
rect 60600 91095 60795 91155
rect 70800 91245 70995 91305
rect 70755 91155 70995 91245
rect 70800 91095 70995 91155
rect 88455 91155 88695 91305
rect 88500 91095 88695 91155
rect 77805 90855 78795 90945
rect 92145 89970 93045 93870
rect 91650 89730 93045 89970
rect 42915 89055 43395 89145
rect 32205 88755 32895 88845
rect 42105 88755 42795 88845
rect 64305 88755 65295 88845
rect 3105 88545 3300 88605
rect 55500 88545 55695 88605
rect 3105 88395 3345 88545
rect 3255 88005 3345 88395
rect 55455 88395 55695 88545
rect 79605 88545 79800 88605
rect 84300 88545 84495 88605
rect 79605 88395 79845 88545
rect 55455 88005 55545 88395
rect 79755 88005 79845 88395
rect 3105 87855 3345 88005
rect 3105 87795 3300 87855
rect 44805 87855 45195 87945
rect 55200 87990 55545 88005
rect 55305 87855 55545 87990
rect 55305 87795 55500 87855
rect 79605 87855 79845 88005
rect 84255 88395 84495 88545
rect 84255 88005 84345 88395
rect 84255 87855 84495 88005
rect 79605 87795 79800 87855
rect 84300 87795 84495 87855
rect 38805 87555 39795 87645
rect 62805 87555 63495 87645
rect 81705 87555 82695 87645
rect -945 85830 450 86070
rect -945 78270 -45 85830
rect 5805 84255 6495 84345
rect 34005 84255 34395 84345
rect 45105 84255 45795 84345
rect 73305 84255 73695 84345
rect 33195 84045 33405 84195
rect 7905 83955 8745 84045
rect 33195 84000 33645 84045
rect 33255 83955 33645 84000
rect 7905 83355 8295 83445
rect 8655 83205 8745 83955
rect 33555 83445 33645 83955
rect 65805 83955 66645 84045
rect 66555 83505 66645 83955
rect 72405 83955 73245 84045
rect 73155 83505 73245 83955
rect 82200 83745 82395 83805
rect 79905 83655 80610 83745
rect 82155 83655 82395 83745
rect 82200 83595 82395 83655
rect 33555 83355 34095 83445
rect 66555 83355 66795 83505
rect 66600 83295 66795 83355
rect 73155 83355 73395 83505
rect 73200 83295 73395 83355
rect 8400 83190 8745 83205
rect 8505 83055 8745 83190
rect 8505 82995 8700 83055
rect 16605 83055 17295 83145
rect 51915 83055 52395 83145
rect 77205 83055 77895 83145
rect 78105 83055 78495 83145
rect 24705 82755 25695 82845
rect 28905 82455 29595 82545
rect 92145 82170 93045 89730
rect 91650 81930 93045 82170
rect 16155 80145 16245 80895
rect 39000 80745 39195 80805
rect 38955 80595 39195 80745
rect 40605 80745 40800 80805
rect 40605 80595 40845 80745
rect 42705 80745 42900 80805
rect 44400 80745 44595 80805
rect 42705 80595 42945 80745
rect 38955 80205 39045 80595
rect 40755 80205 40845 80595
rect 42855 80205 42945 80595
rect 16155 80055 16995 80145
rect 22755 80055 23295 80145
rect 38955 80055 39195 80205
rect 39000 79995 39195 80055
rect 40605 80055 40845 80205
rect 40605 79995 40800 80055
rect 42705 80055 42945 80205
rect 44355 80595 44595 80745
rect 47805 80745 48000 80805
rect 50700 80745 50895 80805
rect 47805 80595 48045 80745
rect 44355 80205 44445 80595
rect 47955 80205 48045 80595
rect 44355 80055 44595 80205
rect 42705 79995 42900 80055
rect 44400 79995 44595 80055
rect 47805 80055 48045 80205
rect 50655 80595 50895 80745
rect 54705 80745 54900 80805
rect 54705 80595 54945 80745
rect 65505 80745 65700 80805
rect 65505 80595 65745 80745
rect 50655 80205 50745 80595
rect 54855 80205 54945 80595
rect 65655 80205 65745 80595
rect 83955 80655 84495 80745
rect 83955 80205 84045 80655
rect 50655 80055 50895 80205
rect 47805 79995 48000 80055
rect 50700 79995 50895 80055
rect 54705 80055 54945 80205
rect 54705 79995 54900 80055
rect 63705 80055 64095 80145
rect 65505 80055 65745 80205
rect 65505 79995 65700 80055
rect 83805 80055 84045 80205
rect 83805 79995 84000 80055
rect 16905 79755 17295 79845
rect 29805 79755 30795 79845
rect 35805 79755 37695 79845
rect 48105 79755 49095 79845
rect 49905 79755 50595 79845
rect 70605 79755 71595 79845
rect 38505 79455 39495 79545
rect -945 78030 450 78270
rect -945 70470 -45 78030
rect 62505 77655 62895 77745
rect 59955 76455 60795 76545
rect 25200 76245 25395 76305
rect 25155 76095 25395 76245
rect 36705 76245 36900 76305
rect 36705 76095 36945 76245
rect 39105 76155 39645 76245
rect 25155 75705 25245 76095
rect 36855 75705 36945 76095
rect 39555 75705 39645 76155
rect 48105 76155 48495 76245
rect 52905 76155 53295 76245
rect 55005 76245 55200 76305
rect 55005 76095 55245 76245
rect 55155 75705 55245 76095
rect 59955 75705 60045 76455
rect 75855 76455 76695 76545
rect 62700 76245 62895 76305
rect 17505 75555 17895 75645
rect 25155 75555 25395 75705
rect 25200 75495 25395 75555
rect 36855 75555 37095 75705
rect 36900 75495 37095 75555
rect 39555 75555 39795 75705
rect 39600 75495 39795 75555
rect 41205 75555 41595 75645
rect 55005 75555 55245 75705
rect 55005 75495 55200 75555
rect 59805 75555 60045 75705
rect 62655 76095 62895 76245
rect 69600 76245 69795 76305
rect 69555 76095 69795 76245
rect 71505 76245 71700 76305
rect 71505 76095 71745 76245
rect 62655 75705 62745 76095
rect 69555 75705 69645 76095
rect 71655 75705 71745 76095
rect 75855 75705 75945 76455
rect 78105 76245 78300 76305
rect 80700 76245 80895 76305
rect 78105 76095 78345 76245
rect 62655 75555 62895 75705
rect 59805 75495 60000 75555
rect 62700 75495 62895 75555
rect 69555 75555 69795 75705
rect 69600 75495 69795 75555
rect 71655 75555 71895 75705
rect 71700 75495 71895 75555
rect 75705 75555 75945 75705
rect 75705 75495 75900 75555
rect 21105 75255 23295 75345
rect 48405 75255 48795 75345
rect 78255 75345 78345 76095
rect 80655 76095 80895 76245
rect 80655 75645 80745 76095
rect 80205 75555 80745 75645
rect 78255 75255 78795 75345
rect 92145 74370 93045 81930
rect 91650 74130 93045 74370
rect 85905 73755 86295 73845
rect 31605 73155 31995 73245
rect 39405 73155 40095 73245
rect 61155 73155 62295 73245
rect 41205 72945 41400 73005
rect 42000 72945 42195 73005
rect 41205 72795 41445 72945
rect 41355 72405 41445 72795
rect 38655 72255 39195 72345
rect 41205 72255 41445 72405
rect 41955 72795 42195 72945
rect 50400 72945 50595 73005
rect 46005 72855 46545 72945
rect 41205 72195 41400 72255
rect 13905 71955 15195 72045
rect 34305 71955 34995 72045
rect 41955 72090 42045 72795
rect 46455 72345 46545 72855
rect 50355 72795 50595 72945
rect 54105 72945 54300 73005
rect 54105 72795 54345 72945
rect 46455 72255 46845 72345
rect 46755 72105 46845 72255
rect 46755 71955 46995 72105
rect 46800 71895 46995 71955
rect 50355 72045 50445 72795
rect 54255 72405 54345 72795
rect 54105 72255 54345 72405
rect 61155 72405 61245 73155
rect 69705 73155 70395 73245
rect 79155 73155 79995 73245
rect 65205 72945 65400 73005
rect 67800 72945 67995 73005
rect 65205 72795 65445 72945
rect 65355 72405 65445 72795
rect 67755 72795 67995 72945
rect 69900 72945 70095 73005
rect 69855 72795 70095 72945
rect 72405 72945 72600 73005
rect 72405 72795 72645 72945
rect 77100 72945 77295 73005
rect 73905 72855 74445 72945
rect 67755 72405 67845 72795
rect 69855 72405 69945 72795
rect 72555 72405 72645 72795
rect 61155 72255 61395 72405
rect 54105 72195 54300 72255
rect 61200 72195 61395 72255
rect 65205 72255 65445 72405
rect 65205 72195 65400 72255
rect 67605 72255 67845 72405
rect 67605 72195 67800 72255
rect 69705 72255 69945 72405
rect 69705 72195 69900 72255
rect 72405 72255 72645 72405
rect 74355 72405 74445 72855
rect 77055 72795 77295 72945
rect 77055 72405 77145 72795
rect 79155 72405 79245 73155
rect 81600 72945 81795 73005
rect 74355 72255 74595 72405
rect 72405 72195 72600 72255
rect 74400 72195 74595 72255
rect 77055 72255 77295 72405
rect 77100 72195 77295 72255
rect 79005 72255 79245 72405
rect 81555 72795 81795 72945
rect 88005 72855 89145 72945
rect 81555 72405 81645 72795
rect 90900 72645 91095 72705
rect 90690 72555 91095 72645
rect 90900 72495 91095 72555
rect 81555 72255 81795 72405
rect 79005 72195 79200 72255
rect 81600 72195 81795 72255
rect 88005 72255 88395 72345
rect 49905 71955 50445 72045
rect 76005 71955 76695 72045
rect 85305 71955 86295 72045
rect 67305 71355 67695 71445
rect -945 70230 450 70470
rect -945 62670 -45 70230
rect 77805 69855 78795 69945
rect 70005 69255 70995 69345
rect 6105 68655 7095 68745
rect 43500 68745 43695 68805
rect 43455 68595 43695 68745
rect 75600 68745 75795 68805
rect 75555 68595 75795 68745
rect 19605 68445 19800 68505
rect 19605 68295 19845 68445
rect 36705 68445 36900 68505
rect 41700 68445 41895 68505
rect 36705 68295 36945 68445
rect 14190 68055 14895 68145
rect 9195 67845 9405 67995
rect 19755 67905 19845 68295
rect 36855 68145 36945 68295
rect 41655 68295 41895 68445
rect 43455 68445 43545 68595
rect 43155 68355 43545 68445
rect 39000 68145 39195 68205
rect 36855 68055 37410 68145
rect 38955 68055 39195 68145
rect 39000 67995 39195 68055
rect 41655 67905 41745 68295
rect 9195 67800 9795 67845
rect 9255 67755 9795 67800
rect 12405 67845 12600 67905
rect 12405 67755 12645 67845
rect 19755 67755 19995 67905
rect 12405 67695 12600 67755
rect 19800 67695 19995 67755
rect 21405 67755 21795 67845
rect 41505 67755 41745 67905
rect 43155 67905 43245 68355
rect 70305 68445 70500 68505
rect 70305 68295 70545 68445
rect 50205 68145 50400 68205
rect 52200 68145 52395 68205
rect 50205 68055 50445 68145
rect 51990 68055 52395 68145
rect 50205 67995 50400 68055
rect 52200 67995 52395 68055
rect 43155 67755 43395 67905
rect 41505 67695 41700 67755
rect 43200 67695 43395 67755
rect 52755 67605 52845 68295
rect 70455 67905 70545 68295
rect 71205 68145 71400 68205
rect 71205 68055 71445 68145
rect 72990 68055 73545 68145
rect 71205 67995 71400 68055
rect 70305 67755 70545 67905
rect 73455 67905 73545 68055
rect 75555 67905 75645 68595
rect 75900 68445 76095 68505
rect 73455 67755 73695 67905
rect 70305 67695 70500 67755
rect 73500 67695 73695 67755
rect 75405 67755 75645 67905
rect 75855 68295 76095 68445
rect 82305 68355 82845 68445
rect 75855 67905 75945 68295
rect 75855 67755 76095 67905
rect 75405 67695 75600 67755
rect 75900 67695 76095 67755
rect 82755 67845 82845 68355
rect 84705 68355 85545 68445
rect 85455 68145 85545 68355
rect 85455 68055 86010 68145
rect 89955 67905 90045 68595
rect 82755 67755 83145 67845
rect 87555 67755 88395 67845
rect 25605 67455 26595 67545
rect 30105 67455 30795 67545
rect 52605 67455 52845 67605
rect 83055 67605 83145 67755
rect 89805 67755 90045 67905
rect 89805 67695 90000 67755
rect 83055 67455 83295 67605
rect 52605 67395 52800 67455
rect 83100 67395 83295 67455
rect 92145 66570 93045 74130
rect 91650 66330 93045 66570
rect 18705 65955 19095 66045
rect 6705 65145 6900 65205
rect 6705 64995 6945 65145
rect 37005 65145 37200 65205
rect 37005 64995 37245 65145
rect 39555 65055 40095 65145
rect 65955 65055 66495 65145
rect 6855 64545 6945 64995
rect 23400 64845 23595 64905
rect 23355 64755 23595 64845
rect 23400 64695 23595 64755
rect 6855 64455 7245 64545
rect 13755 64455 14295 64545
rect 7155 64305 7245 64455
rect 21600 64590 21900 64605
rect 21705 64545 21900 64590
rect 37155 64545 37245 64995
rect 37605 64845 37800 64905
rect 37605 64755 38010 64845
rect 37605 64695 37800 64755
rect 65955 64545 66045 65055
rect 68955 65145 69045 65595
rect 70305 65355 71595 65445
rect 78405 65355 79395 65445
rect 68505 65055 69045 65145
rect 70905 65055 71445 65145
rect 21705 64455 21945 64545
rect 37155 64455 37545 64545
rect 65355 64455 66045 64545
rect 71355 64605 71445 65055
rect 74655 65055 75195 65145
rect 74655 64605 74745 65055
rect 76905 65055 77445 65145
rect 71355 64455 71595 64605
rect 21705 64395 21900 64455
rect 7155 64155 7395 64305
rect 7200 64095 7395 64155
rect 21555 64245 21645 64380
rect 37455 64305 37545 64455
rect 71400 64395 71595 64455
rect 74505 64455 74745 64605
rect 77355 64605 77445 65055
rect 80505 65145 80700 65205
rect 80505 64995 80745 65145
rect 82905 65055 83295 65145
rect 85500 65145 85695 65205
rect 85455 64995 85695 65145
rect 87405 65145 87600 65205
rect 87405 64995 87645 65145
rect 80655 64605 80745 64995
rect 77355 64455 77595 64605
rect 74505 64395 74700 64455
rect 77400 64395 77595 64455
rect 80505 64455 80745 64605
rect 85455 64545 85545 64995
rect 87555 64545 87645 64995
rect 85455 64455 85845 64545
rect 80505 64395 80700 64455
rect 85755 64305 85845 64455
rect 87255 64455 87645 64545
rect 87255 64305 87345 64455
rect 20505 64155 21645 64245
rect 30405 64155 31695 64245
rect 37455 64155 37695 64305
rect 37500 64095 37695 64155
rect 67905 64155 68895 64245
rect 70005 64155 71295 64245
rect 85755 64155 85995 64305
rect 85800 64095 85995 64155
rect 87105 64155 87345 64305
rect 87105 64095 87300 64155
rect -945 62430 450 62670
rect -945 54870 -45 62430
rect 40005 61395 40095 61605
rect 3105 60855 4095 60945
rect 26805 60855 27795 60945
rect 29505 60855 30195 60945
rect 35505 60855 35895 60945
rect 61305 60855 62295 60945
rect 64905 60855 66195 60945
rect 78105 60855 79395 60945
rect 85605 60855 86295 60945
rect 88905 60855 89895 60945
rect 90255 60855 91095 60945
rect 13200 60645 13395 60705
rect 13155 60555 13395 60645
rect 13200 60495 13395 60555
rect 23700 60645 23895 60705
rect 23655 60495 23895 60645
rect 25005 60645 25200 60705
rect 27900 60645 28095 60705
rect 25005 60495 25245 60645
rect 16200 60345 16395 60405
rect 15990 60255 16395 60345
rect 16200 60195 16395 60255
rect 23655 60105 23745 60495
rect 7005 59955 7695 60045
rect 23655 59955 23895 60105
rect 23700 59895 23895 59955
rect 25155 60045 25245 60495
rect 27855 60495 28095 60645
rect 29700 60645 29895 60705
rect 29655 60495 29895 60645
rect 31455 60555 31995 60645
rect 27855 60105 27945 60495
rect 25155 59955 25995 60045
rect 27705 59955 27945 60105
rect 27705 59895 27900 59955
rect 29655 59805 29745 60495
rect 31455 60105 31545 60555
rect 41805 60645 42000 60705
rect 44100 60645 44295 60705
rect 41805 60495 42045 60645
rect 41955 60105 42045 60495
rect 31305 59955 31545 60105
rect 31305 59895 31500 59955
rect 41805 59955 42045 60105
rect 44055 60495 44295 60645
rect 63705 60645 63900 60705
rect 63705 60495 63945 60645
rect 69405 60645 69600 60705
rect 76500 60645 76695 60705
rect 69405 60495 69645 60645
rect 44055 60105 44145 60495
rect 44055 59955 44295 60105
rect 41805 59895 42000 59955
rect 44100 59895 44295 59955
rect 63855 59805 63945 60495
rect 29505 59655 29745 59805
rect 29505 59595 29700 59655
rect 35205 59655 35595 59745
rect 67605 59655 68295 59745
rect 69555 59490 69645 60495
rect 76455 60495 76695 60645
rect 81105 60645 81300 60705
rect 90255 60645 90345 60855
rect 81105 60495 81405 60645
rect 76455 60345 76545 60495
rect 81195 60405 81405 60495
rect 89955 60555 90345 60645
rect 83100 60345 83295 60405
rect 75690 60255 76545 60345
rect 82890 60255 83295 60345
rect 76455 60105 76545 60255
rect 83100 60195 83295 60255
rect 89955 60105 90045 60555
rect 73905 60045 74100 60105
rect 73905 59955 74145 60045
rect 76455 59955 76695 60105
rect 73905 59895 74100 59955
rect 76500 59895 76695 59955
rect 80205 59955 81345 60045
rect 89955 59955 90195 60105
rect 90000 59895 90195 59955
rect 92145 58770 93045 66330
rect 91650 58530 93045 58770
rect 39405 58155 39795 58245
rect 39705 57855 40695 57945
rect 85305 57855 85695 57945
rect 22605 57555 23145 57645
rect 11400 57345 11595 57405
rect 11355 57195 11595 57345
rect 13005 57255 13395 57345
rect 18300 57345 18495 57405
rect 18255 57195 18495 57345
rect 11355 56805 11445 57195
rect 18255 56805 18345 57195
rect 20355 56805 20445 57195
rect 23055 56805 23145 57555
rect 28800 57645 28995 57705
rect 24405 57555 24945 57645
rect 24855 56805 24945 57555
rect 28755 57495 28995 57645
rect 74505 57555 74895 57645
rect 75105 57555 75495 57645
rect 87105 57555 88095 57645
rect 28755 56805 28845 57495
rect 29100 57345 29295 57405
rect 11355 56655 11595 56805
rect 11400 56595 11595 56655
rect 18255 56655 18495 56805
rect 18300 56595 18495 56655
rect 20355 56655 20595 56805
rect 20400 56595 20595 56655
rect 23055 56655 23295 56805
rect 23100 56595 23295 56655
rect 24705 56655 24945 56805
rect 24705 56595 24900 56655
rect 28605 56655 28845 56805
rect 29055 57195 29295 57345
rect 31155 57255 31995 57345
rect 29055 56805 29145 57195
rect 31155 56805 31245 57255
rect 42000 57345 42195 57405
rect 41955 57195 42195 57345
rect 59805 57345 60000 57405
rect 59805 57195 60045 57345
rect 85305 57255 85845 57345
rect 29055 56655 29295 56805
rect 28605 56595 28800 56655
rect 29100 56595 29295 56655
rect 31005 56655 31245 56805
rect 31005 56595 31200 56655
rect 13905 56355 14595 56445
rect 25905 56355 26295 56445
rect 31305 56355 31995 56445
rect 41955 56490 42045 57195
rect 59955 56790 60045 57195
rect 85755 56805 85845 57255
rect 87405 57345 87600 57405
rect 87405 57195 87645 57345
rect 89205 57345 89400 57405
rect 89205 57195 89445 57345
rect 87555 56805 87645 57195
rect 89355 56805 89445 57195
rect 85755 56655 85995 56805
rect 85800 56595 85995 56655
rect 87555 56655 87795 56805
rect 87600 56595 87795 56655
rect 89205 56655 89445 56805
rect 89205 56595 89400 56655
rect 46005 56355 46995 56445
rect 84405 56355 86295 56445
rect 87105 56355 88095 56445
rect -945 54630 450 54870
rect -945 47070 -45 54630
rect 40305 54255 40695 54345
rect 28005 53655 28995 53745
rect 23505 53355 24795 53445
rect 1005 53055 1995 53145
rect 7605 53055 8895 53145
rect 28755 53055 29295 53145
rect 24300 52845 24495 52905
rect 24255 52695 24495 52845
rect 28755 52845 28845 53055
rect 42105 53055 42795 53145
rect 82305 53055 82995 53145
rect 84855 53055 85695 53145
rect 30600 52845 30795 52905
rect 28455 52800 28845 52845
rect 28395 52755 28845 52800
rect 24255 52305 24345 52695
rect 28395 52590 28605 52755
rect 30555 52695 30795 52845
rect 56805 52755 57195 52845
rect 66900 52845 67095 52905
rect 66855 52695 67095 52845
rect 79800 52845 79995 52905
rect 79755 52695 79995 52845
rect 30555 52305 30645 52695
rect 66855 52305 66945 52695
rect 24255 52155 24495 52305
rect 24300 52095 24495 52155
rect 30555 52155 30795 52305
rect 30600 52095 30795 52155
rect 66705 52155 66945 52305
rect 79755 52305 79845 52695
rect 84855 52305 84945 53055
rect 89655 52755 90195 52845
rect 89655 52305 89745 52755
rect 79755 52155 79995 52305
rect 66705 52095 66900 52155
rect 79800 52095 79995 52155
rect 84705 52155 84945 52305
rect 84705 52095 84900 52155
rect 89505 52155 89745 52305
rect 89505 52095 89700 52155
rect 34005 51855 35295 51945
rect 92145 50970 93045 58530
rect 91650 50730 93045 50970
rect 37605 50355 38295 50445
rect 45555 49905 45645 50295
rect 35400 49845 35595 49905
rect 35355 49695 35595 49845
rect 9105 49545 9300 49605
rect 9600 49545 9795 49605
rect 9105 49395 9345 49545
rect 9255 49005 9345 49395
rect 9105 48855 9345 49005
rect 9555 49395 9795 49545
rect 11505 49545 11700 49605
rect 23100 49545 23295 49605
rect 11505 49395 11745 49545
rect 9105 48795 9300 48855
rect 9555 48705 9645 49395
rect 11655 49005 11745 49395
rect 11505 48855 11745 49005
rect 23055 49395 23295 49545
rect 24405 49545 24600 49605
rect 24405 49395 24645 49545
rect 29205 49545 29400 49605
rect 29205 49395 29445 49545
rect 23055 49005 23145 49395
rect 23055 48855 23295 49005
rect 11505 48795 11700 48855
rect 23100 48795 23295 48855
rect 7005 48555 7695 48645
rect 18105 48555 19095 48645
rect 24555 48645 24645 49395
rect 29355 49005 29445 49395
rect 29205 48855 29445 49005
rect 35355 48945 35445 49695
rect 35700 49545 35895 49605
rect 35055 48855 35445 48945
rect 35655 49395 35895 49545
rect 39705 49545 39900 49605
rect 39705 49395 39945 49545
rect 43305 49545 43500 49605
rect 50400 49545 50595 49605
rect 43305 49395 43545 49545
rect 35655 49005 35745 49395
rect 39855 49005 39945 49395
rect 43455 49245 43545 49395
rect 50355 49395 50595 49545
rect 61005 49545 61200 49605
rect 61005 49395 61245 49545
rect 43455 49155 43845 49245
rect 35655 48855 35895 49005
rect 29205 48795 29400 48855
rect 35055 48705 35145 48855
rect 35700 48795 35895 48855
rect 39705 48855 39945 49005
rect 43755 49005 43845 49155
rect 50355 49005 50445 49395
rect 61155 49005 61245 49395
rect 72555 49455 73095 49545
rect 72555 49005 72645 49455
rect 43755 48855 43995 49005
rect 39705 48795 39900 48855
rect 43800 48795 43995 48855
rect 50355 48855 50595 49005
rect 50400 48795 50595 48855
rect 61005 48855 61245 49005
rect 66000 48945 66195 49005
rect 61005 48795 61200 48855
rect 65955 48795 66195 48945
rect 72405 48855 72645 49005
rect 72405 48795 72600 48855
rect 77355 48945 77445 49695
rect 83205 49545 83400 49605
rect 83205 49395 83445 49545
rect 83355 49005 83445 49395
rect 89505 49455 90045 49545
rect 76605 48855 77445 48945
rect 83205 48855 83445 49005
rect 89955 48945 90045 49455
rect 89955 48855 90345 48945
rect 83205 48795 83400 48855
rect 24555 48555 25395 48645
rect 35205 48555 36195 48645
rect 37605 48555 38295 48645
rect 58305 48555 59895 48645
rect 65955 48390 66045 48795
rect 66405 48555 66795 48645
rect 74205 48555 75195 48645
rect 90255 48645 90345 48855
rect 90255 48600 90645 48645
rect 90255 48555 90705 48600
rect 90495 48390 90705 48555
rect 84705 47955 85095 48045
rect -945 46830 450 47070
rect -945 39270 -45 46830
rect 31605 46455 32295 46545
rect 4305 45255 5895 45345
rect 25005 45255 25695 45345
rect 29205 45255 30495 45345
rect 40905 45255 41295 45345
rect 42405 45255 43395 45345
rect 16305 45045 16500 45105
rect 16305 44895 16545 45045
rect 16455 44505 16545 44895
rect 20355 44955 21195 45045
rect 20355 44505 20445 44955
rect 27405 44955 27795 45045
rect 29505 45045 29700 45105
rect 32400 45045 32595 45105
rect 29505 44895 29745 45045
rect 12105 44355 12795 44445
rect 16305 44355 16545 44505
rect 16305 44295 16500 44355
rect 20205 44355 20445 44505
rect 20205 44295 20400 44355
rect 29655 44205 29745 44895
rect 32355 44895 32595 45045
rect 38400 45045 38595 45105
rect 38355 44895 38595 45045
rect 45600 45045 45795 45105
rect 45555 44895 45795 45045
rect 47400 45045 47595 45105
rect 47355 44895 47595 45045
rect 49305 45045 49500 45105
rect 60000 45045 60195 45105
rect 49305 44895 49545 45045
rect 32355 44505 32445 44895
rect 32355 44355 32595 44505
rect 32400 44295 32595 44355
rect 33705 44055 34995 44145
rect 38355 44145 38445 44895
rect 38355 44055 38895 44145
rect 45555 44190 45645 44895
rect 47355 44505 47445 44895
rect 49455 44505 49545 44895
rect 47355 44355 47595 44505
rect 47400 44295 47595 44355
rect 49305 44355 49545 44505
rect 59955 44895 60195 45045
rect 61605 44955 62445 45045
rect 59955 44505 60045 44895
rect 62355 44505 62445 44955
rect 64305 45045 64500 45105
rect 79800 45045 79995 45105
rect 64305 44895 64545 45045
rect 64455 44505 64545 44895
rect 79755 44895 79995 45045
rect 84600 45045 84795 45105
rect 84555 44895 84795 45045
rect 79755 44505 79845 44895
rect 59955 44355 60195 44505
rect 49305 44295 49500 44355
rect 60000 44295 60195 44355
rect 62355 44355 62595 44505
rect 62400 44295 62595 44355
rect 64455 44355 64695 44505
rect 64500 44295 64695 44355
rect 74205 44355 74595 44445
rect 79755 44355 79995 44505
rect 79800 44295 79995 44355
rect 84555 44445 84645 44895
rect 84105 44355 84645 44445
rect 77505 44055 78195 44145
rect 87405 43755 88095 43845
rect 92145 43170 93045 50730
rect 91650 42930 93045 43170
rect 24705 42255 25695 42345
rect 83055 42105 83145 42495
rect 85095 42405 85305 42495
rect 85005 42300 85305 42405
rect 85005 42255 85245 42300
rect 85005 42195 85200 42255
rect 22305 41955 22695 42045
rect 23055 41955 23895 42045
rect 14400 41745 14595 41805
rect 14355 41595 14595 41745
rect 14355 41205 14445 41595
rect 14355 41055 14595 41205
rect 14400 40995 14595 41055
rect 6405 40755 7995 40845
rect 13305 40755 14295 40845
rect 23055 40890 23145 41955
rect 28905 41955 29895 42045
rect 37005 41955 37995 42045
rect 80505 41955 81495 42045
rect 82905 41955 83145 42105
rect 82905 41895 83100 41955
rect 24855 41655 25695 41745
rect 24855 41205 24945 41655
rect 31500 41745 31695 41805
rect 31455 41700 31695 41745
rect 31395 41595 31695 41700
rect 33600 41745 33795 41805
rect 33555 41595 33795 41745
rect 37155 41655 37695 41745
rect 31395 41490 31605 41595
rect 24705 41055 24945 41205
rect 33555 41205 33645 41595
rect 37155 41205 37245 41655
rect 41700 41745 41895 41805
rect 41655 41595 41895 41745
rect 45705 41745 45900 41805
rect 49200 41745 49395 41805
rect 45705 41595 45945 41745
rect 38895 41205 39105 41295
rect 41655 41205 41745 41595
rect 45855 41205 45945 41595
rect 49155 41595 49395 41745
rect 76500 41745 76695 41805
rect 76455 41595 76695 41745
rect 78405 41745 78600 41805
rect 78405 41595 78645 41745
rect 80205 41745 80400 41805
rect 80205 41595 80445 41745
rect 80655 41700 81195 41745
rect 46605 41445 46800 41505
rect 48600 41445 48795 41505
rect 46605 41355 47010 41445
rect 48555 41355 48795 41445
rect 46605 41295 46800 41355
rect 48600 41295 48795 41355
rect 33555 41055 33795 41205
rect 24705 40995 24900 41055
rect 33600 40995 33795 41055
rect 37005 41055 37245 41205
rect 37005 40995 37200 41055
rect 38805 41100 39105 41205
rect 38805 41055 39045 41100
rect 38805 40995 39000 41055
rect 41505 41055 41745 41205
rect 41505 40995 41700 41055
rect 45705 41055 45945 41205
rect 49155 41205 49245 41595
rect 76455 41505 76545 41595
rect 76200 41490 76545 41505
rect 76305 41355 76545 41490
rect 76305 41295 76500 41355
rect 78555 41205 78645 41595
rect 80355 41205 80445 41595
rect 80595 41655 81195 41700
rect 80595 41505 80805 41655
rect 83355 41205 83445 42195
rect 86505 41955 87195 42045
rect 88605 41955 89145 42045
rect 84900 41745 85095 41805
rect 49155 41055 49395 41205
rect 45705 40995 45900 41055
rect 49200 40995 49395 41055
rect 76605 41145 76800 41205
rect 76605 41100 76845 41145
rect 76605 40995 76905 41100
rect 78555 41055 78795 41205
rect 78600 40995 78795 41055
rect 80205 41055 80445 41205
rect 80205 40995 80400 41055
rect 83205 41055 83445 41205
rect 84855 41595 85095 41745
rect 87105 41745 87300 41805
rect 87105 41595 87345 41745
rect 84855 41205 84945 41595
rect 87255 41205 87345 41595
rect 89055 41205 89145 41955
rect 84855 41055 85095 41205
rect 83205 40995 83400 41055
rect 84900 40995 85095 41055
rect 87105 41055 87345 41205
rect 87105 40995 87300 41055
rect 88905 41055 89145 41205
rect 88905 40995 89100 41055
rect 76695 40905 76905 40995
rect 32805 40755 33195 40845
rect 37305 40755 37995 40845
rect 39405 40755 39795 40845
rect 79905 40755 80595 40845
rect 14205 40155 14595 40245
rect -945 39030 450 39270
rect -945 31470 -45 39030
rect 29505 38055 30495 38145
rect 16605 37755 17595 37845
rect 20505 37455 21495 37545
rect 29715 37455 30795 37545
rect 40605 37455 42795 37545
rect 55005 37455 55995 37545
rect 65805 37455 66345 37545
rect 2505 37245 2700 37305
rect 15300 37245 15495 37305
rect 2505 37095 2745 37245
rect 2655 36705 2745 37095
rect 15255 37095 15495 37245
rect 18405 37245 18600 37305
rect 18405 37200 18645 37245
rect 18405 37095 18705 37200
rect 41400 37245 41595 37305
rect 36405 37155 36945 37245
rect 2655 36555 2895 36705
rect 2700 36495 2895 36555
rect 15255 36345 15345 37095
rect 18495 36990 18705 37095
rect 18855 36705 18945 37095
rect 36855 36705 36945 37155
rect 41355 37095 41595 37245
rect 43905 37245 44100 37305
rect 43905 37095 44145 37245
rect 46605 37245 46800 37305
rect 46605 37095 46845 37245
rect 50505 37245 50700 37305
rect 50505 37095 50745 37245
rect 18855 36555 19095 36705
rect 18900 36495 19095 36555
rect 36855 36555 37095 36705
rect 36900 36495 37095 36555
rect 41355 36645 41445 37095
rect 44055 36705 44145 37095
rect 40905 36555 41445 36645
rect 43905 36555 44145 36705
rect 46755 36705 46845 37095
rect 50655 36705 50745 37095
rect 66255 36705 66345 37455
rect 89655 37455 90195 37545
rect 70305 37245 70500 37305
rect 70305 37095 70545 37245
rect 72405 37245 72600 37305
rect 72405 37095 72645 37245
rect 76605 37245 76800 37305
rect 76605 37095 76845 37245
rect 85305 37245 85500 37305
rect 85305 37095 85545 37245
rect 46755 36555 46995 36705
rect 43905 36495 44100 36555
rect 46800 36495 46995 36555
rect 50655 36555 50895 36705
rect 50700 36495 50895 36555
rect 66105 36555 66345 36705
rect 70455 36645 70545 37095
rect 72555 36705 72645 37095
rect 70455 36555 70995 36645
rect 66105 36495 66300 36555
rect 72405 36555 72645 36705
rect 76755 36705 76845 37095
rect 85455 36705 85545 37095
rect 87555 37155 88095 37245
rect 87555 36705 87645 37155
rect 89655 36705 89745 37455
rect 76755 36555 76995 36705
rect 72405 36495 72600 36555
rect 76800 36495 76995 36555
rect 85455 36555 85695 36705
rect 85500 36495 85695 36555
rect 87405 36555 87645 36705
rect 87405 36495 87600 36555
rect 89505 36555 89745 36705
rect 89505 36495 89700 36555
rect 14805 36255 15345 36345
rect 40905 36255 42195 36345
rect 92145 35370 93045 42930
rect 91650 35130 93045 35370
rect 76305 34755 76695 34845
rect 25305 34455 25995 34545
rect 36105 34155 36795 34245
rect 900 33945 1095 34005
rect 855 33795 1095 33945
rect 7605 33945 7800 34005
rect 16800 33945 16995 34005
rect 7605 33795 7845 33945
rect 855 33345 945 33795
rect 3000 33645 3195 33705
rect 2955 33495 3195 33645
rect 2955 33405 3045 33495
rect 855 33255 1245 33345
rect 1155 33105 1245 33255
rect 2805 33255 3045 33405
rect 7755 33405 7845 33795
rect 16755 33795 16995 33945
rect 25605 33945 25800 34005
rect 25605 33795 25845 33945
rect 30600 33945 30795 34005
rect 30555 33795 30795 33945
rect 7755 33255 7995 33405
rect 2805 33195 3000 33255
rect 7800 33195 7995 33255
rect 12705 33255 13095 33345
rect 16755 33345 16845 33795
rect 25755 33405 25845 33795
rect 16455 33255 16845 33345
rect 1155 33075 1500 33105
rect 1155 32955 1395 33075
rect 1200 32895 1395 32955
rect 16455 33045 16545 33255
rect 23505 33255 24195 33345
rect 25755 33255 25995 33405
rect 25800 33195 25995 33255
rect 28155 33345 28245 33795
rect 27855 33255 28245 33345
rect 30555 33405 30645 33795
rect 32655 33405 32745 34095
rect 35805 33945 36000 34005
rect 35805 33795 36045 33945
rect 40605 33945 40800 34005
rect 40605 33795 40845 33945
rect 48405 33945 48600 34005
rect 48405 33795 48645 33945
rect 60405 33945 60600 34005
rect 60900 33945 61095 34005
rect 60405 33795 60645 33945
rect 30555 33255 30795 33405
rect 15705 32955 16545 33045
rect 27855 33045 27945 33255
rect 30600 33195 30795 33255
rect 32655 33255 32895 33405
rect 32700 33195 32895 33255
rect 35955 33345 36045 33795
rect 40755 33390 40845 33795
rect 48555 33405 48645 33795
rect 35955 33255 36495 33345
rect 48405 33255 48645 33405
rect 58155 33345 58245 33795
rect 60555 33405 60645 33795
rect 58155 33255 58545 33345
rect 48405 33195 48600 33255
rect 27405 32955 28395 33045
rect 58455 33045 58545 33255
rect 60405 33255 60645 33405
rect 60855 33795 61095 33945
rect 73005 33855 73395 33945
rect 76005 33855 76845 33945
rect 60855 33405 60945 33795
rect 76755 33405 76845 33855
rect 60855 33255 61095 33405
rect 60405 33195 60600 33255
rect 60900 33195 61095 33255
rect 76755 33255 76995 33405
rect 76800 33195 76995 33255
rect 58455 32955 58995 33045
rect 80205 32655 81195 32745
rect 29805 32355 31095 32445
rect -945 31230 450 31470
rect -945 23670 -45 31230
rect 23805 30255 24795 30345
rect 32505 30255 33195 30345
rect 67305 30255 67995 30345
rect 37305 29955 37695 30045
rect 51405 29955 51795 30045
rect 85605 29955 86595 30045
rect 9705 29655 10095 29745
rect 13305 29745 13500 29805
rect 13305 29595 13545 29745
rect 15705 29655 16095 29745
rect 27705 29655 28995 29745
rect 34305 29655 34995 29745
rect 36705 29655 37695 29745
rect 13455 29445 13545 29595
rect 62805 29655 63495 29745
rect 68805 29655 69345 29745
rect 26100 29445 26295 29505
rect 13455 29355 13845 29445
rect 13755 28905 13845 29355
rect 26055 29295 26295 29445
rect 30105 29445 30300 29505
rect 30105 29295 30345 29445
rect 41205 29445 41400 29505
rect 41700 29445 41895 29505
rect 41205 29295 41445 29445
rect 26055 28905 26145 29295
rect 30255 28905 30345 29295
rect 13605 28755 13845 28905
rect 13605 28695 13800 28755
rect 25905 28755 26145 28905
rect 25905 28695 26100 28755
rect 30105 28755 30345 28905
rect 30105 28695 30300 28755
rect 41355 28605 41445 29295
rect 41655 29295 41895 29445
rect 64905 29445 65100 29505
rect 64905 29295 65145 29445
rect 41655 28905 41745 29295
rect 41655 28755 41895 28905
rect 41700 28695 41895 28755
rect 65055 28890 65145 29295
rect 69255 28905 69345 29655
rect 79155 29655 79695 29745
rect 79155 29445 79245 29655
rect 83505 29655 84495 29745
rect 85605 29655 86295 29745
rect 69105 28755 69345 28905
rect 78855 29355 79245 29445
rect 69105 28695 69300 28755
rect 41355 28455 41595 28605
rect 41400 28395 41595 28455
rect 44655 28500 45495 28545
rect 44595 28455 45495 28500
rect 44595 28305 44805 28455
rect 67605 28455 67995 28545
rect 78855 28545 78945 29355
rect 80805 29445 81000 29505
rect 84000 29445 84195 29505
rect 80805 29295 81045 29445
rect 80955 28905 81045 29295
rect 80805 28755 81045 28905
rect 83955 29295 84195 29445
rect 88005 29355 88545 29445
rect 83955 28845 84045 29295
rect 88455 28905 88545 29355
rect 83955 28800 84345 28845
rect 83955 28755 84405 28800
rect 88455 28755 88695 28905
rect 80805 28695 81000 28755
rect 84195 28605 84405 28755
rect 88500 28695 88695 28755
rect 78855 28455 79695 28545
rect 85905 28455 86595 28545
rect 92145 27570 93045 35130
rect 91650 27330 93045 27570
rect 80505 26655 80895 26745
rect 2805 26145 3000 26205
rect 2805 25995 3045 26145
rect 5205 26055 5595 26145
rect 2955 25605 3045 25995
rect 24255 25605 24345 26595
rect 53805 26355 54795 26445
rect 29055 26055 29595 26145
rect 26355 25605 26445 25995
rect 2955 25455 3195 25605
rect 3000 25395 3195 25455
rect 24255 25455 24495 25605
rect 24300 25395 24495 25455
rect 26205 25455 26445 25605
rect 29055 25545 29145 26055
rect 31500 26145 31695 26205
rect 31455 25995 31695 26145
rect 33600 26145 33795 26205
rect 33555 25995 33795 26145
rect 52395 26145 52605 26295
rect 78705 26355 79095 26445
rect 56700 26145 56895 26205
rect 52155 26100 52605 26145
rect 52155 26055 52545 26100
rect 31455 25605 31545 25995
rect 28755 25455 29145 25545
rect 26205 25395 26400 25455
rect 28755 25245 28845 25455
rect 31305 25455 31545 25605
rect 33555 25605 33645 25995
rect 52155 25605 52245 26055
rect 56655 25995 56895 26145
rect 62100 26145 62295 26205
rect 62055 25995 62295 26145
rect 68205 26145 68400 26205
rect 68205 25995 68445 26145
rect 78405 25995 78645 26175
rect 56655 25605 56745 25995
rect 62055 25605 62145 25995
rect 33555 25455 33795 25605
rect 31305 25395 31500 25455
rect 33600 25395 33795 25455
rect 52155 25455 52395 25605
rect 52200 25395 52395 25455
rect 56655 25455 56895 25605
rect 56700 25395 56895 25455
rect 62055 25455 62295 25605
rect 62100 25395 62295 25455
rect 28305 25155 28845 25245
rect 31005 25155 31995 25245
rect 41205 25155 41595 25245
rect 66705 25155 67095 25245
rect 68355 25245 68445 25995
rect 78555 25605 78645 25995
rect 81855 26055 82395 26145
rect 81855 25605 81945 26055
rect 78555 25455 78795 25605
rect 78600 25395 78795 25455
rect 81705 25455 81945 25605
rect 81705 25395 81900 25455
rect 68355 25155 68895 25245
rect 25305 24855 26595 24945
rect -945 23430 450 23670
rect -945 15870 -45 23430
rect 51705 23055 52395 23145
rect 28305 22155 29595 22245
rect 17205 21855 18495 21945
rect 24405 21855 24795 21945
rect 26205 21855 27195 21945
rect 64005 21855 65595 21945
rect 71205 21855 71895 21945
rect 90705 21855 91095 21945
rect 29400 21645 29595 21705
rect 29355 21495 29595 21645
rect 33105 21645 33300 21705
rect 43500 21645 43695 21705
rect 33105 21495 33345 21645
rect 29355 21105 29445 21495
rect 33255 21105 33345 21495
rect 8805 20955 9195 21045
rect 29355 20955 29595 21105
rect 29400 20895 29595 20955
rect 33105 20955 33345 21105
rect 43455 21495 43695 21645
rect 49305 21645 49500 21705
rect 49305 21495 49545 21645
rect 51405 21645 51600 21705
rect 51405 21495 51645 21645
rect 43455 21105 43545 21495
rect 43455 20955 43695 21105
rect 33105 20895 33300 20955
rect 43500 20895 43695 20955
rect 49455 21045 49545 21495
rect 51555 21105 51645 21495
rect 69255 21555 69795 21645
rect 69255 21105 69345 21555
rect 78105 21555 78645 21645
rect 49155 21000 49545 21045
rect 49095 20955 49545 21000
rect 49095 20805 49305 20955
rect 51405 20955 51645 21105
rect 51405 20895 51600 20955
rect 69105 20955 69345 21105
rect 78555 21105 78645 21555
rect 79905 21645 80100 21705
rect 79905 21495 80145 21645
rect 80055 21105 80145 21495
rect 78555 20955 78795 21105
rect 69105 20895 69300 20955
rect 78600 20895 78795 20955
rect 80055 20955 80295 21105
rect 80100 20895 80295 20955
rect 91005 20955 91695 21045
rect 22305 20655 22995 20745
rect 51705 20655 52395 20745
rect 89205 20355 89895 20445
rect 92145 19770 93045 27330
rect 91650 19530 93045 19770
rect 66705 18555 67095 18645
rect 34305 18345 34500 18405
rect 45300 18345 45495 18405
rect 34305 18195 34545 18345
rect 705 18045 900 18105
rect 705 17895 945 18045
rect 855 17805 945 17895
rect 855 17655 1095 17805
rect 900 17595 1095 17655
rect 34455 17745 34545 18195
rect 45255 18195 45495 18345
rect 54405 18345 54600 18405
rect 54405 18195 54645 18345
rect 55905 18345 56100 18405
rect 56400 18345 56595 18405
rect 55905 18195 56145 18345
rect 45255 17805 45345 18195
rect 54555 17805 54645 18195
rect 34455 17655 35295 17745
rect 45255 17655 45495 17805
rect 45300 17595 45495 17655
rect 54555 17655 54795 17805
rect 54600 17595 54795 17655
rect 8805 17355 9195 17445
rect 18105 17355 18495 17445
rect 56055 17445 56145 18195
rect 56355 18195 56595 18345
rect 82695 18345 82905 18495
rect 82455 18300 82905 18345
rect 82455 18255 82845 18300
rect 56355 17805 56445 18195
rect 56355 17655 56595 17805
rect 56400 17595 56595 17655
rect 82455 17745 82545 18255
rect 82005 17655 82545 17745
rect 56055 17355 56895 17445
rect 58605 17355 59295 17445
rect 78405 17355 79395 17445
rect 91155 17205 91245 17895
rect -945 15630 450 15870
rect -945 8070 -45 15630
rect 47505 15255 47895 15345
rect 32595 14445 32805 14595
rect 31905 14400 32805 14445
rect 31905 14355 32745 14400
rect 76005 14355 76395 14445
rect 1905 14055 3795 14145
rect 15405 14055 16095 14145
rect 18105 14055 19695 14145
rect 22605 14055 23295 14145
rect 38205 14055 39495 14145
rect 62715 14055 63195 14145
rect 64605 14055 65895 14145
rect 85005 14055 85395 14145
rect 23805 13755 24195 13845
rect 29805 13755 30195 13845
rect 60705 13845 60900 13905
rect 76200 13845 76395 13905
rect 60705 13695 60945 13845
rect 60855 13245 60945 13695
rect 76155 13695 76395 13845
rect 78300 13845 78495 13905
rect 78255 13695 78495 13845
rect 82005 13845 82200 13905
rect 82005 13695 82245 13845
rect 76155 13305 76245 13695
rect 78255 13305 78345 13695
rect 82155 13305 82245 13695
rect 60855 13200 61245 13245
rect 60855 13155 61305 13200
rect 76155 13155 76395 13305
rect 61095 13005 61305 13155
rect 76200 13095 76395 13155
rect 78105 13155 78345 13305
rect 78105 13095 78300 13155
rect 82005 13155 82245 13305
rect 82005 13095 82200 13155
rect 49305 12855 49995 12945
rect 92145 11970 93045 19530
rect 91650 11730 93045 11970
rect 28005 10755 28395 10845
rect 44805 10755 45795 10845
rect 58905 10755 59595 10845
rect 64005 10755 64995 10845
rect 73500 10845 73695 10905
rect 73455 10695 73695 10845
rect 19305 10545 19500 10605
rect 19305 10395 19545 10545
rect 25905 10545 26100 10605
rect 25905 10395 26145 10545
rect 19455 10005 19545 10395
rect 19455 9855 19695 10005
rect 19500 9795 19695 9855
rect 26055 9945 26145 10395
rect 30555 10455 31095 10545
rect 30555 10005 30645 10455
rect 33300 10545 33495 10605
rect 33255 10395 33495 10545
rect 44505 10455 45195 10545
rect 73455 10545 73545 10695
rect 87300 10545 87495 10605
rect 73155 10455 73545 10545
rect 33255 10245 33345 10395
rect 32955 10155 33345 10245
rect 32955 10005 33045 10155
rect 47295 10005 47505 10095
rect 47655 10005 47745 10395
rect 26055 9900 26745 9945
rect 26055 9855 26805 9900
rect 26595 9705 26805 9855
rect 30405 9855 30645 10005
rect 30405 9795 30600 9855
rect 32805 9855 33045 10005
rect 32805 9795 33000 9855
rect 47205 9900 47505 10005
rect 47205 9855 47445 9900
rect 47205 9795 47400 9855
rect 55905 9855 56295 9945
rect 56655 9705 56745 10095
rect 73155 10005 73245 10455
rect 87255 10395 87495 10545
rect 87255 10005 87345 10395
rect 73005 9855 73245 10005
rect 73005 9795 73200 9855
rect 87105 9855 87345 10005
rect 87105 9795 87300 9855
rect 23205 9555 25095 9645
rect 57705 9555 59295 9645
rect -945 7830 450 8070
rect -945 270 -45 7830
rect 7005 6255 7395 6345
rect 31905 6255 34095 6345
rect 40905 6255 41895 6345
rect 42105 6255 43095 6345
rect 88005 6255 88695 6345
rect 22755 5955 23895 6045
rect 33000 6045 33195 6105
rect 32955 5895 33195 6045
rect 48405 6045 48600 6105
rect 48900 6045 49095 6105
rect 48405 5895 48645 6045
rect 32955 5445 33045 5895
rect 48555 5505 48645 5895
rect 32655 5400 33045 5445
rect 32595 5355 33045 5400
rect 32595 5205 32805 5355
rect 48405 5355 48645 5505
rect 48855 5895 49095 6045
rect 48405 5295 48600 5355
rect 48855 5205 48945 5895
rect 13305 5055 13995 5145
rect 25605 5055 26895 5145
rect 48600 5190 48945 5205
rect 48705 5055 48945 5190
rect 48705 4995 48900 5055
rect 54405 5055 55095 5145
rect 30405 4755 30795 4845
rect 25305 4455 26295 4545
rect 92145 4170 93045 11730
rect 91650 3930 93045 4170
rect 24405 3555 25095 3645
rect 42705 2955 43695 3045
rect 22305 2655 22995 2745
rect 38100 2745 38295 2805
rect 38055 2595 38295 2745
rect 44505 2745 44700 2805
rect 44505 2595 44745 2745
rect 62205 2745 62400 2805
rect 66600 2745 66795 2805
rect 62205 2595 62445 2745
rect 38055 2205 38145 2595
rect 31605 2055 31995 2145
rect 37905 2055 38145 2205
rect 44655 2205 44745 2595
rect 60000 2445 60195 2505
rect 59955 2355 60195 2445
rect 60000 2295 60195 2355
rect 44655 2055 44895 2205
rect 37905 1995 38100 2055
rect 44700 1995 44895 2055
rect 62355 2145 62445 2595
rect 66555 2595 66795 2745
rect 66555 2205 66645 2595
rect 57705 2055 58545 2145
rect 62355 2055 62745 2145
rect 8805 1755 10095 1845
rect 15105 1755 16395 1845
rect 17490 1695 17505 1800
rect 17805 1755 18795 1845
rect 31305 1755 32895 1845
rect 62655 1845 62745 2055
rect 66405 2055 66645 2205
rect 66405 1995 66600 2055
rect 62655 1755 63195 1845
rect 89805 1755 91095 1845
rect 17295 1545 17505 1695
rect 17295 1500 18495 1545
rect 17355 1455 18495 1500
rect 42105 555 42495 645
rect -945 30 450 270
rect 92145 30 93045 3930
<< m2contact >>
rect 34095 92010 34305 92220
rect 34995 91995 35205 92205
rect 37995 91995 38205 92205
rect 39795 91995 40005 92205
rect 58695 91995 58905 92205
rect 83895 91995 84105 92205
rect 85395 91995 85605 92205
rect 60195 91695 60405 91905
rect 88695 91695 88905 91905
rect 68595 91395 68805 91605
rect 58695 91095 58905 91305
rect 60795 91095 61005 91305
rect 70995 91095 71205 91305
rect 88695 91095 88905 91305
rect 77595 90795 77805 91005
rect 78795 90795 79005 91005
rect 42705 88995 42915 89205
rect 43395 88995 43605 89205
rect 31995 88695 32205 88905
rect 32895 88695 33105 88905
rect 41895 88695 42105 88905
rect 42795 88695 43005 88905
rect 64095 88695 64305 88905
rect 65295 88695 65505 88905
rect 2895 88395 3105 88605
rect 55695 88395 55905 88605
rect 79395 88395 79605 88605
rect 2895 87795 3105 88005
rect 44595 87795 44805 88005
rect 45195 87795 45405 88005
rect 55095 87780 55305 87990
rect 79395 87795 79605 88005
rect 84495 88395 84705 88605
rect 84495 87795 84705 88005
rect 38595 87495 38805 87705
rect 39795 87495 40005 87705
rect 62595 87495 62805 87705
rect 63495 87495 63705 87705
rect 81495 87495 81705 87705
rect 82695 87495 82905 87705
rect 5595 84195 5805 84405
rect 6495 84195 6705 84405
rect 33195 84195 33405 84405
rect 33795 84195 34005 84405
rect 34395 84195 34605 84405
rect 44895 84195 45105 84405
rect 45795 84195 46005 84405
rect 73095 84195 73305 84405
rect 73695 84210 73905 84420
rect 7695 83895 7905 84105
rect 7695 83295 7905 83505
rect 8295 83295 8505 83505
rect 65595 83895 65805 84105
rect 72195 83895 72405 84105
rect 79695 83595 79905 83805
rect 82395 83595 82605 83805
rect 34095 83295 34305 83505
rect 66795 83295 67005 83505
rect 73395 83295 73605 83505
rect 8295 82980 8505 83190
rect 16395 82995 16605 83205
rect 17295 82995 17505 83205
rect 51705 82995 51915 83205
rect 52395 82995 52605 83205
rect 76995 82995 77205 83205
rect 77895 82995 78105 83205
rect 78495 82995 78705 83205
rect 24495 82695 24705 82905
rect 25695 82695 25905 82905
rect 28695 82395 28905 82605
rect 29595 82395 29805 82605
rect 16095 80895 16305 81105
rect 39195 80595 39405 80805
rect 40395 80595 40605 80805
rect 42495 80595 42705 80805
rect 16995 79995 17205 80205
rect 23295 79995 23505 80205
rect 39195 79995 39405 80205
rect 40395 79995 40605 80205
rect 42495 79995 42705 80205
rect 44595 80595 44805 80805
rect 47595 80595 47805 80805
rect 44595 79995 44805 80205
rect 47595 79995 47805 80205
rect 50895 80595 51105 80805
rect 54495 80595 54705 80805
rect 65295 80595 65505 80805
rect 84495 80595 84705 80805
rect 50895 79995 51105 80205
rect 54495 79995 54705 80205
rect 63495 79995 63705 80205
rect 64095 79995 64305 80205
rect 65295 79995 65505 80205
rect 83595 79995 83805 80205
rect 16695 79695 16905 79905
rect 17295 79695 17505 79905
rect 29595 79695 29805 79905
rect 30795 79695 31005 79905
rect 35595 79695 35805 79905
rect 37695 79695 37905 79905
rect 47895 79695 48105 79905
rect 49095 79695 49305 79905
rect 49695 79695 49905 79905
rect 50595 79680 50805 79890
rect 70395 79695 70605 79905
rect 71595 79695 71805 79905
rect 38295 79395 38505 79605
rect 39495 79395 39705 79605
rect 62295 77595 62505 77805
rect 62895 77595 63105 77805
rect 25395 76095 25605 76305
rect 36495 76095 36705 76305
rect 38895 76095 39105 76305
rect 47895 76095 48105 76305
rect 48495 76095 48705 76305
rect 52695 76095 52905 76305
rect 53295 76080 53505 76290
rect 54795 76095 55005 76305
rect 60795 76395 61005 76605
rect 17295 75495 17505 75705
rect 17895 75495 18105 75705
rect 25395 75495 25605 75705
rect 37095 75495 37305 75705
rect 39795 75495 40005 75705
rect 40995 75495 41205 75705
rect 41595 75495 41805 75705
rect 54795 75495 55005 75705
rect 59595 75495 59805 75705
rect 62895 76095 63105 76305
rect 69795 76095 70005 76305
rect 71295 76095 71505 76305
rect 76695 76395 76905 76605
rect 77895 76095 78105 76305
rect 62895 75495 63105 75705
rect 69795 75495 70005 75705
rect 71895 75495 72105 75705
rect 75495 75495 75705 75705
rect 20895 75195 21105 75405
rect 23295 75195 23505 75405
rect 48195 75195 48405 75405
rect 48795 75195 49005 75405
rect 80895 76095 81105 76305
rect 79995 75495 80205 75705
rect 78795 75195 79005 75405
rect 85695 73695 85905 73905
rect 86295 73695 86505 73905
rect 31395 73095 31605 73305
rect 31995 73095 32205 73305
rect 39195 73080 39405 73290
rect 40095 73095 40305 73305
rect 40995 72795 41205 73005
rect 39195 72195 39405 72405
rect 40995 72195 41205 72405
rect 42195 72795 42405 73005
rect 45795 72795 46005 73005
rect 13695 71895 13905 72105
rect 15195 71895 15405 72105
rect 34095 71895 34305 72105
rect 34995 71895 35205 72105
rect 50595 72795 50805 73005
rect 53895 72795 54105 73005
rect 41895 71880 42105 72090
rect 46995 71895 47205 72105
rect 49695 71895 49905 72105
rect 53895 72195 54105 72405
rect 62295 73095 62505 73305
rect 69495 73095 69705 73305
rect 70395 73095 70605 73305
rect 64995 72795 65205 73005
rect 67995 72795 68205 73005
rect 70095 72795 70305 73005
rect 72195 72795 72405 73005
rect 73695 72795 73905 73005
rect 61395 72195 61605 72405
rect 64995 72195 65205 72405
rect 67395 72195 67605 72405
rect 69495 72195 69705 72405
rect 72195 72195 72405 72405
rect 77295 72795 77505 73005
rect 79995 73095 80205 73305
rect 74595 72195 74805 72405
rect 77295 72195 77505 72405
rect 78795 72195 79005 72405
rect 81795 72795 82005 73005
rect 87795 72795 88005 73005
rect 91095 72495 91305 72705
rect 81795 72195 82005 72405
rect 87795 72195 88005 72405
rect 88395 72195 88605 72405
rect 75795 71895 76005 72105
rect 76695 71895 76905 72105
rect 85095 71895 85305 72105
rect 86295 71895 86505 72105
rect 67095 71295 67305 71505
rect 67695 71295 67905 71505
rect 89895 70695 90105 70905
rect 77595 69795 77805 70005
rect 78795 69795 79005 70005
rect 69795 69195 70005 69405
rect 70995 69195 71205 69405
rect 5895 68610 6105 68820
rect 7095 68595 7305 68805
rect 43695 68595 43905 68805
rect 75795 68595 76005 68805
rect 89895 68595 90105 68805
rect 19395 68295 19605 68505
rect 36495 68295 36705 68505
rect 9195 67995 9405 68205
rect 14895 67995 15105 68205
rect 41895 68295 42105 68505
rect 39195 67995 39405 68205
rect 9795 67695 10005 67905
rect 12195 67695 12405 67905
rect 19995 67695 20205 67905
rect 21195 67695 21405 67905
rect 21795 67695 22005 67905
rect 41295 67695 41505 67905
rect 52695 68295 52905 68505
rect 70095 68295 70305 68505
rect 49995 67995 50205 68205
rect 52395 67995 52605 68205
rect 43395 67695 43605 67905
rect 70995 67995 71205 68205
rect 70095 67695 70305 67905
rect 73695 67695 73905 67905
rect 75195 67695 75405 67905
rect 76095 68295 76305 68505
rect 82095 68295 82305 68505
rect 76095 67695 76305 67905
rect 84495 68295 84705 68505
rect 25395 67395 25605 67605
rect 26595 67395 26805 67605
rect 29895 67395 30105 67605
rect 30795 67395 31005 67605
rect 52395 67395 52605 67605
rect 88395 67695 88605 67905
rect 89595 67695 89805 67905
rect 83295 67395 83505 67605
rect 18495 65895 18705 66105
rect 19095 65895 19305 66105
rect 68895 65595 69105 65805
rect 6495 64995 6705 65205
rect 36795 64995 37005 65205
rect 40095 64995 40305 65205
rect 23595 64695 23805 64905
rect 14295 64395 14505 64605
rect 21495 64380 21705 64590
rect 37395 64695 37605 64905
rect 66495 64995 66705 65205
rect 68295 64980 68505 65190
rect 70095 65295 70305 65505
rect 71595 65295 71805 65505
rect 78195 65295 78405 65505
rect 79395 65295 79605 65505
rect 70695 64995 70905 65205
rect 75195 64995 75405 65205
rect 76695 64995 76905 65205
rect 7395 64095 7605 64305
rect 20295 64095 20505 64305
rect 71595 64395 71805 64605
rect 74295 64395 74505 64605
rect 80295 64995 80505 65205
rect 82695 64995 82905 65205
rect 83295 64995 83505 65205
rect 85695 64995 85905 65205
rect 87195 64995 87405 65205
rect 77595 64395 77805 64605
rect 80295 64395 80505 64605
rect 30195 64095 30405 64305
rect 31695 64095 31905 64305
rect 37695 64095 37905 64305
rect 67695 64095 67905 64305
rect 68895 64095 69105 64305
rect 69795 64095 70005 64305
rect 71295 64095 71505 64305
rect 85995 64095 86205 64305
rect 86895 64095 87105 64305
rect 38595 62895 38805 63105
rect 39795 61395 40005 61605
rect 40095 61395 40305 61605
rect 2895 60795 3105 61005
rect 4095 60795 4305 61005
rect 26595 60795 26805 61005
rect 27795 60795 28005 61005
rect 29295 60795 29505 61005
rect 30195 60795 30405 61005
rect 35295 60795 35505 61005
rect 35895 60795 36105 61005
rect 61095 60795 61305 61005
rect 62295 60795 62505 61005
rect 64695 60795 64905 61005
rect 66195 60780 66405 60990
rect 77895 60795 78105 61005
rect 79395 60795 79605 61005
rect 85395 60795 85605 61005
rect 86295 60780 86505 60990
rect 88695 60810 88905 61020
rect 89895 60795 90105 61005
rect 13395 60495 13605 60705
rect 23895 60495 24105 60705
rect 24795 60495 25005 60705
rect 16395 60195 16605 60405
rect 6795 59895 7005 60105
rect 7695 59895 7905 60105
rect 23895 59895 24105 60105
rect 28095 60495 28305 60705
rect 29895 60495 30105 60705
rect 25995 59895 26205 60105
rect 27495 59895 27705 60105
rect 31995 60495 32205 60705
rect 41595 60495 41805 60705
rect 31095 59895 31305 60105
rect 41595 59895 41805 60105
rect 44295 60495 44505 60705
rect 63495 60495 63705 60705
rect 69195 60495 69405 60705
rect 44295 59895 44505 60105
rect 29295 59595 29505 59805
rect 34995 59595 35205 59805
rect 35595 59595 35805 59805
rect 63795 59595 64005 59805
rect 67395 59595 67605 59805
rect 68295 59595 68505 59805
rect 76695 60495 76905 60705
rect 80895 60495 81105 60705
rect 91095 60810 91305 61020
rect 83295 60195 83505 60405
rect 73695 59895 73905 60105
rect 76695 59895 76905 60105
rect 79995 59895 80205 60105
rect 90195 59895 90405 60105
rect 69495 59280 69705 59490
rect 39195 58095 39405 58305
rect 39795 58080 40005 58290
rect 39495 57780 39705 57990
rect 40695 57795 40905 58005
rect 85095 57795 85305 58005
rect 85695 57795 85905 58005
rect 22395 57495 22605 57705
rect 11595 57195 11805 57405
rect 12795 57195 13005 57405
rect 13395 57195 13605 57405
rect 18495 57195 18705 57405
rect 20295 57195 20505 57405
rect 24195 57495 24405 57705
rect 28995 57495 29205 57705
rect 74295 57495 74505 57705
rect 74895 57495 75105 57705
rect 75495 57495 75705 57705
rect 86895 57495 87105 57705
rect 88095 57495 88305 57705
rect 11595 56595 11805 56805
rect 18495 56595 18705 56805
rect 20595 56595 20805 56805
rect 23295 56595 23505 56805
rect 24495 56595 24705 56805
rect 28395 56595 28605 56805
rect 29295 57195 29505 57405
rect 31995 57195 32205 57405
rect 42195 57195 42405 57405
rect 59595 57195 59805 57405
rect 85095 57195 85305 57405
rect 29295 56595 29505 56805
rect 30795 56595 31005 56805
rect 13695 56295 13905 56505
rect 14595 56295 14805 56505
rect 25695 56265 25905 56475
rect 26295 56295 26505 56505
rect 31095 56295 31305 56505
rect 31995 56295 32205 56505
rect 87195 57195 87405 57405
rect 88995 57195 89205 57405
rect 59895 56580 60105 56790
rect 85995 56595 86205 56805
rect 87795 56595 88005 56805
rect 88995 56595 89205 56805
rect 41895 56280 42105 56490
rect 45795 56295 46005 56505
rect 46995 56295 47205 56505
rect 84195 56295 84405 56505
rect 86295 56295 86505 56505
rect 86895 56265 87105 56475
rect 88095 56295 88305 56505
rect 40095 54195 40305 54405
rect 40695 54195 40905 54405
rect 27795 53595 28005 53805
rect 28995 53595 29205 53805
rect 23295 53295 23505 53505
rect 24795 53295 25005 53505
rect 795 52995 1005 53205
rect 1995 52995 2205 53205
rect 7395 52995 7605 53205
rect 8895 52995 9105 53205
rect 24495 52695 24705 52905
rect 29295 52995 29505 53205
rect 41895 52995 42105 53205
rect 42795 52995 43005 53205
rect 82095 52995 82305 53205
rect 82995 52995 83205 53205
rect 28395 52380 28605 52590
rect 30795 52695 31005 52905
rect 56595 52695 56805 52905
rect 57195 52695 57405 52905
rect 67095 52695 67305 52905
rect 79995 52695 80205 52905
rect 24495 52095 24705 52305
rect 30795 52095 31005 52305
rect 66495 52095 66705 52305
rect 85695 52995 85905 53205
rect 90195 52695 90405 52905
rect 79995 52095 80205 52305
rect 84495 52095 84705 52305
rect 89295 52095 89505 52305
rect 33795 51795 34005 52005
rect 35295 51795 35505 52005
rect 37395 50295 37605 50505
rect 38295 50295 38505 50505
rect 45495 50295 45705 50505
rect 35595 49695 35805 49905
rect 45495 49695 45705 49905
rect 77295 49695 77505 49905
rect 8895 49395 9105 49605
rect 8895 48795 9105 49005
rect 9795 49395 10005 49605
rect 11295 49395 11505 49605
rect 11295 48795 11505 49005
rect 23295 49395 23505 49605
rect 24195 49395 24405 49605
rect 28995 49395 29205 49605
rect 23295 48795 23505 49005
rect 6795 48495 7005 48705
rect 7695 48495 7905 48705
rect 9495 48495 9705 48705
rect 17895 48495 18105 48705
rect 19095 48495 19305 48705
rect 28995 48795 29205 49005
rect 35895 49395 36105 49605
rect 39495 49395 39705 49605
rect 43095 49395 43305 49605
rect 50595 49395 50805 49605
rect 60795 49395 61005 49605
rect 35895 48795 36105 49005
rect 39495 48795 39705 49005
rect 73095 49395 73305 49605
rect 43995 48795 44205 49005
rect 50595 48795 50805 49005
rect 60795 48795 61005 49005
rect 66195 48795 66405 49005
rect 72195 48795 72405 49005
rect 76395 48795 76605 49005
rect 82995 49395 83205 49605
rect 89295 49380 89505 49590
rect 82995 48795 83205 49005
rect 25395 48495 25605 48705
rect 34995 48495 35205 48705
rect 36195 48495 36405 48705
rect 37395 48495 37605 48705
rect 38295 48465 38505 48675
rect 58095 48495 58305 48705
rect 59895 48495 60105 48705
rect 66195 48480 66405 48690
rect 66795 48495 67005 48705
rect 73995 48495 74205 48705
rect 75195 48495 75405 48705
rect 65895 48180 66105 48390
rect 90495 48180 90705 48390
rect 84495 47880 84705 48090
rect 85095 47895 85305 48105
rect 31395 46395 31605 46605
rect 32295 46395 32505 46605
rect 4095 45195 4305 45405
rect 5895 45195 6105 45405
rect 24795 45195 25005 45405
rect 25695 45195 25905 45405
rect 28995 45195 29205 45405
rect 30495 45195 30705 45405
rect 40695 45195 40905 45405
rect 41295 45195 41505 45405
rect 42195 45210 42405 45420
rect 43395 45180 43605 45390
rect 16095 44895 16305 45105
rect 21195 44895 21405 45105
rect 27195 44880 27405 45090
rect 27795 44895 28005 45105
rect 29295 44895 29505 45105
rect 11895 44295 12105 44505
rect 12795 44295 13005 44505
rect 16095 44295 16305 44505
rect 19995 44295 20205 44505
rect 32595 44895 32805 45105
rect 38595 44895 38805 45105
rect 45795 44895 46005 45105
rect 47595 44895 47805 45105
rect 49095 44895 49305 45105
rect 32595 44295 32805 44505
rect 29595 43995 29805 44205
rect 33495 43995 33705 44205
rect 34995 43995 35205 44205
rect 38895 43995 39105 44205
rect 47595 44295 47805 44505
rect 49095 44295 49305 44505
rect 60195 44895 60405 45105
rect 61395 44895 61605 45105
rect 64095 44895 64305 45105
rect 79995 44895 80205 45105
rect 84795 44895 85005 45105
rect 60195 44295 60405 44505
rect 62595 44295 62805 44505
rect 64695 44295 64905 44505
rect 73995 44295 74205 44505
rect 74595 44295 74805 44505
rect 79995 44295 80205 44505
rect 83895 44295 84105 44505
rect 45495 43980 45705 44190
rect 77295 43995 77505 44205
rect 78195 43995 78405 44205
rect 87195 43695 87405 43905
rect 88095 43695 88305 43905
rect 82995 42495 83205 42705
rect 85095 42495 85305 42705
rect 24495 42195 24705 42405
rect 25695 42195 25905 42405
rect 83295 42195 83505 42405
rect 84795 42195 85005 42405
rect 22095 41895 22305 42105
rect 22695 41895 22905 42105
rect 14595 41595 14805 41805
rect 14595 40995 14805 41205
rect 6195 40695 6405 40905
rect 7995 40695 8205 40905
rect 13095 40695 13305 40905
rect 14295 40695 14505 40905
rect 23895 41880 24105 42090
rect 28695 41895 28905 42105
rect 29895 41895 30105 42105
rect 36795 41895 37005 42105
rect 37995 41895 38205 42105
rect 80295 41895 80505 42105
rect 81495 41880 81705 42090
rect 82695 41895 82905 42105
rect 25695 41595 25905 41805
rect 31695 41595 31905 41805
rect 33795 41595 34005 41805
rect 31395 41280 31605 41490
rect 24495 40995 24705 41205
rect 37695 41595 37905 41805
rect 41895 41595 42105 41805
rect 45495 41595 45705 41805
rect 38895 41295 39105 41505
rect 49395 41595 49605 41805
rect 76695 41595 76905 41805
rect 78195 41595 78405 41805
rect 79995 41595 80205 41805
rect 46395 41295 46605 41505
rect 48795 41295 49005 41505
rect 33795 40995 34005 41205
rect 36795 40995 37005 41205
rect 38595 40995 38805 41205
rect 41295 40995 41505 41205
rect 45495 40995 45705 41205
rect 76095 41280 76305 41490
rect 81195 41595 81405 41805
rect 80595 41295 80805 41505
rect 86295 41895 86505 42105
rect 87195 41895 87405 42105
rect 88395 41910 88605 42120
rect 49395 40995 49605 41205
rect 76395 40995 76605 41205
rect 78795 40995 79005 41205
rect 79995 40995 80205 41205
rect 82995 40995 83205 41205
rect 85095 41595 85305 41805
rect 86895 41595 87105 41805
rect 85095 40995 85305 41205
rect 86895 40995 87105 41205
rect 88695 40995 88905 41205
rect 22995 40680 23205 40890
rect 32595 40695 32805 40905
rect 33195 40695 33405 40905
rect 37095 40695 37305 40905
rect 37995 40695 38205 40905
rect 39195 40695 39405 40905
rect 39795 40695 40005 40905
rect 76695 40695 76905 40905
rect 79695 40665 79905 40875
rect 80595 40695 80805 40905
rect 13995 40095 14205 40305
rect 14595 40095 14805 40305
rect 29295 37995 29505 38205
rect 30495 37995 30705 38205
rect 16395 37695 16605 37905
rect 17595 37695 17805 37905
rect 20295 37395 20505 37605
rect 21495 37395 21705 37605
rect 29505 37395 29715 37605
rect 30795 37395 31005 37605
rect 40395 37395 40605 37605
rect 42795 37395 43005 37605
rect 54795 37395 55005 37605
rect 55995 37410 56205 37620
rect 65595 37395 65805 37605
rect 2295 37095 2505 37305
rect 15495 37095 15705 37305
rect 18195 37095 18405 37305
rect 18795 37095 19005 37305
rect 36195 37095 36405 37305
rect 2895 36495 3105 36705
rect 14595 36195 14805 36405
rect 18495 36780 18705 36990
rect 41595 37095 41805 37305
rect 43695 37095 43905 37305
rect 46395 37095 46605 37305
rect 50295 37095 50505 37305
rect 19095 36495 19305 36705
rect 37095 36495 37305 36705
rect 40695 36495 40905 36705
rect 43695 36495 43905 36705
rect 70095 37095 70305 37305
rect 72195 37095 72405 37305
rect 76395 37095 76605 37305
rect 85095 37095 85305 37305
rect 46995 36495 47205 36705
rect 50895 36495 51105 36705
rect 65895 36495 66105 36705
rect 70995 36495 71205 36705
rect 72195 36495 72405 36705
rect 88095 37095 88305 37305
rect 90195 37395 90405 37605
rect 76995 36495 77205 36705
rect 85695 36495 85905 36705
rect 87195 36495 87405 36705
rect 89295 36495 89505 36705
rect 40695 36180 40905 36390
rect 42195 36195 42405 36405
rect 76095 34695 76305 34905
rect 76695 34695 76905 34905
rect 25095 34395 25305 34605
rect 25995 34395 26205 34605
rect 32595 34095 32805 34305
rect 35895 34095 36105 34305
rect 36795 34095 37005 34305
rect 1095 33795 1305 34005
rect 7395 33795 7605 34005
rect 3195 33495 3405 33705
rect 2595 33195 2805 33405
rect 16995 33795 17205 34005
rect 25395 33795 25605 34005
rect 28095 33795 28305 34005
rect 30795 33795 31005 34005
rect 7995 33195 8205 33405
rect 12495 33195 12705 33405
rect 13095 33195 13305 33405
rect 1395 32865 1605 33075
rect 15495 32895 15705 33105
rect 23295 33195 23505 33405
rect 24195 33195 24405 33405
rect 25995 33195 26205 33405
rect 35595 33795 35805 34005
rect 40395 33795 40605 34005
rect 48195 33795 48405 34005
rect 58095 33795 58305 34005
rect 60195 33795 60405 34005
rect 27195 32895 27405 33105
rect 30795 33195 31005 33405
rect 32895 33195 33105 33405
rect 36495 33180 36705 33390
rect 40695 33180 40905 33390
rect 48195 33195 48405 33405
rect 28395 32895 28605 33105
rect 60195 33195 60405 33405
rect 61095 33795 61305 34005
rect 72795 33795 73005 34005
rect 73395 33795 73605 34005
rect 75795 33795 76005 34005
rect 61095 33195 61305 33405
rect 76995 33195 77205 33405
rect 58995 32895 59205 33105
rect 79995 32595 80205 32805
rect 81195 32595 81405 32805
rect 29595 32295 29805 32505
rect 31095 32295 31305 32505
rect 23595 30195 23805 30405
rect 24795 30195 25005 30405
rect 32295 30195 32505 30405
rect 33195 30195 33405 30405
rect 67095 30195 67305 30405
rect 67995 30195 68205 30405
rect 37095 29895 37305 30105
rect 37695 29895 37905 30105
rect 51195 29895 51405 30105
rect 51795 29895 52005 30105
rect 85395 29895 85605 30105
rect 86595 29880 86805 30090
rect 9495 29595 9705 29805
rect 10095 29595 10305 29805
rect 13095 29595 13305 29805
rect 15495 29595 15705 29805
rect 16095 29595 16305 29805
rect 27495 29595 27705 29805
rect 28995 29595 29205 29805
rect 34095 29595 34305 29805
rect 34995 29595 35205 29805
rect 36495 29595 36705 29805
rect 37695 29580 37905 29790
rect 62595 29595 62805 29805
rect 63495 29595 63705 29805
rect 68595 29595 68805 29805
rect 26295 29295 26505 29505
rect 29895 29295 30105 29505
rect 40995 29295 41205 29505
rect 13395 28695 13605 28905
rect 25695 28695 25905 28905
rect 29895 28695 30105 28905
rect 41895 29295 42105 29505
rect 64695 29295 64905 29505
rect 41895 28695 42105 28905
rect 79695 29595 79905 29805
rect 83295 29595 83505 29805
rect 84495 29595 84705 29805
rect 85395 29580 85605 29790
rect 86295 29595 86505 29805
rect 64995 28680 65205 28890
rect 68895 28695 69105 28905
rect 41595 28395 41805 28605
rect 45495 28395 45705 28605
rect 67395 28395 67605 28605
rect 67995 28395 68205 28605
rect 80595 29295 80805 29505
rect 80595 28695 80805 28905
rect 84195 29295 84405 29505
rect 87795 29295 88005 29505
rect 88695 28695 88905 28905
rect 79695 28395 79905 28605
rect 84195 28395 84405 28605
rect 85695 28395 85905 28605
rect 86595 28395 86805 28605
rect 44595 28095 44805 28305
rect 24195 26595 24405 26805
rect 80295 26595 80505 26805
rect 80895 26595 81105 26805
rect 2595 25995 2805 26205
rect 4995 25995 5205 26205
rect 5595 25995 5805 26205
rect 52395 26295 52605 26505
rect 53595 26295 53805 26505
rect 54795 26295 55005 26505
rect 26295 25995 26505 26205
rect 3195 25395 3405 25605
rect 24495 25395 24705 25605
rect 25995 25395 26205 25605
rect 29595 25995 29805 26205
rect 31695 25995 31905 26205
rect 33795 25995 34005 26205
rect 78495 26280 78705 26490
rect 79095 26295 79305 26505
rect 28095 25095 28305 25305
rect 31095 25395 31305 25605
rect 56895 25995 57105 26205
rect 62295 25995 62505 26205
rect 67995 25995 68205 26205
rect 78195 25995 78405 26205
rect 33795 25395 34005 25605
rect 52395 25395 52605 25605
rect 56895 25395 57105 25605
rect 62295 25395 62505 25605
rect 30795 25095 31005 25305
rect 31995 25095 32205 25305
rect 40995 25065 41205 25275
rect 41595 25095 41805 25305
rect 66495 25095 66705 25305
rect 67095 25095 67305 25305
rect 82395 25995 82605 26205
rect 78795 25395 79005 25605
rect 81495 25395 81705 25605
rect 68895 25065 69105 25275
rect 25095 24795 25305 25005
rect 26595 24795 26805 25005
rect 85065 23895 85275 24105
rect 51495 22995 51705 23205
rect 52395 22995 52605 23205
rect 88695 22755 88905 22965
rect 28095 22095 28305 22305
rect 29595 22095 29805 22305
rect 16995 21795 17205 22005
rect 18495 21795 18705 22005
rect 24195 21795 24405 22005
rect 24795 21795 25005 22005
rect 25995 21795 26205 22005
rect 27195 21795 27405 22005
rect 63795 21795 64005 22005
rect 65595 21795 65805 22005
rect 70995 21795 71205 22005
rect 71895 21795 72105 22005
rect 90495 21795 90705 22005
rect 91095 21795 91305 22005
rect 29595 21495 29805 21705
rect 32895 21495 33105 21705
rect 8595 20895 8805 21105
rect 9195 20895 9405 21105
rect 29595 20895 29805 21105
rect 32895 20895 33105 21105
rect 43695 21495 43905 21705
rect 49095 21495 49305 21705
rect 51195 21495 51405 21705
rect 43695 20895 43905 21105
rect 69795 21495 70005 21705
rect 77895 21495 78105 21705
rect 51195 20895 51405 21105
rect 68895 20895 69105 21105
rect 79695 21495 79905 21705
rect 78795 20895 79005 21105
rect 80295 20895 80505 21105
rect 90795 20895 91005 21105
rect 91695 20895 91905 21105
rect 22095 20595 22305 20805
rect 22995 20595 23205 20805
rect 49095 20595 49305 20805
rect 51495 20580 51705 20790
rect 52395 20595 52605 20805
rect 88995 20295 89205 20505
rect 89895 20295 90105 20505
rect 66495 18495 66705 18705
rect 67095 18495 67305 18705
rect 82695 18495 82905 18705
rect 34095 18195 34305 18405
rect 495 17895 705 18105
rect 1095 17595 1305 17805
rect 45495 18195 45705 18405
rect 54195 18195 54405 18405
rect 55695 18195 55905 18405
rect 35295 17595 35505 17805
rect 45495 17595 45705 17805
rect 54795 17595 55005 17805
rect 8595 17295 8805 17505
rect 9195 17265 9405 17475
rect 17895 17295 18105 17505
rect 18495 17295 18705 17505
rect 56595 18195 56805 18405
rect 56595 17595 56805 17805
rect 81795 17595 82005 17805
rect 91095 17895 91305 18105
rect 56895 17295 57105 17505
rect 58395 17295 58605 17505
rect 59295 17295 59505 17505
rect 78195 17295 78405 17505
rect 79395 17295 79605 17505
rect 91095 16995 91305 17205
rect 90135 16395 90345 16605
rect 47295 15180 47505 15390
rect 47895 15195 48105 15405
rect 32595 14595 32805 14805
rect 31695 14295 31905 14505
rect 75795 14295 76005 14505
rect 76395 14295 76605 14505
rect 1695 13995 1905 14205
rect 3795 13995 4005 14205
rect 15195 13995 15405 14205
rect 16095 13995 16305 14205
rect 17895 13995 18105 14205
rect 19695 13995 19905 14205
rect 22395 13995 22605 14205
rect 23295 13995 23505 14205
rect 37995 13995 38205 14205
rect 39495 13995 39705 14205
rect 62505 13995 62715 14205
rect 63195 13995 63405 14205
rect 64395 14010 64605 14220
rect 65895 13995 66105 14205
rect 84795 13995 85005 14205
rect 85395 14010 85605 14220
rect 23595 13680 23805 13890
rect 24195 13695 24405 13905
rect 29595 13695 29805 13905
rect 30195 13695 30405 13905
rect 60495 13695 60705 13905
rect 76395 13695 76605 13905
rect 78495 13695 78705 13905
rect 81795 13695 82005 13905
rect 76395 13095 76605 13305
rect 77895 13095 78105 13305
rect 81795 13095 82005 13305
rect 49095 12795 49305 13005
rect 49995 12795 50205 13005
rect 61095 12795 61305 13005
rect 27795 10695 28005 10905
rect 28395 10695 28605 10905
rect 44595 10695 44805 10905
rect 45795 10695 46005 10905
rect 58695 10695 58905 10905
rect 59595 10695 59805 10905
rect 63795 10695 64005 10905
rect 64995 10695 65205 10905
rect 73695 10695 73905 10905
rect 19095 10395 19305 10605
rect 25695 10395 25905 10605
rect 19695 9795 19905 10005
rect 31095 10395 31305 10605
rect 33495 10395 33705 10605
rect 44295 10395 44505 10605
rect 45195 10395 45405 10605
rect 47595 10395 47805 10605
rect 47295 10095 47505 10305
rect 56595 10095 56805 10305
rect 30195 9795 30405 10005
rect 32595 9795 32805 10005
rect 46995 9795 47205 10005
rect 47595 9795 47805 10005
rect 55695 9795 55905 10005
rect 56295 9795 56505 10005
rect 87495 10395 87705 10605
rect 72795 9795 73005 10005
rect 86895 9795 87105 10005
rect 22995 9495 23205 9705
rect 25095 9495 25305 9705
rect 26595 9495 26805 9705
rect 56595 9495 56805 9705
rect 57495 9495 57705 9705
rect 59295 9495 59505 9705
rect 6795 6195 7005 6405
rect 7395 6195 7605 6405
rect 31695 6195 31905 6405
rect 34095 6195 34305 6405
rect 40695 6195 40905 6405
rect 41895 6195 42105 6405
rect 43095 6195 43305 6405
rect 87795 6195 88005 6405
rect 88695 6195 88905 6405
rect 23895 5895 24105 6105
rect 33195 5895 33405 6105
rect 48195 5895 48405 6105
rect 48195 5295 48405 5505
rect 49095 5895 49305 6105
rect 13095 4995 13305 5205
rect 13995 4995 14205 5205
rect 25395 4995 25605 5205
rect 26895 4995 27105 5205
rect 32595 4995 32805 5205
rect 48495 4980 48705 5190
rect 54195 4995 54405 5205
rect 55095 4965 55305 5175
rect 30195 4695 30405 4905
rect 30795 4695 31005 4905
rect 25095 4395 25305 4605
rect 26295 4395 26505 4605
rect 24195 3495 24405 3705
rect 25095 3495 25305 3705
rect 42495 2895 42705 3105
rect 43695 2895 43905 3105
rect 22095 2595 22305 2805
rect 22995 2595 23205 2805
rect 38295 2595 38505 2805
rect 44295 2595 44505 2805
rect 61995 2595 62205 2805
rect 31395 1995 31605 2205
rect 31995 1995 32205 2205
rect 37695 1995 37905 2205
rect 60195 2295 60405 2505
rect 44895 1995 45105 2205
rect 57495 1995 57705 2205
rect 66795 2595 67005 2805
rect 8595 1695 8805 1905
rect 10095 1695 10305 1905
rect 14895 1695 15105 1905
rect 16395 1695 16605 1905
rect 17280 1695 17490 1905
rect 17595 1695 17805 1905
rect 18795 1695 19005 1905
rect 31095 1695 31305 1905
rect 32895 1695 33105 1905
rect 66195 1995 66405 2205
rect 63195 1695 63405 1905
rect 89595 1695 89805 1905
rect 91095 1695 91305 1905
rect 18495 1380 18705 1590
rect 41895 495 42105 705
rect 42495 495 42705 705
<< metal2 >>
rect 50040 94005 50160 94560
rect 72840 94005 72960 94560
rect 1440 91740 1560 92295
rect 3840 91740 3960 92295
rect 4440 91905 4560 93195
rect 2640 91260 2760 91710
rect 5940 91740 6060 92295
rect 7740 91920 7860 92595
rect 4740 91305 4860 91710
rect 8940 91305 9060 91995
rect 9840 91740 9960 93195
rect 11040 91860 11160 92595
rect 11340 92205 11460 92895
rect 11040 91740 11460 91860
rect 11895 91800 12105 91995
rect 11940 91740 12060 91800
rect 1740 88905 1860 91260
rect 2640 91140 3060 91260
rect 1695 88500 1905 88695
rect 1740 88440 1860 88500
rect 2940 88605 3060 91140
rect 4140 88620 4260 91080
rect 5640 89505 5760 91260
rect 5895 88620 6105 88710
rect 1440 87405 1560 87960
rect 1440 84405 1560 87195
rect 240 78705 360 80610
rect 540 75690 660 82695
rect 1440 82305 1560 83460
rect 2040 82905 2160 87960
rect 2640 86805 2760 87960
rect 2940 87405 3060 87795
rect 2340 82260 2460 85695
rect 3240 85005 3360 88395
rect 3840 86805 3960 87960
rect 4440 85605 4560 87780
rect 5040 87705 5160 88410
rect 5640 87405 5760 87960
rect 2805 84060 3000 84105
rect 2805 83940 3060 84060
rect 2805 83895 3000 83940
rect 2205 82140 2460 82260
rect 840 76320 960 81495
rect 2040 80820 2160 82095
rect 1440 79305 1560 80160
rect 2340 80100 2460 80160
rect 2295 79905 2505 80100
rect 2940 79905 3060 81795
rect 3240 80190 3360 80895
rect 3840 80640 3960 81495
rect 4140 81105 4260 84795
rect 5595 84000 5805 84195
rect 5940 84105 6060 87495
rect 7140 87405 7260 91080
rect 8040 90705 8160 91260
rect 11640 90705 11760 91080
rect 12840 91005 12960 91995
rect 13140 91605 13260 92295
rect 13740 91740 13860 93195
rect 53040 93105 53160 93495
rect 16440 91740 16560 92295
rect 8295 88500 8505 88695
rect 8340 88440 8460 88500
rect 8940 88440 9060 89895
rect 9540 89805 9660 90495
rect 11940 89805 12060 90195
rect 12840 90105 12960 90795
rect 14640 90405 14760 91260
rect 15240 89805 15360 91710
rect 9540 89640 9795 89805
rect 9600 89595 9795 89640
rect 6495 84120 6705 84195
rect 5640 83940 5760 84000
rect 4440 83505 4560 83910
rect 7140 83940 7260 85695
rect 7440 84360 7560 88395
rect 9240 87405 9360 87780
rect 7440 84300 7860 84360
rect 7440 84240 7905 84300
rect 7695 84105 7905 84240
rect 4440 82005 4560 83295
rect 7500 83460 7695 83505
rect 5940 82305 6060 83295
rect 6840 82305 6960 83460
rect 7440 83340 7695 83460
rect 7500 83295 7695 83340
rect 8040 83205 8160 83910
rect 8340 83505 8460 87195
rect 4440 80640 4560 81195
rect 4740 79305 4860 80160
rect 1440 76140 1560 76995
rect 1740 75600 1860 75660
rect 1695 75405 1905 75600
rect 2940 73260 3060 78195
rect 5040 77205 5160 79095
rect 5340 78405 5460 82095
rect 6240 80640 6360 81195
rect 7140 80160 7260 82995
rect 8340 81405 8460 82980
rect 8340 80640 8460 81195
rect 8640 81105 8760 84495
rect 9240 84360 9360 85695
rect 9540 84705 9660 89295
rect 16140 89205 16260 91260
rect 17940 89805 18060 92295
rect 20640 91740 20760 92295
rect 21540 91290 21660 92895
rect 24840 91740 24960 92295
rect 25440 91740 25995 91860
rect 26640 91740 26760 92295
rect 18840 91200 18960 91260
rect 18795 91005 19005 91200
rect 10740 87900 10860 87960
rect 10695 87705 10905 87900
rect 11640 87105 11760 87960
rect 9240 84240 9660 84360
rect 9540 83940 9660 84240
rect 10740 83505 10860 86895
rect 12240 85605 12360 88395
rect 11895 84360 12105 84495
rect 11640 84300 12105 84360
rect 11640 84240 12060 84300
rect 11640 83940 11760 84240
rect 12840 83805 12960 84795
rect 9840 82305 9960 83460
rect 13140 82905 13260 87960
rect 13740 87900 13860 87960
rect 13695 87705 13905 87900
rect 14040 82905 14160 83460
rect 14940 81705 15060 88995
rect 17340 88440 18060 88560
rect 18495 88500 18705 88695
rect 18540 88440 18660 88500
rect 15540 87900 15660 87960
rect 15495 87705 15705 87900
rect 16440 85305 16560 87960
rect 15540 83940 15660 84495
rect 16440 83940 16560 85095
rect 17040 84405 17160 88410
rect 17340 85305 17460 88440
rect 20040 88440 20160 90795
rect 20340 90105 20460 91260
rect 20940 90405 21060 91260
rect 20940 89205 21060 90195
rect 20340 87405 20460 87960
rect 17040 83505 17160 84195
rect 17340 84120 17460 85095
rect 18840 85005 18960 87195
rect 18495 84000 18705 84195
rect 18840 84105 18960 84795
rect 18540 83940 18660 84000
rect 9240 80190 9360 80895
rect 10095 80700 10305 80895
rect 10140 80640 10260 80700
rect 11340 80190 11460 81195
rect 12540 80640 12660 81195
rect 5940 79605 6060 80160
rect 4140 74805 4260 75660
rect 2805 73140 3060 73260
rect 1440 71205 1560 72360
rect 2040 72300 2160 72360
rect 1995 72105 2205 72300
rect 240 64860 360 69795
rect 1140 68520 1260 68895
rect 2340 68520 2460 72195
rect 2640 72105 2760 73095
rect 3495 72900 3705 73095
rect 3540 72840 3660 72900
rect 4740 72390 4860 72795
rect 2640 68505 2760 71895
rect 3240 71205 3360 72360
rect 3840 71805 3960 72360
rect 5040 72060 5160 76995
rect 5340 75405 5460 76395
rect 6240 76140 6360 79695
rect 6540 79005 6660 80160
rect 7140 80040 7560 80160
rect 6840 76140 6960 76995
rect 5940 73605 6060 75660
rect 6540 74805 6660 75660
rect 7440 75105 7560 80040
rect 8040 79305 8160 80160
rect 10440 79605 10560 80160
rect 7740 76320 7860 77895
rect 8340 77205 8460 78495
rect 10440 78105 10560 79395
rect 11640 77505 11760 80595
rect 12240 80100 12360 80160
rect 12195 79905 12405 80100
rect 12840 79605 12960 80160
rect 8340 76140 8460 76995
rect 10095 76200 10305 76395
rect 10140 76140 10260 76200
rect 7740 74505 7860 76110
rect 8640 74505 8760 75660
rect 6240 72840 6360 74295
rect 4740 71940 5160 72060
rect 540 65160 660 68310
rect 1440 67005 1560 67860
rect 540 65040 795 65160
rect 2340 65205 2460 68310
rect 2940 68340 3060 70995
rect 3540 68340 3660 68895
rect 2040 65040 2295 65160
rect 240 64740 660 64860
rect 240 54405 360 58995
rect 240 40305 360 54195
rect 540 51705 660 64740
rect 840 60105 960 65010
rect 2640 64605 2760 67095
rect 3540 65040 3660 65595
rect 3840 65505 3960 67860
rect 4440 67305 4560 68295
rect 4740 67905 4860 71940
rect 5040 70905 5160 71595
rect 4440 65505 4560 67095
rect 5040 65205 5160 70695
rect 5940 68820 6060 72180
rect 7140 70305 7260 72810
rect 7440 69405 7560 73395
rect 8295 72900 8505 73095
rect 8340 72840 8460 72900
rect 8040 71205 8160 72360
rect 6240 67005 6360 67860
rect 1740 60540 1860 61095
rect 3840 61005 3960 64560
rect 4740 61305 4860 65010
rect 5640 65040 5760 65595
rect 6300 65160 6495 65205
rect 6240 65040 6495 65160
rect 6300 64995 6495 65040
rect 5940 64500 6060 64560
rect 5895 64305 6105 64500
rect 6540 63660 6660 64395
rect 6840 64005 6960 65295
rect 7140 65160 7260 68595
rect 8340 68520 8460 71895
rect 8640 70905 8760 72360
rect 9240 68205 9360 70095
rect 8040 67005 8160 67680
rect 8640 67005 8760 67860
rect 9540 67605 9660 74895
rect 9840 72405 9960 75660
rect 10440 75600 10560 75660
rect 10395 75405 10605 75600
rect 11340 74505 11460 76110
rect 11640 75405 11760 77295
rect 13740 76560 13860 81195
rect 16140 81105 16260 83280
rect 17340 83205 17460 83910
rect 14040 78705 14160 80610
rect 15540 79605 15660 80160
rect 16140 79605 16260 80580
rect 14640 77505 14760 79395
rect 16440 78105 16560 82995
rect 16740 79905 16860 81495
rect 17640 80640 17760 81195
rect 19140 80820 19260 86595
rect 20640 84060 20760 87495
rect 20340 83940 20760 84060
rect 20040 82905 20160 83460
rect 20940 82905 21060 88410
rect 21240 88005 21360 89595
rect 22440 88440 22560 90495
rect 23040 86805 23160 91260
rect 23640 90105 23760 91710
rect 24540 89205 24660 91260
rect 25740 88440 25860 91080
rect 26040 90405 26160 91710
rect 27540 90705 27660 91260
rect 28140 89505 28260 92295
rect 29940 91740 30060 92895
rect 28740 91290 28860 91710
rect 29640 91200 29760 91260
rect 23340 87405 23460 88410
rect 26040 87840 26460 87960
rect 23340 85860 23460 87195
rect 23040 85740 23460 85860
rect 23040 83505 23160 85740
rect 24195 84000 24405 84195
rect 24240 83940 24360 84000
rect 26040 83940 26160 85995
rect 26340 85905 26460 87840
rect 26640 85305 26760 89295
rect 26940 86205 27060 87795
rect 28140 87405 28260 88410
rect 28440 85860 28560 88995
rect 28740 86805 28860 91080
rect 29595 91005 29805 91200
rect 30540 91005 30660 92595
rect 31140 91740 31260 92895
rect 33540 91740 33660 92895
rect 33840 92205 33960 92595
rect 33840 92055 34095 92205
rect 33900 92010 34095 92055
rect 33900 91995 34200 92010
rect 32640 91305 32760 91710
rect 34995 91800 35205 91995
rect 35040 91740 35160 91800
rect 35640 91740 35760 92595
rect 29340 88440 29460 90195
rect 30840 87705 30960 89895
rect 32040 89505 32160 91260
rect 31695 88860 31905 88995
rect 31695 88800 31995 88860
rect 31740 88740 31995 88800
rect 32040 88440 32160 88695
rect 32895 88560 33105 88695
rect 32895 88500 33360 88560
rect 32940 88440 33360 88500
rect 35940 88560 36060 91260
rect 35940 88440 36360 88560
rect 33540 86205 33660 87960
rect 34140 87405 34260 87960
rect 36240 85905 36360 88440
rect 28440 85740 28695 85860
rect 21840 82605 21960 83460
rect 22440 82905 22560 83460
rect 24840 83490 24960 83895
rect 24495 82605 24705 82695
rect 21840 82005 21960 82395
rect 25440 82305 25560 82695
rect 25695 82605 25905 82695
rect 17340 80100 17460 80160
rect 17040 78705 17160 79995
rect 17295 79905 17505 80100
rect 17340 79305 17460 79695
rect 18840 79305 18960 80160
rect 19440 79605 19560 80160
rect 13740 76440 14160 76560
rect 14040 76140 14160 76440
rect 14640 76140 14760 77295
rect 16440 76320 16560 77295
rect 15240 76140 15960 76260
rect 13140 75405 13260 76095
rect 10395 72900 10605 73095
rect 10440 72840 10560 72900
rect 10740 71805 10860 72360
rect 11040 68805 11160 70995
rect 11340 70905 11460 72360
rect 11640 70005 11760 70395
rect 7140 65040 7560 65160
rect 6540 63540 6960 63660
rect 2895 60720 3105 60795
rect 4095 60600 4305 60795
rect 4140 60540 4260 60600
rect 2040 60000 2160 60060
rect 1995 59805 2205 60000
rect 840 56790 960 57495
rect 1740 57240 1860 58695
rect 2340 57240 2460 58395
rect 2940 57405 3060 60510
rect 5940 60540 6060 61095
rect 2040 53205 2160 56760
rect 2640 56205 2760 56760
rect 840 52275 960 52995
rect 2940 52740 3060 53895
rect 3240 52860 3360 59895
rect 3840 59805 3960 60060
rect 3840 57705 3960 59595
rect 4140 57240 4260 58395
rect 4440 57405 4560 60060
rect 5040 58905 5160 60495
rect 6840 60105 6960 63540
rect 5640 58305 5760 60060
rect 6240 59205 6360 60060
rect 7140 59505 7260 64395
rect 7440 61305 7560 64095
rect 7740 64005 7860 64560
rect 8340 64500 8460 64560
rect 8295 64305 8505 64500
rect 8940 63705 9060 67395
rect 9840 66105 9960 67695
rect 9240 64305 9360 65895
rect 11040 65505 11160 67860
rect 11640 67560 11760 68295
rect 11940 67905 12060 74295
rect 12240 72405 12360 74295
rect 13140 73260 13260 75195
rect 13740 74805 13860 75660
rect 14340 74505 14460 75660
rect 13140 73140 13560 73260
rect 13440 72840 13560 73140
rect 14940 72840 15060 75195
rect 15240 74205 15360 76140
rect 17340 75705 17460 76695
rect 16140 74805 16260 75660
rect 15240 73305 15360 73995
rect 15540 72840 16260 72960
rect 12240 68505 12360 72195
rect 13740 72300 13860 72360
rect 13695 72105 13905 72300
rect 15195 72105 15405 72180
rect 13140 69705 13260 71595
rect 11340 67440 11760 67560
rect 9840 63105 9960 64560
rect 10440 62205 10560 64395
rect 10740 63705 10860 64560
rect 11340 63705 11460 67440
rect 12240 67305 12360 67695
rect 11640 64305 11760 66795
rect 12840 65805 12960 67095
rect 14640 66405 14760 69195
rect 15540 68505 15660 68895
rect 15840 68760 15960 70695
rect 16140 69105 16260 72840
rect 16740 73005 16860 75660
rect 17640 74805 17760 77895
rect 18540 76140 18660 78495
rect 20340 76905 20460 81795
rect 22095 81660 22305 81795
rect 21840 81600 22305 81660
rect 21840 81540 22260 81600
rect 21840 80640 21960 81540
rect 20940 77805 21060 80595
rect 23340 80205 23460 80595
rect 25440 80160 25560 82095
rect 26340 81405 26460 83460
rect 26940 81405 27060 84195
rect 28740 83505 28860 85695
rect 29040 84120 29160 85395
rect 29040 82605 29160 83910
rect 29340 83205 29460 84195
rect 29940 83940 30060 85095
rect 36540 85005 36660 89295
rect 36840 88605 36960 91710
rect 37140 91260 37260 92595
rect 40005 92160 40200 92205
rect 40005 91995 40260 92160
rect 37995 91800 38205 91995
rect 38040 91740 38160 91800
rect 40140 91740 40260 91995
rect 41640 91920 41760 92295
rect 42840 91740 42960 92295
rect 37140 91140 37560 91260
rect 37440 88440 37560 91140
rect 38340 89205 38460 91260
rect 41640 91260 41760 91710
rect 46440 91740 46560 92595
rect 47940 91740 48060 92895
rect 45540 91290 45660 91695
rect 41640 91140 42060 91260
rect 40740 90705 40860 91080
rect 39540 88440 39660 88995
rect 37740 87405 37860 87960
rect 38640 87705 38760 88410
rect 41340 88440 41460 90495
rect 41940 88905 42060 91140
rect 42540 89205 42660 91260
rect 41895 88500 42105 88695
rect 41940 88440 42060 88500
rect 39795 87705 40005 87780
rect 33195 84120 33405 84195
rect 28605 82395 28695 82605
rect 29640 82005 29760 82395
rect 26940 80640 27060 81195
rect 29340 80640 29460 81795
rect 30240 81705 30360 83460
rect 22140 79005 22260 79860
rect 18105 75660 18300 75705
rect 18105 75540 18360 75660
rect 18840 75600 18960 75660
rect 18105 75495 18300 75540
rect 18795 75405 19005 75600
rect 19440 75405 19560 76395
rect 19995 76200 20205 76395
rect 20040 76140 20160 76200
rect 20640 76140 20760 77295
rect 21840 76320 21960 77295
rect 20940 75600 21060 75660
rect 16440 71505 16560 72810
rect 17940 70605 18060 72795
rect 18240 70005 18360 75195
rect 19140 72840 19260 73995
rect 19740 73005 19860 73695
rect 18840 71805 18960 72360
rect 19440 70605 19560 72360
rect 20040 72105 20160 75195
rect 20340 73020 20460 75480
rect 20895 75405 21105 75600
rect 21840 74205 21960 76110
rect 22140 75405 22260 76395
rect 20340 71205 20460 72810
rect 20940 71805 21060 72360
rect 21840 72105 21960 72360
rect 20940 70905 21060 71595
rect 15840 68640 16260 68760
rect 16140 68340 16260 68640
rect 14940 66105 15060 67995
rect 13095 65700 13305 65895
rect 13140 65640 13260 65700
rect 7440 59205 7560 60510
rect 7695 59805 7905 59895
rect 6195 57300 6405 57495
rect 6240 57240 6360 57300
rect 4740 56205 4860 56760
rect 3240 52740 3495 52860
rect 1140 49620 1260 52095
rect 2340 52140 2760 52260
rect 1740 49440 1860 50895
rect 2340 49605 2460 51795
rect 540 44490 660 49395
rect 1440 44940 1560 48780
rect 2040 48405 2160 48960
rect 2640 48360 2760 52140
rect 3540 52005 3660 52695
rect 2940 48660 3060 49695
rect 3495 49500 3705 49695
rect 4140 49620 4260 53595
rect 5040 52740 5160 54195
rect 5340 53805 5460 57195
rect 7740 56790 7860 58095
rect 8940 57705 9060 60060
rect 5640 52740 5760 56295
rect 6540 54405 6660 56760
rect 8940 55905 9060 56760
rect 9240 53205 9360 56595
rect 7395 52920 7605 52995
rect 7995 52800 8205 52995
rect 8895 52800 9105 52995
rect 9540 52920 9660 57495
rect 9840 57405 9960 60060
rect 10440 60000 10860 60060
rect 10440 59940 10905 60000
rect 10695 59805 10905 59940
rect 10905 59640 11160 59760
rect 10140 58905 10260 59295
rect 10440 57240 10560 58995
rect 11040 57405 11160 59640
rect 11340 58860 11460 61095
rect 11640 60540 11760 62895
rect 11940 62805 12060 65295
rect 12840 65040 12960 65595
rect 14340 64605 14460 65895
rect 14940 65040 15060 65895
rect 15540 65040 15660 67695
rect 15840 67305 15960 67860
rect 17040 66405 17160 68595
rect 17340 67005 17460 69495
rect 18195 68400 18405 68595
rect 18240 68340 18360 68400
rect 19440 68505 19560 69795
rect 20340 68340 20460 70680
rect 20940 68340 21060 69495
rect 19740 67905 19860 68310
rect 21840 67905 21960 71895
rect 22440 70305 22560 78495
rect 23040 76605 23160 77895
rect 22995 76200 23205 76395
rect 23040 76140 23160 76200
rect 23640 76140 23760 78795
rect 24240 77505 24360 80160
rect 24840 78705 24960 80160
rect 25140 80040 25560 80160
rect 23340 75405 23460 75660
rect 23340 73605 23460 75195
rect 23640 73260 23760 74895
rect 23940 74805 24060 75480
rect 24840 73905 24960 76110
rect 25140 75105 25260 80040
rect 26640 79005 26760 80160
rect 26340 76320 26460 76695
rect 25605 76260 25800 76305
rect 25605 76140 25860 76260
rect 25605 76095 25800 76140
rect 25440 73605 25560 75495
rect 23340 73140 23760 73260
rect 23340 72840 23460 73140
rect 23940 71505 24060 72795
rect 25740 72405 25860 73995
rect 24540 71805 24660 72360
rect 23340 68520 23460 71295
rect 25140 70305 25260 72360
rect 17640 66705 17760 67680
rect 16440 64590 16560 65295
rect 13440 60705 13560 61995
rect 12240 59205 12360 60060
rect 11340 58740 11760 58860
rect 11340 56790 11460 58395
rect 11640 57405 11760 58740
rect 12540 58305 12660 59460
rect 12195 57300 12405 57495
rect 12840 57405 12960 58695
rect 12240 57240 12360 57300
rect 10140 55905 10260 56580
rect 8040 52740 8160 52800
rect 8940 52740 9060 52800
rect 10140 52905 10260 53295
rect 6540 52305 6660 52710
rect 7140 50460 7260 52260
rect 9240 51960 9360 52260
rect 9840 52200 9960 52260
rect 9795 52005 10005 52200
rect 9240 51840 9660 51960
rect 9540 51660 9660 51840
rect 10140 51660 10260 52095
rect 9540 51540 10260 51660
rect 6840 50340 7260 50460
rect 5640 49620 5760 50295
rect 3540 49440 3660 49500
rect 6240 49440 6360 49995
rect 6840 49305 6960 50340
rect 2940 48540 3360 48660
rect 2640 48240 2895 48360
rect 2640 45120 2760 46695
rect 2040 41640 2160 43395
rect 2640 42405 2760 44910
rect 840 39105 960 41595
rect 1740 41100 1860 41160
rect 1695 40905 1905 41100
rect 2940 41160 3060 48195
rect 3240 45120 3360 48540
rect 3840 48405 3960 48960
rect 4095 45120 4305 45195
rect 4740 44940 4860 47295
rect 5940 46905 6060 48780
rect 6840 48705 6960 49095
rect 7140 47805 7260 49995
rect 8040 49440 8160 50295
rect 8940 49605 9060 51495
rect 10440 51405 10560 54795
rect 11340 53160 11460 53895
rect 11640 53505 11760 56595
rect 12540 56205 12660 56760
rect 11340 53040 11760 53160
rect 11640 52740 11760 53040
rect 12540 52305 12660 52710
rect 7740 48900 7860 48960
rect 7695 48705 7905 48900
rect 9240 48990 9360 49995
rect 8940 48405 9060 48795
rect 9540 48960 9660 51195
rect 10740 50205 10860 51195
rect 11340 51105 11460 52260
rect 12840 52005 12960 56595
rect 13140 55005 13260 58995
rect 13440 57405 13560 57795
rect 13740 57405 13860 62595
rect 14040 57660 14160 64095
rect 16140 61605 16260 63495
rect 16740 62805 16860 66195
rect 18540 66105 18660 67095
rect 19140 66105 19260 67860
rect 19740 66705 19860 67695
rect 20040 66705 20160 67695
rect 21195 67560 21405 67695
rect 20940 67500 21405 67560
rect 20940 67440 21360 67500
rect 17505 65340 17895 65460
rect 17040 64440 17460 64560
rect 17040 63405 17160 64440
rect 17040 62460 17160 63195
rect 16740 62340 17160 62460
rect 16440 60405 16560 61995
rect 14040 57540 14460 57660
rect 14340 57420 14460 57540
rect 14940 57240 15060 58995
rect 16740 58605 16860 62340
rect 17340 60540 17460 63795
rect 17940 63105 18060 64560
rect 18240 62205 18360 64395
rect 18540 63705 18660 65895
rect 19995 65100 20205 65295
rect 20040 65040 20160 65100
rect 20940 64905 21060 67440
rect 22140 67305 22260 67695
rect 22440 66960 22560 67860
rect 22005 66840 22560 66960
rect 21240 64905 21360 66495
rect 23640 64905 23760 65595
rect 19140 63060 19260 64695
rect 19740 64500 19860 64560
rect 20340 64500 20460 64560
rect 19695 64305 19905 64500
rect 20295 64305 20505 64500
rect 23340 64500 23460 64575
rect 19140 62940 19395 63060
rect 17640 59760 17760 60060
rect 17340 59640 17760 59760
rect 13440 56790 13560 57195
rect 14640 56700 14760 56760
rect 14595 56505 14805 56700
rect 13440 54660 13560 55695
rect 13140 54540 13560 54660
rect 13140 51705 13260 54540
rect 13740 52920 13860 56295
rect 15540 55905 15660 58395
rect 17340 58005 17460 59640
rect 16005 56760 16200 56805
rect 16005 56640 16260 56760
rect 16005 56595 16200 56640
rect 16740 56505 16860 56760
rect 17640 56505 17760 58395
rect 14340 53505 14460 53895
rect 14340 52740 14460 53295
rect 14940 52905 15060 55095
rect 13440 51405 13560 52095
rect 14640 52200 14760 52260
rect 14595 52005 14805 52200
rect 11340 50505 11460 50895
rect 10005 49560 10200 49605
rect 10005 49440 10260 49560
rect 10005 49395 10200 49440
rect 11340 49605 11460 50295
rect 12840 49440 12960 50895
rect 13440 49605 13560 51195
rect 9540 48840 9960 48960
rect 3840 43005 3960 44460
rect 3240 41805 3360 42795
rect 4140 42060 4260 43395
rect 3840 41940 4260 42060
rect 3840 41640 3960 41940
rect 2640 41040 3060 41160
rect 240 3705 360 38595
rect 540 35805 660 37695
rect 2340 37305 2460 40095
rect 540 31605 660 33795
rect 540 18105 660 27795
rect 840 27105 960 36195
rect 1440 35805 1560 36660
rect 1740 35205 1860 36495
rect 2640 36405 2760 41040
rect 3240 37905 3360 39495
rect 4140 38505 4260 41160
rect 3240 37140 3360 37695
rect 3840 37320 3960 37995
rect 2895 36405 3105 36495
rect 1140 34005 1260 34995
rect 1740 33840 1860 34395
rect 1140 31305 1260 32895
rect 1440 30405 1560 32865
rect 2040 31905 2160 33360
rect 2940 33360 3060 34995
rect 3540 34020 3660 36660
rect 4440 35805 4560 40095
rect 3840 34605 3960 35595
rect 3900 34260 4095 34305
rect 3840 34095 4095 34260
rect 3240 33900 3495 33960
rect 3195 33840 3495 33900
rect 3195 33705 3405 33840
rect 3840 33840 3960 34095
rect 4440 33840 4560 34995
rect 4740 34305 4860 40695
rect 5040 40305 5160 42195
rect 5340 40905 5460 45195
rect 5895 45000 6105 45195
rect 5940 44940 6060 45000
rect 6540 44940 6660 47295
rect 7440 44505 7560 45795
rect 8895 45000 9105 45195
rect 9540 45105 9660 48495
rect 8940 44940 9060 45000
rect 5940 41640 6060 43095
rect 7740 43005 7860 44910
rect 8640 43605 8760 44280
rect 9240 43905 9360 44460
rect 7440 41190 7560 42195
rect 8340 41820 8460 42495
rect 6840 41040 7395 41160
rect 8040 41100 8160 41160
rect 6195 40905 6405 40980
rect 7995 40905 8205 41100
rect 7740 39105 7860 40395
rect 9540 38505 9660 43995
rect 9840 39405 9960 48840
rect 11100 48960 11295 49005
rect 11040 48840 11295 48960
rect 11100 48795 11295 48840
rect 10740 47805 10860 48495
rect 11640 47505 11760 49410
rect 12540 48900 12660 48960
rect 12495 48705 12705 48900
rect 13740 48105 13860 51495
rect 15240 51105 15360 53295
rect 16140 52740 16260 53895
rect 16740 53505 16860 56295
rect 16740 52740 16860 53295
rect 15540 52200 15960 52260
rect 15495 52140 15960 52200
rect 15495 52005 15705 52140
rect 16440 51705 16560 52260
rect 17340 51105 17460 55695
rect 14940 49440 15060 50295
rect 15540 49440 15660 50295
rect 16740 49905 16860 50295
rect 17340 49905 17460 50295
rect 17340 49440 17460 49695
rect 17640 49605 17760 53895
rect 17940 53505 18060 58995
rect 18240 56790 18360 60060
rect 18840 59505 18960 61395
rect 18540 57405 18660 58995
rect 19140 58605 19260 60510
rect 19440 60105 19560 62895
rect 20040 61005 20160 62595
rect 21540 61605 21660 64380
rect 23295 64305 23505 64500
rect 20040 60540 20160 60795
rect 20640 60540 20760 61395
rect 19140 57240 19260 57795
rect 20340 57405 20460 60060
rect 20940 57660 21060 59295
rect 21240 59205 21360 60495
rect 21540 58305 21660 60795
rect 22140 60720 22260 63495
rect 23940 63405 24060 69495
rect 24240 63405 24360 70095
rect 26040 70005 26160 74295
rect 25740 68520 25860 69195
rect 24840 66405 24960 67860
rect 25440 67800 25560 67860
rect 25395 67605 25605 67800
rect 25395 67305 25605 67395
rect 25140 65040 25260 65895
rect 23040 60540 23160 62295
rect 20940 57540 21360 57660
rect 21240 57240 21360 57540
rect 21840 57240 21960 59295
rect 22440 57705 22560 59880
rect 18540 54105 18660 56595
rect 18840 54705 18960 56580
rect 20040 53505 20160 56595
rect 20340 56205 20460 56880
rect 20640 53805 20760 56595
rect 20940 56205 21060 56760
rect 18840 52920 18960 53295
rect 19440 52740 19560 53295
rect 22440 52860 22560 57180
rect 22740 56790 22860 57795
rect 23040 56205 23160 58095
rect 23340 57405 23460 59895
rect 23640 59505 23760 62595
rect 23940 60705 24060 62880
rect 24540 61560 24660 64395
rect 24840 61905 24960 64560
rect 24540 61440 24960 61560
rect 24840 60705 24960 61440
rect 25140 60060 25260 63795
rect 25440 63705 25560 64560
rect 25740 63360 25860 64395
rect 26040 64005 26160 67395
rect 26340 67305 26460 74895
rect 26640 74805 26760 75495
rect 26940 75405 27060 79695
rect 27240 79605 27360 80160
rect 28140 79905 28260 80610
rect 29040 79605 29160 80160
rect 29640 80100 29760 80160
rect 29595 79905 29805 80100
rect 27240 76305 27360 79395
rect 29040 78705 29160 79395
rect 30240 79005 30360 80610
rect 31140 79905 31260 80160
rect 31005 79740 31260 79905
rect 31005 79695 31200 79740
rect 28740 78105 28860 78495
rect 28140 76140 28260 77895
rect 30240 76140 30360 78195
rect 27840 75600 27960 75660
rect 27795 75405 28005 75600
rect 27240 73020 27360 73395
rect 26940 71160 27060 72360
rect 28440 71760 28560 75495
rect 28740 75405 28860 76110
rect 30840 75705 30960 78795
rect 31140 78405 31260 79395
rect 31740 79005 31860 82995
rect 32040 77805 32160 82395
rect 32340 79605 32460 82695
rect 32940 82605 33060 83460
rect 33540 82905 33660 84195
rect 33840 83505 33960 84195
rect 34395 84000 34605 84195
rect 34440 83940 34560 84000
rect 34740 83400 34860 83460
rect 34140 82905 34260 83295
rect 34695 83205 34905 83400
rect 35340 82905 35460 83460
rect 35940 83205 36060 84195
rect 37395 84000 37605 84195
rect 37440 83940 37560 84000
rect 33240 80640 33360 81495
rect 33840 80640 33960 82395
rect 34740 82005 34860 82680
rect 34140 80805 34260 81195
rect 34740 80820 34860 81795
rect 35940 81660 36060 82395
rect 36540 82305 36660 83460
rect 35940 81540 36360 81660
rect 35340 80640 35460 81195
rect 36240 80205 36360 81540
rect 37140 81060 37260 83460
rect 38040 81105 38160 83910
rect 37140 80940 37560 81060
rect 37440 80820 37560 80940
rect 38340 80760 38460 84195
rect 38940 83940 39060 84495
rect 39240 82605 39360 83460
rect 38040 80640 38760 80760
rect 32940 78705 33060 80160
rect 33540 79005 33660 80160
rect 29340 72840 29460 75195
rect 29640 74805 29760 75660
rect 29040 72300 29160 72360
rect 28305 71640 28560 71760
rect 26940 71040 27360 71160
rect 26940 68340 27060 70695
rect 27240 70605 27360 71040
rect 28140 68505 28260 71595
rect 28740 69405 28860 72180
rect 28995 72105 29205 72300
rect 29805 72240 30060 72360
rect 29040 70305 29160 71895
rect 29940 71805 30060 72240
rect 28440 67905 28560 69195
rect 29940 68340 30060 70995
rect 26595 67605 26805 67695
rect 27840 67305 27960 67860
rect 27240 65040 27360 65595
rect 27840 65040 27960 66195
rect 28140 65205 28260 65895
rect 23940 59205 24060 59895
rect 24240 59760 24360 60060
rect 24840 59940 25260 60060
rect 25440 63240 25860 63360
rect 24240 59640 24660 59760
rect 23940 57240 24060 58395
rect 24240 57705 24360 59295
rect 24540 58605 24660 59640
rect 24540 57405 24660 57795
rect 22140 52740 22560 52860
rect 23040 52740 23160 55095
rect 23340 54105 23460 56595
rect 24240 55605 24360 56760
rect 23295 53505 23505 53580
rect 23640 52920 23760 53295
rect 18540 50760 18660 52260
rect 19140 51705 19260 52260
rect 20640 51360 20760 52260
rect 21240 51705 21360 52260
rect 21840 51705 21960 52095
rect 20640 51240 21060 51360
rect 18540 50640 18960 50760
rect 10695 45000 10905 45195
rect 10740 44940 10860 45000
rect 11340 44940 11460 45795
rect 11940 45105 12060 46095
rect 10140 43905 10260 44895
rect 11700 44460 11895 44505
rect 11040 42705 11160 44460
rect 11640 44340 11895 44460
rect 11700 44295 11895 44340
rect 12240 44205 12360 44910
rect 11595 41700 11805 41895
rect 11640 41640 11760 41700
rect 10140 40005 10260 41595
rect 10740 38805 10860 41160
rect 12240 39405 12360 43095
rect 12540 41805 12660 47895
rect 15240 46905 15360 48960
rect 15840 48405 15960 48960
rect 17940 48900 18060 48960
rect 17895 48705 18105 48900
rect 18540 48960 18660 50295
rect 18840 50205 18960 50640
rect 18540 48840 19260 48960
rect 17895 48405 18105 48495
rect 13740 44940 13860 45495
rect 14340 45105 14460 46695
rect 15240 44940 15360 46095
rect 15900 45060 16095 45105
rect 15840 44940 16095 45060
rect 15900 44895 16095 44940
rect 16440 44505 16560 45195
rect 18240 45060 18360 48795
rect 19305 48495 19395 48705
rect 18240 44940 18660 45060
rect 12795 44205 13005 44295
rect 13440 43305 13560 44460
rect 14640 44340 15060 44460
rect 12795 41700 13005 41895
rect 12840 41640 12960 41700
rect 13440 41640 13560 43095
rect 14640 42405 14760 44340
rect 16140 43905 16260 44295
rect 14640 41805 14760 42195
rect 13140 41100 13260 41160
rect 5940 37140 6060 37695
rect 5640 36360 5760 36660
rect 6240 36600 6360 36660
rect 5340 36240 5760 36360
rect 6195 36405 6405 36600
rect 5340 35205 5460 36240
rect 2940 33240 3360 33360
rect 2640 29505 2760 33195
rect 3240 32205 3360 33240
rect 3540 32805 3660 33180
rect 4140 31905 4260 33360
rect 2340 29340 2595 29460
rect 1440 28005 1560 28860
rect 1740 27705 1860 28395
rect 2040 28005 2160 28860
rect 2640 26205 2760 28695
rect 2940 28605 3060 31695
rect 4440 31005 4560 32895
rect 4440 29520 4560 30195
rect 540 16605 660 17580
rect 540 10905 660 15195
rect 840 15105 960 25995
rect 2940 25590 3060 28395
rect 3240 26205 3360 28695
rect 3540 27105 3660 28860
rect 4140 27705 4260 28860
rect 3840 26040 3960 26595
rect 4740 26505 4860 28695
rect 5040 28005 5160 32595
rect 5340 29505 5460 34095
rect 5640 33390 5760 34395
rect 5940 34005 6060 34995
rect 6840 34305 6960 37095
rect 7140 36660 7260 38295
rect 7140 36540 7560 36660
rect 7140 33840 7260 35595
rect 7440 34005 7560 36540
rect 8040 35805 8160 36660
rect 8640 35205 8760 36795
rect 9240 35805 9360 36660
rect 9840 36405 9960 36660
rect 9840 36240 10095 36405
rect 9900 36195 10095 36240
rect 7740 33390 7860 34095
rect 8640 33840 8760 34995
rect 5895 29400 6105 29595
rect 6540 29520 6660 32895
rect 6840 32505 6960 33360
rect 8040 30405 8160 33195
rect 8940 32805 9060 33360
rect 8940 31905 9060 32595
rect 5940 29340 6060 29400
rect 7395 29400 7605 29595
rect 7440 29340 7560 29400
rect 8940 28890 9060 30795
rect 5640 28800 5760 28860
rect 1440 23805 1560 25560
rect 3405 25560 3600 25605
rect 3405 25440 3660 25560
rect 3405 25395 3600 25440
rect 5040 23505 5160 25995
rect 1740 21540 1860 22695
rect 2340 21540 2460 23295
rect 3240 21540 3360 22695
rect 3840 21540 3960 22395
rect 1440 18705 1560 21060
rect 2040 20505 2160 21060
rect 1740 18240 1860 19695
rect 4140 19005 4260 21060
rect 4740 20505 4860 22395
rect 5040 21090 5160 23295
rect 2940 17790 3060 18795
rect 1140 14205 1260 17595
rect 4740 17760 4860 19980
rect 5340 19905 5460 28695
rect 5595 28605 5805 28800
rect 8340 28305 8460 28860
rect 5805 26160 6000 26205
rect 5805 26040 6060 26160
rect 6540 26040 6660 27495
rect 8340 26505 8460 28095
rect 5805 25995 6000 26040
rect 7440 25590 7560 26295
rect 5640 24705 5760 25395
rect 5940 21540 6060 23895
rect 6240 23805 6360 25380
rect 6540 22905 6660 25095
rect 6240 18420 6360 21060
rect 7140 20205 7260 23295
rect 8340 22005 8460 25560
rect 8940 24105 9060 25395
rect 8340 21540 8460 21795
rect 9240 21105 9360 30195
rect 9495 29505 9705 29595
rect 9840 29520 9960 33795
rect 10140 29805 10260 34095
rect 10440 34005 10560 36495
rect 10740 36405 10860 38280
rect 10740 33840 10860 35595
rect 11040 35505 11160 39195
rect 12540 38505 12660 40995
rect 13095 40905 13305 41100
rect 13740 40605 13860 41160
rect 14340 40905 14460 41595
rect 14595 40905 14805 40995
rect 13740 40305 13860 40395
rect 13740 40140 13995 40305
rect 13800 40095 13995 40140
rect 14805 40095 14895 40305
rect 11340 36105 11460 37695
rect 12240 37140 12360 37695
rect 11940 35505 12060 36660
rect 12540 34605 12660 36660
rect 11295 33900 11505 34095
rect 11340 33840 11460 33900
rect 12540 33405 12660 34080
rect 10440 32805 10560 33195
rect 11040 32805 11160 33360
rect 11640 32205 11760 33180
rect 12840 32805 12960 35895
rect 13140 34305 13260 38895
rect 13440 36105 13560 37995
rect 14040 37140 14160 37695
rect 14640 37140 14760 38295
rect 15540 37305 15660 37995
rect 15840 37320 15960 42495
rect 16140 40305 16260 43695
rect 16440 41805 16560 43980
rect 17340 43305 17460 44460
rect 18540 43560 18660 44940
rect 18240 43440 18660 43560
rect 17040 41640 17160 43095
rect 17595 41700 17805 41895
rect 17640 41640 17760 41700
rect 16740 38205 16860 40980
rect 17340 40305 17460 41160
rect 17595 37905 17805 37995
rect 14340 35205 14460 36660
rect 15240 36405 15360 37110
rect 16440 37140 16560 37695
rect 13740 33840 13860 34995
rect 11805 30360 12000 30405
rect 11805 30300 12060 30360
rect 11805 30195 12105 30300
rect 9690 29400 9705 29505
rect 10440 29340 10560 30195
rect 11895 30105 12105 30195
rect 13140 29805 13260 33195
rect 9540 26205 9660 28695
rect 10740 27705 10860 28860
rect 10740 26040 10860 26895
rect 11340 26220 11460 29295
rect 11640 28305 11760 29595
rect 13440 29505 13560 30495
rect 13740 28905 13860 29895
rect 11940 26505 12060 28695
rect 12540 28305 12660 28860
rect 12840 27405 12960 28395
rect 13140 25590 13260 26295
rect 10440 24705 10560 25560
rect 11940 25500 12060 25560
rect 11895 25305 12105 25500
rect 9540 22140 10695 22260
rect 9540 21720 9660 22140
rect 9795 21600 10005 21795
rect 10395 21600 10605 21795
rect 9840 21540 9960 21600
rect 10440 21540 10560 21600
rect 7440 18240 7560 19395
rect 8040 19305 8160 21060
rect 4140 17640 4860 17760
rect 1440 16005 1560 17580
rect 840 14040 1095 14160
rect 840 13005 960 14040
rect 1695 13800 1905 13995
rect 1740 13740 1860 13800
rect 2340 13740 2460 14895
rect 2940 13905 3060 17580
rect 3795 14205 4005 14295
rect 3195 13800 3405 13995
rect 3240 13740 3360 13800
rect 3840 13740 3960 13995
rect 540 9405 660 10695
rect 840 9990 960 11295
rect 1440 10905 1560 13260
rect 2040 13200 2160 13260
rect 1995 13005 2205 13200
rect 4740 13290 4860 14895
rect 1740 10440 1860 10995
rect 2640 10620 2760 13095
rect 4140 11805 4260 13260
rect 2340 10440 2595 10560
rect 2040 9405 2160 9960
rect 1740 5940 1860 7095
rect 2295 6000 2505 6195
rect 2940 6105 3060 10995
rect 4140 10860 4260 11595
rect 4140 10740 4560 10860
rect 3240 10440 3960 10560
rect 4440 10440 4560 10740
rect 5040 10560 5160 18195
rect 5940 17205 6060 17760
rect 6540 16305 6660 17760
rect 5940 14205 6060 15795
rect 6240 13740 6360 15195
rect 7140 13290 7260 17595
rect 7740 13740 7860 17580
rect 8340 17205 8460 18495
rect 8640 17505 8760 20895
rect 10140 20760 10260 21060
rect 9840 20640 10260 20760
rect 9540 18240 9660 18795
rect 9840 18705 9960 20640
rect 10395 20505 10605 20595
rect 10740 20505 10860 21060
rect 10305 20400 10605 20505
rect 10305 20340 10560 20400
rect 10305 20295 10500 20340
rect 10140 18240 10260 19980
rect 11340 19305 11460 25095
rect 12540 23505 12660 25560
rect 12240 21540 12360 22095
rect 13140 21090 13260 21795
rect 11940 20505 12060 21060
rect 13440 20760 13560 28695
rect 13740 22305 13860 26895
rect 14040 26205 14160 33195
rect 14340 29520 14460 34680
rect 14640 33405 14760 36195
rect 15540 34905 15660 36495
rect 15840 34020 15960 36195
rect 16140 35505 16260 36660
rect 17040 36105 17160 37695
rect 17895 37200 18105 37395
rect 18240 37305 18360 43440
rect 18540 37305 18660 43095
rect 18840 42705 18960 47895
rect 20340 47505 20460 49395
rect 20640 47160 20760 50895
rect 20340 47040 20760 47160
rect 19440 43905 19560 44460
rect 20040 43305 20160 44295
rect 20340 44160 20460 47040
rect 20640 44505 20760 45795
rect 20340 44040 20760 44160
rect 20040 41640 20160 42195
rect 19140 39405 19260 41160
rect 19740 39105 19860 41160
rect 20640 38505 20760 44040
rect 20940 43905 21060 51240
rect 22140 51105 22260 52740
rect 22740 49605 22860 52260
rect 24240 50805 24360 53895
rect 24540 52905 24660 56595
rect 24840 55005 24960 59940
rect 25440 58605 25560 63240
rect 25140 58440 25395 58560
rect 25140 57405 25260 58440
rect 25440 57240 25560 57795
rect 25740 57705 25860 61395
rect 26040 61005 26160 63480
rect 26940 61305 27060 64560
rect 28440 63705 28560 67380
rect 28740 61020 28860 67095
rect 29640 66405 29760 67860
rect 29940 65505 30060 67395
rect 30540 67260 30660 74895
rect 31140 73605 31260 77595
rect 31740 76140 31860 76695
rect 32340 76320 32460 77895
rect 32040 74805 32160 75660
rect 32940 75105 33060 77595
rect 34140 76140 34260 79095
rect 34440 78705 34560 79995
rect 33840 74805 33960 75660
rect 34440 74505 34560 75495
rect 31395 72900 31605 73095
rect 31440 72840 31560 72900
rect 31740 70905 31860 71595
rect 32040 71505 32160 73095
rect 31440 68340 31560 70395
rect 32340 68805 32460 73395
rect 34740 73260 34860 79695
rect 35040 79605 35160 80160
rect 35640 80100 35760 80160
rect 35595 79905 35805 80100
rect 35040 76005 35160 78495
rect 35040 73305 35160 75795
rect 35340 75405 35460 76395
rect 35895 76200 36105 76395
rect 36540 76305 36660 79395
rect 35940 76140 36060 76200
rect 36840 75690 36960 79995
rect 37140 79305 37260 80160
rect 37740 79905 37860 80160
rect 37740 77505 37860 79695
rect 38640 79605 38760 80640
rect 38340 79005 38460 79395
rect 38640 76905 38760 78795
rect 38940 77805 39060 81195
rect 39195 80805 39405 80895
rect 39840 80640 39960 81795
rect 40140 81105 40260 83295
rect 40440 80805 40560 84795
rect 40740 81405 40860 88395
rect 42840 87105 42960 88695
rect 43440 88440 43560 88995
rect 44640 88905 44760 91260
rect 44640 88005 44760 88695
rect 44940 88305 45060 90495
rect 46740 89760 46860 91260
rect 48405 91140 48660 91260
rect 46440 89640 46860 89760
rect 41040 84105 41160 86895
rect 41340 83940 41460 84495
rect 41940 80640 42060 82995
rect 42540 80805 42660 85695
rect 42840 82005 42960 85395
rect 43140 83205 43260 87780
rect 43740 87405 43860 87960
rect 45240 85605 45360 87795
rect 45840 86505 45960 87960
rect 46440 86505 46560 89640
rect 47295 88500 47505 88695
rect 47340 88440 47460 88500
rect 43740 83940 43860 85395
rect 44895 84120 45105 84195
rect 44040 82605 44160 83460
rect 42840 81840 43095 82005
rect 42900 81795 43095 81840
rect 39240 79005 39360 79995
rect 39705 79395 39795 79605
rect 38805 76740 39060 76860
rect 37740 76140 37860 76695
rect 38940 76305 39060 76740
rect 39240 76605 39360 77895
rect 40140 77505 40260 79980
rect 40440 76905 40560 79995
rect 40740 78105 40860 80610
rect 41640 80100 41760 80160
rect 41595 79905 41805 80100
rect 42840 80190 42960 81495
rect 44340 80205 44460 82995
rect 44940 82860 45060 83910
rect 45240 82905 45360 85395
rect 45795 84000 46005 84195
rect 45840 83940 45960 84000
rect 46440 83940 46560 84495
rect 44640 82740 45060 82860
rect 44640 80805 44760 82740
rect 44940 80640 45060 81795
rect 45540 80805 45660 81795
rect 36240 75600 36360 75660
rect 36195 75405 36405 75600
rect 36240 74805 36360 75195
rect 34440 73140 34860 73260
rect 34140 72105 34260 72795
rect 34440 72390 34560 73140
rect 35340 72840 35460 73395
rect 35940 72840 36060 73695
rect 35040 72300 35160 72360
rect 35640 72300 35760 72360
rect 30840 67605 30960 68310
rect 30540 67140 30960 67260
rect 29895 65160 30105 65295
rect 29640 65100 30105 65160
rect 29640 65040 30060 65100
rect 29340 61005 29460 64560
rect 30240 64500 30360 64560
rect 30195 64305 30405 64500
rect 29640 63105 29760 64095
rect 26595 60600 26805 60795
rect 26640 60540 26760 60600
rect 26040 58560 26160 59895
rect 26340 58905 26460 60060
rect 26805 59760 27000 59790
rect 26805 59700 27060 59760
rect 26805 59595 27105 59700
rect 26895 59505 27105 59595
rect 27540 59505 27660 59895
rect 26040 58500 26460 58560
rect 26040 58440 26505 58500
rect 26295 58305 26505 58440
rect 26040 57240 26160 57795
rect 26640 57405 26760 58995
rect 27540 57660 27660 59295
rect 27840 59205 27960 60795
rect 28095 60705 28305 60795
rect 29340 60060 29460 60795
rect 29940 60705 30060 63195
rect 30840 61905 30960 67140
rect 31140 64305 31260 67095
rect 32340 67005 32460 67860
rect 32640 67305 32760 67695
rect 32940 67605 33060 70095
rect 32040 65040 32160 65895
rect 31740 64305 31860 64560
rect 31740 63660 31860 64095
rect 31740 63540 32160 63660
rect 29040 59940 29460 60060
rect 27240 57540 27660 57660
rect 27240 57240 27360 57540
rect 27840 57240 27960 57795
rect 28440 57405 28560 58095
rect 26340 56700 26460 56760
rect 25140 56205 25260 56580
rect 26295 56505 26505 56700
rect 25605 56295 25695 56475
rect 24840 53505 24960 54480
rect 25740 53205 25860 54795
rect 26040 53805 26160 54195
rect 26340 54105 26460 55980
rect 26640 55905 26760 56595
rect 28200 56760 28395 56805
rect 28140 56640 28395 56760
rect 28200 56595 28395 56640
rect 27540 56460 27660 56580
rect 28740 56505 28860 57795
rect 29040 57705 29160 59940
rect 29340 57405 29460 59595
rect 29640 59505 29760 60510
rect 30195 60600 30405 60795
rect 30240 60540 30360 60600
rect 31440 60105 31560 63495
rect 32040 62760 32160 63540
rect 32340 63060 32460 64560
rect 32940 63705 33060 67080
rect 32340 62940 32760 63060
rect 32040 62640 32460 62760
rect 30540 59205 30660 60060
rect 30240 57240 30360 57795
rect 27540 56340 27960 56460
rect 26940 55605 27060 55995
rect 27540 55605 27660 55995
rect 27840 55860 27960 56340
rect 27840 55740 28260 55860
rect 21240 45105 21360 46995
rect 21840 46905 21960 48960
rect 22440 45120 22560 47895
rect 22140 43905 22260 44460
rect 22305 43740 22560 43860
rect 22440 42105 22560 43740
rect 22740 42105 22860 44295
rect 23040 42060 23160 50595
rect 23340 49605 23460 49995
rect 24240 49605 24360 49995
rect 24000 49560 24195 49605
rect 23940 49440 24195 49560
rect 24000 49395 24195 49440
rect 23340 44205 23460 48795
rect 24540 47205 24660 52095
rect 24840 51705 24960 52080
rect 25740 52005 25860 52995
rect 26040 52605 26160 53595
rect 27240 52740 27360 55095
rect 28140 55005 28260 55740
rect 27795 53505 28005 53595
rect 26040 51705 26160 52395
rect 24840 49905 24960 51495
rect 25695 49500 25905 49695
rect 25740 49440 25860 49500
rect 26340 49440 26460 49995
rect 26640 49605 26760 51795
rect 26940 51705 27060 52260
rect 27540 51960 27660 52080
rect 27240 51840 27660 51960
rect 24840 48105 24960 49380
rect 25305 48840 25560 48960
rect 25140 47805 25260 48795
rect 25440 47205 25560 48495
rect 25740 46905 25860 48195
rect 26040 48105 26160 48960
rect 24240 45705 24360 46095
rect 25140 46005 25260 46395
rect 24240 44940 24360 45495
rect 24795 45000 25005 45195
rect 25440 45105 25560 45795
rect 24840 44940 24960 45000
rect 25695 45000 25905 45195
rect 25740 44940 25860 45000
rect 26340 44940 26460 46095
rect 26640 46005 26760 48795
rect 26940 48105 27060 49695
rect 27240 45405 27360 51840
rect 28140 51705 28260 54795
rect 28440 52905 28560 53895
rect 29040 53805 29160 57180
rect 29340 55605 29460 56595
rect 30540 56700 30660 56760
rect 30495 56505 30705 56700
rect 28740 52860 28860 53595
rect 29340 53205 29460 54195
rect 28740 52740 29160 52860
rect 29640 52740 29760 54495
rect 30840 52905 30960 56595
rect 31140 56505 31260 59895
rect 31440 56505 31560 59295
rect 31740 55905 31860 61695
rect 31995 60705 32205 60795
rect 32340 60720 32460 62640
rect 32640 61905 32760 62940
rect 33240 61005 33360 68595
rect 33840 68340 33960 70995
rect 34440 69405 34560 72180
rect 34995 72105 35205 72300
rect 35595 72105 35805 72300
rect 34440 67305 34560 67860
rect 34440 65040 34560 66195
rect 33840 62205 33960 64560
rect 33840 60540 33960 61680
rect 35040 61305 35160 69795
rect 35340 68520 35460 70395
rect 35940 70005 36060 70995
rect 36240 70605 36360 72195
rect 36540 70905 36660 73395
rect 35640 68340 35760 68895
rect 36540 68505 36660 69195
rect 36840 68205 36960 75480
rect 37140 73905 37260 75495
rect 38040 73905 38160 75660
rect 37740 72840 37860 73695
rect 38940 73305 39060 73695
rect 39240 73605 39360 76080
rect 39240 72405 39360 73080
rect 39195 72105 39405 72195
rect 38040 71505 38160 72060
rect 38040 69105 38160 71295
rect 39240 68205 39360 68895
rect 36240 67740 36660 67860
rect 35340 65205 35460 67395
rect 36540 66660 36660 67740
rect 36840 67005 36960 67995
rect 36540 66540 37095 66660
rect 38040 66405 38160 67260
rect 36240 65205 36360 65895
rect 36540 65505 36660 66195
rect 36840 65205 36960 65595
rect 36540 65040 36795 65160
rect 35340 64560 35460 64995
rect 37440 64905 37560 66195
rect 39540 66105 39660 76695
rect 40005 75660 40200 75705
rect 40005 75540 40260 75660
rect 40005 75495 40200 75540
rect 40305 73260 40500 73305
rect 40305 73095 40560 73260
rect 40440 72840 40560 73095
rect 41040 73005 41160 75495
rect 41340 73260 41460 77595
rect 41640 75705 41760 78195
rect 42540 76605 42660 79995
rect 43740 80100 43860 80160
rect 43095 79860 43305 79995
rect 43695 79905 43905 80100
rect 43095 79800 43560 79860
rect 43140 79740 43560 79800
rect 43140 76140 43260 79095
rect 43440 79005 43560 79740
rect 43740 75705 43860 77895
rect 41340 73140 41760 73260
rect 41340 72390 41460 72795
rect 39840 66705 39960 68895
rect 40440 68340 40560 69795
rect 41040 69705 41160 72195
rect 35340 64440 35760 64560
rect 35640 63405 35760 64440
rect 34440 60540 34560 61095
rect 35295 60660 35505 60795
rect 35205 60600 35505 60660
rect 35205 60540 35460 60600
rect 32640 59940 33060 60060
rect 32040 57405 32160 59295
rect 32640 57240 32760 58095
rect 32940 57405 33060 59940
rect 33240 57705 33360 60480
rect 33540 57405 33660 58695
rect 34140 58305 34260 60060
rect 34740 59760 34860 60060
rect 34740 59640 34995 59760
rect 32340 56700 32460 56760
rect 32295 56505 32505 56700
rect 33090 56580 33105 56700
rect 32895 56475 33105 56580
rect 32895 56400 33195 56475
rect 32940 56340 33195 56400
rect 31440 52740 31560 55695
rect 32040 55605 32160 56295
rect 33000 56265 33195 56340
rect 27540 49605 27660 51495
rect 28440 50805 28560 52380
rect 28140 49440 28260 50295
rect 29040 49605 29160 51195
rect 29940 50805 30060 52260
rect 30540 51405 30660 52695
rect 30795 52005 31005 52095
rect 30240 50505 30360 50895
rect 30240 49620 30360 49980
rect 30840 49905 30960 51795
rect 31140 51105 31260 52260
rect 31740 52200 31860 52260
rect 31695 52005 31905 52200
rect 32040 51705 32160 52095
rect 32340 49905 32460 54795
rect 32940 52740 33060 53595
rect 33840 53160 33960 57495
rect 34140 56805 34260 58095
rect 35040 57405 35160 59595
rect 35340 57420 35460 59895
rect 35640 59805 35760 63195
rect 35940 61005 36060 64560
rect 36240 60660 36360 64395
rect 37440 64005 37560 64695
rect 39840 64305 39960 66495
rect 40140 65205 40260 65895
rect 40440 65505 40560 66495
rect 41040 66405 41160 67860
rect 40740 65040 40860 65895
rect 41040 65805 41160 66195
rect 41340 65460 41460 67695
rect 41640 66105 41760 73140
rect 41940 72405 42060 73395
rect 42240 73005 42360 75195
rect 42540 74505 42660 75660
rect 44040 75660 44160 78795
rect 44640 77805 44760 79995
rect 45240 78705 45360 80160
rect 45540 78060 45660 79995
rect 45840 78405 45960 82695
rect 46140 82005 46260 83460
rect 47040 82305 47160 84495
rect 47640 84120 47760 87780
rect 47940 83940 48060 87195
rect 48540 87105 48660 91140
rect 48540 85305 48660 86295
rect 48540 83940 48660 85095
rect 48840 84705 48960 92895
rect 49440 91305 49560 91995
rect 49995 91800 50205 91995
rect 50040 91740 50160 91800
rect 50640 91740 50760 92595
rect 53040 91740 53160 92895
rect 50340 89205 50460 91260
rect 50940 90705 51060 91260
rect 51840 90705 51960 91710
rect 49140 86805 49260 88995
rect 52440 88440 52560 89595
rect 52740 88905 52860 91260
rect 53340 88005 53460 89895
rect 53640 89805 53760 91710
rect 54540 90705 54660 91260
rect 55740 90705 55860 92295
rect 57240 91740 57360 92295
rect 56340 89805 56460 91260
rect 54195 88500 54405 88695
rect 54240 88440 54360 88500
rect 55140 88305 55260 88695
rect 55905 88560 56100 88605
rect 55905 88440 56160 88560
rect 56640 88440 56760 90195
rect 56940 90105 57060 91260
rect 55905 88395 56100 88440
rect 50040 84120 50160 85995
rect 50340 85005 50460 87465
rect 50940 87405 51060 87960
rect 50640 83940 50760 85695
rect 47640 81105 47760 82395
rect 46995 80700 47205 80895
rect 47595 80805 47805 80895
rect 47040 80640 47160 80700
rect 47940 80205 48060 81195
rect 46440 79305 46560 80160
rect 47640 78705 47760 79995
rect 47895 79905 48105 79995
rect 48240 79305 48360 81495
rect 45540 77940 45960 78060
rect 44640 76320 44760 77280
rect 45240 76320 45360 77595
rect 44040 75540 44460 75660
rect 42540 73020 42660 73395
rect 41940 68505 42060 71880
rect 43440 71205 43560 72360
rect 41940 65805 42060 66495
rect 41340 65400 42060 65460
rect 41340 65340 42105 65400
rect 41895 65205 42105 65340
rect 42240 65160 42360 67395
rect 43140 67005 43260 69495
rect 43440 68505 43560 70995
rect 43740 68805 43860 70395
rect 44040 69705 44160 74595
rect 44340 74505 44460 75540
rect 45840 75660 45960 77940
rect 46740 76140 46860 77295
rect 47340 76140 47460 77295
rect 45840 75540 46260 75660
rect 45840 74505 45960 75195
rect 44940 72840 45060 73395
rect 45840 73005 45960 73395
rect 44640 72300 44760 72360
rect 44595 72105 44805 72300
rect 44205 69060 44400 69105
rect 44205 69000 44460 69060
rect 44205 68895 44505 69000
rect 44295 68805 44505 68895
rect 43905 68760 44100 68805
rect 43905 68595 44160 68760
rect 44040 68340 44160 68595
rect 44640 68340 44760 71895
rect 45240 70905 45360 72360
rect 45540 70605 45660 71895
rect 45240 67890 45360 68595
rect 43440 65460 43560 67695
rect 43740 65805 43860 67095
rect 45540 66705 45660 70395
rect 46140 70005 46260 75540
rect 46440 72360 46560 75480
rect 47040 73905 47160 75660
rect 47640 74205 47760 75480
rect 47940 73605 48060 76095
rect 48240 75405 48360 78495
rect 48540 76305 48660 82095
rect 49140 81705 49260 83895
rect 49395 80700 49605 80895
rect 50040 80805 50160 82695
rect 50340 82305 50460 83460
rect 49440 80640 49560 80700
rect 49140 80100 49260 80160
rect 48840 78360 48960 79995
rect 49095 79905 49305 80100
rect 49695 79905 49905 79980
rect 48840 78240 49260 78360
rect 48840 76140 48960 77895
rect 49140 77205 49260 78240
rect 50040 76140 50160 78495
rect 50340 78405 50460 81780
rect 50640 80205 50760 80895
rect 50940 80805 51060 82095
rect 51240 81105 51360 86895
rect 52140 86805 52260 87960
rect 55440 87990 55560 88395
rect 51540 83205 51660 84795
rect 52740 83940 52860 84795
rect 53340 84120 53460 87195
rect 53940 86805 54060 87960
rect 54540 86760 54660 87780
rect 54240 86640 54660 86760
rect 52440 83400 52560 83460
rect 52395 83205 52605 83400
rect 51540 80640 51660 82995
rect 52440 82605 52560 82995
rect 52140 80640 52260 82395
rect 52440 81105 52560 82080
rect 53040 82005 53160 83460
rect 53040 80805 53160 81195
rect 53340 80640 53460 82995
rect 53640 82305 53760 83295
rect 53940 82005 54060 86280
rect 54240 81360 54360 86640
rect 54840 83940 54960 86595
rect 55140 85005 55260 87780
rect 56340 87660 56460 87960
rect 56040 87540 56460 87660
rect 55440 84120 55560 85695
rect 54540 82860 54660 83295
rect 54540 82740 54795 82860
rect 54540 81705 54660 82380
rect 54240 81240 54660 81360
rect 54540 80805 54660 81240
rect 49740 75600 49860 75660
rect 49695 75405 49905 75600
rect 46440 72240 46860 72360
rect 47040 72300 47160 72360
rect 47640 72300 47760 72360
rect 46440 68505 46560 68895
rect 46740 68340 46860 72240
rect 46995 72105 47205 72300
rect 47595 72105 47805 72300
rect 47940 71760 48060 72180
rect 48240 71805 48360 74295
rect 47640 71640 48060 71760
rect 43440 65340 43860 65460
rect 42240 65040 42660 65160
rect 35940 60540 36360 60660
rect 36540 60540 36660 61995
rect 37140 61005 37260 61395
rect 37095 60600 37305 60795
rect 37140 60540 37260 60600
rect 34140 53805 34260 56595
rect 35040 56205 35160 56595
rect 33840 53040 34260 53160
rect 34140 52740 34260 53040
rect 34440 52905 34560 55995
rect 33240 51960 33360 52260
rect 33840 52200 33960 52260
rect 33795 52005 34005 52200
rect 33240 51840 33660 51960
rect 33540 51360 33660 51840
rect 33795 51705 34005 51795
rect 33540 51240 34095 51360
rect 34440 51360 34560 52095
rect 34305 51240 34560 51360
rect 23340 42405 23460 43095
rect 23040 41940 23460 42060
rect 22095 41700 22305 41895
rect 22140 41640 22260 41700
rect 23040 41205 23160 41595
rect 21240 40305 21360 41160
rect 21840 40605 21960 41160
rect 18795 37305 19005 37395
rect 17940 37140 18060 37200
rect 20295 37200 20505 37395
rect 20340 37140 20460 37200
rect 16440 35505 16560 35895
rect 15540 33300 15660 33360
rect 15495 33105 15705 33300
rect 15540 31005 15660 32895
rect 16140 32805 16260 33360
rect 16740 32505 16860 35595
rect 17340 34860 17460 35595
rect 17640 34905 17760 36660
rect 18540 35805 18660 36780
rect 19305 36660 19500 36705
rect 19305 36540 19560 36660
rect 19305 36495 19500 36540
rect 20640 36105 20760 36495
rect 17040 34740 17460 34860
rect 17040 34005 17160 34740
rect 17505 34440 17895 34560
rect 19140 33390 19260 34695
rect 20040 34020 20160 34995
rect 20640 33840 20760 35895
rect 20940 35205 21060 38595
rect 21240 34905 21360 37695
rect 21540 34305 21660 37395
rect 22395 37200 22605 37395
rect 22440 37140 22560 37200
rect 23040 37140 23160 40680
rect 23340 38805 23460 41940
rect 23640 41805 23760 44295
rect 23940 42405 24060 44460
rect 24540 44400 24660 44460
rect 24495 44205 24705 44400
rect 24240 42060 24360 42795
rect 24540 42405 24660 43095
rect 24105 41940 24360 42060
rect 23940 41640 24060 41880
rect 23595 40860 23805 40995
rect 23595 40800 24060 40860
rect 23640 40740 24060 40800
rect 22140 35505 22260 36660
rect 22740 36600 22860 36660
rect 22695 36405 22905 36600
rect 21840 33960 21960 34995
rect 21540 33840 21960 33960
rect 22395 33900 22605 34095
rect 22440 33840 22560 33900
rect 17340 32805 17460 33360
rect 17940 32505 18060 33360
rect 19140 32505 19260 33180
rect 19740 32805 19860 33180
rect 14940 29340 15060 29895
rect 19740 29805 19860 31695
rect 20340 30705 20460 33360
rect 15495 29520 15705 29595
rect 15240 28560 15360 28680
rect 14940 28440 15360 28560
rect 14340 26040 14460 26895
rect 14940 26220 15060 28440
rect 16140 28305 16260 29595
rect 17295 29400 17505 29595
rect 17340 29340 17460 29400
rect 19740 29340 19860 29595
rect 20340 29505 20460 30495
rect 17040 28560 17160 28860
rect 17040 28440 17460 28560
rect 16140 26040 16260 27195
rect 15240 25500 15360 25560
rect 15195 25305 15405 25500
rect 17040 25305 17160 28095
rect 17340 27060 17460 28440
rect 18540 27360 18660 29310
rect 18540 27240 18795 27360
rect 17340 26940 17760 27060
rect 14940 23505 15060 23895
rect 14295 21600 14505 21795
rect 14340 21540 14460 21600
rect 14940 21540 15060 23295
rect 13140 20640 13560 20760
rect 10740 17790 10860 19095
rect 12240 18240 12360 18795
rect 12840 18405 12960 19395
rect 8340 13740 8460 16995
rect 5340 11805 5460 13095
rect 5940 11505 6060 13260
rect 6540 12705 6660 13260
rect 9240 12705 9360 17265
rect 7740 11640 8460 11760
rect 5040 10440 5460 10560
rect 3240 6405 3360 10440
rect 5340 9990 5460 10440
rect 4140 8805 4260 9960
rect 6240 9900 6360 9960
rect 5340 9405 5460 9780
rect 6195 9705 6405 9900
rect 6840 9405 6960 9960
rect 2340 5940 2460 6000
rect 3105 5940 3360 6060
rect 3840 5940 3960 7095
rect 1440 4305 1560 5460
rect 3540 4905 3660 5460
rect 1440 2640 1560 3495
rect 2040 2640 2160 4095
rect 4140 3705 4260 5460
rect 4740 4905 4860 6195
rect 6240 5940 6360 7395
rect 7440 6705 7560 10395
rect 7395 6405 7605 6495
rect 6795 6000 7005 6195
rect 7740 6120 7860 11640
rect 8040 10605 8160 11295
rect 8340 11205 8460 11640
rect 8640 10440 8760 11595
rect 9240 10440 9360 10995
rect 9540 10605 9660 13995
rect 8940 9900 9060 9960
rect 8895 9705 9105 9900
rect 8940 8805 9060 9495
rect 6840 5940 6960 6000
rect 8340 5940 8460 7395
rect 5940 4905 6060 5460
rect 3840 2640 3960 3195
rect 4140 2805 4260 3495
rect 5940 3105 6060 4695
rect 8040 4605 8160 5460
rect 6240 2820 6360 3495
rect 7440 2640 7560 4095
rect 8040 2640 8160 3795
rect 4740 1005 4860 2595
rect 7140 2100 7260 2160
rect 7740 2100 7860 2160
rect 7095 1905 7305 2100
rect 7695 1905 7905 2100
rect 8640 1905 8760 5280
rect 9240 4605 9360 6495
rect 9540 5505 9660 5910
rect 9840 5205 9960 16995
rect 11040 13740 11160 18195
rect 12540 16305 12660 17580
rect 13140 17205 13260 20640
rect 14040 20505 14160 21060
rect 14340 18240 14460 20595
rect 14640 19005 14760 21060
rect 14040 17700 14160 17760
rect 13995 17505 14205 17700
rect 12840 16005 12960 16395
rect 11640 13305 11760 14295
rect 12795 13800 13005 13995
rect 12840 13740 12960 13800
rect 10740 11505 10860 13260
rect 14040 13290 14160 17295
rect 14640 15705 14760 17760
rect 14340 15540 14595 15660
rect 13140 12705 13260 13260
rect 11340 10440 11460 10995
rect 11940 10440 12060 11595
rect 12240 10605 12360 12495
rect 14040 11805 14160 13080
rect 14340 13005 14460 15540
rect 14940 15105 15060 17595
rect 15240 17505 15360 19995
rect 15540 19605 15660 23895
rect 15840 20805 15960 22095
rect 16140 19905 16260 22695
rect 17340 22305 17460 26595
rect 17640 22905 17760 26940
rect 18240 26040 18360 26595
rect 18840 26040 18960 27195
rect 19440 26205 19560 28860
rect 20640 28305 20760 32895
rect 20940 32505 21060 33360
rect 21540 33105 21660 33840
rect 23340 33405 23460 35295
rect 20940 29505 21060 31095
rect 21240 29340 21360 30795
rect 21840 29340 21960 30495
rect 22140 30105 22260 33180
rect 23040 32205 23160 33195
rect 23640 31005 23760 38295
rect 23940 38205 24060 40740
rect 24540 39705 24660 40995
rect 24840 40605 24960 42495
rect 25140 40905 25260 43395
rect 25440 41205 25560 44295
rect 25740 42405 25860 43995
rect 26040 43905 26160 44460
rect 26640 42105 26760 44460
rect 27240 44205 27360 44880
rect 27540 43605 27660 48795
rect 27840 47205 27960 48960
rect 29340 48960 29460 49410
rect 29340 48840 29760 48960
rect 27840 45105 27960 46395
rect 28440 44940 28560 45495
rect 28740 45405 28860 46395
rect 29040 45705 29160 48795
rect 28740 45225 28995 45405
rect 28800 45195 28995 45225
rect 29340 45105 29460 46695
rect 28140 43305 28260 44460
rect 29640 44460 29760 48840
rect 30840 48900 30960 48960
rect 30795 48705 31005 48900
rect 31095 48660 31305 48795
rect 31740 48705 31860 48960
rect 31095 48600 31560 48660
rect 31140 48540 31560 48600
rect 31740 48540 31995 48705
rect 30240 47505 30360 48495
rect 29340 44340 29760 44460
rect 29340 44205 29460 44340
rect 26640 41940 26895 42105
rect 26700 41910 26895 41940
rect 25905 41760 26100 41805
rect 25905 41640 26160 41760
rect 25905 41595 26100 41640
rect 28695 41700 28905 41895
rect 28740 41640 28860 41700
rect 24840 37140 24960 38595
rect 25440 37320 25560 38895
rect 24540 36600 24660 36660
rect 24495 36405 24705 36600
rect 25140 35805 25260 36660
rect 23940 32505 24060 35595
rect 25440 35205 25560 36495
rect 25740 36405 25860 37395
rect 26040 36105 26160 40695
rect 27540 40605 27660 41610
rect 27840 40005 27960 41295
rect 27405 38940 27795 39060
rect 27105 38640 27660 38760
rect 26340 37305 26460 37995
rect 27240 37905 27360 38295
rect 27540 38205 27660 38640
rect 26595 37200 26805 37395
rect 26640 37140 26760 37200
rect 26940 36600 27060 36660
rect 24840 34605 24960 34995
rect 24495 33900 24705 34095
rect 24540 33840 24660 33900
rect 25140 33840 25260 34395
rect 25440 34005 25560 34680
rect 26040 34605 26160 35580
rect 26340 34605 26460 36480
rect 26895 36405 27105 36600
rect 28140 36105 28260 40695
rect 28440 40605 28560 41160
rect 28440 37305 28560 39795
rect 28740 37320 28860 38895
rect 29340 38205 29460 43995
rect 29640 41805 29760 43995
rect 29940 42105 30060 45495
rect 30240 45105 30360 47295
rect 30495 45405 30705 45495
rect 30840 44940 30960 47895
rect 31140 46005 31260 48195
rect 31440 46605 31560 48540
rect 31800 48495 31995 48540
rect 31740 45105 31860 47895
rect 32340 47505 32460 48960
rect 32640 47805 32760 48795
rect 32940 48705 33060 49995
rect 33240 46905 33360 50895
rect 33840 50505 33960 50895
rect 34740 50805 34860 55695
rect 35040 50205 35160 55395
rect 35640 54705 35760 56295
rect 35940 56205 36060 60540
rect 36840 57405 36960 60060
rect 37740 57705 37860 64095
rect 40440 63405 40560 64395
rect 41040 64005 41160 64560
rect 38040 58605 38160 62595
rect 38640 62505 38760 62895
rect 39195 60600 39405 60795
rect 39540 60705 39660 61695
rect 39840 61605 39960 63195
rect 40305 61395 40395 61605
rect 39240 60540 39360 60600
rect 39840 58605 39960 60795
rect 39195 58305 39405 58395
rect 39300 57990 39600 58005
rect 37095 57300 37305 57495
rect 37140 57240 37260 57300
rect 38340 57240 38460 57795
rect 39405 57795 39495 57990
rect 35340 52905 35460 54495
rect 35640 52740 35760 53595
rect 36240 52905 36360 55095
rect 36540 55005 36660 56760
rect 34140 49440 34260 49995
rect 33540 48105 33660 48795
rect 33840 47505 33960 48960
rect 34740 48105 34860 48960
rect 32040 44760 32160 46395
rect 31740 44640 32160 44760
rect 30540 44400 30660 44460
rect 30495 44205 30705 44400
rect 30240 41640 30360 43095
rect 31440 42960 31560 44295
rect 31140 42840 31560 42960
rect 30840 42405 30960 42795
rect 30240 40305 30360 40695
rect 29295 37200 29505 37395
rect 29340 37140 29460 37200
rect 26700 34560 26895 34605
rect 26640 34395 26895 34560
rect 26640 34020 26760 34395
rect 27240 33840 27360 34695
rect 27840 34305 27960 35595
rect 28140 34005 28260 34995
rect 28440 34005 28560 36495
rect 28740 35205 28860 36195
rect 29040 36105 29160 36660
rect 24240 32205 24360 33195
rect 25740 32805 25860 33810
rect 28995 33900 29205 34095
rect 29340 34005 29460 35595
rect 29640 35505 29760 36495
rect 29940 34260 30060 36795
rect 30240 36705 30360 40095
rect 30540 39405 30660 41160
rect 31140 39105 31260 42840
rect 31440 41805 31560 42495
rect 31740 41805 31860 44640
rect 32040 42405 32160 44295
rect 32340 43305 32460 46395
rect 32640 45105 32760 45495
rect 32940 44940 33060 46095
rect 34140 46005 34260 47895
rect 34740 46605 34860 47580
rect 35040 46260 35160 48495
rect 35340 47805 35460 51795
rect 36540 50805 36660 53895
rect 35640 49905 35760 50595
rect 35940 49605 36060 50595
rect 36840 50505 36960 56295
rect 37140 53460 37260 54195
rect 37440 54105 37560 56595
rect 38040 55605 38160 56760
rect 37140 53340 37560 53460
rect 37440 52740 37560 53340
rect 38340 52905 38460 56295
rect 38640 56205 38760 56760
rect 38640 53205 38760 55995
rect 39540 54960 39660 57195
rect 39840 56505 39960 58080
rect 39540 54840 39960 54960
rect 38040 52740 38295 52860
rect 39540 52860 39660 54495
rect 39840 54105 39960 54840
rect 40140 54405 40260 61080
rect 40740 60540 40860 62295
rect 41640 60705 41760 64560
rect 40440 58005 40560 59880
rect 41595 59805 41805 59895
rect 40440 57405 40560 57795
rect 40695 57705 40905 57795
rect 40695 57300 40905 57495
rect 40740 57240 40860 57300
rect 41340 57240 41460 58095
rect 41940 58005 42060 64095
rect 42240 61005 42360 64395
rect 42495 61305 42705 61395
rect 42495 61200 42795 61305
rect 42540 61140 42795 61200
rect 42600 61095 42795 61140
rect 43140 60660 43260 62595
rect 43440 62505 43560 64995
rect 43140 60540 43560 60660
rect 42240 59940 42495 60060
rect 41940 56805 42060 57480
rect 42240 57405 42360 59940
rect 43140 59505 43260 59895
rect 43440 57705 43560 60540
rect 43740 60105 43860 65340
rect 44040 65205 44160 66495
rect 45840 65160 45960 66195
rect 45840 65040 46260 65160
rect 44400 64560 44595 64605
rect 44340 64440 44595 64560
rect 44400 64395 44595 64440
rect 45240 64005 45360 64560
rect 47040 63060 47160 67395
rect 46740 62940 47160 63060
rect 44340 60705 44460 62895
rect 45240 60540 45360 62295
rect 44040 59460 44160 60495
rect 43740 59340 44160 59460
rect 43740 58305 43860 59340
rect 43740 57360 43860 58095
rect 43440 57240 43860 57360
rect 39540 52740 40260 52860
rect 37740 52200 37860 52260
rect 37140 49605 37260 52095
rect 37695 52005 37905 52200
rect 38640 51705 38760 52395
rect 40140 52260 40260 52740
rect 37395 50205 37605 50295
rect 35640 47205 35760 49380
rect 36240 48900 36360 48960
rect 35940 48405 36060 48795
rect 36195 48705 36405 48900
rect 34740 46140 35160 46260
rect 34440 44940 34560 45495
rect 34740 45405 34860 46140
rect 32640 43905 32760 44295
rect 32640 42105 32760 42795
rect 32940 42360 33060 43995
rect 33240 42705 33360 44460
rect 33495 43905 33705 43995
rect 32940 42240 33360 42360
rect 32640 41640 32760 41895
rect 30240 34605 30360 35295
rect 29940 34140 30195 34260
rect 29040 33840 29160 33900
rect 26205 33360 26400 33405
rect 26205 33240 26460 33360
rect 26940 33300 27060 33360
rect 26205 33195 26400 33240
rect 26895 33105 27105 33300
rect 23040 29520 23160 30795
rect 23940 30705 24060 31095
rect 24240 30705 24360 31680
rect 24840 31005 24960 32595
rect 24840 30405 24960 30795
rect 23640 29340 23760 30195
rect 25140 30060 25260 31995
rect 25740 30105 25860 31395
rect 24840 29940 25260 30060
rect 24840 29340 24960 29940
rect 16440 21705 16560 22095
rect 16995 21600 17205 21795
rect 17940 21720 18060 25395
rect 19140 25005 19260 25560
rect 19740 23205 19860 28095
rect 20040 25905 20160 26295
rect 20940 26040 21060 26895
rect 21540 26505 21660 28860
rect 22440 26805 22560 29295
rect 20640 25005 20760 25560
rect 18495 22005 18705 22095
rect 17040 21540 17160 21600
rect 17640 21540 17895 21660
rect 18540 21540 18660 21795
rect 15840 19740 16095 19860
rect 15540 14205 15660 18195
rect 15840 17505 15960 19740
rect 16440 19305 16560 20895
rect 16740 20205 16860 21060
rect 17340 21000 17460 21060
rect 18840 21000 18960 21060
rect 17295 20805 17505 21000
rect 18795 20805 19005 21000
rect 17040 18240 17160 19095
rect 15195 13920 15405 13995
rect 15840 13740 15960 14895
rect 16140 14805 16260 17595
rect 16740 16305 16860 17760
rect 17340 17700 17460 17760
rect 17295 17505 17505 17700
rect 17940 17505 18060 19095
rect 18840 18240 18960 19695
rect 19440 19005 19560 21060
rect 20040 20805 20160 22095
rect 18540 17700 18660 17760
rect 18495 17505 18705 17700
rect 19140 16905 19260 17760
rect 19140 16305 19260 16695
rect 16140 14205 16260 14595
rect 17940 14205 18060 14895
rect 10140 9705 10260 10395
rect 11640 9405 11760 9960
rect 12540 8805 12660 10995
rect 11940 5505 12060 7095
rect 12840 7005 12960 10995
rect 14940 10620 15060 13260
rect 15540 13200 15660 13260
rect 15495 13005 15705 13200
rect 16440 12105 16560 13995
rect 17295 13800 17505 13995
rect 17895 13800 18105 13995
rect 17340 13740 17460 13800
rect 17940 13740 18060 13800
rect 18540 13290 18660 14595
rect 19440 13740 19560 14295
rect 19740 14205 19860 17595
rect 20040 15705 20160 18795
rect 20340 17505 20460 19395
rect 20640 17790 20760 22095
rect 21240 21540 21360 23895
rect 21540 22305 21660 25695
rect 21840 22305 21960 26595
rect 23040 26040 23160 28095
rect 23340 27405 23460 28860
rect 23640 26205 23760 26895
rect 22740 24705 22860 25560
rect 23940 23805 24060 27195
rect 24240 26805 24360 29310
rect 24240 25005 24360 26280
rect 24540 26205 24660 28695
rect 24840 26040 24960 27195
rect 25140 27105 25260 28860
rect 26040 28860 26160 32295
rect 26340 29505 26460 32895
rect 27240 29760 27360 32895
rect 27540 31605 27660 33360
rect 26940 29640 27360 29760
rect 26940 29340 27060 29640
rect 27495 29400 27705 29595
rect 27840 29505 27960 33195
rect 27540 29340 27660 29400
rect 26040 28740 26760 28860
rect 25440 27405 25560 28095
rect 25740 28005 25860 28695
rect 26640 28560 26760 28740
rect 26640 28440 27060 28560
rect 25395 26100 25605 26295
rect 26340 26205 26460 28395
rect 26940 28005 27060 28440
rect 25440 26040 25560 26100
rect 21840 22095 22095 22305
rect 21840 21540 21960 22095
rect 22440 22005 22560 22995
rect 24540 22905 24660 25395
rect 25740 25500 25860 25560
rect 25695 25305 25905 25500
rect 22740 21090 22860 22395
rect 23340 21540 23460 22695
rect 23940 21540 24060 22395
rect 24240 22005 24360 22695
rect 23640 21000 23760 21060
rect 22005 20595 22095 20805
rect 22740 19005 22860 20880
rect 23595 20805 23805 21000
rect 23205 20595 23295 20805
rect 23340 18240 23460 19395
rect 24240 18960 24360 20880
rect 24240 18840 24660 18960
rect 24240 18105 24360 18495
rect 21840 17700 21960 17760
rect 21240 16605 21360 17580
rect 21795 17505 22005 17700
rect 22140 16905 22260 17595
rect 22740 16605 22860 17760
rect 20040 14505 20160 15495
rect 23640 14805 23760 17760
rect 20805 14640 21060 14760
rect 20640 13920 20760 14595
rect 16440 10440 16560 10995
rect 13140 8205 13260 9795
rect 14940 9960 15060 10410
rect 13740 9105 13860 9780
rect 14340 8805 14460 9960
rect 14940 9840 15660 9960
rect 16140 8805 16260 9960
rect 13140 6360 13260 7995
rect 17040 7905 17160 10395
rect 17340 9405 17460 11895
rect 17640 11205 17760 13260
rect 18540 10620 18660 10995
rect 19095 10605 19305 10695
rect 19440 9990 19560 10995
rect 20340 10620 20460 13260
rect 20940 12705 21060 14640
rect 23505 13995 23595 14205
rect 22395 13800 22605 13995
rect 22440 13740 22560 13800
rect 24240 13905 24360 16095
rect 24540 15405 24660 18840
rect 24540 13920 24660 14295
rect 24840 14205 24960 21795
rect 25140 21105 25260 24795
rect 26040 24405 26160 25395
rect 26340 24705 26460 25680
rect 26640 25005 26760 27795
rect 27240 27405 27360 28860
rect 27495 26100 27705 26295
rect 27540 26040 27660 26100
rect 28140 26040 28260 33195
rect 29505 33360 29700 33405
rect 29505 33195 29760 33360
rect 28395 32805 28605 32895
rect 29640 32505 29760 33195
rect 28440 29205 28560 31695
rect 29640 31305 29760 31980
rect 29940 31605 30060 33195
rect 30240 31605 30360 34080
rect 30540 32505 30660 37995
rect 31440 37605 31560 41280
rect 32340 41100 32460 41160
rect 31740 38760 31860 40995
rect 32295 40905 32505 41100
rect 33240 40905 33360 42240
rect 31740 38640 31995 38760
rect 32040 38205 32160 38595
rect 31005 37560 31200 37605
rect 31005 37395 31260 37560
rect 31140 37140 31260 37395
rect 31995 37200 32205 37395
rect 32340 37305 32460 39795
rect 32040 37140 32160 37200
rect 30840 34005 30960 35895
rect 31440 35505 31560 36480
rect 31740 34905 31860 35295
rect 32640 34305 32760 40695
rect 32940 34605 33060 37395
rect 33240 37305 33360 39195
rect 33540 38760 33660 43095
rect 33840 41805 33960 42495
rect 34140 42105 34260 44295
rect 34740 42705 34860 44460
rect 35340 44400 35460 44460
rect 35295 44205 35505 44400
rect 35040 43005 35160 43995
rect 35640 43860 35760 44295
rect 35940 44205 36060 45795
rect 35340 43740 35760 43860
rect 34440 41640 34560 42195
rect 35340 41805 35460 43740
rect 36240 43605 36360 46395
rect 36540 43905 36660 48195
rect 36840 47205 36960 48960
rect 37140 46605 37260 48795
rect 37440 48705 37560 49995
rect 37740 47805 37860 50895
rect 38295 50505 38505 50595
rect 37140 44940 37260 45495
rect 38040 45060 38160 50295
rect 38940 50205 39060 52095
rect 39240 51960 39360 52260
rect 39840 52140 40260 52260
rect 39240 51840 39660 51960
rect 39540 51405 39660 51840
rect 38340 49605 38460 49980
rect 39540 49605 39660 51195
rect 39240 48900 39360 48960
rect 39195 48705 39405 48900
rect 38505 48495 38595 48675
rect 38640 45105 38760 46695
rect 38040 44940 38460 45060
rect 35940 41760 36060 42795
rect 36840 42105 36960 43995
rect 35940 41640 36195 41760
rect 33840 40605 33960 40995
rect 34140 39705 34260 41160
rect 34740 40860 34860 41160
rect 34440 40740 34860 40860
rect 33540 38640 33960 38760
rect 33540 37140 33660 38295
rect 33840 37305 33960 38640
rect 34440 38205 34560 40740
rect 34140 36540 34560 36660
rect 28995 29520 29205 29595
rect 29700 29460 29895 29505
rect 29640 29340 29895 29460
rect 29700 29295 29895 29340
rect 29040 25590 29160 27195
rect 27240 25500 27360 25560
rect 27195 25305 27405 25500
rect 25800 21960 25995 22005
rect 25740 21795 25995 21960
rect 25740 21720 25905 21795
rect 26640 19605 26760 23595
rect 26940 22905 27060 23595
rect 27840 23505 27960 25560
rect 26940 21705 27060 22695
rect 27840 22005 27960 22695
rect 28140 22305 28260 25095
rect 28440 22005 28560 25560
rect 28740 23205 28860 24495
rect 29340 24105 29460 26295
rect 29640 26205 29760 28095
rect 29940 27405 30060 28695
rect 30240 26520 30360 31395
rect 30540 30705 30660 31095
rect 30840 29760 30960 33195
rect 31740 32760 31860 33360
rect 31740 32640 32160 32760
rect 31140 30405 31260 32295
rect 31440 30705 31560 31095
rect 31740 29805 31860 31095
rect 30540 29640 30960 29760
rect 30540 28305 30660 29640
rect 31095 29460 31305 29595
rect 32040 29520 32160 32640
rect 32340 31305 32460 33795
rect 33240 33840 33360 36195
rect 33840 34305 33960 36495
rect 34440 34305 34560 36540
rect 34740 35805 34860 38895
rect 35040 37305 35160 40995
rect 35640 39705 35760 41160
rect 36240 39105 36360 40695
rect 36840 40560 36960 40995
rect 37140 40905 37260 43695
rect 36840 40440 37260 40560
rect 35295 37200 35505 37395
rect 36240 37305 36360 38580
rect 36540 38505 36660 40395
rect 35340 37140 35460 37200
rect 36540 36690 36660 37095
rect 35040 36105 35160 36495
rect 33840 33840 34560 33960
rect 35340 33840 35460 34995
rect 35595 34005 35805 34095
rect 32640 32760 32760 33780
rect 32895 33105 33105 33195
rect 33090 33000 33105 33105
rect 32640 32640 33060 32760
rect 32295 30405 32505 30495
rect 30840 29400 31305 29460
rect 30840 29340 31260 29400
rect 30840 28605 30960 29340
rect 32340 29340 32460 29880
rect 31440 26220 31560 27795
rect 31740 27705 31860 28860
rect 32940 27705 33060 32640
rect 33240 31905 33360 32895
rect 33540 32505 33660 33360
rect 33195 30405 33405 30495
rect 33540 30105 33660 30795
rect 34140 29805 34260 32595
rect 34440 32505 34560 33840
rect 35040 33105 35160 33360
rect 35040 32940 35295 33105
rect 35100 32895 35295 32940
rect 35505 32940 35760 33060
rect 35040 30405 35160 32595
rect 34440 29460 34560 29895
rect 34140 29340 34560 29460
rect 31740 26205 31860 26595
rect 30540 25305 30660 25560
rect 31095 25305 31305 25395
rect 30540 25140 30795 25305
rect 30600 25095 30795 25140
rect 31440 24105 31560 26010
rect 32640 26040 32760 26595
rect 33240 26205 33360 27795
rect 31740 22860 31860 25395
rect 32040 24060 32160 25095
rect 32340 24405 32460 25380
rect 32040 23940 32460 24060
rect 32340 23205 32460 23940
rect 31740 22740 31980 22860
rect 27405 21960 27600 22005
rect 27405 21795 27660 21960
rect 27540 21540 27660 21795
rect 28095 21600 28305 21780
rect 28140 21540 28260 21600
rect 27840 21000 27960 21060
rect 27795 20805 28005 21000
rect 28740 20805 28860 21510
rect 29040 21105 29160 22695
rect 29640 21705 29760 22095
rect 30840 21540 30960 22395
rect 32040 21540 32160 22695
rect 32340 22005 32460 22680
rect 32940 21705 33060 25380
rect 33540 24705 33660 28395
rect 33840 26205 33960 28860
rect 34740 26805 34860 28995
rect 35040 28005 35160 29595
rect 33840 22605 33960 25395
rect 34140 25005 34260 25560
rect 34440 23505 34560 24495
rect 33240 21105 33360 22395
rect 27240 19905 27360 20295
rect 29640 19905 29760 20895
rect 29940 20760 30060 21060
rect 29940 20640 30360 20760
rect 25395 18300 25605 18495
rect 27840 18420 27960 18795
rect 29640 18660 29760 19695
rect 29340 18540 29760 18660
rect 25440 18240 25560 18300
rect 29340 18240 29460 18540
rect 29940 18240 30060 20295
rect 30240 18405 30360 20640
rect 30795 18300 31005 18495
rect 30840 18240 30960 18300
rect 31440 18240 31560 20880
rect 31740 20505 31860 21060
rect 32340 20505 32460 21060
rect 31740 19905 31860 20295
rect 31740 19440 32295 19560
rect 31740 18705 31860 19440
rect 26940 17790 27060 18195
rect 23640 13290 23760 13680
rect 25440 13290 25560 15195
rect 25740 15105 25860 17760
rect 25740 13920 25860 14895
rect 26340 14505 26460 17760
rect 26940 13740 27060 17580
rect 27540 13290 27660 17580
rect 22140 10605 22260 13260
rect 22740 10440 22860 11895
rect 24840 10620 24960 11595
rect 25500 10560 25695 10605
rect 25440 10440 25695 10560
rect 25500 10395 25695 10440
rect 18240 9900 18360 9960
rect 18195 9705 18405 9900
rect 19905 9960 20100 10005
rect 19905 9840 20160 9960
rect 19905 9795 20100 9840
rect 12840 6240 13260 6360
rect 12840 5940 12960 6240
rect 13440 5940 13560 6795
rect 10740 5400 10860 5460
rect 10140 4905 10260 5295
rect 10695 5205 10905 5400
rect 8940 2190 9060 3195
rect 9840 2640 9960 4095
rect 11040 3060 11160 3795
rect 11340 3405 11460 5460
rect 14040 5460 14160 6795
rect 14340 5505 14460 7395
rect 14940 5940 15060 7695
rect 15540 5940 15660 7395
rect 13140 5400 13260 5460
rect 13095 5205 13305 5400
rect 13740 5340 14160 5460
rect 12240 3105 12360 4695
rect 13740 4305 13860 5340
rect 13995 4905 14205 4995
rect 11040 2940 11460 3060
rect 10440 2640 11160 2760
rect 10140 2100 10260 2160
rect 10095 1905 10305 2100
rect 11040 1305 11160 2640
rect 11340 705 11460 2940
rect 12540 2640 12660 3795
rect 13140 2805 13260 3195
rect 13440 1605 13560 3795
rect 13740 2505 13860 4095
rect 14040 2205 14160 4695
rect 15840 4005 15960 5460
rect 14940 2820 15060 3795
rect 16440 3705 16560 7695
rect 17640 7005 17760 7395
rect 16905 6060 17100 6105
rect 16905 5940 17160 6060
rect 17640 5940 17760 6795
rect 18240 6105 18360 7995
rect 16905 5895 17100 5940
rect 19140 5940 19260 6795
rect 16740 4905 16860 5295
rect 16440 3060 16560 3495
rect 16140 2940 16560 3060
rect 16140 2640 16260 2940
rect 16440 2100 16560 2160
rect 14640 1905 14805 1980
rect 16395 1905 16605 2100
rect 17340 1905 17460 2595
rect 17640 1905 17760 3495
rect 18540 2640 18660 4095
rect 19140 2640 19260 4695
rect 19440 3705 19560 5460
rect 20640 4905 20760 7395
rect 21240 7005 21360 9795
rect 22140 9405 22260 10395
rect 26040 10005 26160 12195
rect 26640 11805 26760 13260
rect 27240 11205 27360 11595
rect 27840 10905 27960 16395
rect 28740 16305 28860 18195
rect 28740 15705 28860 16095
rect 28440 13740 28560 14595
rect 28995 13800 29205 13995
rect 29640 13905 29760 17760
rect 32340 17790 32460 18795
rect 32940 18660 33060 20895
rect 33240 18705 33360 20580
rect 34740 20505 34860 23895
rect 35340 23460 35460 32295
rect 35640 31605 35760 32940
rect 35940 30105 36060 34095
rect 36240 32505 36360 34395
rect 36540 33705 36660 34395
rect 36840 34305 36960 40095
rect 37140 37305 37260 40440
rect 37440 40305 37560 43395
rect 37740 41805 37860 42195
rect 38040 42105 38160 43095
rect 38340 42405 38460 44940
rect 38940 44940 39060 47295
rect 39540 46905 39660 48795
rect 39540 44940 39660 45795
rect 39840 45405 39960 52140
rect 40140 49560 40260 49995
rect 40440 49905 40560 56595
rect 41040 54705 41160 56760
rect 44040 56790 44160 58395
rect 44340 57405 44460 59895
rect 45540 59940 45960 60060
rect 45540 58005 45660 59940
rect 46740 58605 46860 62940
rect 47340 60660 47460 68295
rect 47640 67605 47760 71640
rect 48540 68505 48660 72795
rect 48840 69705 48960 75195
rect 49440 74205 49560 74595
rect 49740 73020 49860 73395
rect 49140 70005 49260 70395
rect 48840 68340 48960 69495
rect 48240 66405 48360 67860
rect 49440 66405 49560 71295
rect 49740 68505 49860 71895
rect 50340 71505 50460 75480
rect 50640 73005 50760 79680
rect 50940 78105 51060 79995
rect 51540 77505 51660 79695
rect 51840 79005 51960 80160
rect 52440 78705 52560 79980
rect 54240 79605 54360 79980
rect 51540 76140 51660 77295
rect 52740 76305 52860 77895
rect 54540 77805 54660 79995
rect 50940 74505 51060 76095
rect 53040 75705 53160 77595
rect 53340 76605 53460 76995
rect 53940 76320 54060 76995
rect 54540 76140 54660 77595
rect 54840 76305 54960 82695
rect 51840 73905 51960 75660
rect 52140 74205 52260 74595
rect 50940 72840 51060 73695
rect 51540 72840 51660 73395
rect 52440 72360 52560 74895
rect 53340 74805 53460 76080
rect 53940 73005 54060 74595
rect 51240 71805 51360 72360
rect 51840 71805 51960 72360
rect 52440 72240 52860 72360
rect 49740 67860 49860 68295
rect 50040 68205 50160 70695
rect 52440 68205 52560 68895
rect 52740 68505 52860 72240
rect 53640 71205 53760 72360
rect 53340 69705 53460 70095
rect 53640 69705 53760 70995
rect 53940 68340 54060 72195
rect 54240 71805 54360 72795
rect 54240 68505 54360 70395
rect 49740 67740 50160 67860
rect 47940 63705 48060 64560
rect 48840 64440 49260 64560
rect 49140 64005 49260 64440
rect 48840 61905 48960 62895
rect 47040 60540 47460 60660
rect 47040 58005 47160 60540
rect 49140 60360 49260 63795
rect 49440 61305 49560 65595
rect 49740 61605 49860 67095
rect 50040 65805 50160 67740
rect 51240 66105 51360 67260
rect 50040 60540 50160 61095
rect 50340 61005 50460 64560
rect 50940 60660 51060 64560
rect 51840 63705 51960 65595
rect 52440 65220 52560 67395
rect 53340 67305 53460 67860
rect 53040 65040 53160 65595
rect 53640 65205 53760 66495
rect 52740 61905 52860 64560
rect 53640 63105 53760 64095
rect 53940 62205 54060 65895
rect 54240 64005 54360 67095
rect 54540 65505 54660 75195
rect 54840 74805 54960 75495
rect 55140 75405 55260 82395
rect 56040 82005 56160 87540
rect 56940 86505 57060 86895
rect 57840 86805 57960 93495
rect 56640 82305 56760 83460
rect 57540 80805 57660 83895
rect 57840 83505 57960 85695
rect 58140 84105 58260 93795
rect 58440 91920 58560 92295
rect 58695 91920 58905 91995
rect 60240 91905 60360 92295
rect 58440 91305 58560 91710
rect 58695 90960 58905 91095
rect 59640 91200 59760 91260
rect 59595 91005 59805 91200
rect 58695 90900 59160 90960
rect 58740 90840 59160 90900
rect 59040 88440 59160 90840
rect 59640 88440 59760 88995
rect 59340 87705 59460 87960
rect 60240 87705 60360 90795
rect 60540 89205 60660 91710
rect 61005 91260 61200 91305
rect 61005 91140 61260 91260
rect 61005 91095 61200 91140
rect 62040 91005 62160 91695
rect 62340 90405 62460 91710
rect 63240 90705 63360 91260
rect 64440 91260 64560 92295
rect 65340 91920 65460 93195
rect 65640 93105 65760 93495
rect 65940 91740 66060 92295
rect 64140 91140 64560 91260
rect 63540 90105 63660 90795
rect 63840 90360 63960 91080
rect 64140 90705 64260 91140
rect 63840 90240 64260 90360
rect 62940 89505 63060 89895
rect 62040 88620 62160 88995
rect 64140 88905 64260 90240
rect 64440 88905 64560 90795
rect 65040 90405 65160 91260
rect 63795 88500 64005 88695
rect 63840 88440 63960 88500
rect 58440 83940 58560 85995
rect 59040 85305 59160 86295
rect 59340 85605 59460 87495
rect 61140 87405 61260 87780
rect 61740 87105 61860 87960
rect 62790 87795 62805 87900
rect 62595 87705 62805 87795
rect 63540 87900 63660 87960
rect 63495 87705 63705 87900
rect 65040 87990 65160 89880
rect 65340 88905 65460 89895
rect 65640 88905 65760 91260
rect 65940 88440 66060 90495
rect 66540 90105 66660 93495
rect 71940 91740 72060 92295
rect 68340 91290 68460 91695
rect 66840 89505 66960 91080
rect 67740 90705 67860 91080
rect 66495 88500 66705 88695
rect 66540 88440 66660 88500
rect 67140 87990 67260 89595
rect 67440 89205 67560 90495
rect 68040 88440 68160 88995
rect 68340 88860 68460 91080
rect 68640 90705 68760 91395
rect 68340 88740 68760 88860
rect 68640 88440 68760 88740
rect 69240 88605 69360 88995
rect 69540 87990 69660 89595
rect 64140 87105 64260 87795
rect 66240 87405 66360 87960
rect 65940 87240 66195 87360
rect 57840 80640 57960 82695
rect 58140 82605 58260 83295
rect 58740 82305 58860 83460
rect 59340 82560 59460 83295
rect 59940 82905 60060 85395
rect 60240 84105 60360 84795
rect 60540 84705 60660 86295
rect 60840 83940 60960 86595
rect 63540 83940 63660 85695
rect 65640 84705 65760 86895
rect 65640 84105 65760 84495
rect 59340 82440 59760 82560
rect 58440 80640 58560 81795
rect 59640 81705 59760 82440
rect 59040 80805 59160 81495
rect 60240 81060 60360 83295
rect 60540 82905 60660 83460
rect 61140 82905 61260 83460
rect 62040 82260 62160 83910
rect 62640 83400 62760 83460
rect 62595 83205 62805 83400
rect 63240 82305 63360 83460
rect 62040 82140 62295 82260
rect 60240 80940 60660 81060
rect 59205 80640 59460 80760
rect 60540 80640 60660 80940
rect 56040 79005 56160 80160
rect 55740 77505 55860 78495
rect 56640 78405 56760 80160
rect 57240 79605 57360 80595
rect 58140 79860 58260 80160
rect 57840 79740 58260 79860
rect 57405 77340 57660 77460
rect 55440 73305 55560 76695
rect 56640 76140 56760 76695
rect 57240 76140 57360 77295
rect 57540 76905 57660 77340
rect 55740 75105 55860 75495
rect 56340 75360 56460 75660
rect 56340 75240 56760 75360
rect 56340 73005 56460 74595
rect 56640 74205 56760 75240
rect 56940 75105 57060 75660
rect 57840 75405 57960 79740
rect 58740 79005 58860 79980
rect 59040 78705 59160 79980
rect 58140 76305 58260 78495
rect 59340 78060 59460 80640
rect 61140 79605 61260 81495
rect 59640 78705 59760 79095
rect 59040 77940 59460 78060
rect 58440 76140 58560 76995
rect 59040 76305 59160 77940
rect 59340 76905 59460 77595
rect 59640 76260 59760 78495
rect 59340 76140 59760 76260
rect 58740 75600 58860 75660
rect 58695 75405 58905 75600
rect 57240 74205 57360 74595
rect 56940 72840 57060 73695
rect 54840 71805 54960 72795
rect 55440 70605 55560 72360
rect 54840 65160 54960 70095
rect 55440 68340 55560 70080
rect 56640 67905 56760 70695
rect 55740 66705 55860 67860
rect 55740 65460 55860 65895
rect 55740 65340 56160 65460
rect 56040 65250 56160 65340
rect 54540 65040 54960 65160
rect 54540 62805 54660 65040
rect 54840 63105 54960 64395
rect 55140 64005 55260 64560
rect 50805 60540 51060 60660
rect 49140 60240 49395 60360
rect 44895 57300 45105 57495
rect 44940 57240 45060 57300
rect 41940 55605 42060 56280
rect 40740 50505 40860 54195
rect 41940 53205 42060 55395
rect 42840 53805 42960 56295
rect 43140 54405 43260 56760
rect 45840 56505 45960 57495
rect 43440 55305 43560 56295
rect 41295 52800 41505 52995
rect 41340 52740 41460 52800
rect 41940 52740 42060 52995
rect 42795 52905 43005 52995
rect 43095 52800 43305 52995
rect 43140 52740 43260 52800
rect 43740 52740 43860 54795
rect 44940 52920 45060 55395
rect 41640 51405 41760 52260
rect 41040 49605 41160 50595
rect 40140 49440 40560 49560
rect 40140 46905 40260 48795
rect 40740 48405 40860 48960
rect 40140 45060 40260 46695
rect 40440 45705 40560 47895
rect 40140 44940 40560 45060
rect 40440 44505 40560 44940
rect 39240 44400 39360 44460
rect 39195 44205 39405 44400
rect 37995 41700 38205 41895
rect 38040 41640 38160 41700
rect 38940 41505 39060 43995
rect 39840 43005 39960 44460
rect 40740 43905 40860 45195
rect 41040 45105 41160 48795
rect 41340 46605 41460 49695
rect 41640 48705 41760 50295
rect 42240 49905 42360 51495
rect 42540 50505 42660 52395
rect 44040 51105 44160 52260
rect 43095 49605 43305 49695
rect 43440 48705 43560 50595
rect 44640 50205 44760 51795
rect 44940 51705 45060 52710
rect 45240 50805 45360 53595
rect 45540 50505 45660 55095
rect 45840 52860 45960 54495
rect 46140 53505 46260 57795
rect 47340 57240 47460 59895
rect 49440 59505 49560 60195
rect 52440 60060 52560 61395
rect 50940 58905 51060 59895
rect 47940 58005 48060 58395
rect 47940 57240 48060 57795
rect 48240 57405 48360 58095
rect 48405 57360 48600 57405
rect 48405 57240 48660 57360
rect 48405 57195 48600 57240
rect 46440 56505 46560 57195
rect 47040 56700 47160 56760
rect 46995 56505 47205 56700
rect 47640 56205 47760 56580
rect 47640 54105 47760 54495
rect 47940 54105 48060 55395
rect 48240 53505 48360 56295
rect 49440 56160 49560 58695
rect 51240 58605 51360 59295
rect 52440 59205 52560 59850
rect 52740 58905 52860 60495
rect 54540 59505 54660 59895
rect 49740 56805 49860 57495
rect 51540 57405 51660 58695
rect 51840 56760 51960 58395
rect 49440 56040 49695 56160
rect 50640 56160 50760 56595
rect 52140 56505 52260 58095
rect 52605 57540 53460 57660
rect 53340 57240 53460 57540
rect 50340 56040 50760 56160
rect 49740 55005 49860 55995
rect 50340 55305 50460 56040
rect 45840 52740 46260 52860
rect 47340 52905 47460 53295
rect 48540 52740 48660 53895
rect 48840 52905 48960 54495
rect 41640 47505 41760 48495
rect 41340 45405 41460 46395
rect 42240 45420 42360 47295
rect 42540 46305 42660 46695
rect 41340 44160 41460 44460
rect 41340 44040 41760 44160
rect 41040 42105 41160 42495
rect 40995 41700 41205 41895
rect 41040 41640 41160 41700
rect 37740 38205 37860 40695
rect 37995 40605 38205 40695
rect 38340 40305 38460 41160
rect 38640 40005 38760 40995
rect 39240 40905 39360 41595
rect 39540 40560 39660 41295
rect 41640 41190 41760 44040
rect 41940 43905 42060 44460
rect 41940 41805 42060 43380
rect 42540 41820 42660 44295
rect 42840 43605 42960 47895
rect 43140 46905 43260 48195
rect 43440 45705 43560 47595
rect 43740 46005 43860 49995
rect 44040 48405 44160 48795
rect 43395 45000 43605 45180
rect 43440 44940 43560 45000
rect 44040 44940 44160 47295
rect 44940 46305 45060 48960
rect 44595 45000 44805 45195
rect 44940 45105 45060 46095
rect 44640 44940 44760 45000
rect 43140 43005 43260 44295
rect 44340 43305 44460 44460
rect 45240 43905 45360 48195
rect 45540 48105 45660 49695
rect 46140 49440 46260 49995
rect 46440 49905 46560 52260
rect 47040 51405 47160 52260
rect 47340 51705 47460 52095
rect 46740 49440 46860 50895
rect 47040 50205 47160 51195
rect 46440 48405 46560 48960
rect 45705 47040 46095 47160
rect 45540 44505 45660 45795
rect 45840 45105 45960 46695
rect 47040 46605 47160 47595
rect 47640 46605 47760 52095
rect 47940 51105 48060 51795
rect 48240 51705 48360 52260
rect 48840 51405 48960 52095
rect 49140 52005 49260 54795
rect 52440 54405 52560 56595
rect 53040 54405 53160 56760
rect 53640 56205 53760 56760
rect 54240 54405 54360 58395
rect 54840 57705 54960 61995
rect 55140 58605 55260 61695
rect 55440 60705 55560 63795
rect 55740 62505 55860 64395
rect 55740 60540 55860 62295
rect 56640 62160 56760 62895
rect 56940 62505 57060 71895
rect 57840 71805 57960 72360
rect 57240 68520 57360 69195
rect 58140 69105 58260 72195
rect 58440 68760 58560 75195
rect 58740 70305 58860 73395
rect 59040 70905 59160 73695
rect 59640 73305 59760 75495
rect 59940 73905 60060 79395
rect 60540 77805 60660 78195
rect 60240 76905 60360 77295
rect 60540 76140 60660 77595
rect 60990 76695 61005 76800
rect 60795 76605 61005 76695
rect 61140 76140 61260 76695
rect 61440 76605 61560 81195
rect 62340 80640 62460 82095
rect 63840 80205 63960 82995
rect 64140 80205 64260 83910
rect 65100 80760 65295 80805
rect 65040 80640 65295 80760
rect 65100 80595 65295 80640
rect 65640 80205 65760 82695
rect 65940 81705 66060 87240
rect 68340 85305 68460 87960
rect 66240 81405 66360 85095
rect 67740 83940 67860 84495
rect 68940 83940 69060 85395
rect 69840 84060 69960 90660
rect 70140 88605 70260 90495
rect 71040 89805 71160 91095
rect 72840 90105 72960 91260
rect 73440 90105 73560 91710
rect 74040 90705 74160 93195
rect 74340 93105 74460 94560
rect 76740 93705 76860 94560
rect 74640 91740 74760 92295
rect 75195 91800 75405 91995
rect 75240 91740 75360 91800
rect 71205 89640 71460 89760
rect 70740 88440 70860 89295
rect 71340 88605 71460 89640
rect 71640 87990 71760 89295
rect 71940 88605 72060 89895
rect 74940 89805 75060 91260
rect 72540 88440 72660 88995
rect 72240 86205 72360 87195
rect 69840 83940 70260 84060
rect 66540 82905 66660 83910
rect 66840 82605 66960 83295
rect 68040 82605 68160 83460
rect 69240 83400 69360 83460
rect 69195 83205 69405 83400
rect 68040 81705 68160 82395
rect 68940 80820 69060 82695
rect 69540 82305 69660 82695
rect 69840 81960 69960 83295
rect 70140 82305 70260 83940
rect 70440 82605 70560 84495
rect 71040 83940 71160 85695
rect 72240 84105 72360 85095
rect 69840 81840 70260 81960
rect 61740 77205 61860 79995
rect 63240 79605 63360 80160
rect 64305 80100 64560 80160
rect 64305 80040 64605 80100
rect 63240 78660 63360 79395
rect 63540 79005 63660 79995
rect 64395 79905 64605 80040
rect 67440 80190 67560 80595
rect 65340 79605 65460 79995
rect 63240 78540 63660 78660
rect 62340 77805 62460 78195
rect 62040 76605 62160 77295
rect 60240 74805 60360 75495
rect 60840 73905 60960 75660
rect 60495 72900 60705 73095
rect 61140 73020 61260 75195
rect 61440 74805 61560 75660
rect 61740 73905 61860 74895
rect 62040 74205 62160 75495
rect 62340 73305 62460 76995
rect 62640 73605 62760 77895
rect 63105 77760 63300 77805
rect 63105 77595 63360 77760
rect 62940 76305 63060 77280
rect 63240 76140 63360 77595
rect 63540 76605 63660 78540
rect 65040 78105 65160 78495
rect 63840 76140 63960 77595
rect 64440 76140 64560 77895
rect 65340 76260 65460 79395
rect 66240 79305 66360 80160
rect 66840 79605 66960 80160
rect 65040 76140 65460 76260
rect 65640 76140 65760 78195
rect 66240 77205 66360 79095
rect 66195 76200 66405 76395
rect 66240 76140 66360 76200
rect 62940 74505 63060 75495
rect 62940 73305 63060 73695
rect 60540 72840 60660 72900
rect 62700 72990 63000 73005
rect 62700 72945 62895 72990
rect 62640 72825 62895 72945
rect 61140 72405 61260 72810
rect 62700 72795 62895 72825
rect 63240 72705 63360 74895
rect 64140 74805 64260 75660
rect 64740 74505 64860 75495
rect 61740 72300 61860 72360
rect 59340 70560 59460 71295
rect 59040 70440 59460 70560
rect 58140 68640 58560 68760
rect 58140 68340 58260 68640
rect 56640 62040 57060 62160
rect 56340 60540 56460 61095
rect 56940 60060 57060 62040
rect 57240 61905 57360 68310
rect 57540 65205 57660 67695
rect 57840 67305 57960 67860
rect 58440 67305 58560 67860
rect 59040 67005 59160 70440
rect 59940 70005 60060 70395
rect 60240 68520 60360 72180
rect 59340 67740 59760 67860
rect 59340 66105 59460 67740
rect 57900 64560 58095 64605
rect 57840 64440 58095 64560
rect 57900 64395 58095 64440
rect 57540 61560 57660 64395
rect 58740 64005 58860 64560
rect 56640 59940 57060 60060
rect 57240 61440 57660 61560
rect 54840 56700 54960 56760
rect 54795 56505 55005 56700
rect 50040 52920 50160 54195
rect 50640 52920 50760 54195
rect 54840 54105 54960 56295
rect 55440 55605 55560 56760
rect 49740 52200 49860 52260
rect 49440 50805 49560 52095
rect 49695 52005 49905 52200
rect 47940 45705 48060 49695
rect 48240 48990 48360 49995
rect 48840 49440 48960 50595
rect 48540 46005 48660 48495
rect 48840 46905 48960 47595
rect 47640 45105 47760 45495
rect 45705 44340 45960 44460
rect 43440 41205 43560 42195
rect 44640 41640 44760 42195
rect 45540 41805 45660 43980
rect 39240 40440 39660 40560
rect 41295 40860 41505 40995
rect 39795 40560 40005 40695
rect 41040 40800 41505 40860
rect 41040 40740 41460 40800
rect 39795 40500 40260 40560
rect 39840 40440 40260 40500
rect 37740 37140 37860 37680
rect 38340 37140 38460 39195
rect 37140 34905 37260 36495
rect 37440 35805 37560 36660
rect 38940 35505 39060 39495
rect 39240 37320 39360 40440
rect 39540 37605 39660 40095
rect 40140 39660 40260 40440
rect 41040 40260 41160 40740
rect 40740 40140 41160 40260
rect 40740 40005 40860 40140
rect 40605 39840 40860 40005
rect 40605 39795 40800 39840
rect 40140 39540 40695 39660
rect 40440 38805 40560 39195
rect 41340 39060 41460 40395
rect 41040 38940 41460 39060
rect 40140 37605 40260 38295
rect 40140 37410 40395 37605
rect 39540 37140 39660 37395
rect 40740 37305 40860 37695
rect 40500 36660 40695 36705
rect 39840 35505 39960 36660
rect 40440 36495 40695 36660
rect 37440 33840 37560 35280
rect 36540 32205 36660 33180
rect 37140 31905 37260 33360
rect 36240 29340 36360 31695
rect 37740 31005 37860 31695
rect 38040 31305 38160 33360
rect 38340 31605 38460 32895
rect 38205 31140 38460 31260
rect 36795 30705 37005 30795
rect 36705 30600 37005 30705
rect 36705 30540 36960 30600
rect 36705 30495 36900 30540
rect 36495 29805 36705 29895
rect 36840 29340 36960 30195
rect 37905 29895 37995 30105
rect 37140 29505 37260 29895
rect 38340 29760 38460 31140
rect 38940 29805 39060 34695
rect 40140 33840 40260 34995
rect 40440 34005 40560 36495
rect 40695 36105 40905 36180
rect 40740 33705 40860 34395
rect 40740 32760 40860 33180
rect 41040 33105 41160 38940
rect 41340 36675 41460 37395
rect 41640 37305 41760 40980
rect 42240 40605 42360 41160
rect 41940 38805 42060 39795
rect 42840 39105 42960 40980
rect 43740 40860 43860 41595
rect 43440 40740 43860 40860
rect 43440 40005 43560 40740
rect 44340 40605 44460 41160
rect 42540 37140 42660 37695
rect 42840 37605 42960 38295
rect 43740 37305 43860 40395
rect 44340 40005 44460 40395
rect 44040 37005 44160 38595
rect 44640 37560 44760 40095
rect 45540 37605 45660 40995
rect 45840 38805 45960 44340
rect 46740 43905 46860 44460
rect 47340 44205 47460 44910
rect 49140 45105 49260 47895
rect 49440 44505 49560 48495
rect 49740 47505 49860 48960
rect 50340 45405 50460 52260
rect 51540 52260 51660 52710
rect 53640 52290 53760 53295
rect 56040 53205 56160 57495
rect 56640 57405 56760 59940
rect 57240 57405 57360 61440
rect 58740 60540 58860 61095
rect 59340 60705 59460 65295
rect 59640 64005 59760 66195
rect 59940 64590 60060 67395
rect 60240 66705 60360 67095
rect 60840 66405 60960 70695
rect 61140 65505 61260 71595
rect 61440 70005 61560 72195
rect 61695 72105 61905 72300
rect 62340 68340 62460 69195
rect 62640 68505 62760 71895
rect 62940 70905 63060 72195
rect 63240 70605 63360 72495
rect 63540 71205 63660 74295
rect 64440 72840 64560 73995
rect 65040 73005 65160 76140
rect 64140 71205 64260 72360
rect 65040 71805 65160 72195
rect 62940 67890 63060 69795
rect 64140 69405 64260 70995
rect 65340 70605 65460 75495
rect 65640 71505 65760 74595
rect 65940 73605 66060 75660
rect 66540 73020 66660 75195
rect 66840 74805 66960 78195
rect 67140 73305 67260 78795
rect 67440 76305 67560 78495
rect 67740 76320 67860 77895
rect 68340 76905 68460 77595
rect 68640 77505 68760 80160
rect 67440 73005 67560 75495
rect 67200 72360 67395 72405
rect 67140 72240 67395 72360
rect 67200 72195 67395 72240
rect 66840 71805 66960 72195
rect 67740 71505 67860 73095
rect 68040 73005 68160 75495
rect 68340 74505 68460 75660
rect 68340 73605 68460 74295
rect 69240 74205 69360 81195
rect 70140 80640 70260 81840
rect 71340 81660 71460 83460
rect 71940 82605 72060 83460
rect 71640 82005 71760 82395
rect 72240 81660 72360 83295
rect 72540 82905 72660 84495
rect 72840 82605 72960 85395
rect 73740 84420 73860 88995
rect 74040 85305 74160 88395
rect 74340 87960 74460 88695
rect 74340 87840 75060 87960
rect 73140 82005 73260 84195
rect 74340 83940 74460 85995
rect 71340 81540 72360 81660
rect 70740 80760 70860 81495
rect 72840 81405 72960 81795
rect 70740 80640 71160 80760
rect 70440 80100 70560 80160
rect 70395 79905 70605 80100
rect 69540 75405 69660 77295
rect 69840 76305 69960 78195
rect 70740 76560 70860 79695
rect 71040 78405 71160 80640
rect 71340 79905 71460 81195
rect 72540 80640 72660 81195
rect 71805 79695 71895 79905
rect 70740 76440 71160 76560
rect 71040 76305 71160 76440
rect 71040 76140 71295 76305
rect 71100 76095 71295 76140
rect 69840 73860 69960 75495
rect 70140 74805 70260 75660
rect 71640 75405 71760 77595
rect 72240 76605 72360 80160
rect 73140 79605 73260 80610
rect 73440 79005 73560 83295
rect 73740 78105 73860 82095
rect 74640 81960 74760 83460
rect 75240 82605 75360 87795
rect 76140 85305 76260 93495
rect 76440 87705 76560 90795
rect 76740 90705 76860 91080
rect 77340 90405 77460 91260
rect 77595 91005 77805 91095
rect 77940 91005 78060 93795
rect 78240 91305 78360 91995
rect 79140 91740 79260 92295
rect 78840 91200 78960 91260
rect 78795 91005 79005 91200
rect 78240 90105 78360 90495
rect 76740 88605 76860 89295
rect 78240 88605 78360 89895
rect 78840 88440 78960 88995
rect 79440 88605 79560 91095
rect 77640 87840 78060 87960
rect 75795 84000 76005 84195
rect 75840 83940 75960 84000
rect 76440 83940 76560 86295
rect 76740 84705 76860 86595
rect 77340 86205 77460 86595
rect 77040 83940 77160 85395
rect 77340 84105 77460 84795
rect 74640 81840 75060 81960
rect 74940 80805 75060 81840
rect 75195 81060 75405 81195
rect 75540 81060 75660 82695
rect 75195 81000 75660 81060
rect 75240 80940 75660 81000
rect 75240 80640 75360 80940
rect 74640 80100 74760 80160
rect 74595 79905 74805 80100
rect 75540 80040 75960 80160
rect 74640 78405 74760 78795
rect 74940 77505 75060 79995
rect 72540 76140 72660 76695
rect 70995 75060 71205 75195
rect 70740 75000 71205 75060
rect 70740 74940 71160 75000
rect 70740 74760 70860 74940
rect 70440 74640 70860 74760
rect 69840 73740 70260 73860
rect 69540 73305 69660 73695
rect 68040 71505 68160 72195
rect 65040 69705 65160 70095
rect 64740 68340 65460 68460
rect 62040 67800 62160 67860
rect 61995 67605 62205 67800
rect 62190 67500 62205 67605
rect 62340 65040 62460 67395
rect 64440 67305 64560 68310
rect 64740 67305 64860 68340
rect 60240 61305 60360 62295
rect 61140 61905 61260 64560
rect 57540 60105 57660 60510
rect 57540 57240 57660 58995
rect 57840 57405 57960 59595
rect 58440 58905 58560 60060
rect 59040 58905 59160 60060
rect 56340 56205 56460 57195
rect 56940 56460 57060 56580
rect 56640 56340 57060 56460
rect 55440 52290 55560 52995
rect 56640 52905 56760 56340
rect 57840 55860 57960 56595
rect 57540 55740 57960 55860
rect 51540 52140 51960 52260
rect 50640 49605 50760 51795
rect 50940 50205 51060 52095
rect 51540 49905 51660 51195
rect 51840 49440 51960 52140
rect 52140 49605 52260 50895
rect 52440 48990 52560 49695
rect 50640 48105 50760 48795
rect 50940 47505 51060 48960
rect 52740 48405 52860 52260
rect 53640 51705 53760 52080
rect 56040 51705 56160 52260
rect 53295 49500 53505 49695
rect 53340 49440 53460 49500
rect 54240 49005 54360 49695
rect 55395 49500 55605 49695
rect 55995 49500 56205 49695
rect 55440 49440 55560 49500
rect 56040 49440 56160 49500
rect 56640 48990 56760 52095
rect 56940 50205 57060 52695
rect 57240 49560 57360 52695
rect 57540 51405 57660 55740
rect 58140 53205 58260 57795
rect 59640 57405 59760 61095
rect 60240 60540 60360 61095
rect 60795 60600 61005 60795
rect 61095 60705 61305 60795
rect 60840 60540 60960 60600
rect 61440 59805 61560 63795
rect 62040 63105 62160 64395
rect 59940 57105 60060 59595
rect 61140 57240 61260 57795
rect 61740 57705 61860 61095
rect 62040 60705 62160 62895
rect 62640 61905 62760 64560
rect 62940 62805 63060 64395
rect 63240 61005 63360 67095
rect 65640 66705 65760 67680
rect 63540 62505 63660 66195
rect 64440 65040 64560 65595
rect 63840 63705 63960 64560
rect 64740 61905 64860 64260
rect 62295 60600 62505 60795
rect 62340 60540 62460 60600
rect 63540 60705 63660 61695
rect 64500 60960 64695 61005
rect 64440 60795 64695 60960
rect 64440 60540 64560 60795
rect 62040 57360 62160 59895
rect 62640 58605 62760 60060
rect 63840 60060 63960 60510
rect 65340 60090 65460 61395
rect 63540 59940 63960 60060
rect 63240 58905 63360 59880
rect 61740 57240 62160 57360
rect 58440 55305 58560 56595
rect 58740 54960 58860 56760
rect 60240 56760 60360 57240
rect 63240 56805 63360 58380
rect 60240 56640 60660 56760
rect 59340 56460 59460 56580
rect 58440 54840 58860 54960
rect 59040 56340 59460 56460
rect 58440 54705 58560 54840
rect 58440 52860 58560 54495
rect 59040 52905 59160 56340
rect 59940 55560 60060 56580
rect 59940 55440 60195 55560
rect 58140 52740 58560 52860
rect 60240 52605 60360 55395
rect 58740 51105 58860 52260
rect 60540 52005 60660 56640
rect 60840 55305 60960 56760
rect 61440 55905 61560 56760
rect 61095 52800 61305 52995
rect 62340 52860 62460 54795
rect 61140 52740 61260 52800
rect 62040 52740 62460 52860
rect 56940 49440 57360 49560
rect 46140 37905 46260 43695
rect 47640 43605 47760 44295
rect 47595 42300 47805 42495
rect 47640 42240 47760 42300
rect 48540 41385 48660 43995
rect 46440 40005 46560 41295
rect 48495 41190 48705 41295
rect 48840 40260 48960 41295
rect 49140 40305 49260 44295
rect 49440 41805 49560 43395
rect 49740 42105 49860 45195
rect 50340 43005 50460 44460
rect 50940 43005 51060 44460
rect 50940 41805 51060 42795
rect 48540 40140 48960 40260
rect 46305 37740 46560 37860
rect 44340 37440 44760 37560
rect 42195 36405 42405 36495
rect 42840 35805 42960 36660
rect 43695 36405 43905 36495
rect 42540 34905 42660 35295
rect 42240 33840 42360 34395
rect 44040 34020 44160 36795
rect 41505 33360 41700 33405
rect 41505 33240 41760 33360
rect 41505 33195 41700 33240
rect 40740 32640 41160 32760
rect 37695 29520 37905 29580
rect 37440 29340 37695 29460
rect 37440 28890 37560 29340
rect 38040 29640 38460 29760
rect 38040 29340 38160 29640
rect 35940 28800 36060 28860
rect 35895 28605 36105 28800
rect 38340 28005 38460 28860
rect 35640 25590 35760 27495
rect 35940 26505 36060 27195
rect 36240 26805 36360 27195
rect 36240 26040 36360 26595
rect 36840 26040 36960 27795
rect 36540 25260 36660 25560
rect 36540 25140 36960 25260
rect 35205 23340 35460 23460
rect 32640 18600 33060 18660
rect 32595 18540 33060 18600
rect 32595 18405 32805 18540
rect 32790 18300 32805 18405
rect 33495 18300 33705 18495
rect 34140 18405 34260 20295
rect 34740 19605 34860 20295
rect 35040 18960 35160 23295
rect 36240 21540 36360 22995
rect 36540 22305 36660 22695
rect 34740 18840 35160 18960
rect 33540 18240 33660 18300
rect 34440 17790 34560 18195
rect 31140 17700 31260 17760
rect 30540 16305 30660 17595
rect 31095 17505 31305 17700
rect 29040 13740 29160 13800
rect 29940 13290 30060 14295
rect 30540 13920 30660 16095
rect 31140 13740 31260 14895
rect 31440 14160 31560 15495
rect 31905 14295 31995 14505
rect 31440 14040 31860 14160
rect 31740 13740 31860 14040
rect 29340 11805 29460 12195
rect 29190 11595 29205 11700
rect 28995 11460 29205 11595
rect 28995 11400 29460 11460
rect 29040 11340 29460 11400
rect 27495 10500 27705 10695
rect 27540 10440 27660 10500
rect 23040 9900 23160 9960
rect 22995 9705 23205 9900
rect 22440 9105 22560 9495
rect 24540 9405 24660 9960
rect 25095 9705 25305 9780
rect 26340 9705 26460 10395
rect 26595 9705 26805 9795
rect 20940 5205 21060 6195
rect 22140 4005 22260 4860
rect 18840 2100 18960 2160
rect 18795 1905 19005 2100
rect 14640 1740 14895 1905
rect 14700 1695 14895 1740
rect 18600 1590 18900 1605
rect 18195 1260 18405 1395
rect 18705 1395 18795 1590
rect 19140 1260 19260 1695
rect 18195 1200 19260 1260
rect 18240 1140 19260 1200
rect 20040 705 20160 2610
rect 22140 2190 22260 2595
rect 20640 2100 20760 2160
rect 20595 1905 20805 2100
rect 22440 1305 22560 4395
rect 22740 2190 22860 3495
rect 23040 2805 23160 4095
rect 23640 2640 23760 6495
rect 24240 6105 24360 8295
rect 24840 6120 24960 8595
rect 27240 8205 27360 9960
rect 24105 5940 24360 6105
rect 24105 5895 24300 5940
rect 24240 2805 24360 3495
rect 24540 3405 24660 5460
rect 25440 5205 25560 7395
rect 27840 7305 27960 9780
rect 28440 8805 28560 10695
rect 28740 10605 28860 11295
rect 29340 10440 29460 11340
rect 29940 10440 30060 10995
rect 30240 10560 30360 13695
rect 32340 13290 32460 14595
rect 32595 14505 32805 14595
rect 30840 13200 30960 13260
rect 30795 13005 31005 13200
rect 31140 10605 31260 11895
rect 30240 10440 30660 10560
rect 29640 9105 29760 9960
rect 30240 8205 30360 9795
rect 30540 8505 30660 10440
rect 32340 10440 32460 11895
rect 32940 11805 33060 14895
rect 34440 13905 34560 17580
rect 34740 17505 34860 18840
rect 35940 18705 36060 21060
rect 35040 16605 35160 18495
rect 36240 18240 36360 20595
rect 36840 18660 36960 25140
rect 37140 22005 37260 25395
rect 37440 25005 37560 26895
rect 39240 25590 39360 32295
rect 39540 27105 39660 32595
rect 40140 29520 40260 31395
rect 40740 29340 40860 30195
rect 41040 29505 41160 32640
rect 41340 29205 41460 31095
rect 41640 28860 41760 32895
rect 44340 32205 44460 37440
rect 45705 37440 45960 37560
rect 45840 37140 45960 37440
rect 46440 37305 46560 37740
rect 44640 36105 44760 37095
rect 45540 36600 45660 36660
rect 44640 32505 44760 35295
rect 44940 34905 45060 36495
rect 45495 36405 45705 36600
rect 45540 33840 45660 34695
rect 46140 34020 46260 36165
rect 46740 35505 46860 38895
rect 47205 36660 47400 36705
rect 47205 36540 47460 36660
rect 47205 36495 47400 36540
rect 47040 33840 47160 35595
rect 48240 34005 48360 38595
rect 44940 33405 45060 33810
rect 48000 33360 48195 33405
rect 45840 33300 45960 33360
rect 47340 33300 47460 33360
rect 45795 33105 46005 33300
rect 47295 33105 47505 33300
rect 47940 33240 48195 33360
rect 48000 33195 48195 33240
rect 42105 29460 42300 29505
rect 42105 29340 42360 29460
rect 42795 29400 43005 29595
rect 42840 29340 42960 29400
rect 42105 29295 42300 29340
rect 46740 29340 47460 29460
rect 39540 25605 39660 26295
rect 39840 26205 39960 28695
rect 40440 27105 40560 28860
rect 41340 28740 41760 28860
rect 40740 26805 40860 27495
rect 41340 27405 41460 28740
rect 37440 22005 37560 24795
rect 38640 24705 38760 25560
rect 39240 24705 39360 25380
rect 41640 25305 41760 28395
rect 41940 27105 42060 28695
rect 42540 28005 42660 28860
rect 43140 28800 43260 28860
rect 43095 28605 43305 28800
rect 43740 28605 43860 29310
rect 44790 28365 44805 28500
rect 44595 28305 44805 28365
rect 42840 26040 42960 26595
rect 38595 21600 38805 21795
rect 39495 21600 39705 21795
rect 40140 21720 40260 24795
rect 38640 21540 38760 21600
rect 39540 21540 39660 21600
rect 37140 19005 37260 21480
rect 37740 18705 37860 20295
rect 36840 18540 37260 18660
rect 34140 13740 34395 13860
rect 35040 13740 35160 16080
rect 35340 15705 35460 17595
rect 37140 17760 37260 18540
rect 37695 18300 37905 18495
rect 37740 18240 37860 18300
rect 39240 17760 39360 20295
rect 39840 19605 39960 21060
rect 41040 20505 41160 25065
rect 42240 24705 42360 25380
rect 43140 23205 43260 25560
rect 42495 21600 42705 21795
rect 42540 21540 42660 21600
rect 41340 20805 41460 21510
rect 41100 20160 41295 20205
rect 41040 19995 41295 20160
rect 40140 18240 40260 19695
rect 40695 18300 40905 18495
rect 41040 18405 41160 19995
rect 41940 19605 42060 20595
rect 42240 20205 42360 21060
rect 42840 20205 42960 21060
rect 40740 18240 40860 18300
rect 36840 17640 37260 17760
rect 38040 17700 38160 17760
rect 38640 17700 38760 17760
rect 35640 16005 35760 16395
rect 36840 15405 36960 17640
rect 37995 17505 38205 17700
rect 38595 17505 38805 17700
rect 38940 17640 39360 17760
rect 33840 12405 33960 13260
rect 33840 11205 33960 12195
rect 25140 3705 25260 4395
rect 25740 4305 25860 6795
rect 27240 5940 27360 6795
rect 29640 5940 29760 6495
rect 26040 5205 26160 5910
rect 26940 5400 27060 5460
rect 26895 5205 27105 5400
rect 29940 4905 30060 5460
rect 30540 5205 30660 7695
rect 30840 6120 30960 10395
rect 31440 9900 31560 9960
rect 31395 9705 31605 9900
rect 32040 9105 32160 9960
rect 31695 6000 31905 6195
rect 32640 6060 32760 9795
rect 32940 9705 33060 10995
rect 33240 9990 33360 10695
rect 33705 10560 33900 10605
rect 33705 10440 33960 10560
rect 34440 10440 34560 10995
rect 33705 10395 33900 10440
rect 34140 6405 34260 8295
rect 35340 8205 35460 10995
rect 35640 10605 35760 11295
rect 35940 10440 36060 11895
rect 36540 11760 36660 13695
rect 36840 13305 36960 14295
rect 37740 13740 37860 15795
rect 37995 14205 38205 14295
rect 38340 13920 38460 14595
rect 36240 11640 36660 11760
rect 36240 10905 36360 11640
rect 36540 10440 36660 10995
rect 37140 10605 37260 12195
rect 36240 9405 36360 9960
rect 37440 9405 37560 13260
rect 38940 13005 39060 17640
rect 39540 16005 39660 18195
rect 39495 13800 39705 13995
rect 39540 13740 39660 13800
rect 40140 13740 40260 15795
rect 40440 14805 40560 17760
rect 41340 17505 41460 19395
rect 41340 13290 41460 17295
rect 41640 13860 41760 19095
rect 43140 18960 43260 20895
rect 43440 20805 43560 25380
rect 43740 24105 43860 27495
rect 44940 26805 45060 28395
rect 45240 27705 45360 29310
rect 47340 28905 47460 29340
rect 45840 28605 45960 28860
rect 45705 28440 45960 28605
rect 45705 28395 45900 28440
rect 44940 26040 45060 26595
rect 44040 24705 44160 25995
rect 44640 23505 44760 25560
rect 43905 21660 44100 21705
rect 43905 21540 44160 21660
rect 44595 21600 44805 21795
rect 45540 21705 45660 27795
rect 46140 26040 46260 26895
rect 46440 26505 46560 28860
rect 46740 26805 46860 28095
rect 46740 26040 46860 26595
rect 47340 25005 47460 28095
rect 46140 22005 46260 24195
rect 44640 21540 44760 21600
rect 43905 21495 44100 21540
rect 46095 21600 46305 21795
rect 46140 21540 46260 21600
rect 47640 21705 47760 32595
rect 48240 31605 48360 33195
rect 48540 32805 48660 40140
rect 49140 38205 49260 40095
rect 49440 39105 49560 40995
rect 49740 40905 49860 41160
rect 49740 39705 49860 40695
rect 49740 38160 49860 38595
rect 50040 38505 50160 40995
rect 50640 39705 50760 41160
rect 49740 38040 50160 38160
rect 49395 37200 49605 37395
rect 50040 37320 50160 38040
rect 49440 37140 49560 37200
rect 50340 37305 50460 37995
rect 49740 36600 49860 36660
rect 49695 36405 49905 36600
rect 50640 34905 50760 38895
rect 50940 37320 51060 40995
rect 51240 38205 51360 41895
rect 51540 41805 51660 47895
rect 51840 44490 51960 45495
rect 53040 44940 53160 45795
rect 53940 44490 54060 46395
rect 54840 44940 54960 48495
rect 55740 46905 55860 48960
rect 56940 46605 57060 49440
rect 58140 49440 58260 49995
rect 59040 48990 59160 49695
rect 59940 49440 60060 50295
rect 60840 49605 60960 51195
rect 59640 48900 59760 48960
rect 59595 48705 59805 48900
rect 58095 48360 58305 48495
rect 57705 48300 58305 48360
rect 59895 48405 60105 48495
rect 57705 48240 58260 48300
rect 57540 47205 57660 47595
rect 57240 45120 57360 46095
rect 51840 41640 51960 42795
rect 52140 41100 52260 41160
rect 52095 40905 52305 41100
rect 53340 37605 53460 44460
rect 53640 39105 53760 43995
rect 55140 43005 55260 44460
rect 56040 44340 56295 44460
rect 56040 43605 56160 44340
rect 57240 43305 57360 44910
rect 57540 44460 57660 46995
rect 60840 46905 60960 48795
rect 61140 47805 61260 51795
rect 62640 49905 62760 53595
rect 63240 50805 63360 56280
rect 63540 55905 63660 59940
rect 63840 57405 63960 59595
rect 65040 56640 65460 56760
rect 63540 52905 63660 55695
rect 65340 55005 65460 56640
rect 63840 52740 63960 54195
rect 65040 52260 65160 54495
rect 65640 53805 65760 61095
rect 65940 60705 66060 65295
rect 66240 61305 66360 71295
rect 67140 69105 67260 71295
rect 67440 70005 67560 70695
rect 66840 68520 66960 68895
rect 67440 68340 67560 69795
rect 67740 68805 67860 70695
rect 68040 69405 68160 71295
rect 67140 66405 67260 67860
rect 67740 67740 68160 67860
rect 66840 65205 66960 65895
rect 66705 65040 66960 65205
rect 67440 65040 67560 66795
rect 67740 65805 67860 66495
rect 68040 65805 68160 67740
rect 68340 65505 68460 71895
rect 68640 71805 68760 72360
rect 69240 70305 69360 72360
rect 69540 70905 69660 72195
rect 69840 71505 69960 73395
rect 70140 73005 70260 73740
rect 70440 73305 70560 74640
rect 70740 73305 70860 74295
rect 71040 74205 71160 74595
rect 71640 74205 71760 75195
rect 70740 73110 70995 73305
rect 71940 73005 72060 75495
rect 72840 75105 72960 75660
rect 71940 72840 72195 73005
rect 72000 72795 72195 72840
rect 70140 71805 70260 72480
rect 71040 72060 71160 72360
rect 70740 71940 71160 72060
rect 68640 68505 68760 68895
rect 69240 68340 69360 69780
rect 69795 69405 70005 69495
rect 69540 68805 69660 69195
rect 69900 68460 70095 68505
rect 69840 68340 70095 68460
rect 69900 68295 70095 68340
rect 68805 67860 69000 67905
rect 68805 67740 69060 67860
rect 68805 67695 69000 67740
rect 66705 64995 66900 65040
rect 68340 64605 68460 64980
rect 68640 64605 68760 67095
rect 68940 66705 69060 67395
rect 69240 66405 69360 67095
rect 69540 66705 69660 67860
rect 70440 67890 70560 70695
rect 70740 70605 70860 71940
rect 71040 69405 71160 70395
rect 72240 70305 72360 72195
rect 72540 69360 72660 74595
rect 72795 72960 73005 73095
rect 73740 73005 73860 76395
rect 74040 73605 74160 77295
rect 74895 76560 75105 76695
rect 74640 76500 75105 76560
rect 74640 76440 75060 76500
rect 74640 76140 74760 76440
rect 75240 76140 75360 79695
rect 75540 77805 75660 79395
rect 75840 79005 75960 80040
rect 76140 79305 76260 81795
rect 77040 80805 77160 82995
rect 77340 81705 77460 82395
rect 77340 80640 77460 81495
rect 77640 80805 77760 87495
rect 77940 87405 78060 87840
rect 79440 87405 79560 87795
rect 77940 86505 78060 87195
rect 77940 83205 78060 85095
rect 78540 84405 78660 85695
rect 78840 83940 78960 85395
rect 79140 84105 79260 84795
rect 79440 84705 79560 85995
rect 79740 85605 79860 88410
rect 79740 83805 79860 85395
rect 78405 83340 78660 83460
rect 77940 82305 78060 82680
rect 72795 72900 73260 72960
rect 72840 72840 73260 72900
rect 73140 70305 73260 71595
rect 73440 71505 73560 72180
rect 72240 69300 72660 69360
rect 72195 69240 72660 69300
rect 72195 69105 72405 69240
rect 68895 65505 69105 65595
rect 69240 65160 69360 66195
rect 69540 66105 69660 66495
rect 69840 66405 69960 67395
rect 70140 67305 70260 67695
rect 70440 65505 70560 67680
rect 70095 65220 70305 65295
rect 68940 65040 69360 65160
rect 67140 63705 67260 64560
rect 67740 64500 67860 64560
rect 67695 64305 67905 64500
rect 68940 64305 69060 65040
rect 70740 65205 70860 68595
rect 71040 68205 71160 68880
rect 71040 66405 71160 67995
rect 71940 67140 72360 67260
rect 69840 64500 69960 64560
rect 66195 60600 66405 60780
rect 66240 60540 66360 60600
rect 66840 60540 66960 61695
rect 67740 60060 67860 63195
rect 68340 60540 68460 61695
rect 69240 60705 69360 64395
rect 69795 64305 70005 64500
rect 69540 62205 69660 64095
rect 65940 56505 66060 59895
rect 66240 57420 66360 58995
rect 66540 58605 66660 60060
rect 67140 60000 67560 60060
rect 67140 59940 67605 60000
rect 67740 59940 68160 60060
rect 67395 59805 67605 59940
rect 66240 55905 66360 57210
rect 68040 56760 68160 59940
rect 68505 59700 69060 59760
rect 68505 59640 69105 59700
rect 68895 59505 69105 59640
rect 68340 57405 68460 59280
rect 69240 58305 69360 59895
rect 69540 59805 69660 61680
rect 69840 61605 69960 64095
rect 70140 61905 70260 64095
rect 71040 62505 71160 65880
rect 71340 64305 71460 66795
rect 71640 66105 71760 67095
rect 71940 65760 72060 67140
rect 72240 65805 72360 66795
rect 71640 65700 72060 65760
rect 71595 65640 72060 65700
rect 71595 65505 71805 65640
rect 73440 65220 73560 68595
rect 74040 68340 74160 72795
rect 74340 68805 74460 74595
rect 74940 73020 75060 73995
rect 75540 73905 75660 75495
rect 75840 75405 75960 78195
rect 76140 73005 76260 77895
rect 76440 76305 76560 79995
rect 76740 77505 76860 80160
rect 77040 76560 77160 78495
rect 77940 76905 78060 80895
rect 78240 80805 78360 83280
rect 78705 83160 78900 83205
rect 78705 82995 78960 83160
rect 78540 81105 78660 81795
rect 78840 81405 78960 82995
rect 78495 80700 78705 80895
rect 79095 80700 79305 80895
rect 78540 80640 78660 80700
rect 79140 80640 79260 80700
rect 77805 76740 78060 76905
rect 77805 76695 78000 76740
rect 76905 76440 77160 76560
rect 76740 76140 76860 76395
rect 77295 76200 77505 76395
rect 77895 76305 78105 76395
rect 77340 76140 77460 76200
rect 74640 69105 74760 72195
rect 74940 68760 75060 71895
rect 75240 70905 75360 72360
rect 75840 72300 75960 72360
rect 75795 72105 76005 72300
rect 76140 69960 76260 72195
rect 75840 69840 76260 69960
rect 75840 68805 75960 69840
rect 74640 68640 75060 68760
rect 74640 68340 74760 68640
rect 76140 68505 76260 69495
rect 76440 69405 76560 75495
rect 77040 74505 77160 75660
rect 76740 72390 76860 73695
rect 77340 73005 77460 75195
rect 77640 73305 77760 75480
rect 78240 74805 78360 79095
rect 79740 78405 79860 82395
rect 80040 82005 80160 92895
rect 83895 92205 84105 92295
rect 82305 92040 82695 92160
rect 81495 91800 81705 91995
rect 81540 91740 81660 91800
rect 83295 91800 83505 91995
rect 83895 91905 84105 91995
rect 83340 91740 83460 91800
rect 80640 90105 80760 91095
rect 81240 90705 81360 91260
rect 82140 90405 82260 91095
rect 81240 88440 81360 89895
rect 81540 87900 81660 87960
rect 81495 87705 81705 87900
rect 82140 87405 82260 88410
rect 81840 85605 81960 86595
rect 82140 85905 82260 87195
rect 82440 83805 82560 88995
rect 83040 88620 83160 89295
rect 82740 86505 82860 87495
rect 84240 85560 84360 92595
rect 84540 88605 84660 92295
rect 84840 90705 84960 93495
rect 87240 92205 87360 94560
rect 87840 94005 87960 94560
rect 88735 94440 88860 94560
rect 85395 91800 85605 91995
rect 85440 91740 85560 91800
rect 87540 91740 87660 92595
rect 86340 91200 86460 91260
rect 86295 91005 86505 91200
rect 86040 89805 86160 90495
rect 86940 90105 87060 91395
rect 84840 88440 84960 89295
rect 85440 88440 85560 88995
rect 84540 85860 84660 87795
rect 85140 87105 85260 87780
rect 84540 85740 84960 85860
rect 84240 85440 84660 85560
rect 81240 82800 81360 82860
rect 81195 82605 81405 82800
rect 80040 80205 80160 81195
rect 80340 80805 80460 81195
rect 80895 80700 81105 80895
rect 81540 80820 81660 82695
rect 82440 82560 82560 83280
rect 82740 83205 82860 83895
rect 82440 82440 82860 82560
rect 80940 80640 81060 80700
rect 82440 80640 82560 81795
rect 82740 81060 82860 82440
rect 83040 81405 83160 85395
rect 84240 84105 84360 85095
rect 82740 80940 83160 81060
rect 83040 80640 83160 80940
rect 83640 80805 83760 82995
rect 81240 79305 81360 79980
rect 81240 78705 81360 79095
rect 78840 76320 78960 77895
rect 80640 77805 80760 78195
rect 80940 76305 81060 77595
rect 79140 75360 79260 75660
rect 79005 75240 79260 75360
rect 78495 72900 78705 73095
rect 78840 73005 78960 75195
rect 79740 75105 79860 75660
rect 80040 74805 80160 75495
rect 80340 74505 80460 76110
rect 80640 74805 80760 76110
rect 81840 76305 81960 77295
rect 79995 73305 80205 73395
rect 78540 72840 78660 72900
rect 76695 72105 76905 72180
rect 77040 71805 77160 72795
rect 77340 69705 77460 72195
rect 78240 71205 78360 72360
rect 79140 72390 79260 73095
rect 80040 72840 80160 73095
rect 80640 72840 80760 73995
rect 81240 72390 81360 74895
rect 77640 70005 77760 70995
rect 78240 69705 78360 70395
rect 73740 66705 73860 67695
rect 74940 67800 75060 67860
rect 74895 67605 75105 67800
rect 73740 65040 73860 65895
rect 71340 60090 71460 60495
rect 69840 59940 70260 60060
rect 66840 56700 66960 56760
rect 66795 56505 67005 56700
rect 67740 56640 68160 56760
rect 58140 44940 58260 45495
rect 57540 44340 57960 44460
rect 51105 36660 51300 36705
rect 51105 36540 51360 36660
rect 51105 36495 51300 36540
rect 49140 33105 49260 33795
rect 48240 29340 48360 30195
rect 48840 29520 48960 32295
rect 49740 31905 49860 33360
rect 50940 31005 51060 33810
rect 51240 30105 51360 34095
rect 52140 34005 52260 36495
rect 52440 34305 52560 37395
rect 54240 37140 54360 40095
rect 54540 39705 54660 41160
rect 52740 36405 52860 36795
rect 53340 36105 53460 36660
rect 52740 33960 52860 34695
rect 52440 33840 52860 33960
rect 51840 31305 51960 33360
rect 51840 30360 51960 31095
rect 51840 30240 52260 30360
rect 50340 29520 50460 29895
rect 50640 29340 50760 29895
rect 47940 22005 48060 28680
rect 49440 28605 49560 29310
rect 49440 28005 49560 28395
rect 50940 27405 51060 28860
rect 48840 26220 48960 26595
rect 50040 25605 50160 26895
rect 51840 26205 51960 29895
rect 48540 24405 48660 25560
rect 52140 25590 52260 30240
rect 52740 30105 52860 33195
rect 53040 33105 53160 34395
rect 53940 34305 54060 36660
rect 54840 35205 54960 37395
rect 55140 36705 55260 41160
rect 55440 39705 55560 40980
rect 55740 37260 55860 41595
rect 56040 37620 56160 42795
rect 56340 40305 56460 42195
rect 56640 41805 56760 43095
rect 56340 38205 56460 38895
rect 55440 37140 55860 37260
rect 55440 35160 55560 37140
rect 56640 37140 56760 38295
rect 57540 37305 57660 40980
rect 57840 40605 57960 44340
rect 59040 41640 59160 42195
rect 59640 42105 59760 44940
rect 59940 44505 60060 45795
rect 60240 45105 60360 46395
rect 61440 45105 61560 49695
rect 64440 49620 64560 52260
rect 65040 52140 65460 52260
rect 65340 49605 65460 52140
rect 66240 52200 66360 52260
rect 61740 48405 61860 48780
rect 59940 41760 60060 43395
rect 59640 41640 60060 41760
rect 58140 41205 58260 41610
rect 57540 35205 57660 37095
rect 55440 35040 55860 35160
rect 53340 30705 53460 34095
rect 54240 34020 54360 34995
rect 53640 31605 53760 32895
rect 53940 32805 54060 33360
rect 55740 32505 55860 35040
rect 52740 29340 52860 29895
rect 53295 29400 53505 29595
rect 53340 29340 53460 29400
rect 53940 29340 54060 31095
rect 54540 28890 54660 29595
rect 53040 28305 53160 28680
rect 53640 28005 53760 28860
rect 53805 27840 54060 27960
rect 52395 26220 52605 26295
rect 53595 26205 53805 26295
rect 48840 22605 48960 23895
rect 43005 18840 43260 18960
rect 42840 18240 42960 18795
rect 43740 18420 43860 20895
rect 45105 20940 45360 21060
rect 44340 18240 44460 19995
rect 43740 17790 43860 18210
rect 42540 17700 42660 17760
rect 41940 15405 42060 17595
rect 42495 17505 42705 17700
rect 45240 17505 45360 20940
rect 46440 20505 46560 21060
rect 45540 18405 45660 18795
rect 46440 18705 46560 19395
rect 47040 18360 47160 20295
rect 47340 20205 47460 21510
rect 47895 21600 48105 21795
rect 47940 21540 48060 21600
rect 49140 21705 49260 22695
rect 49440 21105 49560 21795
rect 50040 21705 50160 25080
rect 51240 23505 51360 25395
rect 51540 24660 51660 25560
rect 53940 25590 54060 27840
rect 54840 27105 54960 30495
rect 56040 29460 56160 34995
rect 57840 34005 57960 39795
rect 59040 38160 59160 40395
rect 59340 38505 59460 41160
rect 59940 40005 60060 40995
rect 60240 38205 60360 44295
rect 61440 43305 61560 44295
rect 61740 43605 61860 47295
rect 62040 46305 62160 48960
rect 62040 44805 62160 45495
rect 62340 44205 62460 48195
rect 63240 46605 63360 47595
rect 62640 45060 62760 45795
rect 63540 45705 63660 49395
rect 63840 49005 63960 49410
rect 65040 48900 65160 48960
rect 64740 46305 64860 48795
rect 64995 48705 65205 48900
rect 65340 47205 65460 48795
rect 65640 48405 65760 49695
rect 65940 48705 66060 52095
rect 66195 52005 66405 52200
rect 66240 51105 66360 51795
rect 66540 51705 66660 52095
rect 66240 49005 66360 49995
rect 66840 49905 66960 55695
rect 67440 54705 67560 55995
rect 67740 54105 67860 56640
rect 69540 55905 69660 59280
rect 69840 59205 69960 59940
rect 69840 56205 69960 58995
rect 68040 53505 68160 54495
rect 67140 52905 67260 53295
rect 68040 52740 68160 53295
rect 68340 52905 68460 55695
rect 67140 50205 67260 52095
rect 67740 51105 67860 52260
rect 68340 52140 68760 52260
rect 66840 48900 66960 48960
rect 66795 48705 67005 48900
rect 66105 48690 66300 48705
rect 66105 48495 66195 48690
rect 65940 46005 66060 48180
rect 62640 44940 63060 45060
rect 64140 45105 64260 45495
rect 60540 40605 60660 42495
rect 61440 41805 61560 43095
rect 62640 43005 62760 44295
rect 63840 44400 63960 44460
rect 63795 44205 64005 44400
rect 64140 43305 64260 44295
rect 64440 43905 64560 45795
rect 66240 45405 66360 46695
rect 66540 45105 66660 48495
rect 67440 46905 67560 48960
rect 63840 42405 63960 42795
rect 61695 41700 61905 41895
rect 61740 41640 61860 41700
rect 64140 41805 64260 43095
rect 64740 42660 64860 44295
rect 65040 43905 65160 44460
rect 65640 43905 65760 44460
rect 66195 44160 66405 44295
rect 65940 44100 66405 44160
rect 66540 44340 66795 44460
rect 65940 44040 66360 44100
rect 64440 42540 64860 42660
rect 59040 38040 59460 38160
rect 58740 36105 58860 36660
rect 59340 35805 59460 38040
rect 60240 37560 60360 37995
rect 59940 37440 60360 37560
rect 59940 37140 60060 37440
rect 60495 37200 60705 37395
rect 61140 37305 61260 38595
rect 60540 37140 60660 37200
rect 60840 36600 60960 36660
rect 60795 36405 61005 36600
rect 58140 34005 58260 34395
rect 58995 33900 59205 34095
rect 59040 33840 59160 33900
rect 60240 34005 60360 35595
rect 56640 32205 56760 33360
rect 58140 32505 58260 33480
rect 58440 32160 58560 33195
rect 58740 32805 58860 33360
rect 59040 32505 59160 32895
rect 60240 32805 60360 33195
rect 58005 32040 58560 32160
rect 58740 29805 58860 31695
rect 56040 29340 56460 29460
rect 55740 27705 55860 28680
rect 51540 24540 51960 24660
rect 51495 22905 51705 22995
rect 47040 18240 47460 18360
rect 45705 17760 45900 17805
rect 45705 17640 45960 17760
rect 45705 17595 45900 17640
rect 41640 13740 42060 13860
rect 42540 13740 42660 14595
rect 43440 14505 43560 15495
rect 47040 15105 47160 17595
rect 47340 15705 47460 18240
rect 38340 10440 38460 11295
rect 38640 8205 38760 9960
rect 35340 7305 35460 7995
rect 33195 6105 33405 6195
rect 31740 5940 31860 6000
rect 32340 5940 33060 6060
rect 32940 5490 33060 5940
rect 34095 6000 34305 6195
rect 34140 5940 34260 6000
rect 35640 5505 35760 6495
rect 36840 5940 36960 6495
rect 39240 5505 39360 6495
rect 32790 5280 32805 5400
rect 32595 5205 32805 5280
rect 29940 4740 30195 4905
rect 30000 4695 30195 4740
rect 31005 4695 31095 4905
rect 26505 4395 26595 4605
rect 23940 1605 24060 2160
rect 24840 1605 24960 2895
rect 25440 2640 25560 3195
rect 26040 2820 26160 4395
rect 29940 3405 30060 4095
rect 26340 2100 26460 2160
rect 25740 1005 25860 1980
rect 26295 1905 26505 2100
rect 26940 1305 27060 3195
rect 29040 1605 29160 2595
rect 29340 2190 29460 2895
rect 30240 2640 30360 3795
rect 31440 2205 31560 3195
rect 31740 2190 31860 3795
rect 36540 3705 36660 5460
rect 32595 2700 32805 2895
rect 32640 2640 32760 2700
rect 33240 2640 33360 3195
rect 33840 2190 33960 3495
rect 36405 3240 36795 3360
rect 36495 2700 36705 2895
rect 36540 2640 36660 2700
rect 38340 2805 38460 3795
rect 31095 1905 31305 1980
rect 32040 705 32160 1995
rect 32895 1905 33105 1980
rect 35340 1605 35460 2610
rect 37500 2160 37695 2205
rect 36240 1005 36360 1695
rect 36840 1605 36960 2160
rect 37440 2040 37695 2160
rect 37500 1995 37695 2040
rect 38040 1905 38160 2610
rect 38940 2640 39060 4095
rect 39540 3105 39660 12795
rect 39840 8505 39960 11895
rect 40440 11505 40560 13260
rect 40395 10860 40605 10980
rect 40395 10800 40695 10860
rect 40440 10740 40695 10800
rect 40740 10440 40860 10695
rect 41340 10440 42060 10560
rect 41040 8805 41160 9960
rect 39840 5505 39960 7695
rect 40695 6000 40905 6195
rect 41340 6120 41460 6795
rect 41940 6405 42060 10440
rect 42240 10005 42360 13260
rect 43440 10440 43560 14295
rect 44940 13740 45060 14295
rect 45840 13290 45960 14595
rect 46740 13920 46860 14295
rect 44640 12405 44760 13260
rect 47040 12105 47160 12495
rect 44595 10605 44805 10695
rect 42840 6705 42960 9780
rect 43740 9405 43860 9960
rect 44340 8805 44460 10395
rect 44940 9990 45060 10695
rect 45240 10605 45360 10995
rect 45795 10500 46005 10695
rect 45840 10440 45960 10500
rect 47340 10305 47460 15180
rect 47640 13290 47760 20895
rect 47940 18405 48060 19995
rect 48240 18705 48360 20895
rect 49290 20880 49305 21000
rect 49095 20805 49305 20880
rect 49740 20505 49860 21510
rect 51195 21705 51405 21795
rect 51540 21105 51660 22695
rect 48540 18240 48660 18795
rect 49140 18240 49860 18360
rect 47940 15405 48060 17295
rect 48795 13800 49005 13995
rect 49740 13920 49860 18240
rect 50040 18105 50160 19095
rect 51240 18705 51360 20895
rect 51540 18240 51660 20580
rect 51840 19305 51960 24540
rect 52440 23205 52560 25395
rect 53340 24705 53460 25560
rect 54240 25560 54360 26595
rect 55005 26460 55200 26505
rect 55005 26295 55260 26460
rect 55140 26040 55260 26295
rect 54240 25440 54960 25560
rect 55740 25440 56160 25560
rect 52740 21540 52860 22395
rect 52140 20505 52260 21510
rect 54240 21105 54360 23295
rect 54540 22305 54660 25440
rect 54840 21540 54960 23895
rect 56040 22605 56160 25440
rect 52395 20805 52605 20895
rect 52140 18405 52260 20295
rect 53040 19605 53160 21060
rect 53640 20505 53760 21060
rect 55140 20505 55260 21060
rect 50340 14205 50460 18195
rect 52440 17790 52560 18495
rect 52995 18300 53205 18495
rect 53040 18240 53160 18300
rect 53640 18240 53760 18795
rect 54240 18405 54360 19395
rect 54540 17790 54660 20295
rect 55140 18240 55260 20295
rect 55740 18405 55860 20895
rect 51840 17205 51960 17760
rect 48840 13740 48960 13800
rect 49440 13740 49695 13860
rect 50340 13740 50460 13995
rect 53340 13740 53460 14895
rect 53940 13740 54060 15495
rect 54840 14205 54960 17595
rect 55440 17205 55560 17580
rect 56040 17505 56160 22395
rect 56340 15960 56460 29340
rect 56640 21720 56760 28095
rect 57240 28005 57360 28860
rect 56940 26205 57060 26895
rect 57840 26805 57960 28860
rect 58440 28305 58560 29310
rect 58740 26460 58860 29595
rect 59340 29520 59460 32595
rect 59940 29340 60060 31095
rect 60540 28905 60660 33810
rect 59640 28305 59760 28860
rect 60840 28005 60960 34995
rect 61140 34005 61260 36480
rect 61440 34305 61560 37995
rect 62340 37605 62460 41595
rect 63240 40605 63360 41160
rect 63840 40305 63960 41160
rect 61740 36705 61860 37395
rect 62640 37140 62760 39195
rect 64140 37320 64260 40995
rect 62340 36600 62460 36660
rect 62295 36405 62505 36600
rect 62940 35505 63060 36660
rect 64440 35205 64560 42540
rect 64740 38205 64860 42195
rect 65040 38805 65160 43095
rect 65940 41640 66060 44040
rect 66540 43305 66660 44340
rect 67740 42405 67860 46995
rect 68040 43605 68160 51795
rect 68340 49905 68460 52140
rect 69540 52005 69660 53895
rect 69840 52260 69960 55395
rect 70140 52905 70260 59595
rect 71640 54705 71760 64395
rect 72840 64005 72960 64560
rect 74340 64005 74460 64395
rect 71940 62805 72060 63195
rect 71940 59205 72060 62280
rect 72540 60720 72660 63195
rect 73140 60540 73260 61395
rect 73440 60705 73560 63795
rect 74040 61905 74160 62295
rect 74640 61305 74760 64995
rect 74940 63405 75060 65295
rect 75240 65205 75360 67695
rect 75540 65505 75660 67995
rect 75840 67605 75960 68280
rect 75840 65040 75960 65595
rect 76140 65505 76260 67695
rect 76440 67305 76560 67860
rect 77040 66705 77160 67860
rect 76440 65220 76560 66495
rect 76740 65205 76860 65595
rect 75240 61905 75360 64395
rect 75540 63705 75660 64560
rect 75840 62805 75960 63795
rect 76140 62205 76260 64560
rect 72540 57240 72660 59595
rect 72840 59505 72960 60060
rect 71940 56640 72360 56760
rect 71940 54105 72060 56640
rect 70440 52740 70560 53295
rect 69840 52140 70260 52260
rect 68640 49620 68760 50595
rect 69195 49500 69405 49695
rect 69240 49440 69360 49500
rect 68340 48405 68460 48795
rect 69540 48405 69660 48960
rect 70140 48105 70260 52140
rect 71940 52140 72360 52260
rect 70440 48405 70560 51795
rect 71940 51705 72060 52140
rect 73140 51060 73260 58995
rect 73740 58905 73860 59895
rect 73440 57360 73560 58095
rect 74940 57705 75060 59460
rect 75240 58005 75360 58695
rect 76140 58305 76260 61095
rect 76440 60090 76560 64095
rect 77040 61605 77160 65895
rect 77640 65160 77760 67695
rect 77940 66105 78060 69195
rect 78240 66705 78360 69495
rect 77505 65040 77760 65160
rect 78195 65220 78405 65295
rect 78540 65160 78660 71895
rect 78840 71205 78960 72195
rect 80340 71805 80460 72360
rect 78840 70005 78960 70395
rect 80340 69105 80460 69795
rect 79695 68400 79905 68595
rect 80640 68505 80760 70995
rect 81240 69105 81360 72180
rect 79740 68340 79860 68400
rect 81240 68340 81360 68895
rect 81540 68805 81660 74595
rect 81795 73005 82005 73095
rect 82140 72840 82260 76695
rect 82440 76305 82560 79395
rect 82740 76140 82860 77895
rect 83640 76560 83760 79995
rect 83940 77505 84060 82095
rect 84540 81660 84660 85440
rect 84840 82305 84960 85740
rect 85140 84105 85260 86895
rect 85740 86505 85860 87780
rect 86340 85605 86460 89895
rect 86940 88440 87060 89580
rect 87840 89505 87960 91260
rect 87240 87105 87360 87960
rect 87840 87405 87960 87960
rect 85740 83940 85860 85095
rect 87540 84120 87660 84495
rect 87840 84360 87960 85395
rect 88140 84705 88260 87795
rect 88440 87705 88560 93195
rect 88740 91905 88860 94440
rect 90040 93405 90160 94560
rect 88995 91800 89205 91995
rect 89040 91740 89160 91800
rect 87840 84240 88260 84360
rect 88140 83940 88260 84240
rect 85305 83460 85500 83505
rect 85305 83340 85560 83460
rect 86040 83400 86160 83460
rect 85305 83295 85500 83340
rect 85995 83205 86205 83400
rect 87105 83340 87360 83460
rect 84240 81540 84660 81660
rect 84240 77160 84360 81540
rect 86040 81405 86160 82995
rect 84540 80805 84660 81195
rect 85440 80640 85560 81195
rect 86940 81105 87060 83295
rect 88740 83460 88860 91095
rect 89040 89205 89160 89595
rect 89340 88620 89460 90795
rect 89640 90105 89760 91260
rect 89640 88860 89760 89895
rect 89640 88740 90060 88860
rect 89940 88440 90060 88740
rect 90540 88005 90660 88995
rect 89040 83505 89160 85095
rect 88440 83340 88860 83460
rect 87540 82260 87660 82695
rect 87540 82140 87960 82260
rect 87195 81660 87405 81795
rect 87195 81600 87660 81660
rect 87240 81540 87660 81600
rect 85140 79605 85260 80160
rect 85740 79305 85860 80160
rect 86040 78105 86160 79995
rect 86340 79005 86460 80895
rect 86895 80700 87105 80895
rect 87540 80805 87660 81540
rect 86940 80640 87060 80700
rect 87840 80205 87960 82140
rect 85140 77205 85260 77595
rect 84240 77040 84660 77160
rect 83340 76440 83760 76560
rect 83340 76140 83460 76440
rect 84240 75690 84360 76695
rect 83040 74760 83160 75480
rect 83040 74640 83460 74760
rect 83340 73005 83460 74640
rect 81840 68520 81960 72195
rect 82140 68505 82260 70395
rect 83040 69705 83160 72360
rect 83340 70605 83460 72195
rect 83640 69405 83760 73095
rect 83940 73005 84060 73995
rect 84240 73305 84360 75480
rect 84540 73605 84660 77040
rect 85140 76140 85260 76995
rect 86640 75660 86760 78495
rect 86040 75105 86160 75660
rect 86340 75540 86760 75660
rect 84240 72840 84360 73095
rect 84840 72840 84960 74595
rect 85440 73005 85560 74295
rect 85740 73905 85860 74595
rect 86340 74505 86460 75540
rect 86940 74205 87060 79095
rect 87240 74505 87360 79395
rect 88140 78705 88260 82695
rect 88440 79605 88560 83340
rect 89340 82905 89460 87495
rect 89940 83940 90060 84495
rect 91140 83505 91260 93795
rect 89340 80640 89460 81195
rect 87840 76320 87960 76995
rect 89940 76905 90060 82095
rect 90240 79305 90360 83295
rect 90540 81705 90660 83460
rect 91440 82305 91560 87795
rect 91440 80640 91560 81495
rect 91740 80805 91860 89295
rect 90840 79560 90960 80160
rect 90540 79440 90960 79560
rect 90540 78105 90660 79440
rect 90840 78405 90960 79095
rect 89805 76560 90000 76605
rect 89805 76395 90060 76560
rect 88395 76200 88605 76395
rect 88440 76140 88560 76200
rect 89940 76140 90060 76395
rect 88140 75105 88260 75660
rect 88740 75600 89160 75660
rect 88740 75540 89205 75600
rect 88995 75405 89205 75540
rect 84540 71805 84660 72180
rect 85140 72105 85260 72360
rect 84840 71940 85095 72060
rect 84840 70305 84960 71940
rect 85440 71760 85560 72195
rect 85140 71640 85560 71760
rect 78840 67305 78960 67695
rect 78540 65040 78960 65160
rect 77340 63705 77460 64995
rect 77640 63405 77760 64395
rect 76695 60705 76905 60795
rect 77295 60600 77505 60795
rect 77640 60660 77760 61395
rect 77940 61005 78060 64560
rect 78840 64305 78960 65040
rect 79140 64605 79260 65595
rect 79440 65505 79560 67860
rect 80040 67005 80160 67860
rect 80340 65205 80460 67695
rect 80940 67605 81060 67860
rect 81540 67560 81660 67860
rect 81240 67440 81660 67560
rect 79740 63705 79860 64380
rect 80340 61905 80460 64395
rect 80640 63105 80760 67095
rect 80940 66705 81060 67395
rect 81240 65220 81360 67440
rect 82140 67305 82260 67695
rect 82440 65205 82560 68295
rect 82740 67005 82860 69195
rect 83340 68340 83460 68895
rect 84540 68505 84660 69795
rect 81540 62205 81660 64560
rect 77340 60540 77460 60600
rect 77640 60540 78060 60660
rect 76740 59505 76860 59895
rect 76440 58605 76560 58995
rect 73440 57240 73860 57360
rect 74295 57300 74505 57495
rect 74340 57240 74460 57300
rect 73440 54105 73560 56580
rect 72840 50940 73260 51060
rect 71040 49440 71160 49995
rect 71640 49440 71760 50295
rect 72240 49605 72360 50895
rect 72000 48960 72195 49005
rect 71940 48840 72195 48960
rect 72000 48795 72195 48840
rect 72540 48660 72660 49695
rect 72240 48540 72660 48660
rect 69540 44940 69660 45495
rect 69840 45105 69960 46095
rect 70140 44340 70395 44460
rect 68340 43905 68460 44295
rect 68040 42705 68160 43395
rect 68340 41640 68460 42195
rect 66240 40860 66360 41160
rect 65940 40740 66360 40860
rect 65940 38805 66060 40740
rect 65400 37560 65595 37605
rect 65340 37395 65595 37560
rect 65340 37140 65460 37395
rect 65940 37305 66060 38280
rect 64305 35040 64560 35205
rect 64740 36540 64995 36660
rect 64305 34995 64500 35040
rect 61740 33840 61860 34695
rect 62340 33840 62460 34695
rect 61440 33300 61560 33360
rect 61140 31905 61260 33195
rect 61395 33105 61605 33300
rect 61440 29805 61560 32895
rect 62040 30060 62160 33180
rect 61740 29940 62160 30060
rect 61740 29340 61860 29940
rect 62340 29340 62460 30195
rect 62595 29805 62805 29895
rect 58740 26340 59160 26460
rect 59040 26220 59160 26340
rect 59640 26205 59760 27780
rect 56940 22905 57060 25395
rect 57240 24105 57360 25560
rect 58440 24960 58560 26010
rect 58140 24840 58560 24960
rect 56640 18405 56760 20595
rect 56940 20505 57060 21060
rect 57840 20505 57960 23895
rect 58140 20205 58260 24840
rect 58740 24405 58860 25395
rect 59340 22005 59460 25560
rect 59640 21720 59760 25395
rect 59940 21660 60060 26895
rect 60840 26505 60960 27480
rect 62040 27060 62160 28860
rect 62040 26940 62460 27060
rect 61140 26040 61260 26895
rect 62040 25590 62160 26595
rect 62340 26205 62460 26940
rect 62940 26505 63060 34695
rect 63240 31305 63360 34095
rect 64440 33840 64560 34695
rect 64740 34005 64860 36540
rect 66240 36690 66360 40395
rect 66540 39705 66660 40995
rect 66840 39405 66960 41595
rect 67440 38505 67560 41160
rect 68040 38805 68160 40980
rect 68640 40605 68760 40995
rect 66840 37320 66960 37995
rect 67440 37140 67560 37695
rect 68940 37620 69060 42795
rect 69840 42405 69960 44295
rect 70140 43260 70260 44340
rect 70140 43140 70560 43260
rect 70140 41640 70260 42795
rect 70440 41805 70560 43140
rect 71340 43005 71460 47895
rect 71640 42705 71760 48195
rect 71940 45105 72060 46695
rect 72240 44940 72360 48540
rect 72840 46605 72960 50940
rect 73440 50505 73560 53295
rect 74040 52740 74160 56265
rect 75240 56205 75360 57795
rect 75540 55305 75660 57495
rect 77940 57360 78060 60540
rect 78240 58905 78360 61695
rect 79395 60600 79605 60795
rect 79440 60540 79560 60600
rect 79800 60060 79995 60105
rect 78540 58005 78660 59895
rect 79140 59505 79260 60060
rect 79740 59940 79995 60060
rect 79800 59895 79995 59940
rect 77640 57240 78060 57360
rect 75240 54405 75360 54795
rect 75840 54360 75960 56595
rect 76140 55605 76260 56760
rect 77040 56640 77460 56760
rect 75540 54240 75960 54360
rect 75240 53460 75360 54195
rect 74940 53340 75360 53460
rect 74940 52950 75060 53340
rect 75540 52905 75660 54240
rect 75540 52140 75795 52260
rect 75240 51060 75360 52095
rect 74940 50940 75360 51060
rect 73095 49605 73305 49695
rect 73695 49500 73905 49695
rect 73740 49440 73860 49500
rect 73140 48840 73560 48960
rect 73140 47805 73260 48840
rect 74640 48960 74760 49395
rect 73995 48705 74205 48780
rect 74340 48840 74760 48960
rect 74340 47805 74460 48840
rect 73140 45150 73260 45495
rect 73440 45405 73560 47295
rect 73440 43605 73560 44280
rect 70440 39660 70560 40995
rect 70740 39705 70860 42195
rect 70140 39540 70560 39660
rect 69240 38205 69360 38895
rect 69540 37905 69660 39195
rect 65340 35805 65460 36195
rect 65040 31605 65160 35295
rect 65340 34005 65460 35595
rect 65940 33840 66060 36495
rect 68040 35205 68160 36795
rect 67140 33960 67260 34995
rect 67140 33840 67560 33960
rect 65640 32505 65760 33360
rect 66240 31305 66360 33360
rect 66840 31905 66960 33360
rect 67140 30405 67260 33195
rect 63240 29940 63795 30060
rect 63240 29505 63360 29940
rect 63495 29400 63705 29595
rect 63540 29340 63660 29400
rect 64740 29505 64860 29895
rect 65040 29205 65160 29595
rect 64440 28305 64560 28860
rect 63240 26160 63360 28095
rect 62940 26040 63360 26160
rect 61440 25500 61560 25560
rect 61395 25305 61605 25500
rect 59940 21540 60360 21660
rect 58740 19905 58860 20880
rect 59340 20505 59460 21060
rect 60240 19005 60360 21540
rect 60540 21090 60660 25095
rect 62340 25005 62460 25395
rect 63540 25500 63660 25560
rect 63495 25305 63705 25500
rect 62640 19305 62760 22695
rect 64140 22305 64260 27795
rect 64740 27405 64860 28695
rect 65640 28800 65760 28860
rect 64995 28605 65205 28680
rect 65340 26805 65460 28695
rect 65595 28605 65805 28800
rect 66240 28005 66360 28860
rect 64440 23505 64560 26295
rect 66240 25560 66360 26595
rect 65040 24405 65160 25560
rect 65340 23805 65460 24795
rect 65640 24105 65760 25560
rect 65940 25440 66360 25560
rect 60405 18840 60660 18960
rect 56805 17760 57000 17805
rect 56805 17640 57060 17760
rect 57540 17700 57660 17760
rect 56805 17595 57000 17640
rect 57495 17505 57705 17700
rect 58440 17505 58560 18795
rect 59340 18240 59460 18795
rect 60540 17790 60660 18840
rect 61740 18240 61860 18795
rect 56340 15840 56760 15960
rect 54540 14040 54795 14160
rect 54540 13605 54660 14040
rect 55140 13740 55260 14895
rect 55695 13800 55905 13995
rect 56340 13905 56460 15495
rect 55740 13740 55860 13800
rect 48540 11805 48660 13260
rect 49095 13005 49305 13080
rect 49995 13005 50205 13080
rect 47640 10605 47760 11595
rect 51240 11205 51360 13260
rect 48240 10440 48360 10995
rect 48840 10440 48960 10995
rect 50340 10440 50460 10995
rect 40740 5940 40860 6000
rect 42540 5940 42660 6495
rect 43095 6000 43305 6195
rect 43140 5940 43260 6000
rect 44640 5805 44760 8895
rect 46140 6705 46260 9960
rect 46740 8505 46860 9960
rect 47805 9990 48000 10005
rect 47805 9795 47895 9990
rect 47040 9105 47160 9795
rect 49140 9405 49260 9960
rect 50040 9405 50160 9960
rect 50640 9105 50760 9960
rect 51540 9705 51660 10395
rect 51840 9105 51960 13080
rect 52740 10440 52860 12495
rect 56040 12405 56160 13260
rect 53340 11205 53460 12195
rect 53340 10440 53460 10995
rect 53940 10005 54060 12195
rect 54240 10605 54360 10995
rect 54540 10440 54660 11595
rect 55095 10500 55305 10695
rect 55140 10440 55260 10500
rect 52440 9105 52560 9960
rect 56040 9990 56160 10695
rect 56340 10005 56460 10395
rect 56640 10305 56760 15840
rect 56940 11805 57060 17295
rect 59295 17205 59505 17295
rect 57540 13740 57660 14595
rect 59340 13305 59460 16095
rect 60540 13905 60660 14295
rect 60840 13920 60960 18195
rect 61440 17205 61560 17760
rect 62040 17700 62160 17760
rect 61995 17505 62205 17700
rect 62940 17205 63060 22095
rect 63795 21720 64005 21795
rect 64740 21660 64860 22395
rect 65940 22005 66060 25440
rect 66540 25305 66660 28395
rect 67140 28005 67260 29880
rect 67440 28605 67560 31695
rect 68340 30405 68460 37395
rect 69540 37140 69660 37695
rect 70140 37305 70260 39540
rect 71040 39360 71160 42495
rect 72240 41640 72360 42195
rect 72540 41805 72660 42795
rect 73740 42405 73860 46695
rect 74040 44505 74160 47295
rect 74640 46305 74760 48495
rect 74940 48405 75060 50940
rect 75540 50505 75660 52140
rect 76140 49440 76260 50895
rect 75195 48705 75405 48795
rect 74640 45705 74760 46095
rect 75240 45105 75360 45495
rect 70740 39240 71160 39360
rect 70440 36690 70560 38595
rect 69240 34260 69360 36660
rect 69840 35805 69960 36480
rect 70740 36405 70860 39240
rect 71340 38505 71460 40995
rect 71940 40605 72060 41160
rect 72840 41100 72960 41160
rect 72240 40305 72360 40695
rect 72240 37305 72360 40095
rect 72540 37605 72660 40995
rect 72795 40905 73005 41100
rect 74340 40905 74460 44895
rect 74640 40560 74760 44295
rect 75540 44205 75660 48195
rect 75840 46905 75960 48960
rect 76440 47505 76560 48795
rect 76740 47160 76860 53295
rect 77040 51105 77160 55995
rect 77340 55905 77460 56640
rect 77340 52905 77460 55095
rect 77640 53205 77760 57240
rect 78840 56805 78960 58695
rect 79140 57705 79260 58395
rect 78240 54405 78360 56760
rect 79140 56460 79260 57495
rect 78840 56340 79260 56460
rect 78840 55005 78960 56340
rect 77700 52860 77895 52905
rect 77640 52740 77895 52860
rect 77700 52695 77895 52740
rect 78840 52860 78960 54195
rect 79140 54105 79260 55995
rect 78540 52740 78960 52860
rect 77040 48105 77160 50295
rect 77340 49905 77460 52095
rect 78840 51105 78960 52095
rect 79140 51405 79260 53895
rect 79440 53505 79560 58095
rect 80640 57405 80760 60795
rect 80940 60705 81060 61995
rect 82140 61605 82260 64065
rect 82740 62805 82860 64995
rect 83040 64590 83160 67395
rect 83340 65205 83460 67395
rect 83640 67005 83760 67860
rect 84540 66405 84660 67695
rect 83940 65040 84060 66195
rect 84540 65040 84660 65595
rect 84840 65505 84960 69195
rect 85140 65205 85260 71640
rect 85740 69960 85860 73380
rect 86340 73305 86460 73695
rect 87540 73260 87660 74895
rect 87540 73200 87960 73260
rect 87540 73140 88005 73200
rect 87795 73005 88005 73140
rect 86295 72105 86505 72195
rect 86940 71805 87060 72360
rect 85440 69840 85860 69960
rect 84240 64500 84360 64560
rect 84195 64305 84405 64500
rect 83040 61005 83160 61995
rect 83340 60405 83460 63495
rect 79440 52290 79560 52980
rect 78240 49440 78360 49995
rect 78840 49440 78960 50580
rect 79740 50205 79860 56295
rect 80340 56205 80460 56760
rect 80940 52905 81060 60180
rect 82140 58005 82260 59460
rect 81240 56205 81360 57795
rect 82395 57300 82605 57495
rect 82440 57240 82560 57300
rect 83040 57405 83160 57795
rect 82905 57210 83160 57405
rect 83640 57360 83760 62595
rect 83940 60105 84060 63495
rect 84240 60705 84360 61095
rect 84540 60540 84660 64095
rect 84840 63405 84960 64560
rect 85140 63705 85260 64395
rect 85440 61005 85560 69840
rect 87540 69705 87660 72180
rect 85740 68805 85860 69495
rect 85740 66705 85860 67395
rect 86640 66105 86760 67260
rect 85740 65205 85860 65895
rect 85995 65100 86205 65295
rect 86040 65040 86160 65100
rect 87240 65205 87360 66495
rect 87540 64560 87660 67395
rect 86340 64500 86460 64560
rect 86940 64500 87060 64560
rect 85440 60660 85560 60795
rect 85140 60540 85560 60660
rect 82800 57195 83160 57210
rect 82140 55905 82260 56760
rect 80205 52860 80400 52905
rect 80205 52740 80460 52860
rect 80205 52695 80400 52740
rect 81495 52800 81705 52995
rect 82095 52800 82305 52995
rect 81540 52740 81660 52800
rect 82140 52740 82260 52800
rect 80040 50805 80160 52095
rect 76440 47040 76860 47160
rect 75840 42105 75960 45795
rect 76140 43905 76260 46395
rect 75705 41940 75960 42105
rect 75705 41895 75900 41940
rect 75540 41640 76095 41760
rect 74340 40500 74760 40560
rect 74295 40440 74760 40500
rect 74295 40305 74505 40440
rect 73095 37200 73305 37395
rect 73140 37140 73260 37200
rect 73740 37140 73860 40095
rect 74040 37260 74160 38895
rect 74340 37560 74460 39495
rect 74640 38640 75360 38760
rect 74640 38205 74760 38640
rect 74340 37440 74760 37560
rect 74040 37140 74460 37260
rect 71340 36600 71460 36660
rect 69240 34200 69660 34260
rect 69240 34140 69705 34200
rect 69495 34005 69705 34140
rect 68640 33360 68760 33810
rect 70740 33360 70860 34995
rect 68640 33240 69060 33360
rect 68940 32505 69060 33240
rect 70140 33240 70860 33360
rect 69240 31605 69360 31995
rect 67995 30060 68205 30195
rect 67995 30000 68460 30060
rect 68040 29940 68460 30000
rect 68340 29760 68460 29940
rect 68340 29640 68595 29760
rect 67995 29400 68205 29595
rect 68040 29340 68160 29400
rect 68640 29340 68760 29595
rect 68940 29505 69060 31095
rect 70740 30705 70860 31395
rect 67140 26040 67260 27195
rect 67740 26220 67860 28095
rect 68040 26205 68160 28395
rect 67440 25500 67560 25560
rect 67395 25305 67605 25500
rect 66240 22605 66360 25095
rect 67095 24960 67305 25095
rect 67095 24900 67695 24960
rect 67140 24840 67695 24900
rect 68340 24105 68460 28095
rect 68940 26505 69060 28695
rect 69240 28005 69360 30195
rect 71040 29805 71160 36495
rect 71295 36405 71505 36600
rect 72240 35205 72360 36495
rect 72240 33840 72360 34680
rect 72540 34020 72660 36795
rect 71940 32505 72060 33360
rect 72840 32805 72960 33795
rect 69540 28305 69660 29595
rect 69540 26040 69660 27195
rect 69840 26505 69960 29295
rect 64440 21540 64860 21660
rect 63540 18705 63660 21060
rect 64140 20505 64260 21060
rect 65040 19560 65160 21795
rect 65595 21600 65805 21795
rect 65640 21540 65760 21600
rect 66240 21540 66360 22395
rect 68595 21600 68805 21795
rect 68940 21705 69060 25065
rect 68640 21540 68760 21600
rect 65940 20505 66060 21060
rect 67305 20940 67860 21060
rect 65040 19440 65460 19560
rect 63240 14805 63360 18195
rect 63240 14205 63360 14595
rect 63840 14505 63960 17760
rect 64440 16305 64560 17760
rect 65040 16905 65160 19095
rect 65340 16305 65460 19440
rect 66300 18660 66495 18705
rect 66240 18495 66495 18660
rect 66240 18240 66360 18495
rect 64440 15405 64560 16095
rect 65040 14505 65160 15795
rect 63840 14040 64395 14160
rect 62295 13800 62505 13995
rect 62340 13740 62460 13800
rect 60840 13290 60960 13710
rect 63840 13740 63960 14040
rect 62940 13305 63060 13695
rect 65040 13305 65160 14295
rect 61140 13200 61395 13260
rect 61095 13140 61395 13200
rect 61095 13005 61305 13140
rect 57840 10440 57960 10995
rect 50640 8505 50760 8895
rect 45240 5940 45360 6495
rect 45795 6000 46005 6195
rect 47295 6000 47505 6195
rect 45840 5940 45960 6000
rect 47340 5940 47460 6000
rect 47940 5940 48060 6795
rect 48240 6105 48360 6495
rect 41940 5205 42060 5595
rect 48540 5505 48660 5910
rect 40140 2190 40260 3195
rect 40740 2640 40860 4395
rect 41340 2640 41460 4995
rect 38640 2100 38760 2160
rect 38595 1905 38805 2100
rect 41640 2100 41760 2160
rect 41595 1905 41805 2100
rect 42240 1005 42360 4095
rect 42540 3105 42660 4695
rect 43440 4305 43560 5460
rect 46140 5400 46260 5460
rect 47040 5400 47160 5460
rect 46095 5205 46305 5400
rect 46995 5205 47205 5400
rect 47640 4905 47760 5460
rect 48195 5205 48405 5295
rect 48495 4905 48705 4980
rect 48840 4605 48960 6195
rect 49140 6105 49260 6795
rect 49395 6000 49605 6195
rect 49440 5940 49560 6000
rect 50640 5940 50760 7695
rect 55440 7305 55560 7695
rect 52140 5490 52260 7095
rect 52995 6000 53205 6195
rect 53040 5940 53160 6000
rect 53640 5940 53760 6795
rect 54540 5490 54660 6195
rect 55440 5940 55560 7095
rect 55740 6405 55860 9795
rect 57495 9705 57705 9780
rect 56640 7005 56760 9495
rect 58140 9405 58260 9960
rect 58740 9405 58860 10695
rect 59595 10500 59805 10695
rect 59640 10440 59760 10500
rect 60240 10440 60360 11295
rect 59340 9900 59460 9960
rect 59295 9705 59505 9900
rect 57240 5940 57360 6495
rect 59640 5940 59760 6495
rect 49740 4905 49860 5460
rect 51540 4905 51660 5460
rect 43905 2895 43995 3105
rect 42540 2190 42660 2895
rect 45540 2820 45660 4395
rect 48705 4140 49095 4260
rect 44100 2760 44295 2805
rect 44040 2640 44295 2760
rect 44100 2595 44295 2640
rect 48240 2640 48360 3795
rect 48840 2640 48960 3795
rect 50340 2640 50460 4695
rect 50640 2805 50760 3195
rect 51240 2640 51360 3495
rect 44640 2190 44760 2595
rect 47040 2190 47160 2595
rect 44940 1605 45060 1995
rect 47340 1605 47460 2295
rect 52740 2205 52860 4395
rect 53340 4305 53460 5460
rect 53940 5205 54060 5460
rect 53940 5040 54195 5205
rect 54000 4995 54195 5040
rect 55305 4995 55395 5175
rect 56340 4905 56460 5910
rect 47940 1305 48060 1980
rect 50940 705 51060 1995
rect 51840 705 51960 2160
rect 53040 1905 53160 3495
rect 53340 2805 53460 3195
rect 53640 2640 53760 4395
rect 54840 2805 54960 4695
rect 56940 4005 57060 5460
rect 57540 5400 57660 5460
rect 59340 5400 59460 5460
rect 57495 5205 57705 5400
rect 59295 5205 59505 5400
rect 59040 3240 59160 4695
rect 60540 3405 60660 5895
rect 60840 4905 60960 12195
rect 61140 9990 61260 10995
rect 61440 9105 61560 11595
rect 62040 11205 62160 13260
rect 63540 13200 63660 13260
rect 63495 13005 63705 13200
rect 63840 10905 63960 11295
rect 63840 10440 63960 10695
rect 61740 7905 61860 10095
rect 63300 9960 63495 10005
rect 62340 8805 62460 9960
rect 63240 9840 63495 9960
rect 63300 9795 63495 9840
rect 62340 6705 62460 8595
rect 64440 6120 64560 10695
rect 64740 9990 64860 11595
rect 65340 10905 65460 16095
rect 65640 13905 65760 14595
rect 66105 14160 66300 14205
rect 66105 13995 66360 14160
rect 66240 13740 66360 13995
rect 66540 13860 66660 16995
rect 67140 16905 67260 18495
rect 67440 18405 67560 20595
rect 67695 18300 67905 18495
rect 67740 18240 67860 18300
rect 66840 15960 66960 16695
rect 66840 15840 67260 15960
rect 66540 13740 66960 13860
rect 66840 12105 66960 13740
rect 67140 11205 67260 15840
rect 67440 13905 67560 15195
rect 68040 14160 68160 17580
rect 67740 14040 68160 14160
rect 67740 13740 67860 14040
rect 68340 13740 68460 15795
rect 68940 15705 69060 20895
rect 69240 20505 69360 25395
rect 69840 25005 69960 25560
rect 69540 21090 69660 22095
rect 69840 21705 69960 23595
rect 70140 21960 70260 25395
rect 70440 22305 70560 26595
rect 70740 26505 70860 28860
rect 71040 26040 71160 28695
rect 71340 26505 71460 30795
rect 72540 29340 72660 31995
rect 73140 30405 73260 34095
rect 73440 34005 73560 36660
rect 74340 36105 74460 37140
rect 73740 33840 73860 35595
rect 74640 35505 74760 37440
rect 74940 37305 75060 38295
rect 75240 37560 75360 38640
rect 75840 37605 75960 40995
rect 76140 39105 76260 41280
rect 76440 41205 76560 47040
rect 76740 45405 76860 46395
rect 77340 46305 77460 49380
rect 77940 47805 78060 48960
rect 78540 48405 78660 48960
rect 77505 46140 77760 46260
rect 77205 43995 77295 44205
rect 76740 41805 76860 43695
rect 77040 41640 77160 42795
rect 77340 42105 77460 43395
rect 77640 42705 77760 46140
rect 79140 45405 79260 48195
rect 77940 43305 78060 45195
rect 79140 44940 79260 45195
rect 79740 45120 79860 47595
rect 80640 47460 80760 48195
rect 80940 47805 81060 51195
rect 80640 47340 81060 47460
rect 80040 45105 80160 47295
rect 80340 45360 80460 46995
rect 80940 45705 81060 47340
rect 81240 46305 81360 51495
rect 81840 51405 81960 52260
rect 81540 49605 81660 50895
rect 81840 49440 81960 50595
rect 82440 49920 82560 51795
rect 82740 51105 82860 55995
rect 83040 53205 83160 57195
rect 83340 57240 83760 57360
rect 83940 57240 84060 57795
rect 84540 57240 84660 58095
rect 84840 57705 84960 60060
rect 85140 57405 85260 57795
rect 83340 54105 83460 57240
rect 83640 53805 83760 56595
rect 85440 56760 85560 59895
rect 85740 58005 85860 64395
rect 86295 64305 86505 64500
rect 86895 64305 87105 64500
rect 87240 64440 87660 64560
rect 86040 60705 86160 64095
rect 86940 61905 87060 64095
rect 87240 64005 87360 64440
rect 87840 64260 87960 72195
rect 88140 67605 88260 74295
rect 88440 72405 88560 73995
rect 88440 68505 88560 69795
rect 88740 69405 88860 74895
rect 90240 73905 90360 75660
rect 91140 75105 91260 76110
rect 91440 75405 91560 76695
rect 91740 72960 91860 79995
rect 92040 77805 92160 85395
rect 91605 72840 91860 72960
rect 91140 72060 91260 72495
rect 90840 71940 91260 72060
rect 90840 71505 90960 71940
rect 89940 68805 90060 70695
rect 91440 70005 91560 72795
rect 92040 68805 92160 73395
rect 89940 68340 90660 68460
rect 88440 67305 88560 67695
rect 88740 65505 88860 67680
rect 89340 66405 89460 67860
rect 89040 65040 89160 65595
rect 89640 65205 89760 67695
rect 89940 67005 90060 68340
rect 91440 67305 91560 67860
rect 90240 65040 90360 66195
rect 88140 64305 88260 64995
rect 88740 64500 88860 64560
rect 87540 64140 87960 64260
rect 86340 61305 86460 61695
rect 86295 60600 86505 60780
rect 86940 60720 87060 61380
rect 86340 60540 86460 60600
rect 84195 56505 84405 56580
rect 84840 56205 84960 56760
rect 85140 56640 85560 56760
rect 82995 52905 83205 52995
rect 83295 52800 83505 52995
rect 83340 52740 83460 52800
rect 83940 52740 84060 54795
rect 83040 49605 83160 52095
rect 80340 45300 80760 45360
rect 80340 45240 80805 45300
rect 80595 45105 80805 45240
rect 77640 41640 77760 42180
rect 78240 41805 78360 43995
rect 75240 37440 75660 37560
rect 75540 37140 75660 37440
rect 76440 37305 76560 40680
rect 74940 35205 75060 36495
rect 74040 31605 74160 33360
rect 71640 26040 71760 27495
rect 72540 26205 72660 28395
rect 73140 27405 73260 30195
rect 74640 29805 74760 34095
rect 74940 33960 75060 34995
rect 75240 34305 75360 36660
rect 75840 34005 75960 34995
rect 76140 34905 76260 35895
rect 76440 34905 76560 36495
rect 76740 35805 76860 40695
rect 77940 40605 78060 41160
rect 78540 39405 78660 43095
rect 79740 43005 79860 44910
rect 80940 44940 81060 45495
rect 78840 41805 78960 42195
rect 80040 41805 80160 44295
rect 81240 43605 81360 44295
rect 80340 42105 80460 43095
rect 77040 37305 77160 39195
rect 78840 39060 78960 40995
rect 79140 40860 79260 41160
rect 79140 40740 79695 40860
rect 78540 38940 78960 39060
rect 77640 37140 77760 37695
rect 76695 34905 76905 34995
rect 74940 33840 75360 33960
rect 76140 33360 76260 34095
rect 76440 33705 76560 34695
rect 77040 33960 77160 36495
rect 78240 35760 78360 38295
rect 77940 35640 78360 35760
rect 76740 33840 77160 33960
rect 77340 33840 77460 34695
rect 77940 33840 78060 35640
rect 78540 35460 78660 38940
rect 80040 38505 80160 40995
rect 80340 40605 80460 41580
rect 80640 40905 80760 41295
rect 78840 36405 78960 37995
rect 80640 37305 80760 38295
rect 79740 36600 79860 36660
rect 78240 35340 78660 35460
rect 78240 34305 78360 35340
rect 78840 35205 78960 35595
rect 78540 35040 78795 35160
rect 75840 33240 76260 33360
rect 73440 27360 73560 29595
rect 73440 27240 73860 27360
rect 72795 26100 73005 26295
rect 72840 26040 72960 26100
rect 71340 22905 71460 25560
rect 72540 23505 72660 25395
rect 70140 21840 70560 21960
rect 70440 21540 70560 21840
rect 70995 21600 71205 21795
rect 71040 21540 71160 21600
rect 70140 20205 70260 20880
rect 70740 19605 70860 21060
rect 71640 18450 71760 21495
rect 71940 21105 72060 21795
rect 73440 21540 73560 22395
rect 73740 22005 73860 27240
rect 74040 25560 74160 28395
rect 74340 26205 74460 28695
rect 74640 27405 74760 28860
rect 75240 27405 75360 29595
rect 75540 27360 75660 32595
rect 75840 28605 75960 33240
rect 76740 31605 76860 33840
rect 76995 33105 77205 33195
rect 76140 29505 76260 30795
rect 77640 30105 77760 33360
rect 76395 29400 76605 29595
rect 76440 29340 76560 29400
rect 77640 28560 77760 28860
rect 77640 28440 78060 28560
rect 75540 27240 75960 27360
rect 74640 26805 74760 27195
rect 75840 26205 75960 27240
rect 74040 25440 74460 25560
rect 74040 21705 74160 25095
rect 74340 22905 74460 25440
rect 74640 24705 74760 25560
rect 75540 25500 75660 25560
rect 75495 25305 75705 25500
rect 73740 20505 73860 21060
rect 69540 16605 69660 17760
rect 71940 17205 72060 19995
rect 72240 18405 72360 19395
rect 72405 17760 72600 17805
rect 74040 17760 74160 20895
rect 74340 20805 74460 22380
rect 72405 17640 72660 17760
rect 72405 17595 72600 17640
rect 73605 17640 74160 17760
rect 68640 11805 68760 13080
rect 69240 12405 69360 14895
rect 70140 14505 70260 16695
rect 70440 16305 70560 16695
rect 70740 13740 70860 14295
rect 69540 13305 69660 13710
rect 71340 13305 71460 16095
rect 71640 12705 71760 14595
rect 72540 13740 72660 14895
rect 72240 12705 72360 13260
rect 64995 10560 65205 10695
rect 64995 10500 65460 10560
rect 65040 10440 65460 10500
rect 65640 7905 65760 9960
rect 66840 9405 66960 10395
rect 67740 9900 67860 9960
rect 67140 8805 67260 9795
rect 67695 9705 67905 9900
rect 68640 8205 68760 10995
rect 69540 10440 69660 12495
rect 69240 9405 69360 9960
rect 69840 9900 69960 9960
rect 69795 9705 70005 9900
rect 68940 8505 69060 8895
rect 61440 4005 61560 5460
rect 56040 2640 56160 3195
rect 53940 2100 54060 2160
rect 53895 1905 54105 2100
rect 55440 1605 55560 2295
rect 57540 2205 57660 3195
rect 56340 705 56460 2160
rect 60240 1005 60360 2295
rect 60540 2190 60660 3195
rect 61995 2805 62205 2895
rect 61140 1305 61260 1980
rect 61740 1605 61860 2160
rect 62340 1605 62460 2610
rect 63195 1605 63405 1695
rect 64440 1005 64560 5910
rect 64740 5505 64860 7095
rect 65340 5940 65460 6795
rect 65895 6000 66105 6195
rect 65940 5940 66060 6000
rect 67440 5460 67560 7395
rect 70440 6060 70560 10695
rect 71040 8805 71160 11895
rect 71595 10500 71805 10695
rect 71640 10440 71760 10500
rect 72240 10440 72360 11595
rect 72840 10605 72960 13260
rect 73740 10905 73860 17640
rect 74340 17505 74460 19995
rect 74340 16005 74460 17295
rect 74295 14805 74505 14895
rect 74205 14700 74505 14805
rect 74205 14640 74460 14700
rect 74205 14595 74400 14640
rect 74340 13740 74460 14295
rect 74640 14205 74760 21795
rect 75540 21540 75660 22695
rect 75840 22005 75960 25395
rect 76140 24705 76260 27495
rect 75240 21000 75360 21060
rect 75195 20805 75405 21000
rect 75840 20505 75960 21060
rect 74940 13920 75060 15795
rect 75840 14505 75960 18195
rect 76140 14205 76260 20895
rect 76440 15105 76560 28395
rect 76740 22305 76860 26895
rect 77640 26040 77760 27795
rect 77940 27705 78060 28440
rect 78240 26205 78360 28695
rect 78540 26805 78660 35040
rect 79140 34905 79260 36495
rect 79695 36405 79905 36600
rect 80940 36660 81060 42795
rect 81240 41805 81360 43395
rect 81540 42405 81660 47595
rect 81840 42105 81960 45495
rect 82740 44940 82860 45795
rect 83040 45105 83160 48795
rect 83340 47805 83460 50895
rect 83640 49605 83760 50295
rect 83940 49860 84060 51795
rect 84240 50205 84360 52260
rect 84540 50505 84660 52095
rect 83940 49740 84360 49860
rect 84240 49440 84360 49740
rect 84840 49620 84960 51495
rect 83640 47205 83760 48795
rect 83940 48105 84060 48960
rect 84540 48405 84660 48960
rect 85140 48105 85260 56640
rect 85740 56460 85860 57480
rect 86040 57405 86160 59895
rect 86640 59505 86760 60060
rect 86640 57240 86760 57795
rect 86940 57705 87060 58095
rect 87240 57405 87360 59895
rect 87540 59205 87660 64140
rect 86340 56700 86460 56760
rect 85440 56340 85860 56460
rect 85440 52905 85560 56340
rect 86040 54405 86160 56595
rect 86295 56505 86505 56700
rect 85740 53205 85860 53895
rect 86640 52920 86760 56295
rect 86940 53805 87060 56265
rect 85440 48705 85560 52095
rect 85740 51405 85860 52260
rect 85740 50205 85860 50595
rect 86340 49905 86460 50595
rect 86640 49440 86760 51195
rect 86940 49605 87060 52080
rect 83340 46005 83460 46395
rect 83640 44940 83760 46095
rect 82140 42705 82260 44895
rect 83895 44205 84105 44295
rect 84240 43305 84360 44895
rect 84540 44505 84660 47880
rect 84840 45105 84960 47595
rect 86340 47505 86460 48960
rect 83040 42705 83160 43095
rect 84240 42705 84360 43095
rect 85140 42705 85260 44460
rect 85740 44160 85860 44280
rect 85440 44040 85860 44160
rect 83295 42405 83505 42495
rect 81495 41700 81705 41880
rect 81540 41640 81660 41700
rect 82695 41700 82905 41895
rect 82740 41640 82860 41700
rect 81240 37305 81360 40995
rect 81840 39705 81960 41160
rect 83340 41190 83460 41880
rect 84195 41700 84405 41895
rect 84240 41640 84360 41700
rect 83040 39360 83160 40995
rect 83940 41100 84060 41160
rect 83895 40905 84105 41100
rect 82740 39240 83160 39360
rect 81540 37140 81660 37995
rect 82395 37200 82605 37395
rect 82740 37305 82860 39240
rect 82440 37140 82560 37200
rect 83040 36705 83160 38295
rect 80640 36540 81060 36660
rect 79890 36300 79905 36405
rect 79440 33840 79560 35295
rect 80040 34005 80160 36195
rect 79140 33060 79260 33360
rect 79140 32940 79560 33060
rect 77340 25005 77460 25560
rect 77040 21540 77160 22695
rect 77640 21720 77760 23295
rect 77940 23205 78060 25560
rect 77940 21705 78060 22095
rect 76740 16305 76860 20895
rect 77340 19005 77460 21060
rect 78240 18660 78360 25395
rect 78540 24105 78660 26280
rect 78840 26205 78960 31095
rect 79140 29505 79260 32595
rect 79440 31005 79560 32940
rect 79740 29805 79860 33360
rect 80040 32805 80160 33195
rect 80340 31305 80460 34995
rect 80640 32805 80760 36540
rect 82140 35205 82260 36495
rect 83340 36405 83460 37395
rect 83940 37140 84060 39795
rect 84540 37605 84660 40995
rect 84840 40005 84960 42195
rect 85440 42060 85560 44040
rect 86340 43605 86460 46395
rect 86640 45105 86760 48495
rect 86940 47805 87060 48795
rect 87240 48705 87360 52695
rect 87540 51405 87660 57795
rect 87840 57705 87960 63795
rect 88440 62505 88560 64395
rect 88695 64305 88905 64500
rect 88740 61020 88860 64095
rect 89340 63705 89460 64560
rect 89340 60540 89460 61695
rect 89640 60705 89760 64395
rect 90540 63705 90660 64560
rect 90240 63540 90495 63660
rect 88140 59505 88260 59895
rect 88440 58005 88560 60060
rect 89040 59505 89160 60060
rect 88305 57660 88500 57705
rect 88305 57495 88560 57660
rect 88395 57420 88560 57495
rect 89040 57405 89160 57795
rect 88140 56700 88260 56760
rect 87840 56205 87960 56595
rect 88095 56505 88305 56700
rect 88740 56205 88860 56760
rect 87840 50805 87960 54195
rect 88140 52905 88260 54795
rect 89040 54105 89160 56595
rect 88440 52740 88560 53295
rect 89040 52740 89160 53895
rect 89340 52905 89460 57195
rect 88140 50205 88260 52095
rect 88740 51705 88860 52260
rect 86940 44940 87060 45795
rect 87540 45105 87660 49995
rect 89040 49905 89160 51795
rect 89340 49905 89460 52095
rect 88395 49500 88605 49695
rect 89100 49590 89400 49605
rect 89100 49545 89295 49590
rect 88440 49440 88560 49500
rect 89040 49425 89295 49545
rect 89100 49395 89295 49425
rect 88140 48900 88260 48960
rect 88095 48705 88305 48900
rect 85140 42000 85560 42060
rect 85095 41940 85560 42000
rect 85095 41805 85305 41940
rect 85740 41640 85860 42495
rect 86640 42105 86760 44295
rect 87240 43905 87360 44460
rect 87540 42405 87660 44295
rect 87840 43905 87960 46695
rect 88140 45705 88260 47595
rect 88440 46905 88560 48195
rect 88740 48105 88860 48960
rect 88440 44940 88560 46380
rect 89040 46260 89160 48495
rect 88740 46140 89160 46260
rect 88740 45405 88860 46140
rect 89040 44940 89160 45795
rect 89340 45105 89460 48795
rect 88140 43005 88260 43695
rect 86295 41700 86505 41895
rect 86940 41805 87060 42195
rect 88440 42120 88560 43995
rect 88740 43005 88860 44460
rect 86340 41640 86460 41700
rect 87240 41205 87360 41895
rect 85440 41100 85560 41160
rect 84495 37200 84705 37395
rect 85140 37305 85260 40995
rect 85395 40905 85605 41100
rect 86040 37860 86160 41160
rect 85740 37740 86160 37860
rect 84540 37140 84660 37200
rect 82440 34860 82560 35295
rect 83940 35205 84060 36195
rect 84840 36105 84960 36660
rect 82140 34740 82560 34860
rect 82140 33840 82260 34740
rect 83640 34305 83760 34695
rect 81240 33060 81360 33360
rect 80940 32940 81360 33060
rect 80640 29505 80760 31395
rect 80940 31005 81060 32940
rect 82740 32805 82860 33810
rect 81240 31905 81360 32595
rect 79740 28605 79860 28860
rect 79140 26505 79260 28395
rect 79740 27105 79860 28395
rect 80640 27705 80760 28695
rect 80940 26805 81060 29895
rect 81240 28905 81360 31695
rect 81540 29505 81660 32295
rect 83640 31005 83760 31395
rect 81840 29340 81960 30195
rect 82995 29400 83205 29595
rect 83295 29505 83505 29595
rect 83040 29340 83160 29400
rect 83640 28890 83760 30795
rect 83940 29805 84060 32895
rect 84240 29505 84360 33360
rect 84840 32505 84960 34995
rect 85140 31005 85260 36495
rect 85440 36405 85560 37395
rect 85740 37305 85860 37740
rect 86340 37560 86460 38595
rect 86640 38205 86760 41160
rect 86940 37605 87060 40995
rect 87240 39705 87360 40995
rect 88740 39405 88860 40995
rect 86340 37440 86760 37560
rect 85995 37200 86205 37395
rect 86040 37140 86160 37200
rect 86640 37140 86760 37440
rect 85740 36105 85860 36495
rect 86040 34260 86160 36195
rect 86340 34560 86460 36660
rect 87540 36690 87660 38295
rect 86340 34440 86760 34560
rect 86040 34140 86460 34260
rect 86340 33840 86460 34140
rect 86640 34005 86760 34440
rect 87240 33960 87360 36495
rect 86940 33840 87360 33960
rect 87540 33840 87660 35895
rect 87840 34905 87960 37395
rect 88140 37305 88260 38895
rect 88740 37140 88860 38595
rect 89040 37605 89160 43695
rect 89340 43005 89460 44295
rect 89640 42060 89760 58995
rect 89940 57405 90060 60795
rect 90240 60705 90360 63540
rect 90540 60540 90660 61695
rect 91140 61020 91260 65595
rect 91440 61305 91560 66780
rect 91740 66405 91860 67695
rect 91740 60660 91860 66195
rect 92040 61005 92160 68280
rect 91740 60540 92160 60660
rect 90240 58305 90360 59895
rect 90540 57705 90660 59595
rect 91440 58905 91560 60060
rect 92040 59505 92160 60540
rect 91740 59340 91995 59460
rect 90240 57540 90495 57660
rect 90240 57240 90360 57540
rect 90840 57405 90960 58695
rect 90240 52905 90360 55095
rect 90540 54705 90660 56760
rect 90840 53460 90960 56595
rect 91140 53505 91260 58095
rect 91440 55005 91560 57495
rect 91740 55305 91860 59340
rect 90540 53400 90960 53460
rect 90495 53340 90960 53400
rect 90495 53205 90705 53340
rect 91140 53160 91260 53295
rect 90840 53040 91260 53160
rect 90840 52740 90960 53040
rect 91440 52740 91560 53895
rect 91740 52905 91860 54495
rect 89940 48405 90060 52695
rect 90240 49605 90360 50595
rect 90540 49905 90660 52260
rect 90840 49440 90960 49995
rect 90540 48900 90660 48960
rect 89940 44205 90060 47295
rect 90240 45105 90360 48795
rect 90495 48705 90705 48900
rect 90540 46005 90660 48180
rect 91140 47505 91260 48960
rect 90840 44940 90960 45495
rect 91440 45405 91560 48495
rect 91740 48105 91860 49995
rect 91740 45060 91860 47295
rect 92040 46005 92160 58695
rect 91440 44940 91860 45060
rect 92040 44490 92160 45195
rect 90240 42405 90360 44295
rect 90540 43605 90660 44460
rect 89505 41940 89760 42060
rect 89340 41160 89460 41895
rect 89895 41700 90105 41895
rect 89940 41640 90060 41700
rect 89340 41040 89760 41160
rect 89640 36705 89760 41040
rect 90240 40005 90360 40980
rect 89940 37305 90060 38595
rect 90240 37605 90360 39195
rect 90840 38805 90960 42195
rect 90240 37140 90360 37395
rect 90840 37140 90960 37995
rect 91140 37305 91260 39795
rect 88140 33960 88260 36495
rect 88440 36105 88560 36660
rect 89340 34905 89460 36495
rect 88740 34005 88860 34695
rect 88140 33840 88560 33960
rect 86040 32805 86160 33360
rect 86640 30405 86760 31695
rect 85305 29895 85395 30105
rect 84495 29805 84705 29895
rect 85395 29400 85605 29580
rect 85440 29340 85560 29400
rect 79095 26100 79305 26295
rect 79695 26100 79905 26295
rect 79140 26040 79260 26100
rect 79740 26040 79860 26100
rect 80340 25560 80460 26595
rect 80895 26100 81105 26280
rect 81540 26205 81660 28680
rect 81840 28005 81960 28395
rect 83940 28305 84060 28995
rect 84195 28605 84405 28695
rect 80940 26040 81060 26100
rect 78840 21705 78960 25395
rect 79440 25005 79560 25560
rect 80040 25440 80460 25560
rect 79140 23205 79260 24195
rect 79140 21540 79260 22995
rect 79740 21705 79860 22995
rect 77940 18540 78360 18660
rect 75540 13290 75660 13695
rect 75540 12705 75660 13080
rect 74595 10500 74805 10695
rect 74640 10440 74760 10500
rect 71940 9360 72060 9960
rect 72195 9360 72405 9495
rect 71940 9300 72405 9360
rect 71940 9240 72360 9300
rect 70140 5940 70560 6060
rect 70695 6000 70905 6195
rect 70740 5940 70860 6000
rect 65640 4905 65760 5460
rect 66240 5400 66360 5460
rect 66195 5205 66405 5400
rect 67440 5340 67860 5460
rect 65340 2640 65460 3795
rect 64740 1905 64860 2595
rect 66195 1905 66405 1995
rect 66540 1605 66660 2610
rect 67005 2760 67200 2805
rect 67005 2640 67260 2760
rect 67740 2640 67860 5340
rect 68340 2820 68460 5280
rect 70140 4905 70260 5940
rect 72240 5205 72360 9240
rect 72840 6150 72960 9795
rect 73140 9705 73260 10410
rect 73440 9840 73860 9960
rect 73440 5940 73560 9840
rect 67005 2595 67200 2640
rect 72540 2160 72660 3195
rect 72840 2160 72960 5940
rect 73740 4005 73860 5460
rect 74340 3405 74460 9960
rect 74640 7305 74760 9195
rect 74940 8805 75060 9960
rect 75240 5940 75360 8295
rect 75540 6405 75660 10395
rect 75840 9705 75960 13980
rect 76440 13905 76560 14295
rect 77040 14205 77160 17595
rect 77340 16305 77460 17760
rect 76890 13995 76905 14100
rect 76695 13800 76905 13995
rect 76740 13740 76860 13800
rect 77340 13740 77460 14595
rect 77940 14505 78060 18540
rect 78540 18360 78660 21495
rect 78840 18660 78960 20895
rect 79440 20505 79560 21060
rect 78840 18540 79260 18660
rect 78240 18240 78660 18360
rect 79140 18240 79260 18540
rect 78240 17505 78360 18240
rect 80040 18405 80160 25440
rect 80340 21705 80460 25095
rect 80640 22860 80760 25395
rect 80640 22740 81060 22860
rect 80640 21540 80760 22395
rect 80940 22005 81060 22740
rect 81240 22605 81360 25560
rect 81540 23205 81660 25395
rect 81840 22305 81960 27795
rect 82140 25560 82260 28095
rect 84240 26805 84360 28080
rect 84540 27705 84660 28860
rect 85695 28305 85905 28395
rect 86040 28005 86160 29310
rect 86340 28905 86460 29595
rect 86640 29460 86760 29880
rect 86940 29805 87060 33840
rect 87240 29760 87360 33195
rect 87840 31605 87960 33360
rect 87240 29640 87660 29760
rect 86640 29340 87060 29460
rect 87540 29340 87660 29640
rect 87795 29505 88005 29595
rect 86805 28395 86895 28605
rect 84540 27105 84660 27495
rect 82440 26205 82560 26595
rect 83895 25800 84105 26010
rect 83940 25740 84060 25800
rect 82140 25440 82560 25560
rect 82140 24405 82260 25095
rect 82440 22005 82560 25440
rect 83040 24705 83160 25560
rect 83640 21390 83760 25095
rect 85110 24105 85230 25095
rect 85440 24705 85560 27495
rect 87240 27405 87360 28860
rect 88140 28605 88260 29295
rect 87840 27405 87960 28095
rect 88440 27405 88560 33840
rect 89640 33840 89760 35295
rect 89940 34305 90060 36495
rect 90240 35460 90360 35895
rect 90540 35805 90660 36660
rect 90240 35340 90660 35460
rect 90240 34005 90360 34695
rect 88740 29505 88860 33195
rect 89040 31005 89160 33360
rect 89340 29340 89460 30195
rect 89940 29340 90060 33360
rect 90240 29460 90360 33195
rect 90540 30405 90660 35340
rect 90840 34905 90960 35895
rect 90240 29340 90660 29460
rect 88740 27705 88860 28695
rect 89640 28305 89760 28860
rect 89505 27540 90060 27660
rect 85740 25305 85860 26295
rect 89640 26205 89760 27195
rect 89940 25905 90060 27540
rect 89505 25860 89700 25905
rect 89505 25740 89760 25860
rect 89505 25695 89700 25740
rect 90540 25860 90660 29340
rect 90840 26160 90960 34095
rect 91140 28890 91260 36495
rect 91440 36105 91560 43995
rect 90840 26040 91260 26160
rect 90540 25740 90960 25860
rect 85740 22905 85860 23595
rect 88440 22755 88695 22860
rect 88440 22740 88860 22755
rect 88440 21840 88560 22740
rect 78840 17700 78960 17760
rect 79440 17700 79560 17760
rect 78795 17505 79005 17700
rect 79395 17505 79605 17700
rect 76140 11205 76260 13680
rect 76440 12105 76560 13095
rect 77040 12660 77160 13260
rect 78240 13290 78360 15495
rect 79140 14160 79260 16995
rect 80340 16905 80460 20895
rect 81540 18960 81660 21060
rect 82140 20505 82260 21180
rect 81540 18840 81960 18960
rect 81240 18240 81360 18795
rect 81840 18405 81960 18840
rect 80640 17805 80760 18195
rect 82140 17805 82260 19095
rect 79440 14505 79560 16695
rect 81540 15105 81660 17580
rect 81840 15705 81960 17595
rect 82440 15705 82560 20895
rect 83040 19605 83160 20595
rect 83340 19305 83460 20295
rect 83640 19905 83760 21180
rect 83940 20805 84060 21795
rect 82695 18420 82905 18495
rect 85140 18120 85260 19695
rect 85440 18405 85560 19395
rect 85740 18360 85860 19695
rect 87840 19605 87960 21180
rect 89040 20505 89160 22095
rect 89340 20205 89460 22695
rect 89640 19905 89760 24795
rect 90240 21720 90360 25260
rect 90540 22005 90660 25095
rect 90840 22305 90960 25740
rect 91140 22905 91260 26040
rect 89940 18405 90060 20295
rect 85740 18240 86160 18360
rect 82740 17700 82995 17760
rect 82695 17640 82995 17700
rect 82695 17505 82905 17640
rect 85740 17460 85860 17910
rect 86040 17505 86160 18240
rect 90240 18105 90360 19995
rect 90840 18405 90960 20895
rect 91140 18105 91260 21795
rect 91440 19560 91560 35295
rect 91740 35160 91860 43695
rect 92040 39105 92160 42795
rect 92040 35505 92160 37995
rect 91740 35040 92160 35160
rect 91740 21105 91860 34695
rect 91440 19440 91860 19560
rect 89805 18060 90000 18105
rect 89805 17940 90060 18060
rect 89805 17895 90000 17940
rect 91440 17760 91560 19095
rect 91140 17640 91560 17760
rect 85440 17340 85860 17460
rect 79140 14040 79560 14160
rect 79440 13920 79560 14040
rect 78705 13860 78900 13905
rect 78705 13740 78960 13860
rect 78705 13695 78900 13740
rect 80040 13905 80160 14295
rect 80340 13305 80460 13995
rect 80940 13740 81060 14895
rect 81600 13860 81795 13905
rect 81540 13740 81795 13860
rect 81600 13695 81795 13740
rect 77940 12660 78060 13095
rect 77040 12540 78060 12660
rect 76395 10500 76605 10695
rect 76440 10440 76560 10500
rect 77040 10440 77160 10995
rect 78540 10440 78660 11895
rect 79140 11805 79260 13080
rect 79140 11205 79260 11595
rect 79740 10620 79860 13260
rect 81795 13005 82005 13095
rect 82140 10620 82260 13395
rect 75840 5940 75960 6495
rect 76740 6060 76860 9780
rect 77340 7605 77460 9960
rect 78240 9405 78360 9960
rect 80640 9900 80760 9960
rect 78840 9105 78960 9780
rect 80595 9705 80805 9900
rect 81240 7605 81360 9960
rect 81840 8805 81960 9960
rect 82440 8505 82560 14895
rect 82740 12105 82860 16695
rect 83295 13800 83505 13995
rect 83340 13740 83460 13800
rect 83940 13740 84060 16395
rect 85440 14760 85560 17340
rect 91140 17460 91260 17640
rect 90540 17340 91260 17460
rect 85740 15105 85860 16995
rect 90180 16605 90300 16995
rect 87840 15105 87960 16095
rect 85440 14700 85860 14760
rect 85440 14640 85905 14700
rect 85440 14220 85560 14640
rect 85695 14505 85905 14640
rect 83640 11205 83760 13260
rect 84240 13200 84360 13260
rect 84195 13005 84405 13200
rect 83940 11340 84495 11460
rect 83340 10440 83460 10995
rect 83940 10440 84060 11340
rect 84840 11160 84960 13995
rect 86040 13200 86160 13260
rect 85995 13005 86205 13200
rect 84540 11040 84960 11160
rect 84240 10605 84360 10995
rect 83640 9105 83760 9960
rect 84540 7560 84660 11040
rect 84840 9105 84960 10695
rect 85740 10440 85860 11295
rect 86295 10500 86505 10695
rect 86340 10440 86460 10500
rect 84240 7440 84660 7560
rect 85140 7560 85260 9795
rect 85440 8205 85560 9960
rect 85140 7440 85560 7560
rect 76740 5940 77160 6060
rect 76140 5400 76260 5460
rect 76095 5205 76305 5400
rect 77040 5205 77160 5940
rect 77340 4005 77460 6495
rect 80640 5940 80760 7395
rect 81495 6000 81705 6195
rect 82395 6000 82605 6195
rect 81540 5940 81660 6000
rect 82440 5940 82560 6000
rect 83340 5940 83460 6795
rect 83940 5805 84060 7095
rect 84240 6405 84360 7440
rect 85440 6105 85560 7440
rect 75240 2820 75360 3795
rect 77940 2760 78060 3795
rect 78240 3405 78360 5460
rect 77940 2640 78360 2760
rect 80640 2820 80760 3195
rect 83940 2820 84060 5595
rect 85305 5340 85560 5460
rect 78240 2160 78360 2640
rect 85440 2760 85560 5340
rect 85740 4605 85860 8295
rect 86040 7005 86160 9960
rect 86640 9900 86760 9960
rect 86595 9705 86805 9900
rect 86595 7860 86805 7995
rect 86340 7800 86805 7860
rect 86340 7740 86760 7800
rect 86340 5940 86460 7740
rect 86640 6360 86760 7395
rect 86940 7305 87060 9795
rect 87240 6405 87360 14895
rect 87840 13740 87960 14295
rect 87705 10560 87900 10605
rect 87705 10440 87960 10560
rect 87705 10395 87900 10440
rect 88140 8805 88260 9960
rect 88740 6405 88860 11895
rect 89040 8205 89160 16095
rect 89940 13920 90060 14895
rect 89940 9900 90060 9960
rect 89895 9705 90105 9900
rect 86640 6240 87060 6360
rect 86940 5940 87060 6240
rect 87240 4605 87360 5460
rect 85440 2640 85860 2760
rect 86640 2640 86760 4395
rect 87840 2190 87960 6195
rect 88140 5490 88260 6195
rect 89040 5940 89160 6495
rect 89340 5160 89460 5460
rect 89340 5040 89760 5160
rect 89340 2640 89460 4695
rect 89640 4305 89760 5040
rect 90240 4905 90360 7395
rect 90540 5490 90660 15495
rect 90840 4305 90960 16695
rect 91140 6705 91260 16995
rect 68040 1005 68160 2160
rect 41805 495 41895 705
rect 42705 495 42795 705
rect 70140 -240 70260 2160
rect 75840 -240 75960 2160
rect 81240 -240 81360 2160
rect 83340 -240 83460 2160
rect 69840 -360 70260 -240
rect 75540 -360 75960 -240
rect 80940 -360 81360 -240
rect 83040 -360 83460 -240
rect 85140 -360 85260 2160
rect 87240 -240 87360 2160
rect 89640 2100 89760 2160
rect 89595 1905 89805 2100
rect 91140 1905 91260 6495
rect 91440 6120 91560 17295
rect 91740 7605 91860 19440
rect 92040 16905 92160 35040
rect 92040 4605 92160 16095
rect 86940 -360 87360 -240
<< m3contact >>
rect 49995 93795 50205 94005
rect 58095 93795 58305 94005
rect 72795 93795 73005 94005
rect 52995 93495 53205 93705
rect 57795 93495 58005 93705
rect 4395 93195 4605 93405
rect 9795 93195 10005 93405
rect 13695 93195 13905 93405
rect 1395 92295 1605 92505
rect 3795 92295 4005 92505
rect 2595 91710 2805 91920
rect 3195 91710 3405 91920
rect 7695 92595 7905 92805
rect 5895 92295 6105 92505
rect 4380 91695 4590 91905
rect 4695 91710 4905 91920
rect 5295 91710 5505 91920
rect 8895 91995 9105 92205
rect 7695 91710 7905 91920
rect 11295 92895 11505 93105
rect 10995 92595 11205 92805
rect 10395 91710 10605 91920
rect 13095 92295 13305 92505
rect 11295 91995 11505 92205
rect 11895 91995 12105 92205
rect 12795 91995 13005 92205
rect 1695 88695 1905 88905
rect 2295 88410 2505 88620
rect 3495 91080 3705 91290
rect 4095 91080 4305 91290
rect 4695 91095 4905 91305
rect 6195 91080 6405 91290
rect 7095 91080 7305 91290
rect 5595 89295 5805 89505
rect 5895 88710 6105 88920
rect 3195 88395 3405 88605
rect 4095 88410 4305 88620
rect 4995 88410 5205 88620
rect 5895 88410 6105 88620
rect 6495 88410 6705 88620
rect 1395 87195 1605 87405
rect 1395 84195 1605 84405
rect 1095 83910 1305 84120
rect 495 82695 705 82905
rect 195 80610 405 80820
rect 195 78495 405 78705
rect 2895 87195 3105 87405
rect 2595 86595 2805 86805
rect 2295 85695 2505 85905
rect 1995 82695 2205 82905
rect 1395 82095 1605 82305
rect 1995 82095 2205 82305
rect 4395 87780 4605 87990
rect 3795 86595 4005 86805
rect 4995 87495 5205 87705
rect 6195 87780 6405 87990
rect 5895 87495 6105 87705
rect 5595 87195 5805 87405
rect 4395 85395 4605 85605
rect 3195 84795 3405 85005
rect 4095 84795 4305 85005
rect 2595 83895 2805 84105
rect 3495 83910 3705 84120
rect 3195 83280 3405 83490
rect 795 81495 1005 81705
rect 2895 81795 3105 82005
rect 1995 80610 2205 80820
rect 3795 81495 4005 81705
rect 3195 80895 3405 81105
rect 4395 83910 4605 84120
rect 4995 83910 5205 84120
rect 8895 91095 9105 91305
rect 9495 91080 9705 91290
rect 10095 91080 10305 91290
rect 11595 91080 11805 91290
rect 12195 91080 12405 91290
rect 21495 92895 21705 93105
rect 29895 92895 30105 93105
rect 31095 92895 31305 93105
rect 33495 92895 33705 93105
rect 47895 92895 48105 93105
rect 48795 92895 49005 93105
rect 52995 92895 53205 93105
rect 16395 92295 16605 92505
rect 17895 92295 18105 92505
rect 20595 92295 20805 92505
rect 14295 91710 14505 91920
rect 15195 91710 15405 91920
rect 16995 91710 17205 91920
rect 13095 91395 13305 91605
rect 13995 91080 14205 91290
rect 12795 90795 13005 91005
rect 7995 90495 8205 90705
rect 9495 90495 9705 90705
rect 11595 90495 11805 90705
rect 8895 89895 9105 90105
rect 8295 88695 8505 88905
rect 7395 88395 7605 88605
rect 11895 90195 12105 90405
rect 14595 90195 14805 90405
rect 12795 89895 13005 90105
rect 9795 89595 10005 89805
rect 11895 89595 12105 89805
rect 15195 89595 15405 89805
rect 9495 89295 9705 89505
rect 7095 87195 7305 87405
rect 7095 85695 7305 85905
rect 5895 83895 6105 84105
rect 6495 83910 6705 84120
rect 7995 87780 8205 87990
rect 8595 87780 8805 87990
rect 9195 87780 9405 87990
rect 8295 87195 8505 87405
rect 9195 87195 9405 87405
rect 7995 83910 8205 84120
rect 4395 83295 4605 83505
rect 5295 83280 5505 83490
rect 5895 83295 6105 83505
rect 9195 85695 9405 85905
rect 8595 84495 8805 84705
rect 7095 82995 7305 83205
rect 7995 82995 8205 83205
rect 5295 82095 5505 82305
rect 5895 82095 6105 82305
rect 6795 82095 7005 82305
rect 4395 81795 4605 82005
rect 4395 81195 4605 81405
rect 4095 80895 4305 81105
rect 3195 79980 3405 80190
rect 4095 79980 4305 80190
rect 2295 79695 2505 79905
rect 2895 79695 3105 79905
rect 1395 79095 1605 79305
rect 4680 79095 4890 79305
rect 4995 79095 5205 79305
rect 2895 78195 3105 78405
rect 1395 76995 1605 77205
rect 795 76110 1005 76320
rect 1995 76110 2205 76320
rect 495 75480 705 75690
rect 2295 75480 2505 75690
rect 1695 75195 1905 75405
rect 2595 73095 2805 73305
rect 6195 81195 6405 81405
rect 8295 81195 8505 81405
rect 7695 80610 7905 80820
rect 16695 91080 16905 91290
rect 18495 91710 18705 91920
rect 19995 91710 20205 91920
rect 24795 92295 25005 92505
rect 26595 92295 26805 92505
rect 28095 92295 28305 92505
rect 22095 91710 22305 91920
rect 22695 91710 22905 91920
rect 23595 91710 23805 91920
rect 25995 91710 26205 91920
rect 27195 91710 27405 91920
rect 18795 90795 19005 91005
rect 19995 90795 20205 91005
rect 17895 89595 18105 89805
rect 14895 88995 15105 89205
rect 16095 88995 16305 89205
rect 10995 88410 11205 88620
rect 12195 88395 12405 88605
rect 13395 88410 13605 88620
rect 13995 88410 14205 88620
rect 10695 87495 10905 87705
rect 10695 86895 10905 87105
rect 11595 86895 11805 87105
rect 9495 84495 9705 84705
rect 10095 83910 10305 84120
rect 12195 85395 12405 85605
rect 12795 84795 13005 85005
rect 11895 84495 12105 84705
rect 12195 83910 12405 84120
rect 12795 83595 13005 83805
rect 9195 83280 9405 83490
rect 10695 83295 10905 83505
rect 11295 83280 11505 83490
rect 11895 83280 12105 83490
rect 13695 87495 13905 87705
rect 13695 83910 13905 84120
rect 13095 82695 13305 82905
rect 13995 82695 14205 82905
rect 9795 82095 10005 82305
rect 18495 88695 18705 88905
rect 15795 88410 16005 88620
rect 16995 88410 17205 88620
rect 15495 87495 15705 87705
rect 16395 85095 16605 85305
rect 15495 84495 15705 84705
rect 19395 88410 19605 88620
rect 21495 91080 21705 91290
rect 22395 91080 22605 91290
rect 22395 90495 22605 90705
rect 20895 90195 21105 90405
rect 20295 89895 20505 90105
rect 21195 89595 21405 89805
rect 20895 88995 21105 89205
rect 20895 88410 21105 88620
rect 18195 87780 18405 87990
rect 19695 87780 19905 87990
rect 20595 87495 20805 87705
rect 18795 87195 19005 87405
rect 20295 87195 20505 87405
rect 17295 85095 17505 85305
rect 16995 84195 17205 84405
rect 19095 86595 19305 86805
rect 18795 84795 19005 85005
rect 18495 84195 18705 84405
rect 17295 83910 17505 84120
rect 17895 83910 18105 84120
rect 16095 83280 16305 83490
rect 16995 83295 17205 83505
rect 14895 81495 15105 81705
rect 11295 81195 11505 81405
rect 12495 81195 12705 81405
rect 13695 81195 13905 81405
rect 8595 80895 8805 81105
rect 9195 80895 9405 81105
rect 10095 80895 10305 81105
rect 10695 80610 10905 80820
rect 11595 80595 11805 80805
rect 13095 80610 13305 80820
rect 6195 79695 6405 79905
rect 5895 79395 6105 79605
rect 5295 78195 5505 78405
rect 4995 76995 5205 77205
rect 3795 76110 4005 76320
rect 4395 76110 4605 76320
rect 3495 75480 3705 75690
rect 4095 74595 4305 74805
rect 3495 73095 3705 73305
rect 1695 72810 1905 73020
rect 2295 72195 2505 72405
rect 1995 71895 2205 72105
rect 1395 70995 1605 71205
rect 195 69795 405 70005
rect 1095 68895 1305 69105
rect 4095 72810 4305 73020
rect 4695 72795 4905 73005
rect 2595 71895 2805 72105
rect 495 68310 705 68520
rect 1095 68310 1305 68520
rect 1695 68310 1905 68520
rect 2280 68310 2490 68520
rect 4695 72180 4905 72390
rect 5295 76395 5505 76605
rect 6495 78795 6705 79005
rect 6795 76995 7005 77205
rect 5295 75195 5505 75405
rect 8595 79980 8805 80190
rect 9195 79980 9405 80190
rect 9795 79980 10005 80190
rect 11295 79980 11505 80190
rect 10395 79395 10605 79605
rect 7995 79095 8205 79305
rect 8295 78495 8505 78705
rect 7695 77895 7905 78105
rect 10395 77895 10605 78105
rect 12195 79695 12405 79905
rect 12795 79395 13005 79605
rect 11595 77295 11805 77505
rect 8295 76995 8505 77205
rect 7695 76110 7905 76320
rect 10095 76395 10305 76605
rect 10695 76110 10905 76320
rect 11295 76110 11505 76320
rect 7395 74895 7605 75105
rect 6495 74595 6705 74805
rect 9495 74895 9705 75105
rect 6195 74295 6405 74505
rect 7695 74295 7905 74505
rect 8595 74295 8805 74505
rect 5895 73395 6105 73605
rect 5595 72810 5805 73020
rect 7395 73395 7605 73605
rect 7095 72810 7305 73020
rect 5895 72180 6105 72390
rect 6495 72180 6705 72390
rect 3795 71595 4005 71805
rect 2895 70995 3105 71205
rect 3195 70995 3405 71205
rect 1395 66795 1605 67005
rect 795 65010 1005 65220
rect 1395 65010 1605 65220
rect 2595 68295 2805 68505
rect 3495 68895 3705 69105
rect 4395 68295 4605 68505
rect 3195 67680 3405 67890
rect 2595 67095 2805 67305
rect 195 58995 405 59205
rect 195 54195 405 54405
rect 2295 64995 2505 65205
rect 3495 65595 3705 65805
rect 4995 71595 5205 71805
rect 4995 70695 5205 70905
rect 4695 67695 4905 67905
rect 4395 67095 4605 67305
rect 3795 65295 4005 65505
rect 4395 65295 4605 65505
rect 4095 65010 4305 65220
rect 4680 65010 4890 65220
rect 7095 70095 7305 70305
rect 8295 73095 8505 73305
rect 8895 72810 9105 73020
rect 8295 71895 8505 72105
rect 7995 70995 8205 71205
rect 7395 69195 7605 69405
rect 5895 68295 6105 68505
rect 6495 68310 6705 68520
rect 5595 67680 5805 67890
rect 6195 66795 6405 67005
rect 5595 65595 5805 65805
rect 1695 64380 1905 64590
rect 2595 64395 2805 64605
rect 3195 64380 3405 64590
rect 1695 61095 1905 61305
rect 4995 64995 5205 65205
rect 6795 65295 7005 65505
rect 5295 64380 5505 64590
rect 6495 64395 6705 64605
rect 5895 64095 6105 64305
rect 8595 70695 8805 70905
rect 9195 70095 9405 70305
rect 7695 68310 7905 68520
rect 8295 68310 8505 68520
rect 7995 67680 8205 67890
rect 10395 75195 10605 75405
rect 18795 83895 19005 84105
rect 18195 83280 18405 83490
rect 13995 80610 14205 80820
rect 14595 80610 14805 80820
rect 15195 80610 15405 80820
rect 16095 80580 16305 80790
rect 14895 79980 15105 80190
rect 14595 79395 14805 79605
rect 15495 79395 15705 79605
rect 16095 79395 16305 79605
rect 13995 78495 14205 78705
rect 16695 81495 16905 81705
rect 17595 81195 17805 81405
rect 19695 83910 19905 84120
rect 21195 87795 21405 88005
rect 22095 87780 22305 87990
rect 23595 89895 23805 90105
rect 25095 91080 25305 91290
rect 25695 91080 25905 91290
rect 24495 88995 24705 89205
rect 23295 88410 23505 88620
rect 24195 88410 24405 88620
rect 25095 88410 25305 88620
rect 26895 91080 27105 91290
rect 27495 90495 27705 90705
rect 25995 90195 26205 90405
rect 28695 91710 28905 91920
rect 29295 91710 29505 91920
rect 30495 92595 30705 92805
rect 28695 91080 28905 91290
rect 26595 89295 26805 89505
rect 28095 89295 28305 89505
rect 23895 87780 24105 87990
rect 25395 87780 25605 87990
rect 23295 87195 23505 87405
rect 22995 86595 23205 86805
rect 25995 85995 26205 86205
rect 22095 83910 22305 84120
rect 24195 84195 24405 84405
rect 23595 83910 23805 84120
rect 24795 83895 25005 84105
rect 26295 85695 26505 85905
rect 28395 88995 28605 89205
rect 27195 88410 27405 88620
rect 28095 88410 28305 88620
rect 26895 87795 27105 88005
rect 27495 87780 27705 87990
rect 28095 87195 28305 87405
rect 26895 85995 27105 86205
rect 31695 91710 31905 91920
rect 32595 91710 32805 91920
rect 33795 92595 34005 92805
rect 35595 92595 35805 92805
rect 37095 92595 37305 92805
rect 46395 92595 46605 92805
rect 34095 91695 34305 91905
rect 36795 91710 37005 91920
rect 31395 91080 31605 91290
rect 29595 90795 29805 91005
rect 30495 90795 30705 91005
rect 29295 90195 29505 90405
rect 30795 89895 31005 90105
rect 29895 88410 30105 88620
rect 29595 87780 29805 87990
rect 30195 87780 30405 87990
rect 32595 91095 32805 91305
rect 33795 91080 34005 91290
rect 35295 91080 35505 91290
rect 31995 89295 32205 89505
rect 31695 88995 31905 89205
rect 33795 88410 34005 88620
rect 35295 88410 35505 88620
rect 36495 89295 36705 89505
rect 31695 87780 31905 87990
rect 30795 87495 31005 87705
rect 28695 86595 28905 86805
rect 35595 87780 35805 87990
rect 34095 87195 34305 87405
rect 33495 85995 33705 86205
rect 28695 85695 28905 85905
rect 36195 85695 36405 85905
rect 26595 85095 26805 85305
rect 26895 84195 27105 84405
rect 19995 82695 20205 82905
rect 20895 82695 21105 82905
rect 22995 83295 23205 83505
rect 23895 83280 24105 83490
rect 24795 83280 25005 83490
rect 25695 83280 25905 83490
rect 22395 82695 22605 82905
rect 25395 82695 25605 82905
rect 21795 82395 22005 82605
rect 24495 82395 24705 82605
rect 25695 82395 25905 82605
rect 25395 82095 25605 82305
rect 20295 81795 20505 82005
rect 21780 81795 21990 82005
rect 22095 81795 22305 82005
rect 19095 80610 19305 80820
rect 19695 80610 19905 80820
rect 17895 79980 18105 80190
rect 19395 79395 19605 79605
rect 17295 79095 17505 79305
rect 18795 79095 19005 79305
rect 16995 78495 17205 78705
rect 18495 78495 18705 78705
rect 16395 77895 16605 78105
rect 17595 77895 17805 78105
rect 14595 77295 14805 77505
rect 16395 77295 16605 77505
rect 12195 76110 12405 76320
rect 13095 76095 13305 76305
rect 17295 76695 17505 76905
rect 12495 75480 12705 75690
rect 11595 75195 11805 75405
rect 13095 75195 13305 75405
rect 11295 74295 11505 74505
rect 11880 74295 12090 74505
rect 12195 74295 12405 74505
rect 10395 73095 10605 73305
rect 10995 72810 11205 73020
rect 9795 72195 10005 72405
rect 10695 71595 10905 71805
rect 10995 70995 11205 71205
rect 11295 70695 11505 70905
rect 11595 70395 11805 70605
rect 11595 69795 11805 70005
rect 10995 68595 11205 68805
rect 10095 68310 10305 68520
rect 10695 68310 10905 68520
rect 11595 68295 11805 68505
rect 8895 67395 9105 67605
rect 9495 67395 9705 67605
rect 7995 66795 8205 67005
rect 8595 66795 8805 67005
rect 7995 65010 8205 65220
rect 7095 64395 7305 64605
rect 6795 63795 7005 64005
rect 4695 61095 4905 61305
rect 5895 61095 6105 61305
rect 3795 60795 4005 61005
rect 2295 60510 2505 60720
rect 2895 60510 3105 60720
rect 3495 60510 3705 60720
rect 795 59895 1005 60105
rect 1395 59880 1605 60090
rect 1995 59595 2205 59805
rect 1695 58695 1905 58905
rect 795 57495 1005 57705
rect 2295 58395 2505 58605
rect 4995 60495 5205 60705
rect 3195 59895 3405 60105
rect 2895 57195 3105 57405
rect 795 56580 1005 56790
rect 1395 56580 1605 56790
rect 2595 55995 2805 56205
rect 2895 53895 3105 54105
rect 1995 52680 2205 52890
rect 3795 59595 4005 59805
rect 4095 58395 4305 58605
rect 3795 57495 4005 57705
rect 4995 58695 5205 58905
rect 8295 64095 8505 64305
rect 7695 63795 7905 64005
rect 10395 67680 10605 67890
rect 9195 65895 9405 66105
rect 9795 65895 10005 66105
rect 13695 74595 13905 74805
rect 14895 75195 15105 75405
rect 14295 74295 14505 74505
rect 12795 72810 13005 73020
rect 16395 76110 16605 76320
rect 16095 74595 16305 74805
rect 15195 73995 15405 74205
rect 15195 73095 15405 73305
rect 12195 72195 12405 72405
rect 13095 72180 13305 72390
rect 14595 72180 14805 72390
rect 15195 72180 15405 72390
rect 13095 71595 13305 71805
rect 15795 70695 16005 70905
rect 13095 69495 13305 69705
rect 14595 69195 14805 69405
rect 12195 68295 12405 68505
rect 11895 67695 12105 67905
rect 10995 65295 11205 65505
rect 10095 65010 10305 65220
rect 9195 64095 9405 64305
rect 8895 63495 9105 63705
rect 10395 64395 10605 64605
rect 9795 62895 10005 63105
rect 13395 67395 13605 67605
rect 12195 67095 12405 67305
rect 12795 67095 13005 67305
rect 11595 66795 11805 67005
rect 15495 68895 15705 69105
rect 16395 72810 16605 73020
rect 20895 80595 21105 80805
rect 23295 80595 23505 80805
rect 24495 80610 24705 80820
rect 27495 83910 27705 84120
rect 28095 83910 28305 84120
rect 28995 85395 29205 85605
rect 29895 85095 30105 85305
rect 29295 84195 29505 84405
rect 28995 83910 29205 84120
rect 27795 83280 28005 83490
rect 28695 83295 28905 83505
rect 41595 92295 41805 92505
rect 42795 92295 43005 92505
rect 38595 91710 38805 91920
rect 40995 91710 41205 91920
rect 41595 91710 41805 91920
rect 42195 91710 42405 91920
rect 44295 91710 44505 91920
rect 36795 88395 37005 88605
rect 37695 91080 37905 91290
rect 40695 91080 40905 91290
rect 45495 91695 45705 91905
rect 40695 90495 40905 90705
rect 41295 90495 41505 90705
rect 38295 88995 38505 89205
rect 39495 88995 39705 89205
rect 37995 88410 38205 88620
rect 38595 88410 38805 88620
rect 40095 88410 40305 88620
rect 37095 87780 37305 87990
rect 40695 88395 40905 88605
rect 42495 88995 42705 89205
rect 39195 87780 39405 87990
rect 39795 87780 40005 87990
rect 37695 87195 37905 87405
rect 36495 84795 36705 85005
rect 40395 84795 40605 85005
rect 38895 84495 39105 84705
rect 33495 84195 33705 84405
rect 35895 84195 36105 84405
rect 37395 84195 37605 84405
rect 38295 84195 38505 84405
rect 30795 83910 31005 84120
rect 31995 83910 32205 84120
rect 32595 83910 32805 84120
rect 33195 83910 33405 84120
rect 29295 82995 29505 83205
rect 28395 82395 28605 82605
rect 28995 82395 29205 82605
rect 29280 81795 29490 82005
rect 29595 81795 29805 82005
rect 26295 81195 26505 81405
rect 26895 81195 27105 81405
rect 26295 80610 26505 80820
rect 27495 80610 27705 80820
rect 28095 80610 28305 80820
rect 28695 80610 28905 80820
rect 32295 83280 32505 83490
rect 31695 82995 31905 83205
rect 30195 81495 30405 81705
rect 30195 80610 30405 80820
rect 30795 80610 31005 80820
rect 22095 78795 22305 79005
rect 23595 78795 23805 79005
rect 22395 78495 22605 78705
rect 20895 77595 21105 77805
rect 20595 77295 20805 77505
rect 21795 77295 22005 77505
rect 20295 76695 20505 76905
rect 19395 76395 19605 76605
rect 19995 76395 20205 76605
rect 22095 76395 22305 76605
rect 21195 76110 21405 76320
rect 21795 76110 22005 76320
rect 20295 75480 20505 75690
rect 18195 75195 18405 75405
rect 18795 75195 19005 75405
rect 19395 75195 19605 75405
rect 19995 75195 20205 75405
rect 17595 74595 17805 74805
rect 16695 72795 16905 73005
rect 16995 72810 17205 73020
rect 17895 72795 18105 73005
rect 17295 72180 17505 72390
rect 16395 71295 16605 71505
rect 17895 70395 18105 70605
rect 19095 73995 19305 74205
rect 19695 73695 19905 73905
rect 19695 72795 19905 73005
rect 18795 71595 19005 71805
rect 22095 75195 22305 75405
rect 21795 73995 22005 74205
rect 20295 72810 20505 73020
rect 21195 72810 21405 73020
rect 19995 71895 20205 72105
rect 21795 71895 22005 72105
rect 20895 71595 21105 71805
rect 20295 70995 20505 71205
rect 20295 70680 20505 70890
rect 20895 70695 21105 70905
rect 19395 70395 19605 70605
rect 18195 69795 18405 70005
rect 19395 69795 19605 70005
rect 17295 69495 17505 69705
rect 16095 68895 16305 69105
rect 15495 68295 15705 68505
rect 16995 68595 17205 68805
rect 14595 66195 14805 66405
rect 15495 67695 15705 67905
rect 13095 65895 13305 66105
rect 14295 65895 14505 66105
rect 14895 65895 15105 66105
rect 12795 65595 13005 65805
rect 11895 65295 12105 65505
rect 11595 64095 11805 64305
rect 10695 63495 10905 63705
rect 11295 63495 11505 63705
rect 11595 62895 11805 63105
rect 10395 61995 10605 62205
rect 7395 61095 7605 61305
rect 11295 61095 11505 61305
rect 7395 60510 7605 60720
rect 7995 60510 8205 60720
rect 8595 60510 8805 60720
rect 10095 60510 10305 60720
rect 7095 59295 7305 59505
rect 8295 59880 8505 60090
rect 7695 59595 7905 59805
rect 6195 58995 6405 59205
rect 7395 58995 7605 59205
rect 5595 58095 5805 58305
rect 7695 58095 7905 58305
rect 6195 57495 6405 57705
rect 4395 57195 4605 57405
rect 5295 57195 5505 57405
rect 3795 56580 4005 56790
rect 4695 55995 4905 56205
rect 4995 54195 5205 54405
rect 4095 53595 4305 53805
rect 3495 52695 3705 52905
rect 795 52065 1005 52275
rect 1095 52095 1305 52305
rect 495 51495 705 51705
rect 1395 52065 1605 52275
rect 2295 51795 2505 52005
rect 1695 50895 1905 51105
rect 495 49395 705 49605
rect 1095 49410 1305 49620
rect 2295 49395 2505 49605
rect 1395 48780 1605 48990
rect 1995 48195 2205 48405
rect 3495 51795 3705 52005
rect 2895 49695 3105 49905
rect 3495 49695 3705 49905
rect 8895 57495 9105 57705
rect 9495 57495 9705 57705
rect 8595 57210 8805 57420
rect 5895 56580 6105 56790
rect 5595 56295 5805 56505
rect 5295 53595 5505 53805
rect 7695 56580 7905 56790
rect 8295 56580 8505 56790
rect 9195 56595 9405 56805
rect 8895 55695 9105 55905
rect 6495 54195 6705 54405
rect 6495 52710 6705 52920
rect 7395 52710 7605 52920
rect 7995 52995 8205 53205
rect 9195 52995 9405 53205
rect 10695 59595 10905 59805
rect 10095 59295 10305 59505
rect 10395 58995 10605 59205
rect 10095 58695 10305 58905
rect 9795 57195 10005 57405
rect 16395 67680 16605 67890
rect 15795 67095 16005 67305
rect 18195 68595 18405 68805
rect 18795 68310 19005 68520
rect 19695 68310 19905 68520
rect 20895 69495 21105 69705
rect 22995 77895 23205 78105
rect 22995 76395 23205 76605
rect 24795 78495 25005 78705
rect 24195 77295 24405 77505
rect 24195 76110 24405 76320
rect 24795 76110 25005 76320
rect 23895 75480 24105 75690
rect 23595 74895 23805 75105
rect 23295 73395 23505 73605
rect 23895 74595 24105 74805
rect 26895 79695 27105 79905
rect 26595 78795 26805 79005
rect 26295 76695 26505 76905
rect 26295 76110 26505 76320
rect 25095 74895 25305 75105
rect 24795 73695 25005 73905
rect 25995 75480 26205 75690
rect 26595 75495 26805 75705
rect 26295 74895 26505 75105
rect 25995 74295 26205 74505
rect 25695 73995 25905 74205
rect 25395 73395 25605 73605
rect 23895 72795 24105 73005
rect 24795 72810 25005 73020
rect 22995 72180 23205 72390
rect 24495 71595 24705 71805
rect 23295 71295 23505 71505
rect 23895 71295 24105 71505
rect 22395 70095 22605 70305
rect 25695 72195 25905 72405
rect 24195 70095 24405 70305
rect 25095 70095 25305 70305
rect 23895 69495 24105 69705
rect 22695 68310 22905 68520
rect 23295 68310 23505 68520
rect 17580 67680 17790 67890
rect 17895 67680 18105 67890
rect 18495 67680 18705 67890
rect 17295 66795 17505 67005
rect 18495 67095 18705 67305
rect 17595 66495 17805 66705
rect 16680 66195 16890 66405
rect 16995 66195 17205 66405
rect 16395 65295 16605 65505
rect 12195 64380 12405 64590
rect 15195 64380 15405 64590
rect 15795 64380 16005 64590
rect 16395 64380 16605 64590
rect 13995 64095 14205 64305
rect 11895 62595 12105 62805
rect 13695 62595 13905 62805
rect 13395 61995 13605 62205
rect 11595 60195 11805 60405
rect 12195 58995 12405 59205
rect 11295 58395 11505 58605
rect 10995 57195 11205 57405
rect 13095 58995 13305 59205
rect 12795 58695 13005 58905
rect 12495 58095 12705 58305
rect 12195 57495 12405 57705
rect 10095 56580 10305 56790
rect 10695 56580 10905 56790
rect 11295 56580 11505 56790
rect 10095 55695 10305 55905
rect 10395 54795 10605 55005
rect 10095 53295 10305 53505
rect 9495 52710 9705 52920
rect 10095 52695 10305 52905
rect 5295 52080 5505 52290
rect 6495 52095 6705 52305
rect 5595 50295 5805 50505
rect 7695 52080 7905 52290
rect 10095 52095 10305 52305
rect 8895 51495 9105 51705
rect 9795 51795 10005 52005
rect 6195 49995 6405 50205
rect 4095 49410 4305 49620
rect 5595 49410 5805 49620
rect 7995 50295 8205 50505
rect 7095 49995 7305 50205
rect 6795 49095 7005 49305
rect 2895 48195 3105 48405
rect 2595 46695 2805 46905
rect 1995 44910 2205 45120
rect 2595 44910 2805 45120
rect 495 44280 705 44490
rect 1095 44280 1305 44490
rect 1695 44280 1905 44490
rect 1995 43395 2205 43605
rect 795 41595 1005 41805
rect 1395 41610 1605 41820
rect 2595 42195 2805 42405
rect 195 40095 405 40305
rect 2295 40980 2505 41190
rect 4395 48780 4605 48990
rect 5295 48780 5505 48990
rect 5895 48780 6105 48990
rect 3795 48195 4005 48405
rect 4695 47295 4905 47505
rect 3195 44910 3405 45120
rect 4095 44910 4305 45120
rect 8595 49410 8805 49620
rect 11295 53895 11505 54105
rect 11895 56580 12105 56790
rect 12795 56595 13005 56805
rect 12495 55995 12705 56205
rect 11595 53295 11805 53505
rect 10995 52710 11205 52920
rect 12495 52710 12705 52920
rect 9495 51195 9705 51405
rect 10380 51195 10590 51405
rect 10695 51195 10905 51405
rect 9195 49995 9405 50205
rect 8295 48780 8505 48990
rect 9195 48780 9405 48990
rect 11895 52080 12105 52290
rect 12495 52095 12705 52305
rect 13395 57795 13605 58005
rect 16095 63495 16305 63705
rect 19695 67695 19905 67905
rect 20595 67680 20805 67890
rect 22095 67695 22305 67905
rect 19680 66495 19890 66705
rect 19995 66495 20205 66705
rect 17295 65295 17505 65505
rect 17895 65295 18105 65505
rect 17595 65010 17805 65220
rect 17295 63795 17505 64005
rect 16995 63195 17205 63405
rect 16695 62595 16905 62805
rect 16395 61995 16605 62205
rect 16095 61395 16305 61605
rect 14295 60180 14505 60390
rect 15195 59595 15405 59805
rect 14895 58995 15105 59205
rect 13695 57195 13905 57405
rect 14295 57210 14505 57420
rect 18195 64395 18405 64605
rect 17895 62895 18105 63105
rect 19995 65295 20205 65505
rect 22095 67095 22305 67305
rect 21795 66795 22005 67005
rect 22995 67680 23205 67890
rect 21195 66495 21405 66705
rect 22395 65595 22605 65805
rect 23595 65595 23805 65805
rect 19095 64695 19305 64905
rect 20880 64695 21090 64905
rect 21195 64695 21405 64905
rect 18495 63495 18705 63705
rect 19695 64095 19905 64305
rect 19395 62895 19605 63105
rect 18195 61995 18405 62205
rect 18795 61395 19005 61605
rect 17895 60510 18105 60720
rect 15495 58395 15705 58605
rect 16695 58395 16905 58605
rect 13395 56580 13605 56790
rect 13995 56580 14205 56790
rect 13395 55695 13605 55905
rect 13095 54795 13305 55005
rect 12795 51795 13005 52005
rect 17895 58995 18105 59205
rect 17595 58395 17805 58605
rect 17295 57795 17505 58005
rect 16395 57210 16605 57420
rect 16995 57210 17205 57420
rect 15795 56595 16005 56805
rect 16695 56295 16905 56505
rect 17595 56295 17805 56505
rect 15495 55695 15705 55905
rect 14895 55095 15105 55305
rect 14295 53895 14505 54105
rect 14295 53295 14505 53505
rect 13695 52710 13905 52920
rect 16095 53895 16305 54105
rect 15195 53295 15405 53505
rect 14895 52695 15105 52905
rect 13395 52095 13605 52305
rect 13095 51495 13305 51705
rect 13995 52080 14205 52290
rect 14595 51795 14805 52005
rect 13695 51495 13905 51705
rect 13395 51195 13605 51405
rect 11295 50895 11505 51105
rect 12795 50895 13005 51105
rect 11295 50295 11505 50505
rect 10695 49995 10905 50205
rect 10695 49410 10905 49620
rect 11595 49410 11805 49620
rect 12195 49410 12405 49620
rect 8895 48195 9105 48405
rect 7095 47595 7305 47805
rect 6495 47295 6705 47505
rect 5895 46695 6105 46905
rect 5295 45195 5505 45405
rect 4395 44280 4605 44490
rect 4095 43395 4305 43605
rect 3195 42795 3405 43005
rect 3795 42795 4005 43005
rect 4995 42195 5205 42405
rect 3195 41595 3405 41805
rect 4395 41610 4605 41820
rect 1695 40695 1905 40905
rect 2295 40095 2505 40305
rect 795 38895 1005 39105
rect 195 38595 405 38805
rect 495 37695 705 37905
rect 1095 37110 1305 37320
rect 1995 37110 2205 37320
rect 795 36195 1005 36405
rect 495 35595 705 35805
rect 495 33795 705 34005
rect 495 31395 705 31605
rect 495 27795 705 28005
rect 1695 36495 1905 36705
rect 1395 35595 1605 35805
rect 3495 40980 3705 41190
rect 3195 39495 3405 39705
rect 4695 40695 4905 40905
rect 4395 40095 4605 40305
rect 4095 38295 4305 38505
rect 3795 37995 4005 38205
rect 3195 37695 3405 37905
rect 3795 37110 4005 37320
rect 2580 36195 2790 36405
rect 2895 36195 3105 36405
rect 1095 34995 1305 35205
rect 1695 34995 1905 35205
rect 2895 34995 3105 35205
rect 1695 34395 1905 34605
rect 2295 33810 2505 34020
rect 1395 33180 1605 33390
rect 1095 32895 1305 33105
rect 1095 31095 1305 31305
rect 3795 35595 4005 35805
rect 4395 35595 4605 35805
rect 4395 34995 4605 35205
rect 3795 34395 4005 34605
rect 4095 34095 4305 34305
rect 3495 33810 3705 34020
rect 7395 45795 7605 46005
rect 8895 45195 9105 45405
rect 7695 44910 7905 45120
rect 8295 44910 8505 45120
rect 6195 44280 6405 44490
rect 6795 44280 7005 44490
rect 7395 44295 7605 44505
rect 5895 43095 6105 43305
rect 9495 44895 9705 45105
rect 8595 44280 8805 44490
rect 9495 43995 9705 44205
rect 9195 43695 9405 43905
rect 8595 43395 8805 43605
rect 7695 42795 7905 43005
rect 8295 42495 8505 42705
rect 7395 42195 7605 42405
rect 6495 41610 6705 41820
rect 8295 41610 8505 41820
rect 8895 41610 9105 41820
rect 6195 40980 6405 41190
rect 7395 40980 7605 41190
rect 5295 40695 5505 40905
rect 8595 40980 8805 41190
rect 7695 40395 7905 40605
rect 4995 40095 5205 40305
rect 7695 38895 7905 39105
rect 10395 48780 10605 48990
rect 10695 48495 10905 48705
rect 10695 47595 10905 47805
rect 13395 49395 13605 49605
rect 13095 48780 13305 48990
rect 12495 48495 12705 48705
rect 17295 55695 17505 55905
rect 16695 53295 16905 53505
rect 15495 51795 15705 52005
rect 16395 51495 16605 51705
rect 17595 53895 17805 54105
rect 15195 50895 15405 51105
rect 17295 50895 17505 51105
rect 14895 50295 15105 50505
rect 15495 50295 15705 50505
rect 16695 50295 16905 50505
rect 17295 50295 17505 50505
rect 16695 49695 16905 49905
rect 17295 49695 17505 49905
rect 19095 60510 19305 60720
rect 18795 59295 19005 59505
rect 18495 58995 18705 59205
rect 19995 62595 20205 62805
rect 23295 64095 23505 64305
rect 22095 63495 22305 63705
rect 20595 61395 20805 61605
rect 21495 61395 21705 61605
rect 19995 60795 20205 61005
rect 21495 60795 21705 61005
rect 21195 60495 21405 60705
rect 19395 59895 19605 60105
rect 19095 58395 19305 58605
rect 19095 57795 19305 58005
rect 19695 57210 19905 57420
rect 20895 59295 21105 59505
rect 21195 58995 21405 59205
rect 25995 69795 26205 70005
rect 25695 69195 25905 69405
rect 25095 68310 25305 68520
rect 25695 68310 25905 68520
rect 25995 67395 26205 67605
rect 25395 67095 25605 67305
rect 24795 66195 25005 66405
rect 25095 65895 25305 66105
rect 24495 64395 24705 64605
rect 23880 63195 24090 63405
rect 24195 63195 24405 63405
rect 23895 62880 24105 63090
rect 23595 62595 23805 62805
rect 22995 62295 23205 62505
rect 22095 60510 22305 60720
rect 22395 59880 22605 60090
rect 23295 59895 23505 60105
rect 21795 59295 22005 59505
rect 21495 58095 21705 58305
rect 22995 58095 23205 58305
rect 22695 57795 22905 58005
rect 22395 57180 22605 57390
rect 20295 56880 20505 57090
rect 18195 56580 18405 56790
rect 18795 56580 19005 56790
rect 19395 56580 19605 56790
rect 19995 56595 20205 56805
rect 18795 54495 19005 54705
rect 18495 53895 18705 54105
rect 20295 55995 20505 56205
rect 21495 56580 21705 56790
rect 20895 55995 21105 56205
rect 20595 53595 20805 53805
rect 17895 53295 18105 53505
rect 18795 53295 19005 53505
rect 19395 53295 19605 53505
rect 19995 53295 20205 53505
rect 18795 52710 19005 52920
rect 20895 52710 21105 52920
rect 21495 52710 21705 52920
rect 22695 56580 22905 56790
rect 25095 63795 25305 64005
rect 24795 61695 25005 61905
rect 24495 60510 24705 60720
rect 25695 64395 25905 64605
rect 25395 63495 25605 63705
rect 28095 79695 28305 79905
rect 27195 79395 27405 79605
rect 28995 79395 29205 79605
rect 31095 79395 31305 79605
rect 30195 78795 30405 79005
rect 30795 78795 31005 79005
rect 28680 78495 28890 78705
rect 28995 78495 29205 78705
rect 30195 78195 30405 78405
rect 28095 77895 28305 78105
rect 28695 77895 28905 78105
rect 27180 76095 27390 76305
rect 27495 76110 27705 76320
rect 28695 76110 28905 76320
rect 29295 76110 29505 76320
rect 28395 75495 28605 75705
rect 26895 75195 27105 75405
rect 27795 75195 28005 75405
rect 26595 74595 26805 74805
rect 27195 73395 27405 73605
rect 27195 72810 27405 73020
rect 27795 72180 28005 72390
rect 28095 71595 28305 71805
rect 32295 82695 32505 82905
rect 31995 82395 32205 82605
rect 31695 78795 31905 79005
rect 31095 78195 31305 78405
rect 34995 83910 35205 84120
rect 33795 83295 34005 83505
rect 34695 82995 34905 83205
rect 36795 83910 37005 84120
rect 37995 83910 38205 84120
rect 35895 82995 36105 83205
rect 33495 82695 33705 82905
rect 34095 82695 34305 82905
rect 34695 82680 34905 82890
rect 35295 82695 35505 82905
rect 32895 82395 33105 82605
rect 33795 82395 34005 82605
rect 33195 81495 33405 81705
rect 35895 82395 36105 82605
rect 34695 81795 34905 82005
rect 34095 81195 34305 81405
rect 36495 82095 36705 82305
rect 35295 81195 35505 81405
rect 34095 80595 34305 80805
rect 34695 80610 34905 80820
rect 37995 80895 38205 81105
rect 37395 80610 37605 80820
rect 39795 83910 40005 84120
rect 40095 83295 40305 83505
rect 39195 82395 39405 82605
rect 39795 81795 40005 82005
rect 38895 81195 39105 81405
rect 32295 79395 32505 79605
rect 34395 79995 34605 80205
rect 34095 79095 34305 79305
rect 33495 78795 33705 79005
rect 32895 78495 33105 78705
rect 32295 77895 32505 78105
rect 31095 77595 31305 77805
rect 31995 77595 32205 77805
rect 28695 75195 28905 75405
rect 29295 75195 29505 75405
rect 30795 75495 31005 75705
rect 30495 74895 30705 75105
rect 29595 74595 29805 74805
rect 28695 72180 28905 72390
rect 26895 70695 27105 70905
rect 27195 70395 27405 70605
rect 27495 68310 27705 68520
rect 29595 72180 29805 72390
rect 28995 71895 29205 72105
rect 29895 71595 30105 71805
rect 29895 70995 30105 71205
rect 28995 70095 29205 70305
rect 28380 69195 28590 69405
rect 28695 69195 28905 69405
rect 28095 68295 28305 68505
rect 29295 68310 29505 68520
rect 26595 67695 26805 67905
rect 27195 67680 27405 67890
rect 28395 67695 28605 67905
rect 28395 67380 28605 67590
rect 26295 67095 26505 67305
rect 27795 67095 28005 67305
rect 27795 66195 28005 66405
rect 27195 65595 27405 65805
rect 26595 65010 26805 65220
rect 28095 65895 28305 66105
rect 28095 64995 28305 65205
rect 25995 63795 26205 64005
rect 25995 63480 26205 63690
rect 23595 59295 23805 59505
rect 24195 59295 24405 59505
rect 23895 58995 24105 59205
rect 23895 58395 24105 58605
rect 23295 57195 23505 57405
rect 24495 58395 24705 58605
rect 24495 57795 24705 58005
rect 24495 57195 24705 57405
rect 22995 55995 23205 56205
rect 22995 55095 23205 55305
rect 23595 56580 23805 56790
rect 24195 55395 24405 55605
rect 23295 53895 23505 54105
rect 24195 53895 24405 54105
rect 23295 53580 23505 53790
rect 23595 53295 23805 53505
rect 19095 51495 19305 51705
rect 21795 52095 22005 52305
rect 21195 51495 21405 51705
rect 21795 51495 22005 51705
rect 20595 50895 20805 51105
rect 18495 50295 18705 50505
rect 17595 49395 17805 49605
rect 14595 48780 14805 48990
rect 12495 47895 12705 48105
rect 13695 47895 13905 48105
rect 11595 47295 11805 47505
rect 11895 46095 12105 46305
rect 11295 45795 11505 46005
rect 10695 45195 10905 45405
rect 10095 44895 10305 45105
rect 11880 44895 12090 45105
rect 12195 44910 12405 45120
rect 10095 43695 10305 43905
rect 12195 43995 12405 44205
rect 12195 43095 12405 43305
rect 10995 42495 11205 42705
rect 11595 41895 11805 42105
rect 10095 41595 10305 41805
rect 10995 41610 11205 41820
rect 10095 39795 10305 40005
rect 9795 39195 10005 39405
rect 11295 40980 11505 41190
rect 16995 48780 17205 48990
rect 18195 48795 18405 49005
rect 18795 49995 19005 50205
rect 19395 49410 19605 49620
rect 20295 49395 20505 49605
rect 15795 48195 16005 48405
rect 17895 48195 18105 48405
rect 14295 46695 14505 46905
rect 15195 46695 15405 46905
rect 13695 45495 13905 45705
rect 13095 44910 13305 45120
rect 15195 46095 15405 46305
rect 14295 44895 14505 45105
rect 16395 45195 16605 45405
rect 16995 44910 17205 45120
rect 17595 44910 17805 45120
rect 19695 48780 19905 48990
rect 19395 48495 19605 48705
rect 18795 47895 19005 48105
rect 12795 43995 13005 44205
rect 13995 44280 14205 44490
rect 13395 43095 13605 43305
rect 12795 41895 13005 42105
rect 12495 41595 12705 41805
rect 15495 44280 15705 44490
rect 16395 44295 16605 44505
rect 16395 43980 16605 44190
rect 16095 43695 16305 43905
rect 15795 42495 16005 42705
rect 14595 42195 14805 42405
rect 14295 41595 14505 41805
rect 14895 41610 15105 41820
rect 12495 40995 12705 41205
rect 10995 39195 11205 39405
rect 12195 39195 12405 39405
rect 10695 38595 10905 38805
rect 7095 38295 7305 38505
rect 9495 38295 9705 38505
rect 5895 37695 6105 37905
rect 5295 37110 5505 37320
rect 6795 37095 7005 37305
rect 6195 36195 6405 36405
rect 5295 34995 5505 35205
rect 5895 34995 6105 35205
rect 5595 34395 5805 34605
rect 4695 34095 4905 34305
rect 5295 34095 5505 34305
rect 1995 31695 2205 31905
rect 1395 30195 1605 30405
rect 1695 29310 1905 29520
rect 3495 33180 3705 33390
rect 3495 32595 3705 32805
rect 3195 31995 3405 32205
rect 4695 33180 4905 33390
rect 4395 32895 4605 33105
rect 2895 31695 3105 31905
rect 4095 31695 4305 31905
rect 2595 29295 2805 29505
rect 1695 28395 1905 28605
rect 1395 27795 1605 28005
rect 2595 28695 2805 28905
rect 1995 27795 2205 28005
rect 1695 27495 1905 27705
rect 795 26895 1005 27105
rect 795 25995 1005 26205
rect 1695 26010 1905 26220
rect 2295 26010 2505 26220
rect 4995 32595 5205 32805
rect 4395 30795 4605 31005
rect 4395 30195 4605 30405
rect 3795 29310 4005 29520
rect 4395 29310 4605 29520
rect 3195 28695 3405 28905
rect 2895 28395 3105 28605
rect 495 17580 705 17790
rect 495 16395 705 16605
rect 495 15195 705 15405
rect 4695 28695 4905 28905
rect 4095 27495 4305 27705
rect 3495 26895 3705 27105
rect 3795 26595 4005 26805
rect 3195 25995 3405 26205
rect 10695 38280 10905 38490
rect 7695 37110 7905 37320
rect 9495 37110 9705 37320
rect 10095 37110 10305 37320
rect 8595 36795 8805 37005
rect 7095 35595 7305 35805
rect 6795 34095 7005 34305
rect 5895 33795 6105 34005
rect 6495 33810 6705 34020
rect 7995 35595 8205 35805
rect 10395 36495 10605 36705
rect 10095 36195 10305 36405
rect 9195 35595 9405 35805
rect 8595 34995 8805 35205
rect 7695 34095 7905 34305
rect 10095 34095 10305 34305
rect 9195 33810 9405 34020
rect 9795 33795 10005 34005
rect 5595 33180 5805 33390
rect 6195 33180 6405 33390
rect 6495 32895 6705 33105
rect 5895 29595 6105 29805
rect 5295 29295 5505 29505
rect 7695 33180 7905 33390
rect 6795 32295 7005 32505
rect 8295 33180 8505 33390
rect 8895 32595 9105 32805
rect 8895 31695 9105 31905
rect 8895 30795 9105 31005
rect 7995 30195 8205 30405
rect 7395 29595 7605 29805
rect 6495 29310 6705 29520
rect 7995 29310 8205 29520
rect 5295 28695 5505 28905
rect 9195 30195 9405 30405
rect 4995 27795 5205 28005
rect 4695 26295 4905 26505
rect 4395 26010 4605 26220
rect 1995 25380 2205 25590
rect 2895 25380 3105 25590
rect 4095 25380 4305 25590
rect 1395 23595 1605 23805
rect 2295 23295 2505 23505
rect 4995 23295 5205 23505
rect 1695 22695 1905 22905
rect 3195 22695 3405 22905
rect 3795 22395 4005 22605
rect 4695 22395 4905 22605
rect 3495 20880 3705 21090
rect 1995 20295 2205 20505
rect 1695 19695 1905 19905
rect 1395 18495 1605 18705
rect 4995 20880 5205 21090
rect 4695 20295 4905 20505
rect 4695 19980 4905 20190
rect 2895 18795 3105 19005
rect 4095 18795 4305 19005
rect 2295 18210 2505 18420
rect 3795 18210 4005 18420
rect 795 14895 1005 15105
rect 1395 17580 1605 17790
rect 1995 17580 2205 17790
rect 2895 17580 3105 17790
rect 3495 17580 3705 17790
rect 6195 28680 6405 28890
rect 7695 28680 7905 28890
rect 5595 28395 5805 28605
rect 8895 28680 9105 28890
rect 8295 28095 8505 28305
rect 6495 27495 6705 27705
rect 7395 26295 7605 26505
rect 8295 26295 8505 26505
rect 5595 25395 5805 25605
rect 8595 26010 8805 26220
rect 6195 25380 6405 25590
rect 6795 25380 7005 25590
rect 7395 25380 7605 25590
rect 5595 24495 5805 24705
rect 5895 23895 6105 24105
rect 6495 25095 6705 25305
rect 6195 23595 6405 23805
rect 7095 23295 7305 23505
rect 6495 22695 6705 22905
rect 6495 21510 6705 21720
rect 5295 19695 5505 19905
rect 8895 25395 9105 25605
rect 8895 23895 9105 24105
rect 8295 21795 8505 22005
rect 7695 21510 7905 21720
rect 10695 36195 10905 36405
rect 10695 35595 10905 35805
rect 10395 33795 10605 34005
rect 15195 40980 15405 41190
rect 14595 40695 14805 40905
rect 13695 40395 13905 40605
rect 14895 40095 15105 40305
rect 13095 38895 13305 39105
rect 12495 38295 12705 38505
rect 11295 37695 11505 37905
rect 12195 37695 12405 37905
rect 11295 35895 11505 36105
rect 10995 35295 11205 35505
rect 11895 35295 12105 35505
rect 12795 35895 13005 36105
rect 12495 34395 12705 34605
rect 11295 34095 11505 34305
rect 12495 34080 12705 34290
rect 10395 33195 10605 33405
rect 11595 33180 11805 33390
rect 10395 32595 10605 32805
rect 10995 32595 11205 32805
rect 14595 38295 14805 38505
rect 13395 37995 13605 38205
rect 13995 37695 14205 37905
rect 15495 37995 15705 38205
rect 15195 37110 15405 37320
rect 17895 44280 18105 44490
rect 16995 43095 17205 43305
rect 17295 43095 17505 43305
rect 16395 41595 16605 41805
rect 17595 41895 17805 42105
rect 16695 40980 16905 41190
rect 16095 40095 16305 40305
rect 17295 40095 17505 40305
rect 16695 37995 16905 38205
rect 17595 37995 17805 38205
rect 16995 37695 17205 37905
rect 13395 35895 13605 36105
rect 15795 37110 16005 37320
rect 15495 36495 15705 36705
rect 15195 36195 15405 36405
rect 13695 34995 13905 35205
rect 14295 34995 14505 35205
rect 13095 34095 13305 34305
rect 14295 34680 14505 34890
rect 12795 32595 13005 32805
rect 11595 31995 11805 32205
rect 10395 30195 10605 30405
rect 11595 30195 11805 30405
rect 9480 29295 9690 29505
rect 9795 29310 10005 29520
rect 11895 29895 12105 30105
rect 13395 33180 13605 33390
rect 13995 33195 14205 33405
rect 13395 30495 13605 30705
rect 11595 29595 11805 29805
rect 11295 29295 11505 29505
rect 9495 28695 9705 28905
rect 10095 28680 10305 28890
rect 10695 27495 10905 27705
rect 10695 26895 10905 27105
rect 9495 25995 9705 26205
rect 10095 26010 10305 26220
rect 12195 29310 12405 29520
rect 12795 29310 13005 29520
rect 13695 29895 13905 30105
rect 13395 29295 13605 29505
rect 11895 28695 12105 28905
rect 11595 28095 11805 28305
rect 13095 28680 13305 28890
rect 13695 28695 13905 28905
rect 12795 28395 13005 28605
rect 12495 28095 12705 28305
rect 12795 27195 13005 27405
rect 11895 26295 12105 26505
rect 13095 26295 13305 26505
rect 11295 26010 11505 26220
rect 12195 26010 12405 26220
rect 9795 25380 10005 25590
rect 10995 25380 11205 25590
rect 11295 25095 11505 25305
rect 11895 25095 12105 25305
rect 10395 24495 10605 24705
rect 10695 22095 10905 22305
rect 9795 21795 10005 22005
rect 9495 21510 9705 21720
rect 10395 21795 10605 22005
rect 7095 19995 7305 20205
rect 7395 19395 7605 19605
rect 4995 18195 5205 18405
rect 5595 18210 5805 18420
rect 6195 18210 6405 18420
rect 7995 19095 8205 19305
rect 8295 18495 8505 18705
rect 1395 15795 1605 16005
rect 2295 14895 2505 15105
rect 1095 13995 1305 14205
rect 4695 14895 4905 15105
rect 3795 14295 4005 14505
rect 3195 13995 3405 14205
rect 2895 13695 3105 13905
rect 795 12795 1005 13005
rect 795 11295 1005 11505
rect 495 10695 705 10905
rect 2595 13095 2805 13305
rect 1995 12795 2205 13005
rect 1695 10995 1905 11205
rect 1395 10695 1605 10905
rect 3495 13080 3705 13290
rect 4695 13080 4905 13290
rect 4095 11595 4305 11805
rect 2895 10995 3105 11205
rect 2595 10410 2805 10620
rect 795 9780 1005 9990
rect 1395 9780 1605 9990
rect 495 9195 705 9405
rect 1995 9195 2205 9405
rect 1695 7095 1905 7305
rect 2295 6195 2505 6405
rect 5895 16995 6105 17205
rect 7095 17595 7305 17805
rect 6495 16095 6705 16305
rect 5895 15795 6105 16005
rect 6195 15195 6405 15405
rect 5895 13995 6105 14205
rect 5595 13710 5805 13920
rect 5295 13095 5505 13305
rect 7695 17580 7905 17790
rect 9495 18795 9705 19005
rect 10395 20595 10605 20805
rect 10095 20295 10305 20505
rect 10695 20295 10905 20505
rect 10095 19980 10305 20190
rect 9795 18495 10005 18705
rect 13095 25380 13305 25590
rect 12495 23295 12705 23505
rect 12195 22095 12405 22305
rect 13095 21795 13305 22005
rect 12495 20880 12705 21090
rect 13095 20880 13305 21090
rect 13695 26895 13905 27105
rect 15795 36195 16005 36405
rect 15495 34695 15705 34905
rect 17895 37395 18105 37605
rect 18495 43095 18705 43305
rect 20295 47295 20505 47505
rect 19695 44910 19905 45120
rect 19395 43695 19605 43905
rect 20595 45795 20805 46005
rect 20595 44295 20805 44505
rect 19995 43095 20205 43305
rect 18795 42495 19005 42705
rect 19995 42195 20205 42405
rect 19395 41610 19605 41820
rect 19095 39195 19305 39405
rect 19695 38895 19905 39105
rect 23595 52710 23805 52920
rect 22095 50895 22305 51105
rect 21495 49410 21705 49620
rect 22095 49410 22305 49620
rect 23295 52080 23505 52290
rect 25695 61395 25905 61605
rect 25395 58395 25605 58605
rect 25395 57795 25605 58005
rect 25095 57195 25305 57405
rect 27495 64380 27705 64590
rect 28695 67095 28905 67305
rect 28395 63495 28605 63705
rect 26895 61095 27105 61305
rect 29595 66195 29805 66405
rect 31695 76695 31905 76905
rect 32895 77595 33105 77805
rect 32295 76110 32505 76320
rect 34695 79695 34905 79905
rect 34395 78495 34605 78705
rect 32895 74895 33105 75105
rect 34395 75495 34605 75705
rect 31995 74595 32205 74805
rect 33795 74595 34005 74805
rect 34395 74295 34605 74505
rect 31095 73395 31305 73605
rect 32295 73395 32505 73605
rect 31095 72180 31305 72390
rect 31695 71595 31905 71805
rect 31995 71295 32205 71505
rect 31695 70695 31905 70905
rect 31395 70395 31605 70605
rect 30795 68310 31005 68520
rect 36195 79995 36405 80205
rect 36795 79995 37005 80205
rect 34995 79395 35205 79605
rect 36495 79395 36705 79605
rect 34995 78495 35205 78705
rect 35295 76395 35505 76605
rect 35895 76395 36105 76605
rect 34995 75795 35205 76005
rect 37095 79095 37305 79305
rect 38595 79395 38805 79605
rect 38280 78795 38490 79005
rect 38595 78795 38805 79005
rect 37695 77295 37905 77505
rect 39195 80895 39405 81105
rect 40095 80895 40305 81105
rect 41595 87780 41805 87990
rect 45495 91080 45705 91290
rect 46095 91080 46305 91290
rect 44895 90495 45105 90705
rect 44595 88695 44805 88905
rect 48195 91080 48405 91290
rect 45495 88410 45705 88620
rect 44895 88095 45105 88305
rect 43095 87780 43305 87990
rect 40995 86895 41205 87105
rect 42795 86895 43005 87105
rect 42495 85695 42705 85905
rect 41295 84495 41505 84705
rect 40995 83895 41205 84105
rect 41895 83910 42105 84120
rect 41595 83280 41805 83490
rect 41895 82995 42105 83205
rect 40695 81195 40905 81405
rect 40695 80610 40905 80820
rect 41295 80610 41505 80820
rect 42795 85395 43005 85605
rect 43695 87195 43905 87405
rect 47295 88695 47505 88905
rect 47895 88410 48105 88620
rect 46995 87780 47205 87990
rect 47595 87780 47805 87990
rect 45795 86295 46005 86505
rect 46395 86295 46605 86505
rect 43695 85395 43905 85605
rect 45195 85395 45405 85605
rect 44295 83910 44505 84120
rect 44895 83910 45105 84120
rect 43095 82995 43305 83205
rect 44295 82995 44505 83205
rect 43995 82395 44205 82605
rect 43095 81795 43305 82005
rect 42795 81495 43005 81705
rect 39495 79980 39705 80190
rect 40095 79980 40305 80190
rect 39795 79395 40005 79605
rect 39195 78795 39405 79005
rect 39195 77895 39405 78105
rect 38895 77595 39105 77805
rect 37695 76695 37905 76905
rect 38595 76695 38805 76905
rect 38295 76110 38505 76320
rect 40095 77295 40305 77505
rect 42195 79980 42405 80190
rect 43395 80610 43605 80820
rect 46395 84495 46605 84705
rect 46995 84495 47205 84705
rect 45195 82695 45405 82905
rect 45795 82695 46005 82905
rect 44895 81795 45105 82005
rect 45495 81795 45705 82005
rect 45495 80595 45705 80805
rect 41595 79695 41805 79905
rect 41595 78195 41805 78405
rect 40695 77895 40905 78105
rect 41295 77595 41505 77805
rect 39495 76695 39705 76905
rect 40395 76695 40605 76905
rect 39195 76395 39405 76605
rect 39195 76080 39405 76290
rect 36795 75480 37005 75690
rect 35295 75195 35505 75405
rect 36195 75195 36405 75405
rect 36195 74595 36405 74805
rect 35895 73695 36105 73905
rect 35295 73395 35505 73605
rect 33195 72810 33405 73020
rect 34095 72795 34305 73005
rect 32895 72180 33105 72390
rect 33495 72180 33705 72390
rect 34995 73095 35205 73305
rect 36495 73395 36705 73605
rect 34395 72180 34605 72390
rect 33795 70995 34005 71205
rect 32895 70095 33105 70305
rect 32295 68595 32505 68805
rect 31995 68310 32205 68520
rect 31695 67680 31905 67890
rect 29895 65295 30105 65505
rect 25995 60795 26205 61005
rect 28095 60795 28305 61005
rect 28695 60810 28905 61020
rect 29595 64095 29805 64305
rect 29895 63195 30105 63405
rect 29595 62895 29805 63105
rect 27195 60510 27405 60720
rect 26895 59880 27105 60090
rect 26595 59595 26805 59805
rect 26895 59295 27105 59505
rect 27495 59295 27705 59505
rect 26595 58995 26805 59205
rect 26295 58695 26505 58905
rect 26295 58095 26505 58305
rect 25995 57795 26205 58005
rect 25695 57495 25905 57705
rect 28695 60495 28905 60705
rect 28395 59880 28605 60090
rect 29595 60510 29805 60720
rect 31095 67095 31305 67305
rect 32595 67695 32805 67905
rect 33195 68595 33405 68805
rect 32895 67395 33105 67605
rect 32580 67095 32790 67305
rect 32895 67080 33105 67290
rect 32295 66795 32505 67005
rect 31995 65895 32205 66105
rect 31095 64095 31305 64305
rect 31395 63495 31605 63705
rect 30795 61695 31005 61905
rect 27795 58995 28005 59205
rect 28395 58095 28605 58305
rect 27795 57795 28005 58005
rect 26595 57195 26805 57405
rect 28695 57795 28905 58005
rect 28395 57195 28605 57405
rect 25095 56580 25305 56790
rect 25695 56580 25905 56790
rect 26595 56595 26805 56805
rect 25395 56265 25605 56475
rect 25095 55995 25305 56205
rect 26295 55980 26505 56190
rect 24795 54795 25005 55005
rect 25695 54795 25905 55005
rect 24795 54480 25005 54690
rect 25995 54195 26205 54405
rect 27495 56580 27705 56790
rect 30795 60510 31005 60720
rect 32895 63495 33105 63705
rect 31695 61695 31905 61905
rect 29595 59295 29805 59505
rect 31395 59895 31605 60105
rect 30495 58995 30705 59205
rect 30195 57795 30405 58005
rect 28995 57180 29205 57390
rect 29595 57210 29805 57420
rect 26895 55995 27105 56205
rect 27495 55995 27705 56205
rect 26595 55695 26805 55905
rect 28695 56295 28905 56505
rect 26895 55395 27105 55605
rect 27495 55395 27705 55605
rect 27195 55095 27405 55305
rect 26295 53895 26505 54105
rect 25995 53595 26205 53805
rect 25695 52995 25905 53205
rect 25095 52710 25305 52920
rect 22995 50595 23205 50805
rect 24195 50595 24405 50805
rect 22695 49395 22905 49605
rect 21195 46995 21405 47205
rect 22395 48780 22605 48990
rect 22395 47895 22605 48105
rect 21795 46695 22005 46905
rect 21795 44910 22005 45120
rect 22395 44910 22605 45120
rect 21495 44280 21705 44490
rect 22695 44295 22905 44505
rect 20895 43695 21105 43905
rect 22095 43695 22305 43905
rect 22395 41895 22605 42105
rect 23295 49995 23505 50205
rect 24195 49995 24405 50205
rect 23595 48780 23805 48990
rect 24795 52080 25005 52290
rect 26595 52710 26805 52920
rect 28095 54795 28305 55005
rect 27795 53295 28005 53505
rect 25995 52395 26205 52605
rect 25695 51795 25905 52005
rect 26595 51795 26805 52005
rect 24795 51495 25005 51705
rect 25995 51495 26205 51705
rect 26295 49995 26505 50205
rect 24795 49695 25005 49905
rect 25695 49695 25905 49905
rect 24795 49380 25005 49590
rect 27495 52080 27705 52290
rect 26895 51495 27105 51705
rect 26895 49695 27105 49905
rect 26595 49395 26805 49605
rect 25095 48795 25305 49005
rect 24795 47895 25005 48105
rect 25095 47595 25305 47805
rect 25695 48195 25905 48405
rect 24495 46995 24705 47205
rect 25395 46995 25605 47205
rect 26595 48795 26805 49005
rect 25995 47895 26205 48105
rect 25695 46695 25905 46905
rect 25095 46395 25305 46605
rect 24195 46095 24405 46305
rect 26295 46095 26505 46305
rect 25080 45795 25290 46005
rect 25395 45795 25605 46005
rect 24195 45495 24405 45705
rect 25905 45195 26115 45405
rect 25395 44895 25605 45105
rect 26895 47895 27105 48105
rect 26595 45795 26805 46005
rect 28395 53895 28605 54105
rect 29895 56580 30105 56790
rect 30495 56295 30705 56505
rect 29295 55395 29505 55605
rect 29595 54495 29805 54705
rect 29295 54195 29505 54405
rect 28695 53595 28905 53805
rect 28395 52695 28605 52905
rect 31395 59295 31605 59505
rect 31395 56295 31605 56505
rect 31995 60795 32205 61005
rect 32595 61695 32805 61905
rect 36195 72195 36405 72405
rect 35595 71895 35805 72105
rect 35895 70995 36105 71205
rect 35295 70395 35505 70605
rect 34995 69795 35205 70005
rect 34395 69195 34605 69405
rect 34395 67095 34605 67305
rect 34395 66195 34605 66405
rect 33795 61995 34005 62205
rect 33795 61680 34005 61890
rect 33195 60795 33405 61005
rect 32295 60510 32505 60720
rect 33195 60480 33405 60690
rect 36495 70695 36705 70905
rect 36195 70395 36405 70605
rect 35895 69795 36105 70005
rect 36495 69195 36705 69405
rect 35595 68895 35805 69105
rect 35295 68310 35505 68520
rect 37395 75480 37605 75690
rect 38595 75480 38805 75690
rect 37095 73695 37305 73905
rect 37680 73695 37890 73905
rect 37995 73695 38205 73905
rect 38895 73695 39105 73905
rect 39195 73395 39405 73605
rect 38895 73095 39105 73305
rect 39195 71895 39405 72105
rect 37995 71295 38205 71505
rect 37995 68895 38205 69105
rect 39195 68895 39405 69105
rect 36795 67995 37005 68205
rect 35295 67395 35505 67605
rect 36795 66795 37005 67005
rect 37095 66495 37305 66705
rect 36495 66195 36705 66405
rect 37395 66195 37605 66405
rect 37995 66195 38205 66405
rect 36195 65895 36405 66105
rect 36795 65595 37005 65805
rect 36495 65295 36705 65505
rect 35295 64995 35505 65205
rect 36195 64995 36405 65205
rect 40395 76110 40605 76320
rect 40695 75480 40905 75690
rect 42795 79980 43005 80190
rect 43095 79995 43305 80205
rect 44295 79995 44505 80205
rect 43095 79095 43305 79305
rect 42495 76395 42705 76605
rect 42195 76110 42405 76320
rect 43695 79695 43905 79905
rect 43395 78795 43605 79005
rect 43995 78795 44205 79005
rect 43695 77895 43905 78105
rect 42195 75195 42405 75405
rect 41895 73395 42105 73605
rect 41295 72795 41505 73005
rect 40095 72180 40305 72390
rect 40695 72180 40905 72390
rect 40395 69795 40605 70005
rect 39795 68895 40005 69105
rect 41295 72180 41505 72390
rect 40995 69495 41205 69705
rect 39795 66495 40005 66705
rect 40395 66495 40605 66705
rect 39495 65895 39705 66105
rect 35595 63195 35805 63405
rect 34395 61095 34605 61305
rect 34995 61095 35205 61305
rect 34995 60510 35205 60720
rect 31995 59295 32205 59505
rect 32595 58095 32805 58305
rect 33495 58695 33705 58905
rect 33195 57495 33405 57705
rect 35295 59895 35505 60105
rect 34095 58095 34305 58305
rect 33795 57495 34005 57705
rect 32895 57195 33105 57405
rect 33495 57195 33705 57405
rect 32880 56580 33090 56790
rect 33195 56580 33405 56790
rect 32295 56295 32505 56505
rect 31380 55695 31590 55905
rect 31695 55695 31905 55905
rect 30495 52695 30705 52905
rect 33195 56265 33405 56475
rect 31995 55395 32205 55605
rect 32295 54795 32505 55005
rect 27495 51495 27705 51705
rect 28095 51495 28305 51705
rect 29295 52080 29505 52290
rect 28995 51195 29205 51405
rect 28395 50595 28605 50805
rect 28095 50295 28305 50505
rect 27495 49395 27705 49605
rect 28695 49410 28905 49620
rect 30795 51795 31005 52005
rect 30495 51195 30705 51405
rect 30195 50895 30405 51105
rect 29895 50595 30105 50805
rect 30195 50295 30405 50505
rect 30195 49980 30405 50190
rect 31995 52095 32205 52305
rect 31695 51795 31905 52005
rect 31995 51495 32205 51705
rect 31095 50895 31305 51105
rect 32895 53595 33105 53805
rect 36195 64395 36405 64605
rect 40095 65895 40305 66105
rect 40995 66195 41205 66405
rect 40695 65895 40905 66105
rect 40395 65295 40605 65505
rect 40995 65595 41205 65805
rect 43695 75495 43905 75705
rect 45495 79995 45705 80205
rect 45195 78495 45405 78705
rect 47895 87195 48105 87405
rect 47595 83910 47805 84120
rect 48495 86895 48705 87105
rect 48495 86295 48705 86505
rect 48495 85095 48705 85305
rect 50595 92595 50805 92805
rect 49395 91995 49605 92205
rect 49995 91995 50205 92205
rect 51795 91710 52005 91920
rect 52395 91710 52605 91920
rect 55695 92295 55905 92505
rect 57195 92295 57405 92505
rect 53595 91710 53805 91920
rect 54195 91710 54405 91920
rect 54795 91710 55005 91920
rect 49395 91095 49605 91305
rect 50895 90495 51105 90705
rect 51795 90495 52005 90705
rect 52395 89595 52605 89805
rect 49095 88995 49305 89205
rect 50295 88995 50505 89205
rect 49995 88410 50205 88620
rect 50595 88410 50805 88620
rect 51795 88410 52005 88620
rect 53295 89895 53505 90105
rect 52695 88695 52905 88905
rect 55095 91080 55305 91290
rect 56595 91710 56805 91920
rect 54495 90495 54705 90705
rect 55695 90495 55905 90705
rect 56595 90195 56805 90405
rect 53595 89595 53805 89805
rect 56295 89595 56505 89805
rect 54195 88695 54405 88905
rect 55095 88695 55305 88905
rect 55395 88395 55605 88605
rect 56895 89895 57105 90105
rect 55095 88095 55305 88305
rect 49695 87780 49905 87990
rect 50295 87780 50505 87990
rect 50295 87465 50505 87675
rect 49095 86595 49305 86805
rect 49995 85995 50205 86205
rect 48795 84495 49005 84705
rect 50895 87195 51105 87405
rect 51195 86895 51405 87105
rect 50595 85695 50805 85905
rect 50295 84795 50505 85005
rect 49095 83895 49305 84105
rect 49995 83910 50205 84120
rect 48195 83280 48405 83490
rect 47595 82395 47805 82605
rect 46995 82095 47205 82305
rect 46095 81795 46305 82005
rect 48495 82095 48705 82305
rect 48195 81495 48405 81705
rect 47895 81195 48105 81405
rect 46995 80895 47205 81105
rect 47595 80895 47805 81105
rect 47295 79980 47505 80190
rect 47895 79995 48105 80205
rect 46395 79095 46605 79305
rect 48195 79095 48405 79305
rect 47595 78495 47805 78705
rect 48195 78495 48405 78705
rect 45795 78195 46005 78405
rect 44595 77595 44805 77805
rect 45195 77595 45405 77805
rect 44595 77280 44805 77490
rect 44595 76110 44805 76320
rect 45195 76110 45405 76320
rect 43995 74595 44205 74805
rect 42495 74295 42705 74505
rect 42495 73395 42705 73605
rect 42495 72810 42705 73020
rect 43095 72810 43305 73020
rect 41895 72195 42105 72405
rect 42795 72180 43005 72390
rect 43395 70995 43605 71205
rect 43095 69495 43305 69705
rect 42195 68310 42405 68520
rect 42495 67680 42705 67890
rect 42195 67395 42405 67605
rect 41895 66495 42105 66705
rect 41595 65895 41805 66105
rect 41895 65595 42105 65805
rect 41295 65010 41505 65220
rect 41895 64995 42105 65205
rect 43695 70395 43905 70605
rect 44895 75480 45105 75690
rect 46695 77295 46905 77505
rect 47295 77295 47505 77505
rect 45795 75195 46005 75405
rect 44295 74295 44505 74505
rect 45795 74295 46005 74505
rect 44895 73395 45105 73605
rect 45795 73395 46005 73605
rect 45495 72810 45705 73020
rect 44595 71895 44805 72105
rect 43995 69495 44205 69705
rect 43995 68895 44205 69105
rect 44295 68595 44505 68805
rect 43395 68295 43605 68505
rect 45495 71895 45705 72105
rect 45195 70695 45405 70905
rect 45495 70395 45705 70605
rect 45195 68595 45405 68805
rect 43095 66795 43305 67005
rect 43695 67680 43905 67890
rect 44295 67680 44505 67890
rect 45195 67680 45405 67890
rect 43695 67095 43905 67305
rect 46395 75480 46605 75690
rect 47595 75480 47805 75690
rect 47595 73995 47805 74205
rect 46995 73695 47205 73905
rect 49695 83280 49905 83490
rect 49995 82695 50205 82905
rect 49095 81495 49305 81705
rect 49395 80895 49605 81105
rect 50295 82095 50505 82305
rect 50895 82095 51105 82305
rect 50295 81780 50505 81990
rect 49995 80595 50205 80805
rect 48795 79995 49005 80205
rect 49695 79980 49905 80190
rect 49995 78495 50205 78705
rect 48795 77895 49005 78105
rect 49095 76995 49305 77205
rect 49395 76110 49605 76320
rect 50595 80895 50805 81105
rect 52695 87780 52905 87990
rect 53295 87795 53505 88005
rect 53295 87195 53505 87405
rect 52095 86595 52305 86805
rect 51495 84795 51705 85005
rect 52695 84795 52905 85005
rect 52095 83910 52305 84120
rect 54495 87780 54705 87990
rect 55395 87780 55605 87990
rect 53895 86595 54105 86805
rect 53895 86280 54105 86490
rect 53295 83910 53505 84120
rect 51495 82995 51705 83205
rect 51195 80895 51405 81105
rect 52080 82395 52290 82605
rect 52395 82395 52605 82605
rect 52395 82080 52605 82290
rect 53595 83295 53805 83505
rect 53295 82995 53505 83205
rect 52995 81795 53205 82005
rect 52995 81195 53205 81405
rect 52395 80895 52605 81105
rect 52995 80595 53205 80805
rect 53595 82095 53805 82305
rect 53895 81795 54105 82005
rect 54795 86595 55005 86805
rect 56895 87780 57105 87990
rect 55395 85695 55605 85905
rect 55095 84795 55305 85005
rect 55395 83910 55605 84120
rect 54495 83295 54705 83505
rect 55095 83280 55305 83490
rect 54795 82695 55005 82905
rect 54495 82380 54705 82590
rect 54495 81495 54705 81705
rect 53895 80610 54105 80820
rect 50595 79995 50805 80205
rect 50295 78195 50505 78405
rect 49095 75480 49305 75690
rect 50295 75480 50505 75690
rect 49695 75195 49905 75405
rect 48195 74295 48405 74505
rect 47895 73395 48105 73605
rect 47295 72810 47505 73020
rect 46095 69795 46305 70005
rect 46395 68895 46605 69105
rect 46395 68295 46605 68505
rect 47895 72180 48105 72390
rect 47595 71895 47805 72105
rect 48495 72795 48705 73005
rect 47295 68295 47505 68505
rect 46095 67680 46305 67890
rect 46995 67395 47205 67605
rect 43995 66495 44205 66705
rect 45495 66495 45705 66705
rect 43695 65595 43905 65805
rect 43395 64995 43605 65205
rect 40395 64395 40605 64605
rect 39795 64095 40005 64305
rect 37395 63795 37605 64005
rect 36495 61995 36705 62205
rect 37095 61395 37305 61605
rect 37095 60795 37305 61005
rect 34980 57195 35190 57405
rect 35295 57210 35505 57420
rect 34095 56595 34305 56805
rect 34680 56580 34890 56790
rect 34995 56595 35205 56805
rect 35595 56295 35805 56505
rect 34395 55995 34605 56205
rect 34995 55995 35205 56205
rect 34095 53595 34305 53805
rect 33495 52710 33705 52920
rect 34695 55695 34905 55905
rect 34395 52695 34605 52905
rect 34395 52095 34605 52305
rect 33795 51495 34005 51705
rect 34095 51195 34305 51405
rect 33195 50895 33405 51105
rect 33795 50895 34005 51105
rect 32895 49995 33105 50205
rect 30795 49695 31005 49905
rect 32295 49695 32505 49905
rect 29295 49410 29505 49620
rect 30195 49410 30405 49620
rect 31995 49410 32205 49620
rect 27495 48795 27705 49005
rect 27195 45195 27405 45405
rect 23595 44295 23805 44505
rect 23295 43995 23505 44205
rect 23295 43095 23505 43305
rect 23295 42195 23505 42405
rect 21495 41610 21705 41820
rect 22995 41595 23205 41805
rect 22395 40980 22605 41190
rect 22995 40995 23205 41205
rect 21795 40395 22005 40605
rect 21195 40095 21405 40305
rect 20895 38595 21105 38805
rect 20595 38295 20805 38505
rect 18795 37395 19005 37605
rect 18495 37095 18705 37305
rect 19695 37110 19905 37320
rect 16395 35895 16605 36105
rect 16995 35895 17205 36105
rect 16695 35595 16905 35805
rect 17295 35595 17505 35805
rect 16080 35295 16290 35505
rect 16395 35295 16605 35505
rect 15195 33810 15405 34020
rect 15795 33810 16005 34020
rect 14595 33195 14805 33405
rect 16095 32595 16305 32805
rect 19995 36480 20205 36690
rect 20595 36495 20805 36705
rect 20595 35895 20805 36105
rect 18495 35595 18705 35805
rect 19995 34995 20205 35205
rect 17595 34695 17805 34905
rect 19095 34695 19305 34905
rect 17295 34395 17505 34605
rect 17895 34395 18105 34605
rect 17595 33810 17805 34020
rect 18195 33810 18405 34020
rect 19995 33810 20205 34020
rect 21195 37695 21405 37905
rect 20895 34995 21105 35205
rect 22395 37395 22605 37605
rect 21195 34695 21405 34905
rect 25395 44295 25605 44505
rect 24495 43995 24705 44205
rect 25095 43395 25305 43605
rect 24495 43095 24705 43305
rect 24195 42795 24405 43005
rect 23895 42195 24105 42405
rect 24795 42495 25005 42705
rect 23595 41595 23805 41805
rect 23595 40995 23805 41205
rect 24195 40980 24405 41190
rect 23295 38595 23505 38805
rect 23595 38295 23805 38505
rect 22695 36195 22905 36405
rect 22095 35295 22305 35505
rect 23295 35295 23505 35505
rect 21795 34995 22005 35205
rect 21495 34095 21705 34305
rect 22395 34095 22605 34305
rect 17295 32595 17505 32805
rect 18495 33180 18705 33390
rect 19095 33180 19305 33390
rect 19695 33180 19905 33390
rect 19695 32595 19905 32805
rect 16695 32295 16905 32505
rect 17895 32295 18105 32505
rect 19095 32295 19305 32505
rect 19695 31695 19905 31905
rect 15495 30795 15705 31005
rect 14895 29895 15105 30105
rect 14295 29310 14505 29520
rect 20595 32895 20805 33105
rect 20295 30495 20505 30705
rect 17295 29595 17505 29805
rect 19695 29595 19905 29805
rect 15495 29310 15705 29520
rect 14595 28680 14805 28890
rect 15195 28680 15405 28890
rect 14295 26895 14505 27105
rect 13995 25995 14205 26205
rect 16695 29310 16905 29520
rect 18495 29310 18705 29520
rect 19095 29310 19305 29520
rect 17595 28680 17805 28890
rect 16095 28095 16305 28305
rect 16995 28095 17205 28305
rect 16095 27195 16305 27405
rect 14895 26010 15105 26220
rect 14595 25380 14805 25590
rect 16395 25380 16605 25590
rect 20295 29295 20505 29505
rect 18795 27195 19005 27405
rect 17295 26595 17505 26805
rect 15195 25095 15405 25305
rect 16995 25095 17205 25305
rect 14895 23895 15105 24105
rect 15495 23895 15705 24105
rect 14895 23295 15105 23505
rect 13695 22095 13905 22305
rect 14295 21795 14505 22005
rect 11895 20295 12105 20505
rect 12795 19395 13005 19605
rect 10695 19095 10905 19305
rect 11295 19095 11505 19305
rect 12195 18795 12405 19005
rect 10995 18195 11205 18405
rect 11595 18210 11805 18420
rect 12795 18195 13005 18405
rect 9195 17580 9405 17790
rect 9795 17580 10005 17790
rect 10695 17580 10905 17790
rect 8295 16995 8505 17205
rect 5295 11595 5505 11805
rect 7095 13080 7305 13290
rect 7995 13080 8205 13290
rect 8595 13080 8805 13290
rect 9795 16995 10005 17205
rect 9495 13995 9705 14205
rect 6495 12495 6705 12705
rect 9195 12495 9405 12705
rect 5895 11295 6105 11505
rect 5895 10410 6105 10620
rect 6495 10410 6705 10620
rect 7395 10395 7605 10605
rect 4695 9780 4905 9990
rect 5295 9780 5505 9990
rect 6195 9495 6405 9705
rect 5295 9195 5505 9405
rect 6795 9195 7005 9405
rect 4095 8595 4305 8805
rect 6195 7395 6405 7605
rect 3795 7095 4005 7305
rect 3195 6195 3405 6405
rect 2895 5895 3105 6105
rect 4695 6195 4905 6405
rect 1995 5280 2205 5490
rect 3495 4695 3705 4905
rect 1395 4095 1605 4305
rect 1995 4095 2205 4305
rect 195 3495 405 3705
rect 1395 3495 1605 3705
rect 7395 6495 7605 6705
rect 7995 11295 8205 11505
rect 8595 11595 8805 11805
rect 8295 10995 8505 11205
rect 7995 10395 8205 10605
rect 9195 10995 9405 11205
rect 9495 10395 9705 10605
rect 8295 9780 8505 9990
rect 8895 9495 9105 9705
rect 8895 8595 9105 8805
rect 8295 7395 8505 7605
rect 7695 5910 7905 6120
rect 9195 6495 9405 6705
rect 6495 5280 6705 5490
rect 4695 4695 4905 4905
rect 5895 4695 6105 4905
rect 4095 3495 4305 3705
rect 3795 3195 4005 3405
rect 8595 5280 8805 5490
rect 7995 4395 8205 4605
rect 7395 4095 7605 4305
rect 6195 3495 6405 3705
rect 5895 2895 6105 3105
rect 4095 2595 4305 2805
rect 4695 2595 4905 2805
rect 5595 2610 5805 2820
rect 6195 2610 6405 2820
rect 7995 3795 8205 4005
rect 1695 1980 1905 2190
rect 2295 1980 2505 2190
rect 3495 1980 3705 2190
rect 5295 1980 5505 2190
rect 5895 1980 6105 2190
rect 7095 1695 7305 1905
rect 9495 5910 9705 6120
rect 9495 5295 9705 5505
rect 10395 13710 10605 13920
rect 11895 17580 12105 17790
rect 12495 17580 12705 17790
rect 14295 20595 14505 20805
rect 13995 20295 14205 20505
rect 13695 18210 13905 18420
rect 15195 19995 15405 20205
rect 14595 18795 14805 19005
rect 13995 17295 14205 17505
rect 13095 16995 13305 17205
rect 12795 16395 13005 16605
rect 12495 16095 12705 16305
rect 12795 15795 13005 16005
rect 11595 14295 11805 14505
rect 12795 13995 13005 14205
rect 13395 13710 13605 13920
rect 11595 13095 11805 13305
rect 14895 17595 15105 17805
rect 12495 13080 12705 13290
rect 13995 13080 14205 13290
rect 12195 12495 12405 12705
rect 13095 12495 13305 12705
rect 11895 11595 12105 11805
rect 10695 11295 10905 11505
rect 11295 10995 11505 11205
rect 10095 10395 10305 10605
rect 14595 15495 14805 15705
rect 16095 22695 16305 22905
rect 15795 22095 16005 22305
rect 15795 20595 16005 20805
rect 18195 26595 18405 26805
rect 19995 28680 20205 28890
rect 22095 33180 22305 33390
rect 22680 33180 22890 33390
rect 22995 33195 23205 33405
rect 21495 32895 21705 33105
rect 20895 32295 21105 32505
rect 20895 31095 21105 31305
rect 21195 30795 21405 31005
rect 20895 29295 21105 29505
rect 21795 30495 22005 30705
rect 22995 31995 23205 32205
rect 25695 43995 25905 44205
rect 25995 43695 26205 43905
rect 27195 43995 27405 44205
rect 28395 48780 28605 48990
rect 27795 46995 28005 47205
rect 27795 46395 28005 46605
rect 28695 46395 28905 46605
rect 28395 45495 28605 45705
rect 29295 46695 29505 46905
rect 28995 45495 29205 45705
rect 28995 44895 29205 45105
rect 27495 43395 27705 43605
rect 28695 44280 28905 44490
rect 29895 48780 30105 48990
rect 30195 48495 30405 48705
rect 30795 48495 31005 48705
rect 31095 48795 31305 49005
rect 31095 48195 31305 48405
rect 30795 47895 31005 48105
rect 30195 47295 30405 47505
rect 29895 45495 30105 45705
rect 29295 43995 29505 44205
rect 28095 43095 28305 43305
rect 26895 41895 27105 42105
rect 26595 41610 26805 41820
rect 27495 41610 27705 41820
rect 25395 40995 25605 41205
rect 26295 40980 26505 41190
rect 26895 40980 27105 41190
rect 25095 40695 25305 40905
rect 25980 40695 26190 40905
rect 24795 40395 25005 40605
rect 24495 39495 24705 39705
rect 25395 38895 25605 39105
rect 24795 38595 25005 38805
rect 23895 37995 24105 38205
rect 24195 37110 24405 37320
rect 25695 37395 25905 37605
rect 25395 37110 25605 37320
rect 24495 36195 24705 36405
rect 25395 36495 25605 36705
rect 23895 35595 24105 35805
rect 25095 35595 25305 35805
rect 25695 36195 25905 36405
rect 27795 41295 28005 41505
rect 27495 40395 27705 40605
rect 28095 40695 28305 40905
rect 27795 39795 28005 40005
rect 27195 38895 27405 39105
rect 27795 38895 28005 39105
rect 26895 38595 27105 38805
rect 27195 38295 27405 38505
rect 26295 37995 26505 38205
rect 27495 37995 27705 38205
rect 27195 37695 27405 37905
rect 26595 37395 26805 37605
rect 26295 37095 26505 37305
rect 27195 37110 27405 37320
rect 26295 36480 26505 36690
rect 25995 35895 26205 36105
rect 25995 35580 26205 35790
rect 24795 34995 25005 35205
rect 25395 34995 25605 35205
rect 25395 34680 25605 34890
rect 24795 34395 25005 34605
rect 24495 34095 24705 34305
rect 27495 36480 27705 36690
rect 26895 36195 27105 36405
rect 28395 40395 28605 40605
rect 28395 39795 28605 40005
rect 28695 38895 28905 39105
rect 30495 45495 30705 45705
rect 30195 44895 30405 45105
rect 31995 48495 32205 48705
rect 31695 47895 31905 48105
rect 31095 45795 31305 46005
rect 32595 48795 32805 49005
rect 32895 48495 33105 48705
rect 32595 47595 32805 47805
rect 32295 47295 32505 47505
rect 34995 55395 35205 55605
rect 34695 50595 34905 50805
rect 33795 50295 34005 50505
rect 40995 63795 41205 64005
rect 39795 63195 40005 63405
rect 40395 63195 40605 63405
rect 37995 62595 38205 62805
rect 38595 62295 38805 62505
rect 39495 61695 39705 61905
rect 39195 60795 39405 61005
rect 40695 62295 40905 62505
rect 40395 61395 40605 61605
rect 40095 61080 40305 61290
rect 39795 60795 40005 61005
rect 39495 60495 39705 60705
rect 38595 59880 38805 60090
rect 37995 58395 38205 58605
rect 39195 58395 39405 58605
rect 39795 58395 40005 58605
rect 38295 57795 38505 58005
rect 37095 57495 37305 57705
rect 37695 57495 37905 57705
rect 36795 57195 37005 57405
rect 39195 57780 39405 57990
rect 38895 57210 39105 57420
rect 39495 57195 39705 57405
rect 35895 55995 36105 56205
rect 36195 55095 36405 55305
rect 35280 54495 35490 54705
rect 35595 54495 35805 54705
rect 35595 53595 35805 53805
rect 35295 52695 35505 52905
rect 37395 56595 37605 56805
rect 36795 56295 37005 56505
rect 36495 54795 36705 55005
rect 36495 53895 36705 54105
rect 36195 52695 36405 52905
rect 35895 52080 36105 52290
rect 34095 49995 34305 50205
rect 34995 49995 35205 50205
rect 33495 48795 33705 49005
rect 33495 47895 33705 48105
rect 34095 47895 34305 48105
rect 34695 47895 34905 48105
rect 33795 47295 34005 47505
rect 33195 46695 33405 46905
rect 31995 46395 32205 46605
rect 31695 44895 31905 45105
rect 31080 44280 31290 44490
rect 31395 44295 31605 44505
rect 30495 43995 30705 44205
rect 30195 43095 30405 43305
rect 29595 41595 29805 41805
rect 30795 42795 31005 43005
rect 30795 42195 31005 42405
rect 29895 40980 30105 41190
rect 30195 40695 30405 40905
rect 30195 40095 30405 40305
rect 29295 37395 29505 37605
rect 28380 37095 28590 37305
rect 28695 37110 28905 37320
rect 29895 36795 30105 37005
rect 28395 36495 28605 36705
rect 28095 35895 28305 36105
rect 27795 35595 28005 35805
rect 27195 34695 27405 34905
rect 26295 34395 26505 34605
rect 26895 34395 27105 34605
rect 25695 33810 25905 34020
rect 26595 33810 26805 34020
rect 28095 34995 28305 35205
rect 27780 34095 27990 34305
rect 28695 36195 28905 36405
rect 29595 36495 29805 36705
rect 28995 35895 29205 36105
rect 29295 35595 29505 35805
rect 28695 34995 28905 35205
rect 28995 34095 29205 34305
rect 23895 32295 24105 32505
rect 24795 33180 25005 33390
rect 28395 33795 28605 34005
rect 29595 35295 29805 35505
rect 30495 39195 30705 39405
rect 31395 42495 31605 42705
rect 31995 44295 32205 44505
rect 32895 46095 33105 46305
rect 32595 45495 32805 45705
rect 34695 47580 34905 47790
rect 34695 46395 34905 46605
rect 35580 50595 35790 50805
rect 35895 50595 36105 50805
rect 36495 50595 36705 50805
rect 37095 54195 37305 54405
rect 38295 56295 38505 56505
rect 37995 55395 38205 55605
rect 37395 53895 37605 54105
rect 38595 55995 38805 56205
rect 39795 56295 40005 56505
rect 39495 54495 39705 54705
rect 38595 52995 38805 53205
rect 38295 52695 38505 52905
rect 41295 60510 41505 60720
rect 42195 64395 42405 64605
rect 41895 64095 42105 64305
rect 40395 59880 40605 60090
rect 40995 59880 41205 60090
rect 41595 59595 41805 59805
rect 41295 58095 41505 58305
rect 40395 57795 40605 58005
rect 40695 57495 40905 57705
rect 40395 57195 40605 57405
rect 43095 62595 43305 62805
rect 42495 61395 42705 61605
rect 42795 61095 43005 61305
rect 42195 60795 42405 61005
rect 42795 60510 43005 60720
rect 43395 62295 43605 62505
rect 41895 57795 42105 58005
rect 41895 57480 42105 57690
rect 42495 59880 42705 60090
rect 43095 59895 43305 60105
rect 43095 59295 43305 59505
rect 45795 66195 46005 66405
rect 43995 64995 44205 65205
rect 44595 64395 44805 64605
rect 45195 63795 45405 64005
rect 44295 62895 44505 63105
rect 45195 62295 45405 62505
rect 43995 60495 44205 60705
rect 43695 59895 43905 60105
rect 43995 58395 44205 58605
rect 43695 58095 43905 58305
rect 43395 57495 43605 57705
rect 42795 57210 43005 57420
rect 40395 56595 40605 56805
rect 39795 53895 40005 54105
rect 38595 52395 38805 52605
rect 37095 52095 37305 52305
rect 36795 50295 37005 50505
rect 35595 49380 35805 49590
rect 36495 49410 36705 49620
rect 37695 51795 37905 52005
rect 38895 52095 39105 52305
rect 38595 51495 38805 51705
rect 37695 50895 37905 51105
rect 37395 49995 37605 50205
rect 37095 49395 37305 49605
rect 35295 47595 35505 47805
rect 35895 48195 36105 48405
rect 36495 48195 36705 48405
rect 35595 46995 35805 47205
rect 36195 46395 36405 46605
rect 34095 45795 34305 46005
rect 34395 45495 34605 45705
rect 33495 44910 33705 45120
rect 35895 45795 36105 46005
rect 34695 45195 34905 45405
rect 34995 44910 35205 45120
rect 32895 43995 33105 44205
rect 32595 43695 32805 43905
rect 32295 43095 32505 43305
rect 32595 42795 32805 43005
rect 31995 42195 32205 42405
rect 34095 44295 34305 44505
rect 33495 43695 33705 43905
rect 33495 43095 33705 43305
rect 33195 42495 33405 42705
rect 32595 41895 32805 42105
rect 31395 41595 31605 41805
rect 31995 41610 32205 41820
rect 31095 38895 31305 39105
rect 30195 36495 30405 36705
rect 30195 35295 30405 35505
rect 30195 34395 30405 34605
rect 30195 34080 30405 34290
rect 29295 33795 29505 34005
rect 26295 32895 26505 33105
rect 26895 32895 27105 33105
rect 24795 32595 25005 32805
rect 25695 32595 25905 32805
rect 24195 31995 24405 32205
rect 24195 31680 24405 31890
rect 23895 31095 24105 31305
rect 22995 30795 23205 31005
rect 23595 30795 23805 31005
rect 22095 29895 22305 30105
rect 25995 32295 26205 32505
rect 25095 31995 25305 32205
rect 24795 30795 25005 31005
rect 23880 30495 24090 30705
rect 24195 30495 24405 30705
rect 22395 29295 22605 29505
rect 22995 29310 23205 29520
rect 25695 31395 25905 31605
rect 24195 29310 24405 29520
rect 25695 29895 25905 30105
rect 25395 29310 25605 29520
rect 19695 28095 19905 28305
rect 20595 28095 20805 28305
rect 19395 25995 19605 26205
rect 17895 25395 18105 25605
rect 17595 22695 17805 22905
rect 16395 22095 16605 22305
rect 17295 22095 17505 22305
rect 16395 21495 16605 21705
rect 18495 25380 18705 25590
rect 19095 24795 19305 25005
rect 20895 26895 21105 27105
rect 19995 26295 20205 26505
rect 22995 28095 23205 28305
rect 21795 26595 22005 26805
rect 22395 26595 22605 26805
rect 21495 26295 21705 26505
rect 19995 25695 20205 25905
rect 21495 25695 21705 25905
rect 20595 24795 20805 25005
rect 21195 23895 21405 24105
rect 19695 22995 19905 23205
rect 18495 22095 18705 22305
rect 19995 22095 20205 22305
rect 20595 22095 20805 22305
rect 17895 21510 18105 21720
rect 19095 21510 19305 21720
rect 16395 20895 16605 21105
rect 15495 19395 15705 19605
rect 15495 18195 15705 18405
rect 15195 17295 15405 17505
rect 14895 14895 15105 15105
rect 16095 19695 16305 19905
rect 17295 20595 17505 20805
rect 18795 20595 19005 20805
rect 16695 19995 16905 20205
rect 18795 19695 19005 19905
rect 16395 19095 16605 19305
rect 16995 19095 17205 19305
rect 17895 19095 18105 19305
rect 16395 18210 16605 18420
rect 16095 17595 16305 17805
rect 15795 17295 16005 17505
rect 15795 14895 16005 15105
rect 15495 13995 15705 14205
rect 15195 13710 15405 13920
rect 19995 20595 20205 20805
rect 20295 19395 20505 19605
rect 19395 18795 19605 19005
rect 19995 18795 20205 19005
rect 19395 18210 19605 18420
rect 17295 17295 17505 17505
rect 19695 17595 19905 17805
rect 19095 16695 19305 16905
rect 16695 16095 16905 16305
rect 19095 16095 19305 16305
rect 17895 14895 18105 15105
rect 16095 14595 16305 14805
rect 18495 14595 18705 14805
rect 16395 13995 16605 14205
rect 17295 13995 17505 14205
rect 14295 12795 14505 13005
rect 13995 11595 14205 11805
rect 12480 10995 12690 11205
rect 12795 10995 13005 11205
rect 12195 10395 12405 10605
rect 10995 9780 11205 9990
rect 10095 9495 10305 9705
rect 11595 9195 11805 9405
rect 12495 8595 12705 8805
rect 11895 7095 12105 7305
rect 10395 5910 10605 6120
rect 10995 5910 11205 6120
rect 15495 12795 15705 13005
rect 19395 14295 19605 14505
rect 22395 26010 22605 26220
rect 23295 27195 23505 27405
rect 23895 27195 24105 27405
rect 23595 26895 23805 27105
rect 23595 25995 23805 26205
rect 23295 25380 23505 25590
rect 22695 24495 22905 24705
rect 24495 28695 24705 28905
rect 24195 26280 24405 26490
rect 24795 27195 25005 27405
rect 24495 25995 24705 26205
rect 27780 33195 27990 33405
rect 28095 33195 28305 33405
rect 27495 31395 27705 31605
rect 27795 29295 28005 29505
rect 25395 28095 25605 28305
rect 26295 28395 26505 28605
rect 25695 27795 25905 28005
rect 25395 27195 25605 27405
rect 25095 26895 25305 27105
rect 25395 26295 25605 26505
rect 26580 27795 26790 28005
rect 26895 27795 27105 28005
rect 26295 25680 26505 25890
rect 24195 24795 24405 25005
rect 23895 23595 24105 23805
rect 22395 22995 22605 23205
rect 21495 22095 21705 22305
rect 22095 22095 22305 22305
rect 25095 25380 25305 25590
rect 25695 25095 25905 25305
rect 23295 22695 23505 22905
rect 24180 22695 24390 22905
rect 24495 22695 24705 22905
rect 22695 22395 22905 22605
rect 22395 21795 22605 22005
rect 23895 22395 24105 22605
rect 21495 20880 21705 21090
rect 22695 20880 22905 21090
rect 21795 20595 22005 20805
rect 24195 20880 24405 21090
rect 23295 20595 23505 20805
rect 23595 20595 23805 20805
rect 23295 19395 23505 19605
rect 22695 18795 22905 19005
rect 21495 18210 21705 18420
rect 24195 18495 24405 18705
rect 24195 17895 24405 18105
rect 20595 17580 20805 17790
rect 21195 17580 21405 17790
rect 20295 17295 20505 17505
rect 22095 17595 22305 17805
rect 21795 17295 22005 17505
rect 22095 16695 22305 16905
rect 21195 16395 21405 16605
rect 22695 16395 22905 16605
rect 19995 15495 20205 15705
rect 24195 16095 24405 16305
rect 20595 14595 20805 14805
rect 19995 14295 20205 14505
rect 19995 13710 20205 13920
rect 20595 13710 20805 13920
rect 16995 13080 17205 13290
rect 16395 11895 16605 12105
rect 17295 11895 17505 12105
rect 16395 10995 16605 11205
rect 13395 10410 13605 10620
rect 13995 10410 14205 10620
rect 14895 10410 15105 10620
rect 15795 10410 16005 10620
rect 13095 9795 13305 10005
rect 13695 9780 13905 9990
rect 16995 10395 17205 10605
rect 13695 8895 13905 9105
rect 14295 8595 14505 8805
rect 16095 8595 16305 8805
rect 13095 7995 13305 8205
rect 12795 6795 13005 7005
rect 18495 13080 18705 13290
rect 19695 13080 19905 13290
rect 17595 10995 17805 11205
rect 18495 10995 18705 11205
rect 19395 10995 19605 11205
rect 19095 10695 19305 10905
rect 17895 10410 18105 10620
rect 18495 10410 18705 10620
rect 23595 14595 23805 14805
rect 23595 13995 23805 14205
rect 22995 13710 23205 13920
rect 24495 15195 24705 15405
rect 24495 14295 24705 14505
rect 27195 27195 27405 27405
rect 27495 26295 27705 26505
rect 28695 33180 28905 33390
rect 29295 33195 29505 33405
rect 29895 33195 30105 33405
rect 28395 32595 28605 32805
rect 29595 31980 29805 32190
rect 28395 31695 28605 31905
rect 31695 40995 31905 41205
rect 32295 40695 32505 40905
rect 32295 39795 32505 40005
rect 31995 38595 32205 38805
rect 31995 37995 32205 38205
rect 31395 37395 31605 37605
rect 31995 37395 32205 37605
rect 32295 37095 32505 37305
rect 31395 36480 31605 36690
rect 30795 35895 31005 36105
rect 31380 35295 31590 35505
rect 31695 35295 31905 35505
rect 31695 34695 31905 34905
rect 33195 39195 33405 39405
rect 32895 37395 33105 37605
rect 33795 42495 34005 42705
rect 35595 44295 35805 44505
rect 35295 43995 35505 44205
rect 35895 43995 36105 44205
rect 34995 42795 35205 43005
rect 34695 42495 34905 42705
rect 34395 42195 34605 42405
rect 34095 41895 34305 42105
rect 37095 48795 37305 49005
rect 36795 46995 37005 47205
rect 38295 50595 38505 50805
rect 37995 50295 38205 50505
rect 37695 47595 37905 47805
rect 37095 46395 37305 46605
rect 37095 45495 37305 45705
rect 39495 51195 39705 51405
rect 38295 49980 38505 50190
rect 38895 49995 39105 50205
rect 38295 49395 38505 49605
rect 38895 49410 39105 49620
rect 38595 48780 38805 48990
rect 38595 48465 38805 48675
rect 39195 48495 39405 48705
rect 38895 47295 39105 47505
rect 38595 46695 38805 46905
rect 37695 44280 37905 44490
rect 36795 43995 37005 44205
rect 36495 43695 36705 43905
rect 36195 43395 36405 43605
rect 35895 42795 36105 43005
rect 35295 41595 35505 41805
rect 37095 43695 37305 43905
rect 36195 41610 36405 41820
rect 33795 40395 34005 40605
rect 34995 40995 35205 41205
rect 34095 39495 34305 39705
rect 33495 38295 33705 38505
rect 33195 37095 33405 37305
rect 34695 38895 34905 39105
rect 34395 37995 34605 38205
rect 33795 37095 34005 37305
rect 33795 36495 34005 36705
rect 33195 36195 33405 36405
rect 32895 34395 33105 34605
rect 31395 33810 31605 34020
rect 32280 33795 32490 34005
rect 30495 32295 30705 32505
rect 29880 31395 30090 31605
rect 30195 31395 30405 31605
rect 29595 31095 29805 31305
rect 28995 29310 29205 29520
rect 28395 28995 28605 29205
rect 29295 28680 29505 28890
rect 29595 28095 29805 28305
rect 28995 27195 29205 27405
rect 29295 26295 29505 26505
rect 27195 25095 27405 25305
rect 26295 24495 26505 24705
rect 25995 24195 26205 24405
rect 26580 23595 26790 23805
rect 26895 23595 27105 23805
rect 25695 21510 25905 21720
rect 25095 20895 25305 21105
rect 25995 20880 26205 21090
rect 27795 23295 28005 23505
rect 26895 22695 27105 22905
rect 27795 22695 28005 22905
rect 28995 25380 29205 25590
rect 28695 24495 28905 24705
rect 29895 27195 30105 27405
rect 30495 31095 30705 31305
rect 30495 30495 30705 30705
rect 31095 33180 31305 33390
rect 31380 31095 31590 31305
rect 31695 31095 31905 31305
rect 31395 30495 31605 30705
rect 31095 30195 31305 30405
rect 31095 29595 31305 29805
rect 31695 29595 31905 29805
rect 32595 33780 32805 33990
rect 36495 40980 36705 41190
rect 36195 40695 36405 40905
rect 35595 39495 35805 39705
rect 36495 40395 36705 40605
rect 37395 43395 37605 43605
rect 36195 38895 36405 39105
rect 36195 38580 36405 38790
rect 35295 37395 35505 37605
rect 34995 37095 35205 37305
rect 36795 40095 37005 40305
rect 36495 38295 36705 38505
rect 36495 37095 36705 37305
rect 34995 36495 35205 36705
rect 35895 36480 36105 36690
rect 36495 36480 36705 36690
rect 34995 35895 35205 36105
rect 34695 35595 34905 35805
rect 35295 34995 35505 35205
rect 33795 34095 34005 34305
rect 34395 34095 34605 34305
rect 36180 34395 36390 34605
rect 36495 34395 36705 34605
rect 35595 34095 35805 34305
rect 32880 32895 33090 33105
rect 33195 32895 33405 33105
rect 32295 31095 32505 31305
rect 32295 30495 32505 30705
rect 32295 29880 32505 30090
rect 31395 29310 31605 29520
rect 31995 29310 32205 29520
rect 30795 28395 31005 28605
rect 30495 28095 30705 28305
rect 31395 27795 31605 28005
rect 30195 26310 30405 26520
rect 34095 32595 34305 32805
rect 33495 32295 33705 32505
rect 33195 31695 33405 31905
rect 33495 30795 33705 31005
rect 33195 30495 33405 30705
rect 33495 29895 33705 30105
rect 35295 32895 35505 33105
rect 34995 32595 35205 32805
rect 34395 32295 34605 32505
rect 35295 32295 35505 32505
rect 34995 30195 35205 30405
rect 34395 29895 34605 30105
rect 33495 29310 33705 29520
rect 34695 28995 34905 29205
rect 33495 28395 33705 28605
rect 33195 27795 33405 28005
rect 31695 27495 31905 27705
rect 32895 27495 33105 27705
rect 31695 26595 31905 26805
rect 32595 26595 32805 26805
rect 30195 25995 30405 26205
rect 30795 26010 31005 26220
rect 31395 26010 31605 26220
rect 29895 25380 30105 25590
rect 31095 25095 31305 25305
rect 31995 26010 32205 26220
rect 33195 25995 33405 26205
rect 31695 25395 31905 25605
rect 29295 23895 29505 24105
rect 31395 23895 31605 24105
rect 28695 22995 28905 23205
rect 28995 22695 29205 22905
rect 32295 25380 32505 25590
rect 32895 25380 33105 25590
rect 32295 24195 32505 24405
rect 32295 22995 32505 23205
rect 31980 22695 32190 22905
rect 27780 21795 27990 22005
rect 26895 21495 27105 21705
rect 28095 21780 28305 21990
rect 28395 21795 28605 22005
rect 28695 21510 28905 21720
rect 27195 20880 27405 21090
rect 30795 22395 31005 22605
rect 30195 21510 30405 21720
rect 32295 22680 32505 22890
rect 32295 21795 32505 22005
rect 32595 21510 32805 21720
rect 34995 27795 35205 28005
rect 34695 26595 34905 26805
rect 34395 26010 34605 26220
rect 33495 24495 33705 24705
rect 34695 25380 34905 25590
rect 34095 24795 34305 25005
rect 34395 24495 34605 24705
rect 34695 23895 34905 24105
rect 34395 23295 34605 23505
rect 33195 22395 33405 22605
rect 33795 22395 34005 22605
rect 34095 21510 34305 21720
rect 28995 20895 29205 21105
rect 27795 20595 28005 20805
rect 28695 20595 28905 20805
rect 27195 20295 27405 20505
rect 30495 20880 30705 21090
rect 31395 20880 31605 21090
rect 29895 20295 30105 20505
rect 27195 19695 27405 19905
rect 29595 19695 29805 19905
rect 26595 19395 26805 19605
rect 27795 18795 28005 19005
rect 25395 18495 25605 18705
rect 25995 18210 26205 18420
rect 26895 18195 27105 18405
rect 27795 18210 28005 18420
rect 28695 18195 28905 18405
rect 30795 18495 31005 18705
rect 30195 18195 30405 18405
rect 33195 20895 33405 21105
rect 31695 20295 31905 20505
rect 32295 20295 32505 20505
rect 31695 19695 31905 19905
rect 32295 19395 32505 19605
rect 32295 18795 32505 19005
rect 31695 18495 31905 18705
rect 25395 15195 25605 15405
rect 24795 13995 25005 14205
rect 24495 13710 24705 13920
rect 25695 14895 25905 15105
rect 26895 17580 27105 17790
rect 27495 17580 27705 17790
rect 26295 14295 26505 14505
rect 25695 13710 25905 13920
rect 26295 13710 26505 13920
rect 27795 16395 28005 16605
rect 20895 12495 21105 12705
rect 20295 10410 20505 10620
rect 20895 10410 21105 10620
rect 22695 13080 22905 13290
rect 23595 13080 23805 13290
rect 24795 13080 25005 13290
rect 25395 13080 25605 13290
rect 25995 13080 26205 13290
rect 25995 12195 26205 12405
rect 22695 11895 22905 12105
rect 22095 10395 22305 10605
rect 24795 11595 25005 11805
rect 23295 10410 23505 10620
rect 24795 10410 25005 10620
rect 18795 9780 19005 9990
rect 19395 9780 19605 9990
rect 20595 9780 20805 9990
rect 21195 9795 21405 10005
rect 18195 9495 18405 9705
rect 17295 9195 17505 9405
rect 18195 7995 18405 8205
rect 14895 7695 15105 7905
rect 16395 7695 16605 7905
rect 16995 7695 17205 7905
rect 14295 7395 14505 7605
rect 13395 6795 13605 7005
rect 13995 6795 14205 7005
rect 10095 5295 10305 5505
rect 9795 4995 10005 5205
rect 10695 4995 10905 5205
rect 10095 4695 10305 4905
rect 9195 4395 9405 4605
rect 9795 4095 10005 4305
rect 8895 3195 9105 3405
rect 10995 3795 11205 4005
rect 11895 5295 12105 5505
rect 12495 5280 12705 5490
rect 15495 7395 15705 7605
rect 12195 4695 12405 4905
rect 11295 3195 11505 3405
rect 14295 5295 14505 5505
rect 15195 5280 15405 5490
rect 13995 4695 14205 4905
rect 13695 4095 13905 4305
rect 12495 3795 12705 4005
rect 13395 3795 13605 4005
rect 8895 1980 9105 2190
rect 9495 1980 9705 2190
rect 7695 1695 7905 1905
rect 8385 1695 8595 1905
rect 10995 1095 11205 1305
rect 4695 795 4905 1005
rect 12195 2895 12405 3105
rect 11895 2610 12105 2820
rect 13095 3195 13305 3405
rect 13095 2595 13305 2805
rect 12195 1980 12405 2190
rect 12795 1980 13005 2190
rect 13695 2295 13905 2505
rect 14895 3795 15105 4005
rect 15795 3795 16005 4005
rect 17595 7395 17805 7605
rect 17595 6795 17805 7005
rect 16695 5895 16905 6105
rect 20595 7395 20805 7605
rect 19095 6795 19305 7005
rect 18195 5895 18405 6105
rect 19695 5910 19905 6120
rect 16695 5295 16905 5505
rect 17295 5280 17505 5490
rect 17895 5280 18105 5490
rect 18795 5280 19005 5490
rect 16695 4695 16905 4905
rect 19095 4695 19305 4905
rect 18495 4095 18705 4305
rect 16395 3495 16605 3705
rect 17595 3495 17805 3705
rect 14895 2610 15105 2820
rect 16695 2610 16905 2820
rect 17295 2595 17505 2805
rect 13995 1995 14205 2205
rect 14595 1980 14805 2190
rect 15795 1980 16005 2190
rect 27495 13080 27705 13290
rect 26595 11595 26805 11805
rect 27195 11595 27405 11805
rect 27195 10995 27405 11205
rect 28695 16095 28905 16305
rect 28695 15495 28905 15705
rect 28395 14595 28605 14805
rect 28995 13995 29205 14205
rect 30495 17595 30705 17805
rect 33795 20880 34005 21090
rect 33195 20580 33405 20790
rect 34995 23295 35205 23505
rect 35595 31395 35805 31605
rect 37995 43095 38205 43305
rect 37695 42195 37905 42405
rect 39495 46695 39705 46905
rect 39495 45795 39705 46005
rect 40095 49995 40305 50205
rect 41895 56595 42105 56805
rect 44595 59880 44805 60090
rect 48195 71595 48405 71805
rect 49395 74595 49605 74805
rect 49395 73995 49605 74205
rect 49695 73395 49905 73605
rect 49695 72810 49905 73020
rect 49395 72180 49605 72390
rect 49395 71295 49605 71505
rect 49095 70395 49305 70605
rect 49095 69795 49305 70005
rect 48795 69495 49005 69705
rect 48495 68295 48705 68505
rect 47595 67395 47805 67605
rect 51195 79980 51405 80190
rect 51495 79695 51705 79905
rect 50895 77895 51105 78105
rect 52395 79980 52605 80190
rect 53595 79980 53805 80190
rect 54195 79980 54405 80190
rect 51795 78795 52005 79005
rect 54195 79395 54405 79605
rect 52395 78495 52605 78705
rect 52695 77895 52905 78105
rect 51495 77295 51705 77505
rect 50895 76095 51105 76305
rect 52095 76110 52305 76320
rect 52995 77595 53205 77805
rect 54495 77595 54705 77805
rect 53295 76995 53505 77205
rect 53895 76995 54105 77205
rect 53295 76395 53505 76605
rect 53895 76110 54105 76320
rect 55095 82395 55305 82605
rect 50895 74295 51105 74505
rect 52395 75480 52605 75690
rect 52995 75495 53205 75705
rect 52395 74895 52605 75105
rect 52095 74595 52305 74805
rect 52095 73995 52305 74205
rect 50895 73695 51105 73905
rect 51795 73695 52005 73905
rect 51495 73395 51705 73605
rect 54195 75480 54405 75690
rect 54495 75195 54705 75405
rect 53295 74595 53505 74805
rect 53895 74595 54105 74805
rect 53295 72810 53505 73020
rect 54195 72795 54405 73005
rect 51195 71595 51405 71805
rect 51795 71595 52005 71805
rect 50295 71295 50505 71505
rect 49995 70695 50205 70905
rect 49695 68295 49905 68505
rect 52395 68895 52605 69105
rect 52995 72180 53205 72390
rect 53595 70995 53805 71205
rect 53295 70095 53505 70305
rect 53280 69495 53490 69705
rect 53595 69495 53805 69705
rect 54195 71595 54405 71805
rect 54195 70395 54405 70605
rect 54195 68295 54405 68505
rect 49695 67095 49905 67305
rect 48195 66195 48405 66405
rect 49395 66195 49605 66405
rect 49395 65595 49605 65805
rect 49095 63795 49305 64005
rect 47895 63495 48105 63705
rect 48795 62895 49005 63105
rect 48795 61695 49005 61905
rect 47595 60540 47805 60750
rect 48495 60540 48705 60750
rect 46695 58395 46905 58605
rect 51195 65895 51405 66105
rect 49995 65595 50205 65805
rect 51795 65595 52005 65805
rect 50595 65010 50805 65220
rect 51195 65010 51405 65220
rect 49695 61395 49905 61605
rect 49395 61095 49605 61305
rect 49995 61095 50205 61305
rect 50295 60795 50505 61005
rect 50595 60510 50805 60720
rect 53295 67095 53505 67305
rect 54195 67095 54405 67305
rect 53595 66495 53805 66705
rect 52995 65595 53205 65805
rect 52395 65010 52605 65220
rect 53895 65895 54105 66105
rect 53595 64995 53805 65205
rect 51795 63495 52005 63705
rect 53295 64380 53505 64590
rect 53595 64095 53805 64305
rect 53595 62895 53805 63105
rect 56895 86895 57105 87105
rect 57795 86595 58005 86805
rect 56895 86295 57105 86505
rect 57795 85695 58005 85905
rect 56895 83910 57105 84120
rect 57495 83895 57705 84105
rect 56595 82095 56805 82305
rect 55995 81795 56205 82005
rect 55695 80610 55905 80820
rect 56295 80610 56505 80820
rect 65595 93495 65805 93705
rect 66495 93495 66705 93705
rect 65295 93195 65505 93405
rect 58395 92295 58605 92505
rect 60195 92295 60405 92505
rect 64395 92295 64605 92505
rect 58380 91710 58590 91920
rect 58695 91710 58905 91920
rect 59295 91710 59505 91920
rect 59895 91710 60105 91920
rect 60495 91710 60705 91920
rect 61395 91710 61605 91920
rect 58395 91095 58605 91305
rect 58995 91080 59205 91290
rect 59595 90795 59805 91005
rect 60195 90795 60405 91005
rect 59595 88995 59805 89205
rect 58695 87780 58905 87990
rect 61980 91695 62190 91905
rect 62295 91710 62505 91920
rect 62895 91710 63105 91920
rect 63495 91710 63705 91920
rect 61995 90795 62205 91005
rect 63795 91080 64005 91290
rect 65595 92895 65805 93105
rect 65895 92295 66105 92505
rect 65295 91710 65505 91920
rect 63495 90795 63705 91005
rect 63195 90495 63405 90705
rect 62295 90195 62505 90405
rect 64395 90795 64605 91005
rect 64095 90495 64305 90705
rect 62895 89895 63105 90105
rect 63495 89895 63705 90105
rect 62895 89295 63105 89505
rect 60495 88995 60705 89205
rect 61995 88995 62205 89205
rect 64995 90195 65205 90405
rect 64980 89880 65190 90090
rect 65295 89895 65505 90105
rect 63795 88695 64005 88905
rect 64395 88695 64605 88905
rect 61395 88410 61605 88620
rect 61995 88410 62205 88620
rect 63195 88410 63405 88620
rect 61095 87780 61305 87990
rect 59295 87495 59505 87705
rect 60195 87495 60405 87705
rect 58995 86295 59205 86505
rect 58395 85995 58605 86205
rect 58095 83895 58305 84105
rect 61095 87195 61305 87405
rect 62580 87795 62790 88005
rect 62895 87780 63105 87990
rect 64095 87795 64305 88005
rect 65895 90495 66105 90705
rect 65595 88695 65805 88905
rect 73995 93195 74205 93405
rect 71895 92295 72105 92505
rect 67395 91710 67605 91920
rect 68295 91695 68505 91905
rect 72495 91710 72705 91920
rect 73395 91710 73605 91920
rect 66795 91080 67005 91290
rect 67695 91080 67905 91290
rect 68295 91080 68505 91290
rect 66495 89895 66705 90105
rect 67380 90495 67590 90705
rect 67695 90495 67905 90705
rect 67095 89595 67305 89805
rect 66795 89295 67005 89505
rect 66495 88695 66705 88905
rect 67395 88995 67605 89205
rect 67995 88995 68205 89205
rect 68595 90495 68805 90705
rect 69495 89595 69705 89805
rect 69195 88995 69405 89205
rect 69195 88395 69405 88605
rect 64995 87780 65205 87990
rect 65595 87780 65805 87990
rect 67095 87780 67305 87990
rect 67695 87780 67905 87990
rect 61695 86895 61905 87105
rect 64095 86895 64305 87105
rect 65595 86895 65805 87105
rect 60795 86595 61005 86805
rect 60495 86295 60705 86505
rect 59295 85395 59505 85605
rect 59895 85395 60105 85605
rect 58995 85095 59205 85305
rect 58995 83910 59205 84120
rect 57780 83295 57990 83505
rect 58095 83295 58305 83505
rect 57795 82695 58005 82905
rect 57180 80595 57390 80805
rect 57495 80595 57705 80805
rect 58095 82395 58305 82605
rect 59295 83295 59505 83505
rect 60195 84795 60405 85005
rect 60495 84495 60705 84705
rect 60195 83895 60405 84105
rect 63495 85695 63705 85905
rect 61395 83910 61605 84120
rect 61995 83910 62205 84120
rect 62895 83910 63105 84120
rect 65595 84495 65805 84705
rect 64095 83910 64305 84120
rect 64695 83910 64905 84120
rect 65295 83910 65505 84120
rect 60195 83295 60405 83505
rect 59895 82695 60105 82905
rect 58695 82095 58905 82305
rect 58395 81795 58605 82005
rect 58995 81495 59205 81705
rect 59595 81495 59805 81705
rect 60495 82695 60705 82905
rect 61095 82695 61305 82905
rect 62595 82995 62805 83205
rect 63795 82995 64005 83205
rect 62295 82095 62505 82305
rect 63195 82095 63405 82305
rect 61095 81495 61305 81705
rect 58995 80595 59205 80805
rect 55995 78795 56205 79005
rect 55695 78495 55905 78705
rect 58680 79980 58890 80190
rect 58995 79980 59205 80190
rect 57195 79395 57405 79605
rect 56595 78195 56805 78405
rect 55695 77295 55905 77505
rect 57195 77295 57405 77505
rect 55395 76695 55605 76905
rect 56595 76695 56805 76905
rect 55095 75195 55305 75405
rect 54795 74595 55005 74805
rect 55995 76110 56205 76320
rect 57495 76695 57705 76905
rect 55695 75495 55905 75705
rect 55695 74895 55905 75105
rect 56295 74595 56505 74805
rect 55395 73095 55605 73305
rect 54795 72795 55005 73005
rect 55695 72810 55905 73020
rect 58695 78795 58905 79005
rect 58095 78495 58305 78705
rect 58995 78495 59205 78705
rect 60195 79980 60405 80190
rect 61395 81195 61605 81405
rect 59895 79395 60105 79605
rect 61095 79395 61305 79605
rect 59595 79095 59805 79305
rect 59595 78495 59805 78705
rect 58395 76995 58605 77205
rect 58095 76095 58305 76305
rect 59295 77595 59505 77805
rect 59295 76695 59505 76905
rect 58995 76095 59205 76305
rect 57795 75195 58005 75405
rect 58380 75195 58590 75405
rect 58695 75195 58905 75405
rect 56895 74895 57105 75105
rect 57195 74595 57405 74805
rect 56595 73995 56805 74205
rect 57195 73995 57405 74205
rect 56895 73695 57105 73905
rect 56295 72795 56505 73005
rect 57495 72810 57705 73020
rect 54795 71595 55005 71805
rect 55995 72180 56205 72390
rect 57195 72180 57405 72390
rect 56895 71895 57105 72105
rect 56595 70695 56805 70905
rect 55395 70395 55605 70605
rect 54795 70095 55005 70305
rect 54495 65295 54705 65505
rect 55395 70080 55605 70290
rect 55995 68310 56205 68520
rect 56595 67695 56805 67905
rect 55695 66495 55905 66705
rect 55695 65895 55905 66105
rect 54195 63795 54405 64005
rect 55395 65010 55605 65220
rect 55995 65040 56205 65250
rect 54795 64395 55005 64605
rect 55695 64395 55905 64605
rect 55080 63795 55290 64005
rect 55395 63795 55605 64005
rect 54795 62895 55005 63105
rect 54495 62595 54705 62805
rect 53895 61995 54105 62205
rect 54795 61995 55005 62205
rect 52695 61695 52905 61905
rect 52395 61395 52605 61605
rect 49395 60195 49605 60405
rect 47295 59895 47505 60105
rect 45495 57795 45705 58005
rect 46095 57795 46305 58005
rect 46995 57795 47205 58005
rect 44895 57495 45105 57705
rect 45795 57495 46005 57705
rect 44295 57195 44505 57405
rect 42495 56580 42705 56790
rect 42795 56295 43005 56505
rect 41895 55395 42105 55605
rect 40995 54495 41205 54705
rect 43995 56580 44205 56790
rect 44595 56580 44805 56790
rect 45195 56580 45405 56790
rect 43395 56295 43605 56505
rect 44895 55395 45105 55605
rect 43395 55095 43605 55305
rect 43695 54795 43905 55005
rect 43095 54195 43305 54405
rect 42795 53595 43005 53805
rect 41295 52995 41505 53205
rect 42795 52695 43005 52905
rect 43095 52995 43305 53205
rect 45495 55095 45705 55305
rect 45195 53595 45405 53805
rect 44295 52710 44505 52920
rect 44895 52710 45105 52920
rect 42495 52395 42705 52605
rect 42195 51495 42405 51705
rect 41595 51195 41805 51405
rect 40995 50595 41205 50805
rect 40695 50295 40905 50505
rect 40395 49695 40605 49905
rect 41595 50295 41805 50505
rect 41295 49695 41505 49905
rect 40995 49395 41205 49605
rect 40095 48795 40305 49005
rect 40995 48795 41205 49005
rect 40695 48195 40905 48405
rect 40395 47895 40605 48105
rect 40095 46695 40305 46905
rect 39795 45195 40005 45405
rect 40395 45495 40605 45705
rect 39195 43995 39405 44205
rect 38295 42195 38505 42405
rect 40395 44295 40605 44505
rect 43395 52080 43605 52290
rect 44595 51795 44805 52005
rect 43995 50895 44205 51105
rect 43395 50595 43605 50805
rect 42495 50295 42705 50505
rect 42195 49695 42405 49905
rect 43095 49695 43305 49905
rect 42495 49410 42705 49620
rect 42195 48780 42405 48990
rect 42795 48780 43005 48990
rect 44895 51495 45105 51705
rect 45195 50595 45405 50805
rect 45795 54495 46005 54705
rect 46395 57195 46605 57405
rect 50295 59880 50505 60090
rect 50895 59895 51105 60105
rect 52695 60495 52905 60705
rect 53295 60540 53505 60750
rect 54195 60540 54405 60750
rect 49395 59295 49605 59505
rect 51495 59850 51705 60060
rect 52395 59850 52605 60060
rect 51195 59295 51405 59505
rect 49395 58695 49605 58905
rect 50895 58695 51105 58905
rect 47895 58395 48105 58605
rect 48195 58095 48405 58305
rect 47895 57795 48105 58005
rect 48195 57195 48405 57405
rect 47595 56580 47805 56790
rect 46395 56295 46605 56505
rect 48195 56295 48405 56505
rect 47595 55995 47805 56205
rect 47895 55395 48105 55605
rect 47595 54495 47805 54705
rect 47580 53895 47790 54105
rect 47895 53895 48105 54105
rect 52395 58995 52605 59205
rect 54495 59895 54705 60105
rect 54495 59295 54705 59505
rect 51495 58695 51705 58905
rect 52695 58695 52905 58905
rect 51195 58395 51405 58605
rect 49695 57495 49905 57705
rect 51795 58395 52005 58605
rect 54195 58395 54405 58605
rect 51495 57195 51705 57405
rect 49695 56595 49905 56805
rect 50280 56550 50490 56760
rect 50595 56595 50805 56805
rect 52095 58095 52305 58305
rect 49695 55995 49905 56205
rect 51195 56550 51405 56760
rect 51795 56550 52005 56760
rect 52395 57495 52605 57705
rect 52695 57210 52905 57420
rect 52395 56595 52605 56805
rect 52095 56295 52305 56505
rect 50295 55095 50505 55305
rect 49095 54795 49305 55005
rect 49695 54795 49905 55005
rect 48795 54495 49005 54705
rect 48495 53895 48705 54105
rect 46095 53295 46305 53505
rect 47295 53295 47505 53505
rect 48195 53295 48405 53505
rect 46695 52710 46905 52920
rect 47295 52695 47505 52905
rect 47895 52710 48105 52920
rect 48795 52695 49005 52905
rect 43695 49995 43905 50205
rect 44595 49995 44805 50205
rect 46095 49995 46305 50205
rect 41595 48495 41805 48705
rect 43395 48495 43605 48705
rect 43095 48195 43305 48405
rect 42795 47895 43005 48105
rect 41595 47295 41805 47505
rect 42195 47295 42405 47505
rect 41295 46395 41505 46605
rect 42495 46695 42705 46905
rect 42495 46095 42705 46305
rect 40995 44895 41205 45105
rect 41595 44910 41805 45120
rect 42195 44895 42405 45105
rect 40695 43695 40905 43905
rect 39795 42795 40005 43005
rect 40995 42495 41205 42705
rect 40995 41895 41205 42105
rect 39195 41595 39405 41805
rect 40395 41610 40605 41820
rect 37695 40695 37905 40905
rect 37395 40095 37605 40305
rect 37995 40395 38205 40605
rect 38295 40095 38505 40305
rect 39495 41295 39705 41505
rect 40095 40980 40305 41190
rect 40695 40980 40905 41190
rect 42495 44295 42705 44505
rect 41895 43695 42105 43905
rect 41895 43380 42105 43590
rect 43395 47595 43605 47805
rect 43095 46695 43305 46905
rect 44595 49410 44805 49620
rect 44295 48780 44505 48990
rect 43995 48195 44205 48405
rect 43995 47295 44205 47505
rect 43695 45795 43905 46005
rect 43395 45495 43605 45705
rect 45195 48195 45405 48405
rect 44895 46095 45105 46305
rect 44595 45195 44805 45405
rect 44895 44895 45105 45105
rect 43095 44295 43305 44505
rect 42795 43395 43005 43605
rect 43695 44280 43905 44490
rect 47280 52095 47490 52305
rect 47595 52095 47805 52305
rect 47295 51495 47505 51705
rect 46995 51195 47205 51405
rect 46695 50895 46905 51105
rect 46395 49695 46605 49905
rect 46995 49995 47205 50205
rect 46995 48780 47205 48990
rect 46395 48195 46605 48405
rect 45495 47895 45705 48105
rect 46995 47595 47205 47805
rect 45495 46995 45705 47205
rect 46095 46995 46305 47205
rect 45795 46695 46005 46905
rect 45495 45795 45705 46005
rect 47895 51795 48105 52005
rect 48795 52095 49005 52305
rect 48195 51495 48405 51705
rect 53595 55995 53805 56205
rect 55095 61695 55305 61905
rect 56595 62895 56805 63105
rect 55695 62295 55905 62505
rect 55395 60495 55605 60705
rect 58095 72195 58305 72405
rect 57795 71595 58005 71805
rect 57195 69195 57405 69405
rect 58095 68895 58305 69105
rect 58995 73695 59205 73905
rect 58695 73395 58905 73605
rect 60495 78195 60705 78405
rect 60495 77595 60705 77805
rect 60195 77295 60405 77505
rect 60195 76695 60405 76905
rect 60780 76695 60990 76905
rect 61095 76695 61305 76905
rect 62895 80610 63105 80820
rect 64995 83280 65205 83490
rect 65595 82695 65805 82905
rect 66195 87195 66405 87405
rect 68895 87780 69105 87990
rect 69495 87780 69705 87990
rect 68895 85395 69105 85605
rect 66195 85095 66405 85305
rect 68295 85095 68505 85305
rect 65895 81495 66105 81705
rect 67695 84495 67905 84705
rect 66495 83910 66705 84120
rect 67095 83910 67305 84120
rect 69495 83910 69705 84120
rect 70095 90495 70305 90705
rect 72195 91080 72405 91290
rect 77895 93795 78105 94005
rect 76095 93495 76305 93705
rect 76695 93495 76905 93705
rect 74295 92895 74505 93105
rect 74595 92295 74805 92505
rect 75195 91995 75405 92205
rect 73995 90495 74205 90705
rect 71895 89895 72105 90105
rect 72795 89895 73005 90105
rect 73395 89895 73605 90105
rect 70995 89595 71205 89805
rect 70695 89295 70905 89505
rect 70095 88395 70305 88605
rect 71595 89295 71805 89505
rect 71295 88395 71505 88605
rect 75495 91080 75705 91290
rect 74895 89595 75105 89805
rect 72495 88995 72705 89205
rect 73695 88995 73905 89205
rect 71895 88395 72105 88605
rect 73095 88410 73305 88620
rect 70395 87780 70605 87990
rect 70995 87780 71205 87990
rect 71595 87780 71805 87990
rect 72195 87780 72405 87990
rect 72795 87780 73005 87990
rect 72195 87195 72405 87405
rect 72195 85995 72405 86205
rect 70995 85695 71205 85905
rect 70395 84495 70605 84705
rect 66495 82695 66705 82905
rect 67395 83280 67605 83490
rect 69795 83295 70005 83505
rect 69195 82995 69405 83205
rect 68895 82695 69105 82905
rect 69495 82695 69705 82905
rect 66795 82395 67005 82605
rect 67995 82395 68205 82605
rect 67995 81495 68205 81705
rect 66195 81195 66405 81405
rect 69495 82095 69705 82305
rect 72795 85395 73005 85605
rect 72195 85095 72405 85305
rect 71595 83910 71805 84120
rect 72495 84495 72705 84705
rect 70395 82395 70605 82605
rect 70095 82095 70305 82305
rect 69195 81195 69405 81405
rect 66495 80610 66705 80820
rect 67395 80595 67605 80805
rect 68295 80610 68505 80820
rect 68895 80610 69105 80820
rect 61680 79995 61890 80205
rect 61995 79980 62205 80190
rect 62595 79980 62805 80190
rect 63795 79995 64005 80205
rect 63195 79395 63405 79605
rect 64695 79980 64905 80190
rect 65595 79995 65805 80205
rect 64395 79695 64605 79905
rect 65295 79395 65505 79605
rect 63495 78795 63705 79005
rect 62295 78195 62505 78405
rect 62595 77895 62805 78105
rect 61995 77295 62205 77505
rect 61695 76995 61905 77205
rect 62295 76995 62505 77205
rect 61395 76395 61605 76605
rect 61995 76395 62205 76605
rect 61695 76110 61905 76320
rect 60195 75495 60405 75705
rect 60195 74595 60405 74805
rect 61095 75195 61305 75405
rect 59895 73695 60105 73905
rect 60795 73695 61005 73905
rect 59595 73095 59805 73305
rect 60495 73095 60705 73305
rect 59895 72810 60105 73020
rect 61995 75495 62205 75705
rect 61695 74895 61905 75105
rect 61395 74595 61605 74805
rect 61995 73995 62205 74205
rect 61695 73695 61905 73905
rect 62895 77280 63105 77490
rect 64995 78495 65205 78705
rect 64395 77895 64605 78105
rect 64995 77895 65205 78105
rect 63795 77595 64005 77805
rect 63495 76395 63705 76605
rect 67395 79980 67605 80190
rect 67995 79980 68205 80190
rect 66795 79395 67005 79605
rect 66195 79095 66405 79305
rect 65595 78195 65805 78405
rect 67095 78795 67305 79005
rect 66795 78195 67005 78405
rect 66195 76995 66405 77205
rect 66195 76395 66405 76605
rect 63495 75480 63705 75690
rect 63195 74895 63405 75105
rect 62895 74295 63105 74505
rect 62895 73695 63105 73905
rect 62595 73395 62805 73605
rect 62895 73095 63105 73305
rect 61095 72810 61305 73020
rect 61995 72810 62205 73020
rect 62895 72780 63105 72990
rect 64695 75495 64905 75705
rect 64095 74595 64305 74805
rect 63495 74295 63705 74505
rect 64695 74295 64905 74505
rect 63195 72495 63405 72705
rect 59595 72180 59805 72390
rect 60195 72180 60405 72390
rect 61095 72195 61305 72405
rect 59295 71295 59505 71505
rect 58995 70695 59205 70905
rect 58695 70095 58905 70305
rect 57195 68310 57405 68520
rect 56895 62295 57105 62505
rect 56295 61095 56505 61305
rect 55995 59880 56205 60090
rect 57495 67695 57705 67905
rect 57795 67095 58005 67305
rect 58395 67095 58605 67305
rect 59895 70395 60105 70605
rect 59895 69795 60105 70005
rect 61095 71595 61305 71805
rect 60795 70695 61005 70905
rect 60195 68310 60405 68520
rect 58995 66795 59205 67005
rect 59895 67395 60105 67605
rect 59595 66195 59805 66405
rect 59295 65895 59505 66105
rect 59295 65295 59505 65505
rect 57495 64995 57705 65205
rect 57495 64395 57705 64605
rect 58095 64395 58305 64605
rect 57195 61695 57405 61905
rect 58695 63795 58905 64005
rect 55095 58395 55305 58605
rect 54795 57495 55005 57705
rect 55995 57495 56205 57705
rect 55095 57210 55305 57420
rect 54795 56295 55005 56505
rect 49995 54195 50205 54405
rect 50595 54195 50805 54405
rect 52395 54195 52605 54405
rect 52995 54195 53205 54405
rect 54195 54195 54405 54405
rect 55395 55395 55605 55605
rect 54795 53895 55005 54105
rect 53595 53295 53805 53505
rect 49995 52710 50205 52920
rect 50595 52710 50805 52920
rect 51495 52710 51705 52920
rect 52395 52710 52605 52920
rect 52995 52710 53205 52920
rect 49395 52095 49605 52305
rect 49095 51795 49305 52005
rect 48795 51195 49005 51405
rect 47895 50895 48105 51105
rect 49695 51795 49905 52005
rect 48795 50595 49005 50805
rect 49395 50595 49605 50805
rect 48195 49995 48405 50205
rect 47895 49695 48105 49905
rect 46995 46395 47205 46605
rect 47595 46395 47805 46605
rect 49395 49410 49605 49620
rect 48195 48780 48405 48990
rect 49095 48780 49305 48990
rect 48495 48495 48705 48705
rect 49395 48495 49605 48705
rect 49095 47895 49305 48105
rect 48795 47595 49005 47805
rect 48795 46695 49005 46905
rect 48495 45795 48705 46005
rect 47580 45495 47790 45705
rect 47895 45495 48105 45705
rect 46395 44910 46605 45120
rect 47295 44910 47505 45120
rect 45495 44295 45705 44505
rect 45195 43695 45405 43905
rect 44295 43095 44505 43305
rect 43095 42795 43305 43005
rect 43395 42195 43605 42405
rect 44595 42195 44805 42405
rect 42495 41610 42705 41820
rect 43695 41595 43905 41805
rect 45195 41610 45405 41820
rect 41595 40980 41805 41190
rect 38595 39795 38805 40005
rect 38895 39495 39105 39705
rect 38295 39195 38505 39405
rect 37695 37995 37905 38205
rect 37695 37680 37905 37890
rect 37095 37095 37305 37305
rect 37995 36480 38205 36690
rect 37395 35595 37605 35805
rect 39495 40095 39705 40305
rect 41295 40395 41505 40605
rect 40395 39795 40605 40005
rect 40695 39495 40905 39705
rect 40395 39195 40605 39405
rect 40395 38595 40605 38805
rect 40095 38295 40305 38505
rect 40695 37695 40905 37905
rect 39495 37395 39705 37605
rect 39195 37110 39405 37320
rect 40095 37110 40305 37320
rect 40695 37095 40905 37305
rect 37395 35280 37605 35490
rect 38895 35295 39105 35505
rect 39795 35295 40005 35505
rect 37095 34695 37305 34905
rect 40095 34995 40305 35205
rect 38895 34695 39105 34905
rect 36495 33495 36705 33705
rect 36195 32295 36405 32505
rect 36495 31995 36705 32205
rect 36195 31695 36405 31905
rect 37095 31695 37305 31905
rect 37695 31695 37905 31905
rect 35895 29895 36105 30105
rect 38295 32895 38505 33105
rect 38295 31395 38505 31605
rect 37995 31095 38205 31305
rect 36795 30795 37005 31005
rect 37695 30795 37905 31005
rect 36495 30495 36705 30705
rect 36795 30195 37005 30405
rect 36495 29895 36705 30105
rect 37995 29895 38205 30105
rect 40695 35895 40905 36105
rect 40695 34395 40905 34605
rect 40695 33495 40905 33705
rect 39495 33180 39705 33390
rect 39495 32595 39705 32805
rect 41295 37395 41505 37605
rect 42795 40980 43005 41190
rect 43395 40995 43605 41205
rect 42195 40395 42405 40605
rect 41895 39795 42105 40005
rect 44895 40980 45105 41190
rect 43695 40395 43905 40605
rect 44295 40395 44505 40605
rect 43395 39795 43605 40005
rect 42795 38895 43005 39105
rect 41895 38595 42105 38805
rect 42795 38295 43005 38505
rect 42495 37695 42705 37905
rect 44595 40095 44805 40305
rect 44295 39795 44505 40005
rect 43995 38595 44205 38805
rect 43395 37095 43605 37305
rect 46095 44280 46305 44490
rect 47895 44910 48105 45120
rect 48495 44910 48705 45120
rect 49695 47295 49905 47505
rect 50895 52095 51105 52305
rect 58695 61095 58905 61305
rect 57495 60510 57705 60720
rect 58095 60510 58305 60720
rect 60195 67095 60405 67305
rect 60195 66495 60405 66705
rect 60795 66195 61005 66405
rect 62295 72180 62505 72390
rect 62895 72195 63105 72405
rect 61695 71895 61905 72105
rect 62595 71895 62805 72105
rect 61395 69795 61605 70005
rect 62295 69195 62505 69405
rect 61695 68310 61905 68520
rect 62895 70695 63105 70905
rect 64395 73995 64605 74205
rect 65295 75495 65505 75705
rect 64695 72180 64905 72390
rect 64995 71595 65205 71805
rect 63495 70995 63705 71205
rect 64095 70995 64305 71205
rect 63195 70395 63405 70605
rect 62895 69795 63105 70005
rect 62595 68295 62805 68505
rect 65595 74595 65805 74805
rect 66495 75195 66705 75405
rect 65895 73395 66105 73605
rect 66795 74595 67005 74805
rect 67395 78495 67605 78705
rect 67695 77895 67905 78105
rect 68295 77595 68505 77805
rect 68595 77295 68805 77505
rect 68295 76695 68505 76905
rect 67380 76095 67590 76305
rect 67695 76110 67905 76320
rect 68595 76110 68805 76320
rect 67395 75495 67605 75705
rect 67995 75495 68205 75705
rect 67095 73095 67305 73305
rect 66495 72810 66705 73020
rect 67695 73095 67905 73305
rect 67395 72795 67605 73005
rect 66195 72180 66405 72390
rect 66795 72195 67005 72405
rect 66795 71595 67005 71805
rect 68295 74295 68505 74505
rect 70695 81495 70905 81705
rect 72195 83295 72405 83505
rect 71580 82395 71790 82605
rect 71895 82395 72105 82605
rect 71595 81795 71805 82005
rect 72495 82695 72705 82905
rect 74295 88695 74505 88905
rect 73995 88395 74205 88605
rect 75495 88410 75705 88620
rect 75195 87795 75405 88005
rect 74295 85995 74505 86205
rect 73995 85095 74205 85305
rect 72795 82395 73005 82605
rect 73695 83895 73905 84105
rect 72780 81795 72990 82005
rect 73095 81795 73305 82005
rect 71295 81195 71505 81405
rect 72480 81195 72690 81405
rect 72795 81195 73005 81405
rect 69795 79980 70005 80190
rect 70695 79695 70905 79905
rect 69795 78195 70005 78405
rect 69495 77295 69705 77505
rect 71895 80610 72105 80820
rect 73095 80610 73305 80820
rect 71295 79695 71505 79905
rect 71895 79695 72105 79905
rect 70995 78195 71205 78405
rect 71595 77595 71805 77805
rect 70395 76110 70605 76320
rect 69495 75195 69705 75405
rect 69195 73995 69405 74205
rect 69495 73695 69705 73905
rect 70695 75480 70905 75690
rect 73095 79395 73305 79605
rect 73995 83280 74205 83490
rect 73695 82095 73905 82305
rect 73395 78795 73605 79005
rect 76995 91710 77205 91920
rect 76695 91080 76905 91290
rect 76395 90795 76605 91005
rect 76695 90495 76905 90705
rect 77595 91095 77805 91305
rect 84795 93495 85005 93705
rect 79995 92895 80205 93105
rect 79095 92295 79305 92505
rect 78195 91995 78405 92205
rect 78195 91095 78405 91305
rect 79395 91095 79605 91305
rect 77895 90795 78105 91005
rect 78195 90495 78405 90705
rect 77295 90195 77505 90405
rect 78195 89895 78405 90105
rect 76695 89295 76905 89505
rect 76695 88395 76905 88605
rect 77295 88410 77505 88620
rect 78795 88995 79005 89205
rect 78195 88395 78405 88605
rect 79695 88410 79905 88620
rect 76995 87780 77205 87990
rect 76395 87495 76605 87705
rect 77595 87495 77805 87705
rect 76695 86595 76905 86805
rect 77295 86595 77505 86805
rect 76395 86295 76605 86505
rect 76095 85095 76305 85305
rect 75795 84195 76005 84405
rect 77295 85995 77505 86205
rect 76995 85395 77205 85605
rect 76695 84495 76905 84705
rect 77295 84795 77505 85005
rect 77295 83895 77505 84105
rect 76095 83280 76305 83490
rect 76695 83280 76905 83490
rect 75495 82695 75705 82905
rect 75195 82395 75405 82605
rect 74295 80610 74505 80820
rect 75195 81195 75405 81405
rect 76095 81795 76305 82005
rect 74895 80595 75105 80805
rect 74895 79995 75105 80205
rect 74595 79695 74805 79905
rect 74595 78795 74805 79005
rect 74595 78195 74805 78405
rect 73695 77895 73905 78105
rect 75195 79695 75405 79905
rect 73995 77295 74205 77505
rect 74895 77295 75105 77505
rect 72495 76695 72705 76905
rect 72195 76395 72405 76605
rect 73695 76395 73905 76605
rect 73095 76110 73305 76320
rect 70995 75195 71205 75405
rect 71595 75195 71805 75405
rect 70095 74595 70305 74805
rect 68295 73395 68505 73605
rect 69795 73395 70005 73605
rect 68295 72810 68505 73020
rect 68895 72810 69105 73020
rect 67995 72195 68205 72405
rect 68295 71895 68505 72105
rect 65595 71295 65805 71505
rect 66195 71295 66405 71505
rect 67995 71295 68205 71505
rect 65295 70395 65505 70605
rect 64995 70095 65205 70305
rect 64995 69495 65205 69705
rect 64095 69195 64305 69405
rect 63795 68310 64005 68520
rect 64395 68310 64605 68520
rect 62895 67680 63105 67890
rect 63495 67680 63705 67890
rect 61980 67395 62190 67605
rect 62295 67395 62505 67605
rect 61095 65295 61305 65505
rect 60795 65010 61005 65220
rect 61395 65010 61605 65220
rect 65595 67680 65805 67890
rect 63195 67095 63405 67305
rect 64380 67095 64590 67305
rect 64695 67095 64905 67305
rect 59895 64380 60105 64590
rect 60495 64380 60705 64590
rect 59595 63795 59805 64005
rect 60195 62295 60405 62505
rect 61995 64395 62205 64605
rect 61395 63795 61605 64005
rect 61095 61695 61305 61905
rect 59595 61095 59805 61305
rect 60195 61095 60405 61305
rect 59295 60495 59505 60705
rect 57495 59895 57705 60105
rect 57795 59595 58005 59805
rect 57495 58995 57705 59205
rect 56280 57195 56490 57405
rect 56595 57195 56805 57405
rect 57195 57195 57405 57405
rect 58395 58695 58605 58905
rect 58995 58695 59205 58905
rect 58095 57795 58305 58005
rect 57795 57195 58005 57405
rect 56895 56580 57105 56790
rect 57795 56595 58005 56805
rect 56295 55995 56505 56205
rect 55395 52995 55605 53205
rect 55995 52995 56205 53205
rect 54495 52710 54705 52920
rect 56295 52710 56505 52920
rect 56895 52695 57105 52905
rect 50595 51795 50805 52005
rect 51495 51195 51705 51405
rect 50895 49995 51105 50205
rect 51495 49695 51705 49905
rect 51195 49410 51405 49620
rect 52095 52080 52305 52290
rect 52095 50895 52305 51105
rect 52395 49695 52605 49905
rect 52095 49395 52305 49605
rect 50595 47895 50805 48105
rect 51495 48780 51705 48990
rect 52395 48780 52605 48990
rect 53595 52080 53805 52290
rect 54795 52080 55005 52290
rect 55395 52080 55605 52290
rect 56595 52095 56805 52305
rect 53595 51495 53805 51705
rect 55995 51495 56205 51705
rect 53295 49695 53505 49905
rect 54195 49695 54405 49905
rect 55395 49695 55605 49905
rect 55995 49695 56205 49905
rect 53595 48780 53805 48990
rect 54195 48795 54405 49005
rect 56895 49995 57105 50205
rect 58995 57210 59205 57420
rect 60795 60795 61005 61005
rect 61095 60495 61305 60705
rect 60495 59880 60705 60090
rect 61995 62895 62205 63105
rect 61695 61095 61905 61305
rect 59895 59595 60105 59805
rect 61395 59595 61605 59805
rect 61095 57795 61305 58005
rect 60195 57240 60405 57450
rect 62895 64395 63105 64605
rect 62895 62595 63105 62805
rect 62595 61695 62805 61905
rect 65595 66495 65805 66705
rect 63495 66195 63705 66405
rect 64395 65595 64605 65805
rect 65895 65295 66105 65505
rect 63795 63495 64005 63705
rect 63495 62295 63705 62505
rect 63495 61695 63705 61905
rect 64695 61695 64905 61905
rect 63195 60795 63405 61005
rect 61995 60495 62205 60705
rect 62895 60510 63105 60720
rect 65295 61395 65505 61605
rect 63795 60510 64005 60720
rect 61995 59895 62205 60105
rect 61695 57495 61905 57705
rect 63195 59880 63405 60090
rect 65595 61095 65805 61305
rect 63195 58695 63405 58905
rect 62595 58395 62805 58605
rect 63195 58380 63405 58590
rect 62295 57240 62505 57450
rect 59895 56895 60105 57105
rect 58395 56595 58605 56805
rect 58395 55095 58605 55305
rect 59295 56580 59505 56790
rect 58395 54495 58605 54705
rect 58095 52995 58305 53205
rect 60195 55395 60405 55605
rect 58995 52695 59205 52905
rect 60195 52395 60405 52605
rect 57495 51195 57705 51405
rect 59295 52050 59505 52260
rect 63195 56595 63405 56805
rect 63195 56280 63405 56490
rect 61395 55695 61605 55905
rect 60795 55095 61005 55305
rect 62295 54795 62505 55005
rect 61095 52995 61305 53205
rect 62595 53595 62805 53805
rect 60495 51795 60705 52005
rect 61095 51795 61305 52005
rect 60795 51195 61005 51405
rect 58695 50895 58905 51105
rect 59895 50295 60105 50505
rect 58095 49995 58305 50205
rect 55095 48780 55305 48990
rect 54795 48495 55005 48705
rect 52695 48195 52905 48405
rect 51495 47895 51705 48105
rect 50895 47295 51105 47505
rect 49695 45195 49905 45405
rect 50295 45195 50505 45405
rect 47295 43995 47505 44205
rect 46095 43695 46305 43905
rect 46695 43695 46905 43905
rect 45795 38595 46005 38805
rect 48195 44280 48405 44490
rect 48795 44280 49005 44490
rect 49395 44295 49605 44505
rect 48495 43995 48705 44205
rect 47595 43395 47805 43605
rect 47595 42495 47805 42705
rect 48495 40980 48705 41190
rect 49395 43395 49605 43605
rect 50595 44910 50805 45120
rect 50295 42795 50505 43005
rect 50895 42795 51105 43005
rect 49695 41895 49905 42105
rect 50295 41610 50505 41820
rect 51195 41895 51405 42105
rect 50895 41595 51105 41805
rect 46395 39795 46605 40005
rect 46695 38895 46905 39105
rect 46095 37695 46305 37905
rect 43995 36795 44205 37005
rect 41295 36465 41505 36675
rect 41880 36465 42090 36675
rect 42195 36495 42405 36705
rect 43695 36195 43905 36405
rect 42795 35595 43005 35805
rect 42495 35295 42705 35505
rect 42495 34695 42705 34905
rect 42195 34395 42405 34605
rect 43395 33810 43605 34020
rect 43995 33810 44205 34020
rect 41295 33195 41505 33405
rect 43695 33180 43905 33390
rect 40995 32895 41205 33105
rect 41595 32895 41805 33105
rect 39195 32295 39405 32505
rect 37080 29295 37290 29505
rect 37695 29310 37905 29520
rect 38895 29595 39105 29805
rect 38595 29310 38805 29520
rect 36495 28680 36705 28890
rect 37395 28680 37605 28890
rect 35895 28395 36105 28605
rect 36795 27795 37005 28005
rect 38295 27795 38505 28005
rect 35595 27495 35805 27705
rect 35880 27195 36090 27405
rect 36195 27195 36405 27405
rect 36195 26595 36405 26805
rect 35895 26295 36105 26505
rect 37395 26895 37605 27105
rect 35595 25380 35805 25590
rect 37095 25395 37305 25605
rect 34095 20295 34305 20505
rect 34695 20295 34905 20505
rect 33180 18495 33390 18705
rect 33495 18495 33705 18705
rect 32580 18195 32790 18405
rect 32895 18210 33105 18420
rect 34695 19395 34905 19605
rect 36195 22995 36405 23205
rect 35595 21510 35805 21720
rect 36495 22695 36705 22905
rect 36495 22095 36705 22305
rect 34395 18195 34605 18405
rect 31695 17580 31905 17790
rect 32295 17580 32505 17790
rect 33195 17580 33405 17790
rect 33795 17580 34005 17790
rect 34395 17580 34605 17790
rect 31095 17295 31305 17505
rect 30495 16095 30705 16305
rect 29895 14295 30105 14505
rect 31395 15495 31605 15705
rect 31095 14895 31305 15105
rect 30495 13710 30705 13920
rect 32895 14895 33105 15105
rect 32295 14595 32505 14805
rect 31995 14295 32205 14505
rect 28695 13080 28905 13290
rect 29295 13080 29505 13290
rect 29895 13080 30105 13290
rect 29295 12195 29505 12405
rect 28980 11595 29190 11805
rect 29295 11595 29505 11805
rect 28695 11295 28905 11505
rect 27495 10695 27705 10905
rect 26295 10395 26505 10605
rect 26895 10410 27105 10620
rect 23595 9780 23805 9990
rect 22395 9495 22605 9705
rect 22095 9195 22305 9405
rect 25095 9780 25305 9990
rect 25995 9795 26205 10005
rect 26595 9795 26805 10005
rect 26295 9495 26505 9705
rect 24495 9195 24705 9405
rect 22395 8895 22605 9105
rect 24795 8595 25005 8805
rect 24195 8295 24405 8505
rect 21195 6795 21405 7005
rect 23595 6495 23805 6705
rect 20895 6195 21105 6405
rect 22095 5910 22305 6120
rect 21195 5595 21405 5805
rect 20895 4995 21105 5205
rect 20595 4695 20805 4905
rect 22395 4395 22605 4605
rect 22095 3795 22305 4005
rect 19395 3495 19605 3705
rect 19995 2610 20205 2820
rect 20895 2610 21105 2820
rect 21495 2610 21705 2820
rect 18195 1980 18405 2190
rect 19095 1695 19305 1905
rect 13395 1395 13605 1605
rect 18195 1395 18405 1605
rect 18795 1380 19005 1590
rect 21195 1980 21405 2190
rect 22095 1980 22305 2190
rect 20595 1695 20805 1905
rect 22995 4095 23205 4305
rect 22695 3495 22905 3705
rect 27795 9780 28005 9990
rect 27195 7995 27405 8205
rect 25395 7395 25605 7605
rect 24795 5910 25005 6120
rect 28695 10395 28905 10605
rect 29895 10995 30105 11205
rect 32595 14295 32805 14505
rect 31395 13080 31605 13290
rect 32295 13080 32505 13290
rect 30795 12795 31005 13005
rect 31095 11895 31305 12105
rect 32295 11895 32505 12105
rect 28995 9780 29205 9990
rect 29595 8895 29805 9105
rect 28395 8595 28605 8805
rect 30795 10395 31005 10605
rect 31695 10410 31905 10620
rect 33495 13710 33705 13920
rect 36195 20595 36405 20805
rect 34995 18495 35205 18705
rect 35895 18495 36105 18705
rect 34695 17295 34905 17505
rect 35595 18210 35805 18420
rect 38295 26010 38505 26220
rect 40095 31395 40305 31605
rect 40695 30195 40905 30405
rect 40095 29310 40305 29520
rect 41295 31095 41505 31305
rect 41295 28995 41505 29205
rect 39795 28695 40005 28905
rect 45495 37395 45705 37605
rect 44595 37095 44805 37305
rect 45195 37110 45405 37320
rect 44895 36495 45105 36705
rect 44595 35895 44805 36105
rect 44595 35295 44805 35505
rect 46095 36480 46305 36690
rect 45495 36195 45705 36405
rect 46095 36165 46305 36375
rect 44895 34695 45105 34905
rect 45495 34695 45705 34905
rect 44895 33810 45105 34020
rect 48195 38595 48405 38805
rect 47595 37110 47805 37320
rect 46995 35595 47205 35805
rect 46695 35295 46905 35505
rect 46095 33810 46305 34020
rect 47595 33810 47805 34020
rect 44895 33195 45105 33405
rect 45795 32895 46005 33105
rect 47295 32895 47505 33105
rect 47595 32595 47805 32805
rect 44595 32295 44805 32505
rect 44295 31995 44505 32205
rect 42795 29595 43005 29805
rect 43695 29310 43905 29520
rect 44295 29310 44505 29520
rect 45195 29310 45405 29520
rect 46095 29310 46305 29520
rect 39495 26895 39705 27105
rect 39495 26295 39705 26505
rect 40695 27495 40905 27705
rect 40395 26895 40605 27105
rect 41295 27195 41505 27405
rect 40695 26595 40905 26805
rect 39795 25995 40005 26205
rect 40395 26010 40605 26220
rect 37995 25380 38205 25590
rect 37395 24795 37605 25005
rect 39180 25380 39390 25590
rect 39495 25395 39705 25605
rect 40095 25380 40305 25590
rect 40995 25380 41205 25590
rect 44595 28680 44805 28890
rect 43095 28395 43305 28605
rect 43695 28395 43905 28605
rect 44580 28365 44790 28575
rect 44895 28395 45105 28605
rect 42495 27795 42705 28005
rect 43695 27495 43905 27705
rect 41895 26895 42105 27105
rect 42795 26595 43005 26805
rect 42195 25380 42405 25590
rect 40095 24795 40305 25005
rect 38595 24495 38805 24705
rect 39195 24495 39405 24705
rect 37080 21795 37290 22005
rect 37395 21795 37605 22005
rect 38595 21795 38805 22005
rect 37095 21480 37305 21690
rect 37695 21510 37905 21720
rect 39495 21795 39705 22005
rect 40095 21510 40305 21720
rect 37995 20880 38205 21090
rect 37695 20295 37905 20505
rect 39195 20295 39405 20505
rect 37095 18795 37305 19005
rect 34995 16395 35205 16605
rect 34995 16080 35205 16290
rect 34395 13695 34605 13905
rect 35895 17580 36105 17790
rect 36495 17580 36705 17790
rect 37695 18495 37905 18705
rect 38295 18210 38505 18420
rect 42195 24495 42405 24705
rect 43395 25380 43605 25590
rect 43095 22995 43305 23205
rect 42495 21795 42705 22005
rect 41295 21510 41505 21720
rect 41895 21510 42105 21720
rect 41295 20595 41505 20805
rect 41895 20595 42105 20805
rect 40995 20295 41205 20505
rect 41295 19995 41505 20205
rect 40095 19695 40305 19905
rect 39795 19395 40005 19605
rect 39495 18195 39705 18405
rect 40695 18495 40905 18705
rect 43095 20895 43305 21105
rect 42195 19995 42405 20205
rect 42795 19995 43005 20205
rect 41295 19395 41505 19605
rect 41895 19395 42105 19605
rect 40995 18195 41205 18405
rect 35595 16395 35805 16605
rect 35595 15795 35805 16005
rect 35295 15495 35505 15705
rect 37995 17295 38205 17505
rect 38595 17295 38805 17505
rect 37695 15795 37905 16005
rect 36795 15195 37005 15405
rect 36795 14295 37005 14505
rect 35895 13710 36105 13920
rect 36495 13695 36705 13905
rect 35595 13080 35805 13290
rect 33795 12195 34005 12405
rect 32895 11595 33105 11805
rect 35895 11895 36105 12105
rect 35595 11295 35805 11505
rect 32895 10995 33105 11205
rect 33795 10995 34005 11205
rect 34395 10995 34605 11205
rect 35295 10995 35505 11205
rect 30495 8295 30705 8505
rect 30195 7995 30405 8205
rect 30495 7695 30705 7905
rect 27795 7095 28005 7305
rect 25695 6795 25905 7005
rect 27195 6795 27405 7005
rect 25995 5910 26205 6120
rect 26595 5910 26805 6120
rect 29595 6495 29805 6705
rect 27795 5910 28005 6120
rect 28995 5910 29205 6120
rect 27495 5280 27705 5490
rect 29295 5280 29505 5490
rect 25995 4995 26205 5205
rect 31395 9495 31605 9705
rect 31995 8895 32205 9105
rect 30795 5910 31005 6120
rect 33195 10695 33405 10905
rect 33195 9780 33405 9990
rect 34095 9780 34305 9990
rect 34695 9780 34905 9990
rect 32895 9495 33105 9705
rect 34095 8295 34305 8505
rect 35595 10395 35805 10605
rect 38295 14595 38505 14805
rect 37995 14295 38205 14505
rect 38295 13710 38505 13920
rect 36795 13095 37005 13305
rect 37095 12195 37305 12405
rect 36495 10995 36705 11205
rect 36195 10695 36405 10905
rect 37095 10395 37305 10605
rect 36795 9780 37005 9990
rect 37995 13080 38205 13290
rect 39495 15795 39705 16005
rect 40095 15795 40305 16005
rect 41595 19095 41805 19305
rect 41295 17295 41505 17505
rect 40395 14595 40605 14805
rect 42795 18795 43005 19005
rect 45495 27795 45705 28005
rect 45195 27495 45405 27705
rect 44895 26595 45105 26805
rect 43995 25995 44205 26205
rect 43995 24495 44205 24705
rect 43695 23895 43905 24105
rect 44595 23295 44805 23505
rect 44595 21795 44805 22005
rect 46095 26895 46305 27105
rect 47295 28695 47505 28905
rect 46695 28095 46905 28305
rect 47295 28095 47505 28305
rect 46695 26595 46905 26805
rect 46395 26295 46605 26505
rect 46395 25380 46605 25590
rect 47295 24795 47505 25005
rect 46095 24195 46305 24405
rect 46095 21795 46305 22005
rect 45495 21495 45705 21705
rect 46695 21510 46905 21720
rect 47280 21510 47490 21720
rect 49095 40095 49305 40305
rect 49995 40995 50205 41205
rect 49695 40695 49905 40905
rect 49695 39495 49905 39705
rect 49395 38895 49605 39105
rect 49695 38595 49905 38805
rect 49095 37995 49305 38205
rect 50895 40995 51105 41205
rect 50595 39495 50805 39705
rect 50595 38895 50805 39105
rect 49995 38295 50205 38505
rect 49395 37395 49605 37605
rect 50295 37995 50505 38205
rect 49995 37110 50205 37320
rect 49095 36480 49305 36690
rect 49695 36195 49905 36405
rect 53895 46395 54105 46605
rect 52995 45795 53205 46005
rect 51795 45495 52005 45705
rect 52395 44910 52605 45120
rect 56595 48780 56805 48990
rect 55695 46695 55905 46905
rect 57495 49410 57705 49620
rect 58995 49695 59205 49905
rect 60495 49410 60705 49620
rect 57795 48780 58005 48990
rect 58395 48780 58605 48990
rect 58995 48780 59205 48990
rect 60195 48780 60405 48990
rect 59595 48495 59805 48705
rect 57495 48195 57705 48405
rect 59895 48195 60105 48405
rect 57495 47595 57705 47805
rect 57495 46995 57705 47205
rect 56895 46395 57105 46605
rect 57195 46095 57405 46305
rect 55395 44910 55605 45120
rect 57195 44910 57405 45120
rect 51795 44280 52005 44490
rect 52695 44280 52905 44490
rect 51795 42795 52005 43005
rect 51495 41595 51705 41805
rect 52395 41610 52605 41820
rect 52695 40980 52905 41190
rect 52095 40695 52305 40905
rect 51195 37995 51405 38205
rect 53895 44280 54105 44490
rect 54495 44280 54705 44490
rect 53595 43995 53805 44205
rect 56295 44250 56505 44460
rect 55995 43395 56205 43605
rect 64695 59880 64905 60090
rect 65295 59880 65505 60090
rect 63795 57195 64005 57405
rect 64095 56550 64305 56760
rect 63495 55695 63705 55905
rect 65295 54795 65505 55005
rect 64995 54495 65205 54705
rect 63795 54195 64005 54405
rect 63495 52695 63705 52905
rect 67380 70695 67590 70905
rect 67695 70695 67905 70905
rect 67395 69795 67605 70005
rect 66780 68895 66990 69105
rect 67095 68895 67305 69105
rect 66795 68310 67005 68520
rect 67995 69195 68205 69405
rect 67695 68595 67905 68805
rect 67395 66795 67605 67005
rect 67095 66195 67305 66405
rect 66795 65895 67005 66105
rect 67695 66495 67905 66705
rect 67680 65595 67890 65805
rect 67995 65595 68205 65805
rect 68595 71595 68805 71805
rect 70995 74595 71205 74805
rect 70695 74295 70905 74505
rect 70995 73995 71205 74205
rect 71595 73995 71805 74205
rect 70995 73095 71205 73305
rect 70695 72810 70905 73020
rect 71295 72810 71505 73020
rect 72195 75480 72405 75690
rect 72795 74895 73005 75105
rect 72495 74595 72705 74805
rect 70095 72480 70305 72690
rect 71595 72180 71805 72390
rect 70095 71595 70305 71805
rect 69795 71295 70005 71505
rect 69495 70695 69705 70905
rect 70395 70695 70605 70905
rect 69195 70095 69405 70305
rect 69195 69780 69405 69990
rect 68595 68895 68805 69105
rect 68595 68295 68805 68505
rect 69795 69495 70005 69705
rect 69495 69195 69705 69405
rect 69495 68595 69705 68805
rect 68595 67695 68805 67905
rect 68895 67395 69105 67605
rect 68595 67095 68805 67305
rect 68295 65295 68505 65505
rect 69195 67095 69405 67305
rect 68895 66495 69105 66705
rect 70680 70395 70890 70605
rect 70995 70395 71205 70605
rect 72195 70095 72405 70305
rect 72795 73095 73005 73305
rect 74895 76695 75105 76905
rect 75495 79395 75705 79605
rect 77295 82395 77505 82605
rect 77295 81495 77505 81705
rect 76995 80595 77205 80805
rect 78495 87780 78705 87990
rect 79095 87780 79305 87990
rect 77895 87195 78105 87405
rect 79395 87195 79605 87405
rect 77895 86295 78105 86505
rect 79395 85995 79605 86205
rect 78495 85695 78705 85905
rect 77895 85095 78105 85305
rect 78795 85395 79005 85605
rect 78495 84195 78705 84405
rect 79095 84795 79305 85005
rect 79695 85395 79905 85605
rect 79395 84495 79605 84705
rect 79095 83895 79305 84105
rect 78195 83280 78405 83490
rect 77895 82680 78105 82890
rect 77895 82095 78105 82305
rect 77895 80895 78105 81105
rect 77595 80595 77805 80805
rect 76395 79995 76605 80205
rect 76095 79095 76305 79305
rect 75795 78795 76005 79005
rect 75795 78195 76005 78405
rect 75495 77595 75705 77805
rect 74895 75480 75105 75690
rect 74295 74595 74505 74805
rect 73995 73395 74205 73605
rect 73995 72795 74205 73005
rect 73395 72180 73605 72390
rect 73095 71595 73305 71805
rect 73395 71295 73605 71505
rect 73095 70095 73305 70305
rect 70995 68880 71205 69090
rect 72195 68895 72405 69105
rect 70695 68595 70905 68805
rect 69795 67395 70005 67605
rect 69495 66495 69705 66705
rect 69195 66195 69405 66405
rect 68895 65295 69105 65505
rect 70395 67680 70605 67890
rect 70095 67095 70305 67305
rect 69795 66195 70005 66405
rect 69495 65895 69705 66105
rect 70395 65295 70605 65505
rect 68280 64395 68490 64605
rect 68595 64395 68805 64605
rect 69495 65010 69705 65220
rect 70095 65010 70305 65220
rect 73395 68595 73605 68805
rect 71595 67095 71805 67305
rect 71295 66795 71505 67005
rect 70995 66195 71205 66405
rect 70995 65880 71205 66090
rect 69195 64395 69405 64605
rect 67095 63495 67305 63705
rect 67695 63195 67905 63405
rect 66795 61695 67005 61905
rect 66195 61095 66405 61305
rect 65895 60495 66105 60705
rect 65895 59895 66105 60105
rect 68295 61695 68505 61905
rect 68895 60510 69105 60720
rect 70395 64380 70605 64590
rect 69495 64095 69705 64305
rect 70095 64095 70305 64305
rect 69495 61995 69705 62205
rect 69495 61680 69705 61890
rect 66195 58995 66405 59205
rect 66495 58395 66705 58605
rect 66195 57210 66405 57420
rect 67395 57210 67605 57420
rect 65895 56295 66105 56505
rect 68595 59880 68805 60090
rect 69195 59895 69405 60105
rect 68295 59280 68505 59490
rect 68895 59295 69105 59505
rect 71595 65895 71805 66105
rect 72195 66795 72405 67005
rect 72195 65595 72405 65805
rect 74895 73995 75105 74205
rect 76095 77895 76305 78105
rect 75795 75195 76005 75405
rect 75495 73695 75705 73905
rect 74895 72810 75105 73020
rect 75495 72810 75705 73020
rect 76995 78495 77205 78705
rect 76695 77295 76905 77505
rect 78495 81795 78705 82005
rect 79695 82395 79905 82605
rect 78795 81195 79005 81405
rect 78495 80895 78705 81105
rect 78195 80595 78405 80805
rect 79095 80895 79305 81105
rect 78795 79980 79005 80190
rect 78195 79095 78405 79305
rect 77595 76695 77805 76905
rect 77295 76395 77505 76605
rect 76395 76095 76605 76305
rect 77895 76395 78105 76605
rect 76395 75495 76605 75705
rect 76095 72795 76305 73005
rect 74895 71895 75105 72105
rect 74595 68895 74805 69105
rect 74295 68595 74505 68805
rect 76095 72195 76305 72405
rect 75195 70695 75405 70905
rect 76095 69495 76305 69705
rect 77595 75480 77805 75690
rect 77295 75195 77505 75405
rect 76995 74295 77205 74505
rect 76695 73695 76905 73905
rect 84195 92595 84405 92805
rect 83895 92295 84105 92505
rect 81495 91995 81705 92205
rect 82095 91995 82305 92205
rect 82695 91995 82905 92205
rect 83295 91995 83505 92205
rect 80895 91710 81105 91920
rect 82395 91710 82605 91920
rect 83895 91695 84105 91905
rect 80595 91095 80805 91305
rect 82095 91095 82305 91305
rect 81195 90495 81405 90705
rect 82695 91080 82905 91290
rect 83595 91080 83805 91290
rect 82095 90195 82305 90405
rect 80595 89895 80805 90105
rect 81195 89895 81405 90105
rect 80595 88410 80805 88620
rect 82995 89295 83205 89505
rect 82395 88995 82605 89205
rect 82095 88410 82305 88620
rect 80895 87780 81105 87990
rect 82095 87195 82305 87405
rect 81795 86595 82005 86805
rect 82095 85695 82305 85905
rect 81795 85395 82005 85605
rect 82995 88410 83205 88620
rect 83595 88410 83805 88620
rect 83295 87780 83505 87990
rect 82695 86295 82905 86505
rect 82995 85395 83205 85605
rect 84495 92295 84705 92505
rect 87795 93795 88005 94005
rect 88395 93195 88605 93405
rect 87495 92595 87705 92805
rect 87195 91995 87405 92205
rect 85995 91710 86205 91920
rect 86895 91395 87105 91605
rect 85695 91080 85905 91290
rect 86295 90795 86505 91005
rect 84795 90495 85005 90705
rect 85995 90495 86205 90705
rect 86295 89895 86505 90105
rect 86895 89895 87105 90105
rect 85995 89595 86205 89805
rect 84795 89295 85005 89505
rect 85395 88995 85605 89205
rect 85095 87780 85305 87990
rect 85695 87780 85905 87990
rect 85095 86895 85305 87105
rect 82695 83895 82905 84105
rect 82395 83280 82605 83490
rect 81495 82695 81705 82905
rect 81195 82395 81405 82605
rect 79995 81795 80205 82005
rect 79980 81195 80190 81405
rect 80295 81195 80505 81405
rect 80895 80895 81105 81105
rect 80295 80595 80505 80805
rect 82695 82995 82905 83205
rect 82395 81795 82605 82005
rect 81495 80610 81705 80820
rect 84195 85095 84405 85305
rect 83595 83910 83805 84120
rect 84195 83895 84405 84105
rect 83895 83280 84105 83490
rect 83595 82995 83805 83205
rect 82995 81195 83205 81405
rect 83895 82095 84105 82305
rect 83595 80595 83805 80805
rect 79995 79995 80205 80205
rect 80595 79980 80805 80190
rect 81195 79980 81405 80190
rect 82695 79980 82905 80190
rect 83295 79980 83505 80190
rect 82395 79395 82605 79605
rect 81195 79095 81405 79305
rect 81195 78495 81405 78705
rect 79695 78195 79905 78405
rect 80595 78195 80805 78405
rect 78795 77895 79005 78105
rect 80580 77595 80790 77805
rect 80895 77595 81105 77805
rect 78795 76110 79005 76320
rect 79395 76110 79605 76320
rect 80280 76110 80490 76320
rect 80595 76110 80805 76320
rect 81795 77295 82005 77505
rect 78195 74595 78405 74805
rect 77595 73095 77805 73305
rect 78495 73095 78705 73305
rect 76995 72795 77205 73005
rect 77895 72810 78105 73020
rect 79695 74895 79905 75105
rect 79995 74595 80205 74805
rect 81195 76110 81405 76320
rect 82095 76695 82305 76905
rect 81795 76095 82005 76305
rect 81495 75480 81705 75690
rect 81195 74895 81405 75105
rect 80595 74595 80805 74805
rect 80295 74295 80505 74505
rect 80595 73995 80805 74205
rect 79995 73395 80205 73605
rect 79095 73095 79305 73305
rect 78795 72795 79005 73005
rect 76695 72180 76905 72390
rect 76995 71595 77205 71805
rect 77595 72180 77805 72390
rect 81495 74595 81705 74805
rect 78495 71895 78705 72105
rect 77595 70995 77805 71205
rect 78195 70995 78405 71205
rect 78195 70395 78405 70605
rect 77295 69495 77505 69705
rect 78195 69495 78405 69705
rect 76395 69195 76605 69405
rect 77895 69195 78105 69405
rect 75795 68280 76005 68490
rect 76695 68310 76905 68520
rect 77295 68310 77505 68520
rect 75495 67995 75705 68205
rect 74295 67680 74505 67890
rect 74895 67395 75105 67605
rect 73695 66495 73905 66705
rect 73695 65895 73905 66105
rect 71895 65010 72105 65220
rect 72495 65010 72705 65220
rect 73395 65010 73605 65220
rect 74895 65295 75105 65505
rect 74595 64995 74805 65205
rect 70995 62295 71205 62505
rect 70095 61695 70305 61905
rect 69795 61395 70005 61605
rect 70395 60510 70605 60720
rect 71295 60495 71505 60705
rect 69495 59595 69705 59805
rect 69195 58095 69405 58305
rect 68295 57195 68505 57405
rect 66795 56295 67005 56505
rect 67395 55995 67605 56205
rect 66195 55695 66405 55905
rect 66795 55695 67005 55905
rect 65595 53595 65805 53805
rect 65595 52710 65805 52920
rect 63195 50595 63405 50805
rect 61395 49695 61605 49905
rect 62595 49695 62805 49905
rect 61095 47595 61305 47805
rect 60795 46695 61005 46905
rect 60195 46395 60405 46605
rect 59895 45795 60105 46005
rect 58095 45495 58305 45705
rect 58995 44940 59205 45150
rect 59595 44940 59805 45150
rect 56595 43095 56805 43305
rect 57195 43095 57405 43305
rect 55095 42795 55305 43005
rect 55995 42795 56205 43005
rect 54195 41610 54405 41820
rect 54795 41610 55005 41820
rect 55695 41595 55905 41805
rect 54195 40095 54405 40305
rect 53595 38895 53805 39105
rect 52395 37395 52605 37605
rect 53295 37395 53505 37605
rect 50895 37110 51105 37320
rect 51795 37110 52005 37320
rect 52095 36495 52305 36705
rect 50595 34695 50805 34905
rect 51195 34095 51405 34305
rect 49095 33795 49305 34005
rect 50295 33810 50505 34020
rect 50895 33810 51105 34020
rect 49095 32895 49305 33105
rect 48495 32595 48705 32805
rect 48795 32295 49005 32505
rect 48195 31395 48405 31605
rect 48195 30195 48405 30405
rect 49695 31695 49905 31905
rect 50895 30795 51105 31005
rect 53595 37110 53805 37320
rect 54495 39495 54705 39705
rect 52695 36795 52905 37005
rect 52695 36195 52905 36405
rect 53295 35895 53505 36105
rect 52695 34695 52905 34905
rect 52395 34095 52605 34305
rect 52095 33795 52305 34005
rect 52995 34395 53205 34605
rect 52695 33195 52905 33405
rect 51795 31095 52005 31305
rect 50280 29895 50490 30105
rect 50595 29895 50805 30105
rect 48795 29310 49005 29520
rect 49395 29310 49605 29520
rect 50295 29310 50505 29520
rect 51195 29310 51405 29520
rect 47895 28680 48105 28890
rect 48495 28680 48705 28890
rect 49395 28395 49605 28605
rect 49395 27795 49605 28005
rect 50895 27195 51105 27405
rect 49995 26895 50205 27105
rect 48795 26595 49005 26805
rect 48795 26010 49005 26220
rect 50895 26010 51105 26220
rect 51795 25995 52005 26205
rect 49395 25380 49605 25590
rect 49995 25395 50205 25605
rect 50595 25380 50805 25590
rect 51195 25395 51405 25605
rect 55395 40980 55605 41190
rect 55395 39495 55605 39705
rect 56295 42195 56505 42405
rect 56595 41595 56805 41805
rect 57195 41610 57405 41820
rect 56895 40980 57105 41190
rect 57495 40980 57705 41190
rect 56295 40095 56505 40305
rect 56295 38895 56505 39105
rect 56595 38295 56805 38505
rect 56295 37995 56505 38205
rect 55095 36495 55305 36705
rect 54195 34995 54405 35205
rect 54795 34995 55005 35205
rect 55995 37095 56205 37305
rect 58995 42195 59205 42405
rect 58095 41610 58305 41820
rect 60495 44910 60705 45120
rect 61095 44910 61305 45120
rect 62295 49410 62505 49620
rect 62895 49410 63105 49620
rect 63480 49395 63690 49605
rect 63795 49410 64005 49620
rect 64395 49410 64605 49620
rect 65895 52095 66105 52305
rect 65595 49695 65805 49905
rect 61695 48780 61905 48990
rect 61695 48195 61905 48405
rect 61695 47295 61905 47505
rect 59895 44295 60105 44505
rect 59895 43395 60105 43605
rect 59595 41895 59805 42105
rect 58095 40995 58305 41205
rect 58695 40980 58905 41190
rect 57795 40395 58005 40605
rect 58995 40395 59205 40605
rect 57795 39795 58005 40005
rect 57495 37095 57705 37305
rect 56295 36480 56505 36690
rect 56895 36480 57105 36690
rect 53295 34095 53505 34305
rect 53895 34095 54105 34305
rect 52995 32895 53205 33105
rect 54195 33810 54405 34020
rect 54795 33840 55005 34050
rect 53595 32895 53805 33105
rect 53895 32595 54105 32805
rect 55995 34995 56205 35205
rect 57495 34995 57705 35205
rect 55695 32295 55905 32505
rect 53595 31395 53805 31605
rect 53895 31095 54105 31305
rect 53295 30495 53505 30705
rect 52695 29895 52905 30105
rect 53295 29595 53505 29805
rect 54795 30495 55005 30705
rect 54495 29595 54705 29805
rect 52995 28680 53205 28890
rect 52995 28095 53205 28305
rect 54495 28680 54705 28890
rect 53595 27795 53805 28005
rect 52395 26010 52605 26220
rect 52995 26010 53205 26220
rect 53595 25995 53805 26205
rect 49995 25080 50205 25290
rect 48495 24195 48705 24405
rect 48795 23895 49005 24105
rect 49095 22695 49305 22905
rect 48795 22395 49005 22605
rect 47895 21795 48105 22005
rect 43395 20595 43605 20805
rect 42195 18210 42405 18420
rect 44295 20880 44505 21090
rect 44895 20880 45105 21090
rect 44295 19995 44505 20205
rect 43695 18210 43905 18420
rect 41895 17595 42105 17805
rect 43095 17580 43305 17790
rect 43695 17580 43905 17790
rect 44595 17580 44805 17790
rect 45795 20880 46005 21090
rect 46395 20295 46605 20505
rect 46995 20295 47205 20505
rect 46395 19395 46605 19605
rect 45495 18795 45705 19005
rect 46395 18495 46605 18705
rect 46095 18210 46305 18420
rect 46695 18210 46905 18420
rect 47595 21495 47805 21705
rect 48795 21510 49005 21720
rect 49395 21795 49605 22005
rect 49680 21510 49890 21720
rect 52095 25380 52305 25590
rect 55395 29310 55605 29520
rect 59895 40995 60105 41205
rect 59895 39795 60105 40005
rect 59295 38295 59505 38505
rect 60795 44280 61005 44490
rect 61395 44295 61605 44505
rect 62595 48780 62805 48990
rect 62295 48195 62505 48405
rect 61995 46095 62205 46305
rect 61995 45495 62205 45705
rect 61995 44595 62205 44805
rect 63195 47595 63405 47805
rect 63195 46395 63405 46605
rect 62595 45795 62805 46005
rect 65295 49395 65505 49605
rect 63795 48795 64005 49005
rect 64695 48795 64905 49005
rect 65295 48795 65505 49005
rect 64995 48495 65205 48705
rect 66195 51795 66405 52005
rect 66495 51495 66705 51705
rect 66195 50895 66405 51105
rect 66195 49995 66405 50205
rect 67395 54495 67605 54705
rect 68595 56580 68805 56790
rect 70695 59880 70905 60090
rect 71295 59880 71505 60090
rect 70095 59595 70305 59805
rect 69795 58995 70005 59205
rect 69795 55995 70005 56205
rect 68295 55695 68505 55905
rect 69495 55695 69705 55905
rect 67995 54495 68205 54705
rect 67695 53895 67905 54105
rect 67095 53295 67305 53505
rect 67995 53295 68205 53505
rect 67395 52710 67605 52920
rect 69795 55395 70005 55605
rect 69495 53895 69705 54105
rect 68295 52695 68505 52905
rect 67095 52095 67305 52305
rect 67995 51795 68205 52005
rect 67695 50895 67905 51105
rect 67095 49995 67305 50205
rect 66795 49695 67005 49905
rect 67095 49410 67305 49620
rect 65895 48495 66105 48705
rect 66495 48495 66705 48705
rect 65595 48195 65805 48405
rect 65295 46995 65505 47205
rect 64695 46095 64905 46305
rect 66195 46695 66405 46905
rect 64395 45795 64605 46005
rect 65895 45795 66105 46005
rect 63495 45495 63705 45705
rect 64095 45495 64305 45705
rect 63495 44910 63705 45120
rect 62295 43995 62505 44205
rect 61695 43395 61905 43605
rect 61395 43095 61605 43305
rect 60495 42495 60705 42705
rect 63195 44280 63405 44490
rect 64095 44295 64305 44505
rect 63795 43995 64005 44205
rect 66195 45195 66405 45405
rect 65295 44910 65505 45120
rect 65895 44910 66105 45120
rect 67695 46995 67905 47205
rect 67395 46695 67605 46905
rect 66495 44895 66705 45105
rect 64395 43695 64605 43905
rect 64095 43095 64305 43305
rect 62595 42795 62805 43005
rect 63795 42795 64005 43005
rect 63795 42195 64005 42405
rect 61695 41895 61905 42105
rect 61395 41595 61605 41805
rect 62295 41595 62505 41805
rect 62895 41610 63105 41820
rect 63495 41610 63705 41820
rect 66195 44295 66405 44505
rect 64995 43695 65205 43905
rect 65595 43695 65805 43905
rect 64995 43095 65205 43305
rect 64095 41595 64305 41805
rect 61095 40980 61305 41190
rect 60495 40395 60705 40605
rect 61095 38595 61305 38805
rect 58395 37110 58605 37320
rect 58695 35895 58905 36105
rect 60195 37995 60405 38205
rect 60495 37395 60705 37605
rect 61395 37995 61605 38205
rect 61095 37095 61305 37305
rect 60195 36480 60405 36690
rect 61095 36480 61305 36690
rect 60795 36195 61005 36405
rect 59295 35595 59505 35805
rect 60195 35595 60405 35805
rect 58095 34395 58305 34605
rect 58995 34095 59205 34305
rect 57795 33795 58005 34005
rect 59595 33810 59805 34020
rect 60795 34995 61005 35205
rect 60495 33810 60705 34020
rect 58095 33480 58305 33690
rect 57495 33150 57705 33360
rect 58395 33195 58605 33405
rect 58095 32295 58305 32505
rect 56595 31995 56805 32205
rect 57795 31995 58005 32205
rect 59295 33180 59505 33390
rect 59895 33180 60105 33390
rect 58695 32595 58905 32805
rect 59295 32595 59505 32805
rect 60195 32595 60405 32805
rect 58995 32295 59205 32505
rect 58695 31695 58905 31905
rect 58695 29595 58905 29805
rect 55695 28680 55905 28890
rect 55695 27495 55905 27705
rect 54795 26895 55005 27105
rect 54195 26595 54405 26805
rect 51195 23295 51405 23505
rect 51495 22695 51705 22905
rect 51195 21795 51405 22005
rect 47595 20895 47805 21105
rect 48180 20895 48390 21105
rect 47295 19995 47505 20205
rect 46395 17580 46605 17790
rect 46995 17595 47205 17805
rect 42495 17295 42705 17505
rect 45195 17295 45405 17505
rect 43395 15495 43605 15705
rect 41895 15195 42105 15405
rect 42495 14595 42705 14805
rect 47295 15495 47505 15705
rect 46995 14895 47205 15105
rect 45795 14595 46005 14805
rect 43395 14295 43605 14505
rect 44895 14295 45105 14505
rect 39795 13080 40005 13290
rect 38895 12795 39105 13005
rect 39495 12795 39705 13005
rect 38295 11295 38505 11505
rect 38895 10410 39105 10620
rect 37995 9780 38205 9990
rect 36195 9195 36405 9405
rect 37395 9195 37605 9405
rect 35295 7995 35505 8205
rect 38595 7995 38805 8205
rect 35295 7095 35505 7305
rect 35595 6495 35805 6705
rect 36795 6495 37005 6705
rect 39195 6495 39405 6705
rect 33195 6195 33405 6405
rect 33495 5910 33705 6120
rect 36195 5910 36405 6120
rect 38595 5910 38805 6120
rect 31395 5280 31605 5490
rect 31995 5280 32205 5490
rect 32580 5280 32790 5490
rect 32895 5280 33105 5490
rect 33795 5280 34005 5490
rect 34395 5280 34605 5490
rect 35595 5295 35805 5505
rect 30495 4995 30705 5205
rect 31095 4695 31305 4905
rect 25995 4395 26205 4605
rect 26595 4395 26805 4605
rect 25695 4095 25905 4305
rect 24495 3195 24705 3405
rect 25395 3195 25605 3405
rect 24795 2895 25005 3105
rect 24195 2595 24405 2805
rect 22695 1980 22905 2190
rect 23295 1980 23505 2190
rect 29895 4095 30105 4305
rect 30195 3795 30405 4005
rect 31695 3795 31905 4005
rect 26895 3195 27105 3405
rect 29895 3195 30105 3405
rect 25995 2610 26205 2820
rect 25695 1980 25905 2190
rect 23895 1395 24105 1605
rect 24795 1395 25005 1605
rect 22395 1095 22605 1305
rect 26295 1695 26505 1905
rect 29295 2895 29505 3105
rect 27795 2610 28005 2820
rect 28395 2610 28605 2820
rect 28995 2595 29205 2805
rect 27495 1980 27705 2190
rect 28095 1980 28305 2190
rect 31395 3195 31605 3405
rect 30795 2610 31005 2820
rect 29295 1980 29505 2190
rect 29895 1980 30105 2190
rect 30495 1980 30705 2190
rect 31095 1980 31305 2190
rect 37095 5280 37305 5490
rect 38295 5280 38505 5490
rect 39195 5295 39405 5505
rect 38895 4095 39105 4305
rect 38295 3795 38505 4005
rect 33795 3495 34005 3705
rect 36495 3495 36705 3705
rect 33195 3195 33405 3405
rect 32595 2895 32805 3105
rect 31695 1980 31905 2190
rect 36195 3195 36405 3405
rect 36795 3195 37005 3405
rect 36495 2895 36705 3105
rect 34395 2610 34605 2820
rect 35295 2610 35505 2820
rect 37095 2610 37305 2820
rect 37995 2610 38205 2820
rect 28995 1395 29205 1605
rect 26895 1095 27105 1305
rect 25695 795 25905 1005
rect 32295 1980 32505 2190
rect 32895 1980 33105 2190
rect 33795 1980 34005 2190
rect 34695 1980 34905 2190
rect 36195 1695 36405 1905
rect 35295 1395 35505 1605
rect 39795 11895 40005 12105
rect 41295 13080 41505 13290
rect 40395 11295 40605 11505
rect 40395 10980 40605 11190
rect 40695 10695 40905 10905
rect 40395 9780 40605 9990
rect 40995 8595 41205 8805
rect 39795 8295 40005 8505
rect 39795 7695 40005 7905
rect 41295 6795 41505 7005
rect 44295 13710 44505 13920
rect 46695 14295 46905 14505
rect 46695 13710 46905 13920
rect 43995 13080 44205 13290
rect 45795 13080 46005 13290
rect 46395 13080 46605 13290
rect 46995 12495 47205 12705
rect 44595 12195 44805 12405
rect 46995 11895 47205 12105
rect 45195 10995 45405 11205
rect 44895 10695 45105 10905
rect 44595 10395 44805 10605
rect 42195 9795 42405 10005
rect 42795 9780 43005 9990
rect 43695 9195 43905 9405
rect 46395 10410 46605 10620
rect 47895 19995 48105 20205
rect 48495 20880 48705 21090
rect 49080 20880 49290 21090
rect 49395 20895 49605 21105
rect 49995 21495 50205 21705
rect 50595 21510 50805 21720
rect 50295 20880 50505 21090
rect 50895 20880 51105 21090
rect 51495 20895 51705 21105
rect 49695 20295 49905 20505
rect 49995 19095 50205 19305
rect 48495 18795 48705 19005
rect 48195 18495 48405 18705
rect 47895 18195 48105 18405
rect 48195 17580 48405 17790
rect 48795 17580 49005 17790
rect 47895 17295 48105 17505
rect 48795 13995 49005 14205
rect 51195 18495 51405 18705
rect 50295 18195 50505 18405
rect 50895 18210 51105 18420
rect 52695 25380 52905 25590
rect 53895 25380 54105 25590
rect 53295 24495 53505 24705
rect 54195 23295 54405 23505
rect 52695 22395 52905 22605
rect 52095 21510 52305 21720
rect 53295 21510 53505 21720
rect 54795 23895 55005 24105
rect 54495 22095 54705 22305
rect 55995 22395 56205 22605
rect 55395 21510 55605 21720
rect 52395 20895 52605 21105
rect 52095 20295 52305 20505
rect 51795 19095 52005 19305
rect 54195 20895 54405 21105
rect 55695 20895 55905 21105
rect 53595 20295 53805 20505
rect 54495 20295 54705 20505
rect 55095 20295 55305 20505
rect 52995 19395 53205 19605
rect 54195 19395 54405 19605
rect 53595 18795 53805 19005
rect 52395 18495 52605 18705
rect 52995 18495 53205 18705
rect 52095 18195 52305 18405
rect 49995 17895 50205 18105
rect 51195 17580 51405 17790
rect 52395 17580 52605 17790
rect 53295 17580 53505 17790
rect 53895 17580 54105 17790
rect 54495 17580 54705 17790
rect 51795 16995 52005 17205
rect 53895 15495 54105 15705
rect 53295 14895 53505 15105
rect 50295 13995 50505 14205
rect 49695 13710 49905 13920
rect 50895 13710 51105 13920
rect 55395 17580 55605 17790
rect 55995 17295 56205 17505
rect 55395 16995 55605 17205
rect 56895 29310 57105 29520
rect 57495 29310 57705 29520
rect 58395 29310 58605 29520
rect 56595 28095 56805 28305
rect 57195 27795 57405 28005
rect 56895 26895 57105 27105
rect 58395 28095 58605 28305
rect 57795 26595 58005 26805
rect 59895 31095 60105 31305
rect 59295 29310 59505 29520
rect 60495 28695 60705 28905
rect 59595 28095 59805 28305
rect 63195 40395 63405 40605
rect 64095 40995 64305 41205
rect 63795 40095 64005 40305
rect 62595 39195 62805 39405
rect 61695 37395 61905 37605
rect 62295 37395 62505 37605
rect 63195 37110 63405 37320
rect 64095 37110 64305 37320
rect 61695 36495 61905 36705
rect 62295 36195 62505 36405
rect 62895 35295 63105 35505
rect 64695 42195 64905 42405
rect 66795 44250 67005 44460
rect 66495 43095 66705 43305
rect 70695 56580 70905 56790
rect 72195 64380 72405 64590
rect 73995 64380 74205 64590
rect 72795 63795 73005 64005
rect 73395 63795 73605 64005
rect 74295 63795 74505 64005
rect 71895 63195 72105 63405
rect 72495 63195 72705 63405
rect 71895 62595 72105 62805
rect 71895 62280 72105 62490
rect 73095 61395 73305 61605
rect 72495 60510 72705 60720
rect 73995 62295 74205 62505
rect 73995 61695 74205 61905
rect 75795 67395 76005 67605
rect 75795 65595 76005 65805
rect 75495 65295 75705 65505
rect 76395 67095 76605 67305
rect 77595 67695 77805 67905
rect 76395 66495 76605 66705
rect 76995 66495 77205 66705
rect 76095 65295 76305 65505
rect 76995 65895 77205 66105
rect 76695 65595 76905 65805
rect 76395 65010 76605 65220
rect 75195 64395 75405 64605
rect 74895 63195 75105 63405
rect 75795 63795 76005 64005
rect 75495 63495 75705 63705
rect 75795 62595 76005 62805
rect 76395 64095 76605 64305
rect 76095 61995 76305 62205
rect 75195 61695 75405 61905
rect 74595 61095 74805 61305
rect 76095 61095 76305 61305
rect 73395 60495 73605 60705
rect 72495 59595 72705 59805
rect 71895 58995 72105 59205
rect 72795 59295 73005 59505
rect 73095 58995 73305 59205
rect 71595 54495 71805 54705
rect 71895 53895 72105 54105
rect 70395 53295 70605 53505
rect 70095 52695 70305 52905
rect 71295 52740 71505 52950
rect 69495 51795 69705 52005
rect 68595 50595 68805 50805
rect 68295 49695 68505 49905
rect 69195 49695 69405 49905
rect 68595 49410 68805 49620
rect 68295 48795 68505 49005
rect 68895 48780 69105 48990
rect 68295 48195 68505 48405
rect 69495 48195 69705 48405
rect 70395 51795 70605 52005
rect 71895 51495 72105 51705
rect 72195 50895 72405 51105
rect 73695 58695 73905 58905
rect 73395 58095 73605 58305
rect 75195 58695 75405 58905
rect 77295 64995 77505 65205
rect 78195 66495 78405 66705
rect 77895 65895 78105 66105
rect 78195 65010 78405 65220
rect 79095 72180 79305 72390
rect 79695 72180 79905 72390
rect 81195 72180 81405 72390
rect 80295 71595 80505 71805
rect 78795 70995 79005 71205
rect 80595 70995 80805 71205
rect 78795 70395 79005 70605
rect 80295 69795 80505 70005
rect 80295 68895 80505 69105
rect 79695 68595 79905 68805
rect 79095 68310 79305 68520
rect 81195 68895 81405 69105
rect 80595 68295 80805 68505
rect 81795 73095 82005 73305
rect 82695 77895 82905 78105
rect 82395 76095 82605 76305
rect 85695 86295 85905 86505
rect 86895 89580 87105 89790
rect 87795 89295 88005 89505
rect 87495 88410 87705 88620
rect 88095 87795 88305 88005
rect 87795 87195 88005 87405
rect 87195 86895 87405 87105
rect 86295 85395 86505 85605
rect 87795 85395 88005 85605
rect 85695 85095 85905 85305
rect 85095 83895 85305 84105
rect 87495 84495 87705 84705
rect 91095 93795 91305 94005
rect 89995 93195 90205 93405
rect 88995 91995 89205 92205
rect 88395 87495 88605 87705
rect 88095 84495 88305 84705
rect 86295 83910 86505 84120
rect 87495 83910 87705 84120
rect 85095 83295 85305 83505
rect 86895 83295 87105 83505
rect 85995 82995 86205 83205
rect 84795 82095 85005 82305
rect 83895 77295 84105 77505
rect 84495 81195 84705 81405
rect 85395 81195 85605 81405
rect 85995 81195 86205 81405
rect 84795 80610 85005 80820
rect 87795 83280 88005 83490
rect 89295 90795 89505 91005
rect 88995 89595 89205 89805
rect 88995 88995 89205 89205
rect 89595 89895 89805 90105
rect 90495 88995 90705 89205
rect 89295 88410 89505 88620
rect 89595 87780 89805 87990
rect 90495 87795 90705 88005
rect 89295 87495 89505 87705
rect 88995 85095 89205 85305
rect 87495 82695 87705 82905
rect 88095 82695 88305 82905
rect 87195 81795 87405 82005
rect 86295 80895 86505 81105
rect 86895 80895 87105 81105
rect 85095 79395 85305 79605
rect 85995 79995 86205 80205
rect 85695 79095 85905 79305
rect 87495 80595 87705 80805
rect 87195 79980 87405 80190
rect 87795 79995 88005 80205
rect 87195 79395 87405 79605
rect 86895 79095 87105 79305
rect 86295 78795 86505 79005
rect 86595 78495 86805 78705
rect 85995 77895 86205 78105
rect 85095 77595 85305 77805
rect 84195 76695 84405 76905
rect 82995 75480 83205 75690
rect 83595 75480 83805 75690
rect 84195 75480 84405 75690
rect 82695 72810 82905 73020
rect 83895 73995 84105 74205
rect 83595 73095 83805 73305
rect 83295 72795 83505 73005
rect 81495 68595 81705 68805
rect 82395 72180 82605 72390
rect 82095 70395 82305 70605
rect 81795 68310 82005 68520
rect 83295 72195 83505 72405
rect 83295 70395 83505 70605
rect 82995 69495 83205 69705
rect 85095 76995 85305 77205
rect 85695 76110 85905 76320
rect 85395 75480 85605 75690
rect 85995 74895 86205 75105
rect 84795 74595 85005 74805
rect 85695 74595 85905 74805
rect 84495 73395 84705 73605
rect 84195 73095 84405 73305
rect 83895 72795 84105 73005
rect 85395 74295 85605 74505
rect 86295 74295 86505 74505
rect 88995 83295 89205 83505
rect 89895 84495 90105 84705
rect 91695 89295 91905 89505
rect 91395 87795 91605 88005
rect 90195 83295 90405 83505
rect 89295 82695 89505 82905
rect 89895 82095 90105 82305
rect 89295 81195 89505 81405
rect 88995 79980 89205 80190
rect 88395 79395 88605 79605
rect 88095 78495 88305 78705
rect 87795 76995 88005 77205
rect 91095 83295 91305 83505
rect 91395 82095 91605 82305
rect 90495 81495 90705 81705
rect 91395 81495 91605 81705
rect 91995 85395 92205 85605
rect 91695 80595 91905 80805
rect 91695 79995 91905 80205
rect 90195 79095 90405 79305
rect 90795 79095 91005 79305
rect 90795 78195 91005 78405
rect 90495 77895 90705 78105
rect 89895 76695 90105 76905
rect 91395 76695 91605 76905
rect 88395 76395 88605 76605
rect 89595 76395 89805 76605
rect 87795 76110 88005 76320
rect 90495 76110 90705 76320
rect 91095 76110 91305 76320
rect 89595 75480 89805 75690
rect 88995 75195 89205 75405
rect 87495 74895 87705 75105
rect 88095 74895 88305 75105
rect 88695 74895 88905 75105
rect 87195 74295 87405 74505
rect 86895 73995 87105 74205
rect 85695 73380 85905 73590
rect 85395 72795 85605 73005
rect 84495 72180 84705 72390
rect 85395 72195 85605 72405
rect 84495 71595 84705 71805
rect 84795 70095 85005 70305
rect 84495 69795 84705 70005
rect 82695 69195 82905 69405
rect 83595 69195 83805 69405
rect 82395 68295 82605 68505
rect 78795 67695 79005 67905
rect 78795 67095 79005 67305
rect 79095 65595 79305 65805
rect 77295 63495 77505 63705
rect 77595 63195 77805 63405
rect 76995 61395 77205 61605
rect 77595 61395 77805 61605
rect 76695 60795 76905 61005
rect 77295 60795 77505 61005
rect 80295 67695 80505 67905
rect 79995 66795 80205 67005
rect 79995 65010 80205 65220
rect 80895 67395 81105 67605
rect 82095 67695 82305 67905
rect 80595 67095 80805 67305
rect 79095 64395 79305 64605
rect 79695 64380 79905 64590
rect 78795 64095 79005 64305
rect 79695 63495 79905 63705
rect 80895 66495 81105 66705
rect 82095 67095 82305 67305
rect 81195 65010 81405 65220
rect 81795 65010 82005 65220
rect 83295 68895 83505 69105
rect 84195 68310 84405 68520
rect 84795 69195 85005 69405
rect 82995 67395 83205 67605
rect 82695 66795 82905 67005
rect 82395 64995 82605 65205
rect 80595 62895 80805 63105
rect 82095 64380 82305 64590
rect 82095 64065 82305 64275
rect 80895 61995 81105 62205
rect 81495 61995 81705 62205
rect 78195 61695 78405 61905
rect 80295 61695 80505 61905
rect 76395 59880 76605 60090
rect 76995 59880 77205 60090
rect 76695 59295 76905 59505
rect 76395 58995 76605 59205
rect 76395 58395 76605 58605
rect 76095 58095 76305 58305
rect 75195 57795 75405 58005
rect 73395 56580 73605 56790
rect 73995 56580 74205 56790
rect 73995 56265 74205 56475
rect 73395 53895 73605 54105
rect 73395 53295 73605 53505
rect 71595 50295 71805 50505
rect 70995 49995 71205 50205
rect 72495 49695 72705 49905
rect 72195 49395 72405 49605
rect 71295 48780 71505 48990
rect 70395 48195 70605 48405
rect 71595 48195 71805 48405
rect 70095 47895 70305 48105
rect 71295 47895 71505 48105
rect 69795 46095 70005 46305
rect 69495 45495 69705 45705
rect 68595 44940 68805 45150
rect 69795 44895 70005 45105
rect 68295 44295 68505 44505
rect 69795 44295 70005 44505
rect 68295 43695 68505 43905
rect 67995 43395 68205 43605
rect 68895 42795 69105 43005
rect 67995 42495 68205 42705
rect 67695 42195 67905 42405
rect 68295 42195 68505 42405
rect 66795 41595 67005 41805
rect 67695 41610 67905 41820
rect 65595 40980 65805 41190
rect 66495 40995 66705 41205
rect 66195 40395 66405 40605
rect 64995 38595 65205 38805
rect 65895 38595 66105 38805
rect 65895 38280 66105 38490
rect 64695 37995 64905 38205
rect 65895 37095 66105 37305
rect 64095 34995 64305 35205
rect 61695 34695 61905 34905
rect 62295 34695 62505 34905
rect 62895 34695 63105 34905
rect 64395 34695 64605 34905
rect 61395 34095 61605 34305
rect 61995 33180 62205 33390
rect 61395 32895 61605 33105
rect 61095 31695 61305 31905
rect 62295 30195 62505 30405
rect 61395 29595 61605 29805
rect 62595 29895 62805 30105
rect 61395 28680 61605 28890
rect 59595 27780 59805 27990
rect 60795 27795 61005 28005
rect 57495 26010 57705 26220
rect 58395 26010 58605 26220
rect 58995 26010 59205 26220
rect 60795 27480 61005 27690
rect 59895 26895 60105 27105
rect 57795 25380 58005 25590
rect 59595 25995 59805 26205
rect 58695 25395 58905 25605
rect 57195 23895 57405 24105
rect 57795 23895 58005 24105
rect 56895 22695 57105 22905
rect 56595 21510 56805 21720
rect 57195 21510 57405 21720
rect 56595 20595 56805 20805
rect 56895 20295 57105 20505
rect 57795 20295 58005 20505
rect 58695 24195 58905 24405
rect 59595 25395 59805 25605
rect 59295 21795 59505 22005
rect 58995 21510 59205 21720
rect 59595 21510 59805 21720
rect 61095 26895 61305 27105
rect 60795 26295 61005 26505
rect 60495 26010 60705 26220
rect 61995 26595 62205 26805
rect 63195 34095 63405 34305
rect 63795 33810 64005 34020
rect 64995 36480 65205 36690
rect 65595 36480 65805 36690
rect 66495 39495 66705 39705
rect 66795 39195 67005 39405
rect 67995 40980 68205 41190
rect 68595 40995 68805 41205
rect 68595 40395 68805 40605
rect 67995 38595 68205 38805
rect 67395 38295 67605 38505
rect 66795 37995 67005 38205
rect 67395 37695 67605 37905
rect 66795 37110 67005 37320
rect 70395 44250 70605 44460
rect 70095 42795 70305 43005
rect 69795 42195 70005 42405
rect 69495 41610 69705 41820
rect 71295 42795 71505 43005
rect 71895 46695 72105 46905
rect 71895 44895 72105 45105
rect 75195 55995 75405 56205
rect 76395 57210 76605 57420
rect 80595 60795 80805 61005
rect 78795 60510 79005 60720
rect 78495 59895 78705 60105
rect 78195 58695 78405 58905
rect 79095 59295 79305 59505
rect 78795 58695 79005 58905
rect 78495 57795 78705 58005
rect 75795 56595 76005 56805
rect 75495 55095 75705 55305
rect 75195 54795 75405 55005
rect 75195 54195 75405 54405
rect 76995 55995 77205 56205
rect 76095 55395 76305 55605
rect 74895 52740 75105 52950
rect 76695 53295 76905 53505
rect 75495 52695 75705 52905
rect 75180 52095 75390 52305
rect 73395 50295 73605 50505
rect 73095 49695 73305 49905
rect 73695 49695 73905 49905
rect 74595 49395 74805 49605
rect 73995 48780 74205 48990
rect 74595 48495 74805 48705
rect 73095 47595 73305 47805
rect 74295 47595 74505 47805
rect 73395 47295 73605 47505
rect 73995 47295 74205 47505
rect 72795 46395 73005 46605
rect 73095 45495 73305 45705
rect 73695 46695 73905 46905
rect 73395 45195 73605 45405
rect 73095 44940 73305 45150
rect 73395 44280 73605 44490
rect 73395 43395 73605 43605
rect 72495 42795 72705 43005
rect 70995 42495 71205 42705
rect 71595 42495 71805 42705
rect 70695 42195 70905 42405
rect 70395 41595 70605 41805
rect 69795 40980 70005 41190
rect 70395 40995 70605 41205
rect 69495 39195 69705 39405
rect 69195 38895 69405 39105
rect 69195 37995 69405 38205
rect 69495 37695 69705 37905
rect 68295 37395 68505 37605
rect 68895 37410 69105 37620
rect 67995 36795 68205 37005
rect 65295 36195 65505 36405
rect 65295 35595 65505 35805
rect 64995 35295 65205 35505
rect 64695 33795 64905 34005
rect 64095 33180 64305 33390
rect 65295 33795 65505 34005
rect 66195 36480 66405 36690
rect 67095 36480 67305 36690
rect 67095 34995 67305 35205
rect 67995 34995 68205 35205
rect 66495 33810 66705 34020
rect 65595 32295 65805 32505
rect 64995 31395 65205 31605
rect 67095 33195 67305 33405
rect 66795 31695 67005 31905
rect 63195 31095 63405 31305
rect 66195 31095 66405 31305
rect 67395 31695 67605 31905
rect 63795 29895 64005 30105
rect 64695 29895 64905 30105
rect 63705 29595 63915 29805
rect 63195 29295 63405 29505
rect 64095 29310 64305 29520
rect 67095 29880 67305 30090
rect 64995 29595 65205 29805
rect 65895 29310 66105 29520
rect 66495 29310 66705 29520
rect 64995 28995 65205 29205
rect 63795 28680 64005 28890
rect 64695 28695 64905 28905
rect 63195 28095 63405 28305
rect 64395 28095 64605 28305
rect 62895 26295 63105 26505
rect 64095 27795 64305 28005
rect 60795 25380 61005 25590
rect 61995 25380 62205 25590
rect 60495 25095 60705 25305
rect 61395 25095 61605 25305
rect 58695 20880 58905 21090
rect 58095 19995 58305 20205
rect 59295 20295 59505 20505
rect 58695 19695 58905 19905
rect 62595 25380 62805 25590
rect 63495 25095 63705 25305
rect 62295 24795 62505 25005
rect 62595 22695 62805 22905
rect 61095 21510 61305 21720
rect 61995 21510 62205 21720
rect 60495 20880 60705 21090
rect 61395 20880 61605 21090
rect 65295 28695 65505 28905
rect 64995 28395 65205 28605
rect 64695 27195 64905 27405
rect 65595 28395 65805 28605
rect 66495 28395 66705 28605
rect 66195 27795 66405 28005
rect 65295 26595 65505 26805
rect 66195 26595 66405 26805
rect 64395 26295 64605 26505
rect 65295 26010 65505 26220
rect 65295 24795 65505 25005
rect 64995 24195 65205 24405
rect 65595 23895 65805 24105
rect 65295 23595 65505 23805
rect 64395 23295 64605 23505
rect 64695 22395 64905 22605
rect 62895 22095 63105 22305
rect 64095 22095 64305 22305
rect 62595 19095 62805 19305
rect 58395 18795 58605 19005
rect 59295 18795 59505 19005
rect 60195 18795 60405 19005
rect 57195 18210 57405 18420
rect 57795 18210 58005 18420
rect 59895 18210 60105 18420
rect 61695 18795 61905 19005
rect 60795 18195 61005 18405
rect 62295 18210 62505 18420
rect 58995 17580 59205 17790
rect 59595 17580 59805 17790
rect 60495 17580 60705 17790
rect 57495 17295 57705 17505
rect 56295 15495 56505 15705
rect 55095 14895 55305 15105
rect 54795 13995 55005 14205
rect 55695 13995 55905 14205
rect 56295 13695 56505 13905
rect 54495 13395 54705 13605
rect 47595 13080 47805 13290
rect 49095 13080 49305 13290
rect 49995 13080 50205 13290
rect 50595 13080 50805 13290
rect 47595 11595 47805 11805
rect 48495 11595 48705 11805
rect 51795 13080 52005 13290
rect 52995 13080 53205 13290
rect 53595 13080 53805 13290
rect 55395 13080 55605 13290
rect 48195 10995 48405 11205
rect 48795 10995 49005 11205
rect 50295 10995 50505 11205
rect 51195 10995 51405 11205
rect 50895 10410 51105 10620
rect 51495 10395 51705 10605
rect 44895 9780 45105 9990
rect 45495 9780 45705 9990
rect 44595 8895 44805 9105
rect 44295 8595 44505 8805
rect 42495 6495 42705 6705
rect 42795 6495 43005 6705
rect 41295 5910 41505 6120
rect 47895 9780 48105 9990
rect 48495 9780 48705 9990
rect 49095 9195 49305 9405
rect 49995 9195 50205 9405
rect 51495 9495 51705 9705
rect 52695 12495 52905 12705
rect 53295 12195 53505 12405
rect 53895 12195 54105 12405
rect 55995 12195 56205 12405
rect 53295 10995 53505 11205
rect 54495 11595 54705 11805
rect 54195 10995 54405 11205
rect 54195 10395 54405 10605
rect 55095 10695 55305 10905
rect 55995 10695 56205 10905
rect 52995 9780 53205 9990
rect 53895 9795 54105 10005
rect 54795 9780 55005 9990
rect 55395 9780 55605 9990
rect 56295 10395 56505 10605
rect 59295 16995 59505 17205
rect 59295 16095 59505 16305
rect 57495 14595 57705 14805
rect 58095 13710 58305 13920
rect 60495 14295 60705 14505
rect 59895 13710 60105 13920
rect 61995 17295 62205 17505
rect 63795 21510 64005 21720
rect 68895 37095 69105 37305
rect 70695 39495 70905 39705
rect 72195 42195 72405 42405
rect 71595 41610 71805 41820
rect 75795 52050 76005 52260
rect 76095 50895 76305 51105
rect 75495 50295 75705 50505
rect 75495 49410 75705 49620
rect 75195 48795 75405 49005
rect 74895 48195 75105 48405
rect 75495 48195 75705 48405
rect 74595 46095 74805 46305
rect 74595 45495 74805 45705
rect 75195 45495 75405 45705
rect 74295 44895 74505 45105
rect 74880 44910 75090 45120
rect 75195 44895 75405 45105
rect 73695 42195 73905 42405
rect 72495 41595 72705 41805
rect 71295 40995 71505 41205
rect 70395 38595 70605 38805
rect 69795 36480 70005 36690
rect 70395 36480 70605 36690
rect 72495 40995 72705 41205
rect 72195 40695 72405 40905
rect 71895 40395 72105 40605
rect 72195 40095 72405 40305
rect 71295 38295 71505 38505
rect 71595 37110 71805 37320
rect 73695 40950 73905 41160
rect 72795 40695 73005 40905
rect 74295 40695 74505 40905
rect 76395 47295 76605 47505
rect 77295 55695 77505 55905
rect 77295 55095 77505 55305
rect 79095 58395 79305 58605
rect 79395 58095 79605 58305
rect 79095 57495 79305 57705
rect 78795 56595 79005 56805
rect 79095 55995 79305 56205
rect 78795 54795 79005 55005
rect 78195 54195 78405 54405
rect 78795 54195 79005 54405
rect 77595 52995 77805 53205
rect 77295 52695 77505 52905
rect 77895 52695 78105 52905
rect 79095 53895 79305 54105
rect 77295 52095 77505 52305
rect 78795 52095 79005 52305
rect 76995 50895 77205 51105
rect 76995 50295 77205 50505
rect 84495 67695 84705 67905
rect 83595 66795 83805 67005
rect 83895 66195 84105 66405
rect 84495 66195 84705 66405
rect 84495 65595 84705 65805
rect 84795 65295 85005 65505
rect 86295 73095 86505 73305
rect 88095 74295 88305 74505
rect 86595 72810 86805 73020
rect 87195 72810 87405 73020
rect 86295 72195 86505 72405
rect 87495 72180 87705 72390
rect 86895 71595 87105 71805
rect 85095 64995 85305 65205
rect 82995 64380 83205 64590
rect 83595 64380 83805 64590
rect 84195 64095 84405 64305
rect 84495 64095 84705 64305
rect 83295 63495 83505 63705
rect 83895 63495 84105 63705
rect 82695 62595 82905 62805
rect 82995 61995 83205 62205
rect 82095 61395 82305 61605
rect 82995 60795 83205 61005
rect 83595 62595 83805 62805
rect 80895 60180 81105 60390
rect 80595 57195 80805 57405
rect 79695 56295 79905 56505
rect 79395 53295 79605 53505
rect 79395 52980 79605 53190
rect 79395 52080 79605 52290
rect 79095 51195 79305 51405
rect 78795 50895 79005 51105
rect 78795 50580 79005 50790
rect 78195 49995 78405 50205
rect 77295 49380 77505 49590
rect 80295 55995 80505 56205
rect 81195 57795 81405 58005
rect 82095 57795 82305 58005
rect 82995 57795 83205 58005
rect 82395 57495 82605 57705
rect 81795 57210 82005 57420
rect 82695 57210 82905 57420
rect 84195 61095 84405 61305
rect 84195 60495 84405 60705
rect 85095 64395 85305 64605
rect 85095 63495 85305 63705
rect 84795 63195 85005 63405
rect 85695 69495 85905 69705
rect 87495 69495 87705 69705
rect 85695 68595 85905 68805
rect 85695 67395 85905 67605
rect 87495 67395 87705 67605
rect 85695 66495 85905 66705
rect 87195 66495 87405 66705
rect 85695 65895 85905 66105
rect 86595 65895 86805 66105
rect 85995 65295 86205 65505
rect 86595 65010 86805 65220
rect 85695 64395 85905 64605
rect 83895 59895 84105 60105
rect 84495 58095 84705 58305
rect 83895 57795 84105 58005
rect 81195 55995 81405 56205
rect 82695 55995 82905 56205
rect 82095 55695 82305 55905
rect 81495 52995 81705 53205
rect 80895 52695 81105 52905
rect 80595 52080 80805 52290
rect 81195 51495 81405 51705
rect 80895 51195 81105 51405
rect 79995 50595 80205 50805
rect 79695 49995 79905 50205
rect 79695 49410 79905 49620
rect 76995 47895 77205 48105
rect 75795 46695 76005 46905
rect 76095 46395 76305 46605
rect 75795 45795 76005 46005
rect 75495 43995 75705 44205
rect 76095 43695 76305 43905
rect 75495 41895 75705 42105
rect 76095 41595 76305 41805
rect 75795 40995 76005 41205
rect 73695 40095 73905 40305
rect 74295 40095 74505 40305
rect 72495 37395 72705 37605
rect 73095 37395 73305 37605
rect 74295 39495 74505 39705
rect 73995 38895 74205 39105
rect 74895 38295 75105 38505
rect 74595 37995 74805 38205
rect 72495 36795 72705 37005
rect 70695 36195 70905 36405
rect 69795 35595 70005 35805
rect 70695 34995 70905 35205
rect 68595 33810 68805 34020
rect 69495 33795 69705 34005
rect 69195 33150 69405 33360
rect 68895 32295 69105 32505
rect 69195 31995 69405 32205
rect 69195 31395 69405 31605
rect 70695 31395 70905 31605
rect 68895 31095 69105 31305
rect 68295 30195 68505 30405
rect 67995 29595 68205 29805
rect 70695 30495 70905 30705
rect 69195 30195 69405 30405
rect 68895 29295 69105 29505
rect 68295 28680 68505 28890
rect 67695 28095 67905 28305
rect 67095 27795 67305 28005
rect 67095 27195 67305 27405
rect 67695 26010 67905 26220
rect 68295 28095 68505 28305
rect 66195 25095 66405 25305
rect 67395 25095 67605 25305
rect 67695 24795 67905 25005
rect 71895 36480 72105 36690
rect 71295 36195 71505 36405
rect 72195 34995 72405 35205
rect 72195 34680 72405 34890
rect 71595 33810 71805 34020
rect 73095 34095 73305 34305
rect 72495 33810 72705 34020
rect 72795 32595 73005 32805
rect 71895 32295 72105 32505
rect 72495 31995 72705 32205
rect 71295 30795 71505 31005
rect 69495 29595 69705 29805
rect 70995 29595 71205 29805
rect 69795 29295 70005 29505
rect 70395 29310 70605 29520
rect 69495 28095 69705 28305
rect 69195 27795 69405 28005
rect 69495 27195 69705 27405
rect 68895 26295 69105 26505
rect 70395 26595 70605 26805
rect 69795 26295 70005 26505
rect 68880 25380 69090 25590
rect 69195 25395 69405 25605
rect 68295 23895 68505 24105
rect 66195 22395 66405 22605
rect 64995 21795 65205 22005
rect 65895 21795 66105 22005
rect 64095 20295 64305 20505
rect 68595 21795 68805 22005
rect 67995 21510 68205 21720
rect 68895 21495 69105 21705
rect 66495 20880 66705 21090
rect 67095 20895 67305 21105
rect 68295 20880 68505 21090
rect 67395 20595 67605 20805
rect 65895 20295 66105 20505
rect 64995 19095 65205 19305
rect 63495 18495 63705 18705
rect 63195 18195 63405 18405
rect 64095 18210 64305 18420
rect 61395 16995 61605 17205
rect 62895 16995 63105 17205
rect 63195 14595 63405 14805
rect 64995 16695 65205 16905
rect 65895 17580 66105 17790
rect 66495 17580 66705 17790
rect 66495 16995 66705 17205
rect 64395 16095 64605 16305
rect 65295 16095 65505 16305
rect 64995 15795 65205 16005
rect 64395 15195 64605 15405
rect 63795 14295 64005 14505
rect 64995 14295 65205 14505
rect 62295 13995 62505 14205
rect 60795 13710 61005 13920
rect 61695 13710 61905 13920
rect 57795 13080 58005 13290
rect 58395 13080 58605 13290
rect 59295 13095 59505 13305
rect 62895 13695 63105 13905
rect 64395 13695 64605 13905
rect 60195 13080 60405 13290
rect 60780 13080 60990 13290
rect 61395 13080 61605 13290
rect 60795 12195 61005 12405
rect 56895 11595 57105 11805
rect 60195 11295 60405 11505
rect 57795 10995 58005 11205
rect 57195 10410 57405 10620
rect 46995 8895 47205 9105
rect 50595 8895 50805 9105
rect 51795 8895 52005 9105
rect 52395 8895 52605 9105
rect 46695 8295 46905 8505
rect 50595 8295 50805 8505
rect 50595 7695 50805 7905
rect 55395 7695 55605 7905
rect 47895 6795 48105 7005
rect 49095 6795 49305 7005
rect 45195 6495 45405 6705
rect 46095 6495 46305 6705
rect 45795 6195 46005 6405
rect 47295 6195 47505 6405
rect 48195 6495 48405 6705
rect 48795 6195 49005 6405
rect 48495 5910 48705 6120
rect 41895 5595 42105 5805
rect 44595 5595 44805 5805
rect 39795 5295 40005 5505
rect 40395 5280 40605 5490
rect 40995 5280 41205 5490
rect 42795 5280 43005 5490
rect 41295 4995 41505 5205
rect 41895 4995 42105 5205
rect 40695 4395 40905 4605
rect 40095 3195 40305 3405
rect 39495 2895 39705 3105
rect 42495 4695 42705 4905
rect 42195 4095 42405 4305
rect 39195 1980 39405 2190
rect 40095 1980 40305 2190
rect 40995 1980 41205 2190
rect 37995 1695 38205 1905
rect 38595 1695 38805 1905
rect 41595 1695 41805 1905
rect 36795 1395 37005 1605
rect 45495 5280 45705 5490
rect 46095 4995 46305 5205
rect 46995 4995 47205 5205
rect 48495 5295 48705 5505
rect 48195 4995 48405 5205
rect 47595 4695 47805 4905
rect 48495 4695 48705 4905
rect 49395 6195 49605 6405
rect 52095 7095 52305 7305
rect 55395 7095 55605 7305
rect 51195 5910 51405 6120
rect 53595 6795 53805 7005
rect 52995 6195 53205 6405
rect 54495 6195 54705 6405
rect 55995 9780 56205 9990
rect 57495 9780 57705 9990
rect 59895 9780 60105 9990
rect 58095 9195 58305 9405
rect 58695 9195 58905 9405
rect 56595 6795 56805 7005
rect 57195 6495 57405 6705
rect 59595 6495 59805 6705
rect 55695 6195 55905 6405
rect 56295 5910 56505 6120
rect 57795 5910 58005 6120
rect 58995 5910 59205 6120
rect 50895 5280 51105 5490
rect 52095 5280 52305 5490
rect 49695 4695 49905 4905
rect 50295 4695 50505 4905
rect 51495 4695 51705 4905
rect 45495 4395 45705 4605
rect 48795 4395 49005 4605
rect 43395 4095 43605 4305
rect 43995 2895 44205 3105
rect 48495 4095 48705 4305
rect 49095 4095 49305 4305
rect 48195 3795 48405 4005
rect 48795 3795 49005 4005
rect 43395 2610 43605 2820
rect 44595 2595 44805 2805
rect 45495 2610 45705 2820
rect 46095 2610 46305 2820
rect 46995 2595 47205 2805
rect 52695 4395 52905 4605
rect 51195 3495 51405 3705
rect 50595 3195 50805 3405
rect 50595 2595 50805 2805
rect 42495 1980 42705 2190
rect 43095 1980 43305 2190
rect 43695 1980 43905 2190
rect 44595 1980 44805 2190
rect 47295 2295 47505 2505
rect 45195 1980 45405 2190
rect 45795 1980 46005 2190
rect 46995 1980 47205 2190
rect 54495 5280 54705 5490
rect 55095 5280 55305 5490
rect 55395 4995 55605 5205
rect 60495 5895 60705 6105
rect 54795 4695 55005 4905
rect 56295 4695 56505 4905
rect 53595 4395 53805 4605
rect 53295 4095 53505 4305
rect 52995 3495 53205 3705
rect 47895 1980 48105 2190
rect 48495 1980 48705 2190
rect 50895 1995 51105 2205
rect 44895 1395 45105 1605
rect 47295 1395 47505 1605
rect 47895 1095 48105 1305
rect 36195 795 36405 1005
rect 42195 795 42405 1005
rect 52695 1995 52905 2205
rect 53295 3195 53505 3405
rect 53295 2595 53505 2805
rect 54195 2610 54405 2820
rect 57495 4995 57705 5205
rect 59895 5280 60105 5490
rect 59295 4995 59505 5205
rect 58995 4695 59205 4905
rect 56895 3795 57105 4005
rect 55995 3195 56205 3405
rect 57495 3195 57705 3405
rect 61395 11595 61605 11805
rect 61095 10995 61305 11205
rect 61095 9780 61305 9990
rect 62895 13095 63105 13305
rect 64095 13080 64305 13290
rect 64995 13095 65205 13305
rect 63495 12795 63705 13005
rect 64695 11595 64905 11805
rect 63795 11295 64005 11505
rect 61995 10995 62205 11205
rect 64395 10695 64605 10905
rect 62895 10425 63105 10635
rect 61695 10095 61905 10305
rect 61395 8895 61605 9105
rect 63495 9795 63705 10005
rect 62295 8595 62505 8805
rect 61695 7695 61905 7905
rect 62295 6495 62505 6705
rect 65595 14595 65805 14805
rect 65595 13695 65805 13905
rect 67695 18495 67905 18705
rect 67395 18195 67605 18405
rect 67995 17580 68205 17790
rect 66780 16695 66990 16905
rect 67095 16695 67305 16905
rect 65895 13080 66105 13290
rect 66795 11895 67005 12105
rect 67395 15195 67605 15405
rect 68295 15795 68505 16005
rect 67395 13695 67605 13905
rect 70095 25395 70305 25605
rect 69795 24795 70005 25005
rect 69795 23595 70005 23805
rect 69495 22095 69705 22305
rect 70995 28695 71205 28905
rect 70695 26295 70905 26505
rect 71895 29310 72105 29520
rect 74295 35895 74505 36105
rect 73695 35595 73905 35805
rect 76695 46395 76905 46605
rect 80295 48780 80505 48990
rect 78495 48195 78705 48405
rect 79095 48195 79305 48405
rect 80595 48195 80805 48405
rect 77895 47595 78105 47805
rect 77295 46095 77505 46305
rect 76695 45195 76905 45405
rect 76995 44910 77205 45120
rect 76995 43995 77205 44205
rect 76695 43695 76905 43905
rect 77295 43395 77505 43605
rect 76995 42795 77205 43005
rect 79695 47595 79905 47805
rect 77895 45195 78105 45405
rect 79095 45195 79305 45405
rect 79995 47295 80205 47505
rect 80895 47595 81105 47805
rect 79695 44910 79905 45120
rect 80295 46995 80505 47205
rect 82395 51795 82605 52005
rect 81795 51195 82005 51405
rect 81495 50895 81705 51105
rect 81795 50595 82005 50805
rect 81495 49395 81705 49605
rect 85395 59895 85605 60105
rect 84795 57495 85005 57705
rect 83595 56595 83805 56805
rect 83295 53895 83505 54105
rect 84195 56580 84405 56790
rect 86295 64095 86505 64305
rect 88395 73995 88605 74205
rect 88395 69795 88605 70005
rect 91395 75195 91605 75405
rect 91095 74895 91305 75105
rect 90195 73695 90405 73905
rect 91395 72795 91605 73005
rect 92040 77595 92250 77805
rect 91995 73395 92205 73605
rect 90795 71295 91005 71505
rect 88695 69195 88905 69405
rect 91395 69795 91605 70005
rect 91995 68595 92205 68805
rect 88395 68295 88605 68505
rect 88995 68310 89205 68520
rect 88095 67395 88305 67605
rect 88695 67680 88905 67890
rect 88395 67095 88605 67305
rect 89295 66195 89505 66405
rect 88995 65595 89205 65805
rect 88695 65295 88905 65505
rect 88095 64995 88305 65205
rect 91095 68310 91305 68520
rect 91995 68280 92205 68490
rect 90795 67680 91005 67890
rect 91695 67695 91905 67905
rect 91395 67095 91605 67305
rect 89895 66795 90105 67005
rect 91395 66780 91605 66990
rect 90195 66195 90405 66405
rect 89595 64995 89805 65205
rect 91095 65595 91305 65805
rect 88395 64395 88605 64605
rect 87195 63795 87405 64005
rect 86295 61695 86505 61905
rect 86895 61695 87105 61905
rect 86895 61380 87105 61590
rect 86295 61095 86505 61305
rect 85995 60495 86205 60705
rect 86895 60510 87105 60720
rect 85995 59895 86205 60105
rect 85695 57480 85905 57690
rect 84795 55995 85005 56205
rect 83895 54795 84105 55005
rect 83595 53595 83805 53805
rect 82995 52695 83205 52905
rect 83295 52995 83505 53205
rect 82995 52095 83205 52305
rect 82695 50895 82905 51105
rect 82395 49710 82605 49920
rect 83595 52080 83805 52290
rect 83895 51795 84105 52005
rect 83295 50895 83505 51105
rect 82395 49395 82605 49605
rect 82095 48780 82305 48990
rect 82695 48780 82905 48990
rect 81495 47595 81705 47805
rect 81195 46095 81405 46305
rect 80895 45495 81105 45705
rect 78495 44280 78705 44490
rect 77895 43095 78105 43305
rect 77595 42495 77805 42705
rect 77595 42180 77805 42390
rect 77295 41895 77505 42105
rect 78495 43095 78705 43305
rect 77295 40980 77505 41190
rect 76395 40680 76605 40890
rect 76095 38895 76305 39105
rect 74895 37095 75105 37305
rect 75795 37395 76005 37605
rect 76095 37110 76305 37320
rect 74895 36495 75105 36705
rect 74595 35295 74805 35505
rect 74895 34995 75105 35205
rect 74595 34095 74805 34305
rect 73995 31395 74205 31605
rect 73095 30195 73305 30405
rect 72195 28680 72405 28890
rect 72495 28395 72705 28605
rect 71595 27495 71805 27705
rect 71295 26295 71505 26505
rect 75795 36480 76005 36690
rect 76395 36495 76605 36705
rect 76095 35895 76305 36105
rect 75795 34995 76005 35205
rect 75195 34095 75405 34305
rect 77895 40395 78105 40605
rect 80595 44895 80805 45105
rect 79695 42795 79905 43005
rect 78795 42195 79005 42405
rect 78795 41595 79005 41805
rect 79395 41610 79605 41820
rect 80295 44280 80505 44490
rect 81195 44295 81405 44505
rect 81195 43395 81405 43605
rect 80295 43095 80505 43305
rect 80895 42795 81105 43005
rect 80295 41580 80505 41790
rect 76995 39195 77205 39405
rect 78495 39195 78705 39405
rect 79695 40980 79905 41190
rect 78195 38295 78405 38505
rect 77595 37695 77805 37905
rect 76995 37095 77205 37305
rect 76695 35595 76905 35805
rect 76695 34995 76905 35205
rect 76395 34695 76605 34905
rect 76095 34095 76305 34305
rect 75495 33180 75705 33390
rect 77295 36480 77505 36690
rect 77295 34695 77505 34905
rect 80295 40395 80505 40605
rect 79995 38295 80205 38505
rect 80595 38295 80805 38505
rect 78795 37995 79005 38205
rect 79395 37110 79605 37320
rect 79995 37110 80205 37320
rect 80595 37095 80805 37305
rect 79095 36495 79305 36705
rect 78795 36195 79005 36405
rect 78795 35595 79005 35805
rect 78195 34095 78405 34305
rect 76395 33495 76605 33705
rect 75495 32595 75705 32805
rect 73395 29595 73605 29805
rect 74595 29595 74805 29805
rect 75195 29595 75405 29805
rect 73095 27195 73305 27405
rect 73995 29310 74205 29520
rect 74295 28695 74505 28905
rect 73995 28395 74205 28605
rect 72795 26295 73005 26505
rect 72495 25995 72705 26205
rect 71895 25380 72105 25590
rect 72495 25395 72705 25605
rect 72495 23295 72705 23505
rect 71295 22695 71505 22905
rect 73395 22395 73605 22605
rect 70395 22095 70605 22305
rect 71595 21495 71805 21705
rect 69495 20880 69705 21090
rect 70095 20880 70305 21090
rect 69195 20295 69405 20505
rect 70095 19995 70305 20205
rect 70695 19395 70905 19605
rect 72795 21510 73005 21720
rect 74595 27195 74805 27405
rect 75195 27195 75405 27405
rect 76995 32895 77205 33105
rect 76695 31395 76905 31605
rect 76095 30795 76305 31005
rect 77595 29895 77805 30105
rect 76395 29595 76605 29805
rect 76095 29295 76305 29505
rect 77895 29310 78105 29520
rect 76695 28680 76905 28890
rect 75795 28395 76005 28605
rect 76395 28395 76605 28605
rect 78195 28695 78405 28905
rect 76095 27495 76305 27705
rect 74595 26595 74805 26805
rect 74295 25995 74505 26205
rect 75795 25995 76005 26205
rect 73995 25095 74205 25305
rect 73695 21795 73905 22005
rect 75795 25395 76005 25605
rect 75495 25095 75705 25305
rect 74595 24495 74805 24705
rect 74295 22695 74505 22905
rect 75495 22695 75705 22905
rect 74295 22380 74505 22590
rect 73995 21495 74205 21705
rect 71895 20895 72105 21105
rect 73095 20880 73305 21090
rect 73995 20895 74205 21105
rect 73695 20295 73905 20505
rect 71895 19995 72105 20205
rect 70095 18210 70305 18420
rect 70695 18240 70905 18450
rect 71595 18240 71805 18450
rect 72195 19395 72405 19605
rect 72195 18195 72405 18405
rect 72195 17595 72405 17805
rect 74595 21795 74805 22005
rect 74295 20595 74505 20805
rect 74295 19995 74505 20205
rect 73395 17550 73605 17760
rect 71895 16995 72105 17205
rect 70080 16695 70290 16905
rect 70395 16695 70605 16905
rect 69495 16395 69705 16605
rect 68895 15495 69105 15705
rect 69195 14895 69405 15105
rect 67995 13080 68205 13290
rect 68595 13080 68805 13290
rect 70395 16095 70605 16305
rect 71295 16095 71505 16305
rect 70095 14295 70305 14505
rect 70695 14295 70905 14505
rect 69495 13710 69705 13920
rect 70095 13710 70305 13920
rect 72495 14895 72705 15105
rect 71595 14595 71805 14805
rect 69495 13095 69705 13305
rect 70395 13080 70605 13290
rect 71295 13095 71505 13305
rect 73095 13710 73305 13920
rect 69495 12495 69705 12705
rect 71595 12495 71805 12705
rect 72195 12495 72405 12705
rect 69195 12195 69405 12405
rect 68595 11595 68805 11805
rect 67095 10995 67305 11205
rect 68595 10995 68805 11205
rect 65295 10695 65505 10905
rect 65895 10410 66105 10620
rect 66795 10395 67005 10605
rect 67395 10410 67605 10620
rect 64695 9780 64905 9990
rect 66195 9780 66405 9990
rect 67095 9795 67305 10005
rect 66795 9195 67005 9405
rect 67695 9495 67905 9705
rect 67095 8595 67305 8805
rect 70995 11895 71205 12105
rect 70395 10695 70605 10905
rect 69795 9495 70005 9705
rect 69195 9195 69405 9405
rect 68895 8895 69105 9105
rect 68895 8295 69105 8505
rect 68595 7995 68805 8205
rect 65595 7695 65805 7905
rect 67395 7395 67605 7605
rect 64695 7095 64905 7305
rect 61695 5910 61905 6120
rect 63195 5910 63405 6120
rect 63795 5910 64005 6120
rect 64395 5910 64605 6120
rect 60795 4695 61005 4905
rect 62895 5280 63105 5490
rect 63495 5280 63705 5490
rect 61395 3795 61605 4005
rect 60495 3195 60705 3405
rect 54795 2595 55005 2805
rect 56595 2610 56805 2820
rect 55395 2295 55605 2505
rect 54495 1980 54705 2190
rect 52995 1695 53205 1905
rect 53895 1695 54105 1905
rect 55395 1395 55605 1605
rect 56895 1980 57105 2190
rect 61995 2895 62205 3105
rect 61395 2610 61605 2820
rect 62295 2610 62505 2820
rect 63195 2610 63405 2820
rect 63795 2610 64005 2820
rect 60495 1980 60705 2190
rect 61095 1980 61305 2190
rect 62895 1980 63105 2190
rect 63495 1980 63705 2190
rect 61695 1395 61905 1605
rect 62295 1395 62505 1605
rect 63195 1395 63405 1605
rect 61095 1095 61305 1305
rect 65295 6795 65505 7005
rect 65895 6195 66105 6405
rect 66495 5910 66705 6120
rect 64695 5295 64905 5505
rect 67995 5910 68205 6120
rect 72195 11595 72405 11805
rect 71595 10695 71805 10905
rect 74295 17295 74505 17505
rect 74295 15795 74505 16005
rect 74295 14895 74505 15105
rect 73995 14595 74205 14805
rect 74295 14295 74505 14505
rect 76095 24495 76305 24705
rect 75795 21795 76005 22005
rect 75195 20595 75405 20805
rect 76095 20895 76305 21105
rect 75795 20295 76005 20505
rect 75795 18195 76005 18405
rect 75195 17580 75405 17790
rect 74895 15795 75105 16005
rect 74595 13995 74805 14205
rect 77595 27795 77805 28005
rect 76695 26895 76905 27105
rect 77895 27495 78105 27705
rect 78795 34995 79005 35205
rect 80295 36480 80505 36690
rect 82695 45795 82905 46005
rect 81795 45495 82005 45705
rect 81495 42195 81705 42405
rect 82095 44895 82305 45105
rect 83595 50295 83805 50505
rect 84795 51495 85005 51705
rect 84495 50295 84705 50505
rect 84195 49995 84405 50205
rect 83595 49395 83805 49605
rect 84795 49410 85005 49620
rect 83595 48795 83805 49005
rect 83295 47595 83505 47805
rect 84495 48195 84705 48405
rect 87195 59895 87405 60105
rect 86595 59295 86805 59505
rect 86895 58095 87105 58305
rect 86595 57795 86805 58005
rect 85995 57195 86205 57405
rect 88095 64095 88305 64305
rect 87795 63795 88005 64005
rect 87495 58995 87705 59205
rect 87495 57795 87705 58005
rect 86895 56580 87105 56790
rect 86595 56295 86805 56505
rect 85995 54195 86205 54405
rect 85695 53895 85905 54105
rect 86895 53595 87105 53805
rect 85395 52695 85605 52905
rect 85995 52710 86205 52920
rect 86595 52710 86805 52920
rect 87195 52695 87405 52905
rect 85395 52095 85605 52305
rect 86295 52080 86505 52290
rect 86895 52080 87105 52290
rect 85695 51195 85905 51405
rect 86595 51195 86805 51405
rect 85695 50595 85905 50805
rect 86295 50595 86505 50805
rect 85695 49995 85905 50205
rect 86295 49695 86505 49905
rect 85995 49410 86205 49620
rect 86895 49395 87105 49605
rect 85395 48495 85605 48705
rect 83895 47895 84105 48105
rect 83595 46995 83805 47205
rect 83295 46395 83505 46605
rect 83595 46095 83805 46305
rect 83295 45795 83505 46005
rect 82995 44895 83205 45105
rect 84195 44895 84405 45105
rect 83295 44280 83505 44490
rect 83895 43995 84105 44205
rect 84795 47595 85005 47805
rect 86895 48795 87105 49005
rect 86595 48495 86805 48705
rect 86295 47295 86505 47505
rect 86295 46395 86505 46605
rect 85395 44910 85605 45120
rect 84495 44295 84705 44505
rect 82995 43095 83205 43305
rect 84195 43095 84405 43305
rect 85695 44280 85905 44490
rect 82095 42495 82305 42705
rect 83295 42495 83505 42705
rect 84195 42495 84405 42705
rect 81795 41895 82005 42105
rect 82095 41610 82305 41820
rect 83295 41880 83505 42090
rect 84195 41895 84405 42105
rect 81195 40995 81405 41205
rect 82395 40980 82605 41190
rect 81795 39495 82005 39705
rect 83295 40980 83505 41190
rect 84495 40995 84705 41205
rect 83895 40695 84105 40905
rect 83895 39795 84105 40005
rect 81495 37995 81705 38205
rect 81195 37095 81405 37305
rect 82395 37395 82605 37605
rect 82995 38295 83205 38505
rect 82695 37095 82905 37305
rect 83295 37395 83505 37605
rect 79680 36195 79890 36405
rect 79995 36195 80205 36405
rect 79395 35295 79605 35505
rect 79095 34695 79305 34905
rect 80295 34995 80505 35205
rect 79995 33795 80205 34005
rect 79095 32595 79305 32805
rect 78795 31095 79005 31305
rect 78495 26595 78705 26805
rect 77295 24795 77505 25005
rect 77595 23295 77805 23505
rect 76995 22695 77205 22905
rect 76695 22095 76905 22305
rect 78195 25395 78405 25605
rect 77895 22995 78105 23205
rect 77895 22095 78105 22305
rect 77595 21510 77805 21720
rect 76695 20895 76905 21105
rect 77295 18795 77505 19005
rect 79395 30795 79605 31005
rect 79995 33195 80205 33405
rect 81780 36480 81990 36690
rect 82095 36495 82305 36705
rect 82995 36495 83205 36705
rect 88695 64095 88905 64305
rect 88395 62295 88605 62505
rect 89595 64395 89805 64605
rect 89295 63495 89505 63705
rect 89295 61695 89505 61905
rect 88695 60495 88905 60705
rect 89595 60495 89805 60705
rect 88095 59895 88305 60105
rect 88095 59295 88305 59505
rect 88995 59295 89205 59505
rect 89595 58995 89805 59205
rect 88395 57795 88605 58005
rect 88995 57795 89205 58005
rect 87795 57495 88005 57705
rect 88395 57210 88605 57420
rect 89295 57195 89505 57405
rect 87795 55995 88005 56205
rect 88695 55995 88905 56205
rect 88095 54795 88305 55005
rect 87795 54195 88005 54405
rect 87495 51195 87705 51405
rect 88995 53895 89205 54105
rect 88395 53295 88605 53505
rect 88095 52695 88305 52905
rect 89295 52695 89505 52905
rect 88095 52095 88305 52305
rect 87795 50595 88005 50805
rect 88995 51795 89205 52005
rect 88695 51495 88905 51705
rect 87495 49995 87705 50205
rect 88095 49995 88305 50205
rect 87195 48495 87405 48705
rect 86895 47595 87105 47805
rect 86895 45795 87105 46005
rect 86595 44895 86805 45105
rect 88395 49695 88605 49905
rect 88980 49695 89190 49905
rect 89295 49695 89505 49905
rect 88095 48495 88305 48705
rect 88395 48195 88605 48405
rect 88095 47595 88305 47805
rect 87795 46695 88005 46905
rect 87495 44895 87705 45105
rect 86595 44295 86805 44505
rect 86295 43395 86505 43605
rect 85695 42495 85905 42705
rect 87495 44295 87705 44505
rect 89295 48795 89505 49005
rect 88995 48495 89205 48705
rect 88695 47895 88905 48105
rect 88395 46695 88605 46905
rect 88395 46380 88605 46590
rect 88095 45495 88305 45705
rect 88995 45795 89205 46005
rect 88695 45195 88905 45405
rect 89295 44895 89505 45105
rect 88395 43995 88605 44205
rect 87795 43695 88005 43905
rect 88095 42795 88305 43005
rect 86895 42195 87105 42405
rect 87495 42195 87705 42405
rect 86595 41895 86805 42105
rect 89295 44295 89505 44505
rect 88995 43695 89205 43905
rect 88695 42795 88905 43005
rect 87795 41610 88005 41820
rect 88395 41595 88605 41805
rect 84795 39795 85005 40005
rect 84495 37395 84705 37605
rect 85395 40695 85605 40905
rect 86295 38595 86505 38805
rect 85395 37395 85605 37605
rect 84195 36480 84405 36690
rect 83295 36195 83505 36405
rect 83895 36195 84105 36405
rect 82395 35295 82605 35505
rect 82095 34995 82305 35205
rect 85095 36495 85305 36705
rect 84795 35895 85005 36105
rect 83895 34995 84105 35205
rect 84795 34995 85005 35205
rect 81495 33810 81705 34020
rect 83595 34695 83805 34905
rect 83595 34095 83805 34305
rect 82695 33810 82905 34020
rect 83295 33810 83505 34020
rect 83895 33810 84105 34020
rect 81795 33180 82005 33390
rect 80595 32595 80805 32805
rect 80595 31395 80805 31605
rect 80295 31095 80505 31305
rect 79080 29295 79290 29505
rect 79395 29310 79605 29520
rect 79995 29310 80205 29520
rect 83595 33180 83805 33390
rect 83895 32895 84105 33105
rect 82695 32595 82905 32805
rect 81495 32295 81705 32505
rect 81195 31695 81405 31905
rect 80895 30795 81105 31005
rect 80895 29895 81105 30105
rect 80295 28680 80505 28890
rect 79095 28395 79305 28605
rect 80595 27495 80805 27705
rect 79695 26895 79905 27105
rect 83595 31395 83805 31605
rect 83595 30795 83805 31005
rect 81795 30195 82005 30405
rect 81495 29295 81705 29505
rect 82995 29595 83205 29805
rect 82395 29310 82605 29520
rect 83295 29295 83505 29505
rect 81180 28695 81390 28905
rect 83895 29595 84105 29805
rect 84795 32295 85005 32505
rect 85995 37395 86205 37605
rect 87195 40995 87405 41205
rect 86595 37995 86805 38205
rect 88095 40980 88305 41190
rect 87195 39495 87405 39705
rect 88695 39195 88905 39405
rect 88095 38895 88305 39105
rect 87495 38295 87705 38505
rect 85695 37095 85905 37305
rect 86895 37395 87105 37605
rect 85395 36195 85605 36405
rect 85995 36195 86205 36405
rect 85695 35895 85905 36105
rect 86895 36480 87105 36690
rect 87795 37395 88005 37605
rect 86595 33795 86805 34005
rect 87495 36480 87705 36690
rect 87495 35895 87705 36105
rect 88695 38595 88905 38805
rect 89295 42795 89505 43005
rect 89295 41895 89505 42105
rect 90495 63495 90705 63705
rect 90495 61695 90705 61905
rect 90195 60495 90405 60705
rect 91695 66195 91905 66405
rect 91395 61095 91605 61305
rect 91095 60495 91305 60705
rect 91995 60795 92205 61005
rect 90795 59880 91005 60090
rect 90495 59595 90705 59805
rect 90195 58095 90405 58305
rect 90795 58695 91005 58905
rect 91395 58695 91605 58905
rect 89895 57195 90105 57405
rect 90495 57495 90705 57705
rect 91095 58095 91305 58305
rect 90795 57195 91005 57405
rect 90195 55095 90405 55305
rect 90795 56595 91005 56805
rect 90495 54495 90705 54705
rect 91395 57495 91605 57705
rect 91995 59295 92205 59505
rect 91995 58695 92205 58905
rect 91695 55095 91905 55305
rect 91395 54795 91605 55005
rect 91695 54495 91905 54705
rect 91395 53895 91605 54105
rect 91095 53295 91305 53505
rect 90495 52995 90705 53205
rect 89895 52695 90105 52905
rect 91695 52695 91905 52905
rect 90195 50595 90405 50805
rect 91095 52080 91305 52290
rect 90795 49995 91005 50205
rect 91695 49995 91905 50205
rect 90495 49695 90705 49905
rect 90195 49395 90405 49605
rect 90195 48795 90405 49005
rect 89895 48195 90105 48405
rect 89895 47295 90105 47505
rect 90495 48495 90705 48705
rect 91395 48495 91605 48705
rect 91095 47295 91305 47505
rect 90495 45795 90705 46005
rect 90795 45495 91005 45705
rect 90195 44895 90405 45105
rect 91695 47895 91905 48105
rect 91695 47295 91905 47505
rect 91395 45195 91605 45405
rect 91995 45795 92205 46005
rect 91995 45195 92205 45405
rect 90195 44295 90405 44505
rect 89895 43995 90105 44205
rect 91095 44280 91305 44490
rect 91995 44280 92205 44490
rect 91395 43995 91605 44205
rect 90495 43395 90705 43605
rect 90195 42195 90405 42405
rect 90795 42195 91005 42405
rect 89895 41895 90105 42105
rect 88995 37395 89205 37605
rect 90195 40980 90405 41190
rect 90195 39795 90405 40005
rect 90195 39195 90405 39405
rect 89895 38595 90105 38805
rect 91095 39795 91305 40005
rect 90795 38595 91005 38805
rect 90795 37995 91005 38205
rect 89895 37095 90105 37305
rect 91095 37095 91305 37305
rect 88095 36495 88305 36705
rect 87795 34695 88005 34905
rect 88995 36480 89205 36690
rect 89595 36495 89805 36705
rect 89895 36495 90105 36705
rect 88395 35895 88605 36105
rect 89595 35295 89805 35505
rect 88695 34695 88905 34905
rect 89295 34695 89505 34905
rect 85995 32595 86205 32805
rect 86595 31695 86805 31905
rect 85095 30795 85305 31005
rect 86595 30195 86805 30405
rect 84495 29895 84705 30105
rect 85095 29895 85305 30105
rect 84795 29310 85005 29520
rect 85995 29310 86205 29520
rect 83895 28995 84105 29205
rect 81495 28680 81705 28890
rect 82095 28680 82305 28890
rect 82695 28680 82905 28890
rect 83595 28680 83805 28890
rect 78795 25995 79005 26205
rect 79695 26295 79905 26505
rect 80895 26280 81105 26490
rect 81795 28395 82005 28605
rect 84195 28695 84405 28905
rect 82095 28095 82305 28305
rect 83880 28095 84090 28305
rect 81795 27795 82005 28005
rect 81495 25995 81705 26205
rect 78495 23895 78705 24105
rect 79395 24795 79605 25005
rect 79095 24195 79305 24405
rect 79095 22995 79305 23205
rect 79695 22995 79905 23205
rect 78480 21495 78690 21705
rect 78795 21495 79005 21705
rect 76995 17595 77205 17805
rect 76695 16095 76905 16305
rect 76395 14895 76605 15105
rect 75780 13980 75990 14190
rect 76095 13995 76305 14205
rect 74895 13710 75105 13920
rect 75495 13695 75705 13905
rect 74595 13080 74805 13290
rect 75495 13080 75705 13290
rect 75495 12495 75705 12705
rect 74595 10695 74805 10905
rect 72780 10395 72990 10605
rect 73095 10410 73305 10620
rect 73995 10410 74205 10620
rect 72495 9780 72705 9990
rect 72195 9495 72405 9705
rect 70995 8595 71205 8805
rect 70695 6195 70905 6405
rect 71595 5940 71805 6150
rect 66195 4995 66405 5205
rect 65595 4695 65805 4905
rect 65295 3795 65505 4005
rect 64695 2595 64905 2805
rect 65895 2610 66105 2820
rect 66495 2610 66705 2820
rect 65595 1980 65805 2190
rect 64695 1695 64905 1905
rect 66195 1695 66405 1905
rect 68295 5280 68505 5490
rect 68895 5250 69105 5460
rect 75495 10395 75705 10605
rect 73095 9495 73305 9705
rect 72795 5940 73005 6150
rect 72195 4995 72405 5205
rect 70095 4695 70305 4905
rect 72495 3195 72705 3405
rect 68295 2610 68505 2820
rect 69495 2610 69705 2820
rect 67395 1980 67605 2190
rect 73695 3795 73905 4005
rect 74595 9195 74805 9405
rect 74895 8595 75105 8805
rect 75195 8295 75405 8505
rect 74595 7095 74805 7305
rect 77295 16095 77505 16305
rect 77295 14595 77505 14805
rect 76680 13995 76890 14205
rect 76995 13995 77205 14205
rect 76095 13680 76305 13890
rect 79395 20295 79605 20505
rect 79680 18210 79890 18420
rect 80595 25395 80805 25605
rect 80295 25095 80505 25305
rect 80595 22395 80805 22605
rect 80295 21495 80505 21705
rect 81495 22995 81705 23205
rect 81195 22395 81405 22605
rect 84195 28080 84405 28290
rect 85095 28680 85305 28890
rect 85695 28095 85905 28305
rect 87195 33195 87405 33405
rect 86895 29595 87105 29805
rect 87795 31395 88005 31605
rect 87795 29595 88005 29805
rect 88095 29295 88305 29505
rect 86295 28695 86505 28905
rect 86895 28395 87105 28605
rect 85995 27795 86205 28005
rect 84495 27495 84705 27705
rect 85395 27495 85605 27705
rect 84495 26895 84705 27105
rect 82395 26595 82605 26805
rect 84195 26595 84405 26805
rect 82695 26010 82905 26220
rect 83295 26010 83505 26220
rect 83895 26010 84105 26220
rect 84795 25710 85005 25920
rect 82095 25095 82305 25305
rect 82095 24195 82305 24405
rect 81795 22095 82005 22305
rect 83595 25095 83805 25305
rect 85065 25095 85275 25305
rect 82995 24495 83205 24705
rect 80895 21795 81105 22005
rect 82395 21795 82605 22005
rect 81195 21510 81405 21720
rect 88095 28395 88305 28605
rect 87795 28095 88005 28305
rect 88695 33795 88905 34005
rect 90195 35895 90405 36105
rect 91095 36495 91305 36705
rect 90795 35895 91005 36105
rect 90495 35595 90705 35805
rect 90195 34695 90405 34905
rect 89895 34095 90105 34305
rect 90195 33795 90405 34005
rect 88695 33195 88905 33405
rect 88995 30795 89205 31005
rect 89295 30195 89505 30405
rect 88695 29295 88905 29505
rect 90195 33195 90405 33405
rect 90795 34695 91005 34905
rect 90795 34095 91005 34305
rect 90495 30195 90705 30405
rect 88995 28680 89205 28890
rect 89595 28095 89805 28305
rect 88695 27495 88905 27705
rect 89295 27495 89505 27705
rect 87195 27195 87405 27405
rect 87795 27195 88005 27405
rect 88395 27195 88605 27405
rect 89595 27195 89805 27405
rect 85695 26295 85905 26505
rect 89595 25995 89805 26205
rect 87795 25680 88005 25890
rect 89295 25695 89505 25905
rect 89895 25695 90105 25905
rect 91695 43695 91905 43905
rect 91395 35895 91605 36105
rect 91395 35295 91605 35505
rect 91095 28680 91305 28890
rect 85695 25095 85905 25305
rect 89595 24795 89805 25005
rect 85395 24495 85605 24705
rect 85695 23595 85905 23805
rect 85695 22695 85905 22905
rect 83895 21795 84105 22005
rect 89295 22695 89505 22905
rect 88995 22095 89205 22305
rect 82095 21180 82305 21390
rect 82995 21180 83205 21390
rect 83595 21180 83805 21390
rect 79995 18195 80205 18405
rect 78795 17295 79005 17505
rect 79605 17295 79815 17505
rect 79095 16995 79305 17205
rect 78195 15495 78405 15705
rect 77895 14295 78105 14505
rect 77595 13080 77805 13290
rect 80895 20880 81105 21090
rect 81195 18795 81405 19005
rect 82395 20895 82605 21105
rect 82095 20295 82305 20505
rect 82095 19095 82305 19305
rect 80595 18195 80805 18405
rect 81795 18195 82005 18405
rect 80595 17595 80805 17805
rect 81495 17580 81705 17790
rect 82095 17595 82305 17805
rect 79395 16695 79605 16905
rect 80295 16695 80505 16905
rect 82995 20595 83205 20805
rect 83295 20295 83505 20505
rect 82995 19395 83205 19605
rect 85995 21210 86205 21420
rect 87795 21180 88005 21390
rect 83895 20595 84105 20805
rect 83595 19695 83805 19905
rect 85095 19695 85305 19905
rect 85695 19695 85905 19905
rect 83295 19095 83505 19305
rect 82695 18210 82905 18420
rect 83295 18210 83505 18420
rect 85395 19395 85605 19605
rect 85395 18195 85605 18405
rect 89295 19995 89505 20205
rect 90495 25095 90705 25305
rect 91095 22695 91305 22905
rect 90795 22095 91005 22305
rect 90195 21510 90405 21720
rect 90495 20880 90705 21090
rect 89595 19695 89805 19905
rect 87795 19395 88005 19605
rect 90195 19995 90405 20205
rect 84195 17910 84405 18120
rect 85095 17910 85305 18120
rect 85695 17910 85905 18120
rect 82995 17580 83205 17790
rect 82695 17295 82905 17505
rect 89895 18195 90105 18405
rect 90795 18195 91005 18405
rect 91995 42795 92205 43005
rect 91995 38895 92205 39105
rect 91995 37995 92205 38205
rect 91995 35295 92205 35505
rect 91695 34695 91905 34905
rect 91395 19095 91605 19305
rect 88095 17880 88305 18090
rect 89595 17895 89805 18105
rect 90195 17895 90405 18105
rect 82695 16695 82905 16905
rect 81795 15495 82005 15705
rect 82395 15495 82605 15705
rect 80895 14895 81105 15105
rect 81495 14895 81705 15105
rect 82395 14895 82605 15105
rect 79395 14295 79605 14505
rect 79995 14295 80205 14505
rect 79395 13710 79605 13920
rect 80295 13995 80505 14205
rect 79995 13695 80205 13905
rect 82095 13395 82305 13605
rect 78195 13080 78405 13290
rect 79095 13080 79305 13290
rect 76395 11895 76605 12105
rect 78495 11895 78705 12105
rect 76095 10995 76305 11205
rect 76995 10995 77205 11205
rect 76395 10695 76605 10905
rect 79095 11595 79305 11805
rect 79095 10995 79305 11205
rect 80295 13095 80505 13305
rect 81195 13080 81405 13290
rect 81795 12795 82005 13005
rect 79095 10410 79305 10620
rect 79695 10410 79905 10620
rect 80895 10410 81105 10620
rect 81495 10410 81705 10620
rect 82095 10410 82305 10620
rect 76695 9780 76905 9990
rect 75795 9495 76005 9705
rect 75795 6495 76005 6705
rect 75495 6195 75705 6405
rect 76395 5910 76605 6120
rect 78795 9780 79005 9990
rect 78195 9195 78405 9405
rect 80595 9495 80805 9705
rect 78795 8895 79005 9105
rect 81795 8595 82005 8805
rect 83895 16395 84105 16605
rect 83295 13995 83505 14205
rect 85995 17295 86205 17505
rect 91395 17295 91605 17505
rect 85695 16995 85905 17205
rect 90135 16995 90345 17205
rect 90795 16695 91005 16905
rect 87795 16095 88005 16305
rect 88995 16095 89205 16305
rect 85695 14895 85905 15105
rect 87195 14895 87405 15105
rect 87795 14895 88005 15105
rect 85695 14295 85905 14505
rect 82695 11895 82905 12105
rect 84195 12795 84405 13005
rect 83280 10995 83490 11205
rect 83595 10995 83805 11205
rect 84495 11295 84705 11505
rect 84195 10995 84405 11205
rect 85395 13695 85605 13905
rect 85995 12795 86205 13005
rect 85695 11295 85905 11505
rect 84195 10395 84405 10605
rect 82995 9780 83205 9990
rect 83595 8895 83805 9105
rect 82395 8295 82605 8505
rect 77295 7395 77505 7605
rect 80595 7395 80805 7605
rect 81195 7395 81405 7605
rect 84795 10695 85005 10905
rect 86295 10695 86505 10905
rect 85095 9795 85305 10005
rect 84795 8895 85005 9105
rect 85695 8295 85905 8505
rect 85395 7995 85605 8205
rect 77295 6495 77505 6705
rect 75495 5280 75705 5490
rect 76095 4995 76305 5205
rect 76995 4995 77205 5205
rect 77895 5910 78105 6120
rect 83895 7095 84105 7305
rect 83295 6795 83505 7005
rect 81495 6195 81705 6405
rect 82395 6195 82605 6405
rect 84195 6195 84405 6405
rect 85395 5895 85605 6105
rect 83895 5595 84105 5805
rect 75195 3795 75405 4005
rect 77295 3795 77505 4005
rect 77895 3795 78105 4005
rect 74295 3195 74505 3405
rect 73695 2640 73905 2850
rect 75195 2610 75405 2820
rect 78795 5250 79005 5460
rect 78195 3195 78405 3405
rect 80595 3195 80805 3405
rect 79395 2640 79605 2850
rect 85095 5250 85305 5460
rect 80595 2610 80805 2820
rect 82695 2610 82905 2820
rect 83895 2610 84105 2820
rect 86595 9495 86805 9705
rect 86595 7995 86805 8205
rect 85995 6795 86205 7005
rect 86595 7395 86805 7605
rect 86895 7095 87105 7305
rect 87795 14295 88005 14505
rect 88695 11895 88905 12105
rect 88095 8595 88305 8805
rect 90495 15495 90705 15705
rect 89895 14895 90105 15105
rect 89895 13710 90105 13920
rect 89595 10410 89805 10620
rect 89895 9495 90105 9705
rect 88995 7995 89205 8205
rect 90195 7395 90405 7605
rect 88995 6495 89205 6705
rect 87195 6195 87405 6405
rect 88095 6195 88305 6405
rect 86595 5280 86805 5490
rect 85695 4395 85905 4605
rect 86595 4395 86805 4605
rect 87195 4395 87405 4605
rect 89595 5910 89805 6120
rect 88095 5280 88305 5490
rect 88695 5280 88905 5490
rect 89295 4695 89505 4905
rect 90495 5280 90705 5490
rect 90195 4695 90405 4905
rect 91095 6495 91305 6705
rect 89595 4095 89805 4305
rect 90795 4095 91005 4305
rect 66495 1395 66705 1605
rect 60195 795 60405 1005
rect 64395 795 64605 1005
rect 67995 795 68205 1005
rect 11295 495 11505 705
rect 19995 495 20205 705
rect 31995 495 32205 705
rect 41595 495 41805 705
rect 42795 495 43005 705
rect 50895 495 51105 705
rect 51795 495 52005 705
rect 56295 495 56505 705
rect 70995 1950 71205 2160
rect 71895 1950 72105 2160
rect 72480 1950 72690 2160
rect 72795 1950 73005 2160
rect 76695 1950 76905 2160
rect 77595 1950 77805 2160
rect 78195 1950 78405 2160
rect 87795 1980 88005 2190
rect 88995 1980 89205 2190
rect 91995 16695 92205 16905
rect 91995 16095 92205 16305
rect 91695 7395 91905 7605
rect 91395 5910 91605 6120
rect 91995 4395 92205 4605
<< metal3 >>
rect 50205 93840 58095 93960
rect 73005 93840 77895 93960
rect 88005 93840 91095 93960
rect 53205 93540 57795 93660
rect 58005 93540 65595 93660
rect 66705 93540 74460 93660
rect 4605 93240 9795 93360
rect 10005 93240 13695 93360
rect 65505 93240 73995 93360
rect 74340 93360 74460 93540
rect 76305 93540 76695 93660
rect 77040 93540 84795 93660
rect 77040 93360 77160 93540
rect 74340 93240 77160 93360
rect 88605 93240 89995 93360
rect 11505 92940 21495 93060
rect 21705 92940 29895 93060
rect 30105 92940 31095 93060
rect 33705 92940 35760 93060
rect 35640 92805 35760 92940
rect 48105 92940 48795 93060
rect 49005 92940 52995 93060
rect 65805 92940 74295 93060
rect 74505 92940 79995 93060
rect 7905 92640 10995 92760
rect 30705 92640 33795 92760
rect 35805 92640 37095 92760
rect 46605 92640 50595 92760
rect 84405 92640 87495 92760
rect 1605 92340 3795 92460
rect 4005 92340 5895 92460
rect 13305 92340 16395 92460
rect 18105 92340 20595 92460
rect 25005 92340 26595 92460
rect 26805 92340 28095 92460
rect 41805 92340 42795 92460
rect 55905 92340 57195 92460
rect 58605 92340 60195 92460
rect 64605 92340 65895 92460
rect 66105 92340 71895 92460
rect 72105 92340 74595 92460
rect 79305 92340 83895 92460
rect 84705 92340 87360 92460
rect 87240 92205 87360 92340
rect 9105 92040 11295 92160
rect 12105 92040 12795 92160
rect 49605 92040 49995 92160
rect 75405 92040 78195 92160
rect 81705 92040 82095 92160
rect 82905 92040 83295 92160
rect 87405 92040 88995 92160
rect 2805 91755 3195 91875
rect 3840 91740 4380 91860
rect 3840 91560 3960 91740
rect 4905 91755 5295 91875
rect 7905 91740 9660 91860
rect 3540 91440 3960 91560
rect 9540 91560 9660 91740
rect 14505 91755 15195 91875
rect 17205 91740 18495 91860
rect 21240 91740 22095 91860
rect 9540 91440 10260 91560
rect 3540 91290 3660 91440
rect 4305 91140 4695 91260
rect 6405 91125 7095 91245
rect 10140 91290 10260 91440
rect 9105 91140 9495 91260
rect 10440 91260 10560 91710
rect 12540 91440 13095 91560
rect 10440 91140 11595 91260
rect 12540 91260 12660 91440
rect 12405 91140 12660 91260
rect 14205 91140 16695 91260
rect 20040 91260 20160 91710
rect 18540 91140 20160 91260
rect 18540 90960 18660 91140
rect 13005 90840 18660 90960
rect 19005 90840 19995 90960
rect 21240 90960 21360 91740
rect 22905 91755 23595 91875
rect 26205 91755 27195 91875
rect 28905 91755 29295 91875
rect 31905 91755 32595 91875
rect 37005 91755 38595 91875
rect 41205 91755 41595 91875
rect 44505 91740 45495 91860
rect 21705 91125 22395 91245
rect 25305 91125 25695 91245
rect 25905 91140 26895 91260
rect 28905 91125 31395 91245
rect 32805 91140 33795 91260
rect 34140 91260 34260 91695
rect 34140 91140 35295 91260
rect 35505 91140 37695 91260
rect 42240 91260 42360 91710
rect 52005 91755 52395 91875
rect 53805 91755 54195 91875
rect 55005 91740 56595 91860
rect 56805 91755 58380 91875
rect 58905 91755 59295 91875
rect 60105 91755 60495 91875
rect 61605 91740 61980 91860
rect 62505 91755 62895 91875
rect 63705 91740 65295 91860
rect 55140 91440 59460 91560
rect 40905 91140 42360 91260
rect 45705 91125 46095 91245
rect 48405 91140 49395 91260
rect 55140 91290 55260 91440
rect 58605 91140 58995 91260
rect 59340 91260 59460 91440
rect 59340 91140 63795 91260
rect 20205 90840 21360 90960
rect 29805 90840 30495 90960
rect 59805 90840 60195 90960
rect 62205 90840 63495 90960
rect 65040 90960 65160 91740
rect 67605 91740 68295 91860
rect 72705 91755 73395 91875
rect 75540 91740 76995 91860
rect 75540 91290 75660 91740
rect 83040 91740 83895 91860
rect 80940 91305 81060 91710
rect 82440 91305 82560 91710
rect 83040 91560 83160 91740
rect 67005 91125 67695 91245
rect 68505 91125 72195 91245
rect 76905 91140 77595 91260
rect 78405 91140 79395 91260
rect 80805 91140 81060 91305
rect 80805 91095 81000 91140
rect 82305 91140 82560 91305
rect 82740 91440 83160 91560
rect 86040 91560 86160 91710
rect 86040 91440 86895 91560
rect 82740 91290 82860 91440
rect 82305 91095 82500 91140
rect 83805 91140 85695 91260
rect 64605 90840 65160 90960
rect 76605 90840 77895 90960
rect 86505 90840 89295 90960
rect 8205 90540 9495 90660
rect 11805 90540 22395 90660
rect 22605 90540 27495 90660
rect 27705 90540 40695 90660
rect 40905 90540 41295 90660
rect 45105 90540 50895 90660
rect 51105 90540 51795 90660
rect 54705 90540 55695 90660
rect 63405 90540 64095 90660
rect 66105 90540 67380 90660
rect 67905 90540 68595 90660
rect 68805 90540 70095 90660
rect 74205 90540 76695 90660
rect 78405 90540 81195 90660
rect 85005 90540 85995 90660
rect 12105 90240 14595 90360
rect 14805 90240 20895 90360
rect 26205 90240 29295 90360
rect 56805 90240 62295 90360
rect 62505 90240 64995 90360
rect 65205 90240 77295 90360
rect 77505 90240 82095 90360
rect 9105 89940 12795 90060
rect 20505 89940 23595 90060
rect 31005 89940 53295 90060
rect 57105 89940 62895 90060
rect 63705 89940 64980 90060
rect 65505 89940 66495 90060
rect 72105 89940 72795 90060
rect 73605 89940 78195 90060
rect 80805 89940 81195 90060
rect 86505 89940 86895 90060
rect 87105 89940 89595 90060
rect 10005 89640 11895 89760
rect 15405 89640 17895 89760
rect 18105 89640 21195 89760
rect 52605 89640 53595 89760
rect 53805 89640 56295 89760
rect 56505 89640 67095 89760
rect 69705 89640 70995 89760
rect 71205 89640 74895 89760
rect 86205 89640 86895 89760
rect 87105 89640 88995 89760
rect 5805 89340 9495 89460
rect 26805 89340 28095 89460
rect 32205 89340 36495 89460
rect 63105 89340 66795 89460
rect 70905 89340 71595 89460
rect 72240 89340 76695 89460
rect 15105 89040 16095 89160
rect 21105 89040 24495 89160
rect 28605 89040 31695 89160
rect 38505 89040 39495 89160
rect 39705 89040 42495 89160
rect 49305 89040 50295 89160
rect 59805 89040 60495 89160
rect 60705 89040 61995 89160
rect 62205 89040 66660 89160
rect 1905 88740 5895 88860
rect 66540 88905 66660 89040
rect 67605 89040 67995 89160
rect 72240 89160 72360 89340
rect 83205 89340 84795 89460
rect 88005 89340 91695 89460
rect 69405 89040 72360 89160
rect 72705 89040 73695 89160
rect 73905 89040 78795 89160
rect 82605 89040 85395 89160
rect 89205 89040 90495 89160
rect 6105 88740 8295 88860
rect 17040 88740 18495 88860
rect 17040 88620 17160 88740
rect 44805 88740 47295 88860
rect 47505 88740 50460 88860
rect 2340 87960 2460 88410
rect 3405 88440 4095 88560
rect 5205 88455 5895 88575
rect 6705 88440 7395 88560
rect 11205 88440 12195 88560
rect 12405 88440 13395 88560
rect 16005 88455 16995 88575
rect 19605 88455 20895 88575
rect 23505 88455 24195 88575
rect 28305 88455 29895 88575
rect 34005 88440 35295 88560
rect 35505 88440 36795 88560
rect 14040 88260 14160 88410
rect 25140 88260 25260 88410
rect 27240 88260 27360 88410
rect 37005 88440 37860 88560
rect 14040 88140 15060 88260
rect 25140 88140 27360 88260
rect 2340 87840 4395 87960
rect 6405 87840 7995 87960
rect 8205 87840 8460 87960
rect 5205 87540 5895 87660
rect 8340 87660 8460 87840
rect 8805 87825 9195 87945
rect 14940 87960 15060 88140
rect 27240 88005 27360 88140
rect 14940 87840 18195 87960
rect 18405 87840 19695 87960
rect 21405 87840 22095 87960
rect 24105 87840 25395 87960
rect 27105 87840 27360 88005
rect 27105 87795 27300 87840
rect 27705 87840 29595 87960
rect 30405 87840 31695 87960
rect 35805 87840 37095 87960
rect 37740 87960 37860 88440
rect 38205 88455 38595 88575
rect 40305 88440 40695 88560
rect 45705 88440 47460 88560
rect 37740 87840 39195 87960
rect 40005 87840 41595 87960
rect 44895 87945 45105 88095
rect 43305 87825 46995 87945
rect 47340 87960 47460 88440
rect 48105 88440 49860 88560
rect 49740 87990 49860 88440
rect 50340 88560 50460 88740
rect 52905 88740 53460 88860
rect 50340 88440 50595 88560
rect 53340 88560 53460 88740
rect 54405 88740 55095 88860
rect 64005 88740 64395 88860
rect 65805 88740 66360 88860
rect 53340 88440 55395 88560
rect 47340 87840 47595 87960
rect 8340 87540 10695 87660
rect 13905 87540 15495 87660
rect 20805 87540 30795 87660
rect 50040 87675 50160 88410
rect 51840 87960 51960 88410
rect 62205 88440 63060 88560
rect 52740 88140 55095 88260
rect 52740 87990 52860 88140
rect 61440 88260 61560 88410
rect 61440 88200 62745 88260
rect 61440 88140 62805 88200
rect 62595 88005 62805 88140
rect 50505 87840 51960 87960
rect 53505 87840 54495 87960
rect 55605 87825 56895 87945
rect 58905 87840 61095 87960
rect 62790 87900 62805 88005
rect 62940 87990 63060 88440
rect 66240 88560 66360 88740
rect 66705 88740 74295 88860
rect 66240 88440 69195 88560
rect 63240 87960 63360 88410
rect 70305 88560 70500 88605
rect 71100 88560 71295 88605
rect 70305 88395 70560 88560
rect 63240 87840 64095 87960
rect 70440 87990 70560 88395
rect 71040 88395 71295 88560
rect 72105 88440 72960 88560
rect 71040 87990 71160 88395
rect 72840 87990 72960 88440
rect 73305 88440 73995 88560
rect 75540 88005 75660 88410
rect 76905 88560 77100 88605
rect 76905 88395 77160 88560
rect 77505 88440 78060 88560
rect 65205 87825 65595 87945
rect 67305 87825 67695 87945
rect 69105 87825 69495 87945
rect 71805 87825 72195 87945
rect 75405 87840 75660 88005
rect 77040 87990 77160 88395
rect 75405 87795 75600 87840
rect 77940 87960 78060 88440
rect 78405 88440 79260 88560
rect 79140 87990 79260 88440
rect 79905 88455 80595 88575
rect 82305 88455 82995 88575
rect 85740 88440 87495 88560
rect 77940 87840 78495 87960
rect 81105 87840 83295 87960
rect 83640 87960 83760 88410
rect 85740 87990 85860 88440
rect 89340 88260 89460 88410
rect 88140 88200 89460 88260
rect 88095 88140 89460 88200
rect 88095 88005 88305 88140
rect 83640 87840 85095 87960
rect 89805 87840 90495 87960
rect 90705 87840 91395 87960
rect 50040 87495 50295 87675
rect 59505 87540 60195 87660
rect 76605 87540 77595 87660
rect 88605 87540 89295 87660
rect 1605 87240 2895 87360
rect 3105 87240 5595 87360
rect 7305 87240 8295 87360
rect 8505 87240 9195 87360
rect 19005 87240 20295 87360
rect 23505 87240 28095 87360
rect 28305 87240 34095 87360
rect 37905 87240 43695 87360
rect 48105 87240 50895 87360
rect 51105 87240 53295 87360
rect 61305 87240 66195 87360
rect 66405 87240 72195 87360
rect 78105 87240 79395 87360
rect 82305 87240 87795 87360
rect 10905 86940 11595 87060
rect 41205 86940 42795 87060
rect 48705 86940 51195 87060
rect 57105 86940 61695 87060
rect 61905 86940 64095 87060
rect 65805 86940 73860 87060
rect 2805 86640 3795 86760
rect 10740 86760 10860 86895
rect 4005 86640 10860 86760
rect 19305 86640 22995 86760
rect 23205 86640 28695 86760
rect 49305 86640 52095 86760
rect 54105 86640 54795 86760
rect 55005 86640 57795 86760
rect 58005 86640 60795 86760
rect 73740 86760 73860 86940
rect 85305 86940 87195 87060
rect 73740 86640 76695 86760
rect 77505 86640 81795 86760
rect 46005 86340 46395 86460
rect 46605 86340 48495 86460
rect 54105 86340 56895 86460
rect 59205 86340 60495 86460
rect 76605 86340 77895 86460
rect 82905 86340 85695 86460
rect 26205 86040 26895 86160
rect 27105 86040 33495 86160
rect 50205 86040 58395 86160
rect 72405 86040 74295 86160
rect 74505 86040 77295 86160
rect 79605 86040 83460 86160
rect 2505 85740 7095 85860
rect 7305 85740 9195 85860
rect 26505 85740 28695 85860
rect 36405 85740 42495 85860
rect 50805 85740 55395 85860
rect 58005 85740 63495 85860
rect 63705 85740 70995 85860
rect 78705 85740 82095 85860
rect 83340 85860 83460 86040
rect 83340 85740 91860 85860
rect 91740 85605 91860 85740
rect 4605 85440 12195 85560
rect 29205 85440 42795 85560
rect 43005 85440 43695 85560
rect 45405 85440 59295 85560
rect 60105 85440 68895 85560
rect 73005 85440 76995 85560
rect 79005 85440 79695 85560
rect 82005 85440 82995 85560
rect 83205 85440 86295 85560
rect 86505 85440 87795 85560
rect 91740 85440 91995 85605
rect 91800 85395 91995 85440
rect 16605 85140 17295 85260
rect 26805 85140 29895 85260
rect 48705 85140 58995 85260
rect 66405 85140 68295 85260
rect 72405 85140 73995 85260
rect 76305 85140 77895 85260
rect 84405 85140 85695 85260
rect 85905 85140 88995 85260
rect 3405 84840 4095 84960
rect 13005 84840 18795 84960
rect 36705 84840 40395 84960
rect 50505 84840 51495 84960
rect 52905 84840 55095 84960
rect 76140 84960 76260 85095
rect 60405 84840 76260 84960
rect 77505 84840 79095 84960
rect 8805 84540 9495 84660
rect 12105 84540 15495 84660
rect 37440 84540 38895 84660
rect 37440 84405 37560 84540
rect 39540 84540 41295 84660
rect 1605 84240 3060 84360
rect 1305 83940 2595 84060
rect 2940 83460 3060 84240
rect 17205 84240 18495 84360
rect 24405 84240 26895 84360
rect 27840 84240 29295 84360
rect 3705 83955 4395 84075
rect 5040 83760 5160 83910
rect 6105 84060 6300 84105
rect 6105 83895 6360 84060
rect 6705 83955 7995 84075
rect 8205 83940 10095 84060
rect 12405 83940 13695 84060
rect 17505 83955 17895 84075
rect 22305 83940 23595 84060
rect 23805 83940 24795 84060
rect 5040 83640 5760 83760
rect 5640 83505 5760 83640
rect 2940 83340 3195 83460
rect 4605 83340 5295 83460
rect 5640 83340 5895 83505
rect 5700 83295 5895 83340
rect 6240 83460 6360 83895
rect 11940 83640 12795 83760
rect 6240 83340 9195 83460
rect 11940 83490 12060 83640
rect 10905 83340 11295 83460
rect 16305 83340 16995 83460
rect 18840 83460 18960 83895
rect 18405 83340 18960 83460
rect 19740 83460 19860 83910
rect 27840 84060 27960 84240
rect 31995 84240 33495 84360
rect 31995 84120 32205 84240
rect 33705 84240 34260 84360
rect 27705 83940 27960 84060
rect 28305 83955 28995 84075
rect 31005 83940 31995 84060
rect 32805 83955 33195 84075
rect 34140 84060 34260 84240
rect 36105 84240 37395 84360
rect 39540 84360 39660 84540
rect 46605 84540 46995 84660
rect 47205 84540 48795 84660
rect 60705 84540 65595 84660
rect 67905 84540 70395 84660
rect 72705 84540 75360 84660
rect 38505 84240 39660 84360
rect 75240 84360 75360 84540
rect 76905 84540 79395 84660
rect 87705 84540 88095 84660
rect 88305 84540 89895 84660
rect 75240 84240 75795 84360
rect 76005 84240 78495 84360
rect 34140 83940 34995 84060
rect 37005 83955 37995 84075
rect 40005 83940 40260 84060
rect 29040 83760 29160 83910
rect 20940 83640 29160 83760
rect 20940 83460 21060 83640
rect 40140 83505 40260 83940
rect 44505 83955 44895 84075
rect 47805 83955 49095 84075
rect 40995 83760 41205 83895
rect 40995 83700 41760 83760
rect 41040 83640 41760 83700
rect 19740 83340 21060 83460
rect 23205 83340 23895 83460
rect 25005 83325 25695 83445
rect 28005 83340 28695 83460
rect 32505 83340 33795 83460
rect 41640 83490 41760 83640
rect 41940 83205 42060 83910
rect 49305 83955 49995 84075
rect 57105 83940 57495 84060
rect 48405 83340 49560 83460
rect 7305 83040 7995 83160
rect 29505 83040 31695 83160
rect 34905 83040 35895 83160
rect 43305 83040 44295 83160
rect 49440 83160 49560 83340
rect 52140 83460 52260 83910
rect 53340 83760 53460 83910
rect 55440 83760 55560 83910
rect 53340 83700 53760 83760
rect 54540 83700 55560 83760
rect 53340 83640 53805 83700
rect 49905 83340 52260 83460
rect 53595 83505 53805 83640
rect 54495 83640 55560 83700
rect 54495 83505 54705 83640
rect 58140 83505 58260 83895
rect 59040 83505 59160 83910
rect 61605 83955 61995 84075
rect 64305 83955 64695 84075
rect 66705 83955 67095 84075
rect 71340 83940 71595 84060
rect 60240 83505 60360 83895
rect 55305 83340 57780 83460
rect 59040 83340 59295 83505
rect 59100 83295 59295 83340
rect 62940 83460 63060 83910
rect 62940 83340 64995 83460
rect 65340 83460 65460 83910
rect 69540 83505 69660 83910
rect 65340 83340 67395 83460
rect 69540 83340 69795 83505
rect 69600 83295 69795 83340
rect 49440 83040 51495 83160
rect 52140 83040 53295 83160
rect 705 82740 1995 82860
rect 13305 82740 13995 82860
rect 14205 82740 19995 82860
rect 20205 82740 20895 82860
rect 22605 82740 25395 82860
rect 32505 82740 33495 82860
rect 34305 82740 34695 82860
rect 34905 82740 35295 82860
rect 45405 82740 45795 82860
rect 52140 82860 52260 83040
rect 62805 83040 63795 83160
rect 71340 83160 71460 83940
rect 75540 83940 77295 84060
rect 73740 83760 73860 83895
rect 75540 83760 75660 83940
rect 79305 83940 81060 84060
rect 72240 83700 75660 83760
rect 72195 83640 75660 83700
rect 80940 83760 81060 83940
rect 82905 83940 83595 84060
rect 84000 84060 84195 84105
rect 83940 83895 84195 84060
rect 87240 83940 87495 84060
rect 80940 83640 81360 83760
rect 72195 83505 72405 83640
rect 74205 83340 76095 83460
rect 76905 83325 78195 83445
rect 81240 83460 81360 83640
rect 83940 83490 84060 83895
rect 85140 83505 85260 83895
rect 81240 83340 82395 83460
rect 86340 83460 86460 83910
rect 86340 83340 86895 83460
rect 69405 83040 71460 83160
rect 82905 83040 83595 83160
rect 87240 83160 87360 83940
rect 88005 83340 88995 83460
rect 90405 83340 91095 83460
rect 86205 83040 87360 83160
rect 50205 82740 52260 82860
rect 55005 82740 57795 82860
rect 60105 82740 60495 82860
rect 61305 82740 65595 82860
rect 65805 82740 66495 82860
rect 66705 82740 68895 82860
rect 69705 82740 72495 82860
rect 75705 82740 77895 82860
rect 81705 82740 87495 82860
rect 88305 82740 89295 82860
rect 22005 82440 24495 82560
rect 25905 82440 28395 82560
rect 29205 82440 31995 82560
rect 33105 82440 33795 82560
rect 34005 82440 35895 82560
rect 39405 82440 43995 82560
rect 47805 82440 52080 82560
rect 52605 82440 54495 82560
rect 55305 82440 58095 82560
rect 67005 82440 67995 82560
rect 70605 82440 71580 82560
rect 72105 82440 72795 82560
rect 75405 82440 77295 82560
rect 79905 82440 81195 82560
rect 1605 82140 1995 82260
rect 5505 82140 5895 82260
rect 6105 82140 6795 82260
rect 7005 82140 9795 82260
rect 25605 82140 36495 82260
rect 47205 82140 48495 82260
rect 50505 82140 50895 82260
rect 3105 81840 4395 81960
rect 20505 81840 21780 81960
rect 22305 81840 29280 81960
rect 29805 81840 34695 81960
rect 40005 81840 42060 81960
rect 1005 81540 3795 81660
rect 15105 81540 16695 81660
rect 30405 81540 33195 81660
rect 41940 81660 42060 81840
rect 43305 81840 44895 81960
rect 45105 81840 45495 81960
rect 46305 81840 50295 81960
rect 50940 81960 51060 82095
rect 52605 82140 53595 82260
rect 53805 82140 56595 82260
rect 58905 82140 62295 82260
rect 63405 82140 69495 82260
rect 70305 82140 73695 82260
rect 78105 82140 82560 82260
rect 82440 82005 82560 82140
rect 84105 82140 84795 82260
rect 90105 82140 91395 82260
rect 50940 81840 52995 81960
rect 53205 81840 53895 81960
rect 56205 81840 58395 81960
rect 71805 81840 72780 81960
rect 73305 81840 76095 81960
rect 78705 81840 79995 81960
rect 82605 81840 87195 81960
rect 41940 81540 42795 81660
rect 48405 81540 49095 81660
rect 54705 81540 58995 81660
rect 59805 81540 61095 81660
rect 63240 81540 65895 81660
rect 4605 81240 6195 81360
rect 8505 81240 11295 81360
rect 11505 81240 12495 81360
rect 13905 81240 17595 81360
rect 26505 81240 26895 81360
rect 34305 81240 35295 81360
rect 39105 81240 40695 81360
rect 48105 81240 52995 81360
rect 63240 81360 63360 81540
rect 68205 81540 70695 81660
rect 77505 81540 90495 81660
rect 90705 81540 91395 81660
rect 91605 81540 92760 81660
rect 61605 81240 63360 81360
rect 66405 81240 69195 81360
rect 71505 81240 72480 81360
rect 73005 81240 75195 81360
rect 79005 81240 79980 81360
rect 80505 81240 82995 81360
rect 84705 81240 85395 81360
rect 86205 81240 89295 81360
rect 3405 80940 4095 81060
rect 8805 80940 9195 81060
rect 9405 80940 10095 81060
rect 38205 80940 39195 81060
rect 47205 80940 47595 81060
rect 49605 80940 50595 81060
rect 51405 81060 51600 81105
rect 51405 80895 51660 81060
rect 78105 80940 78495 81060
rect 79305 80940 80895 81060
rect 86505 80940 86895 81060
rect 405 80655 1995 80775
rect 6240 80640 7695 80760
rect 3405 80025 4095 80145
rect 6240 79905 6360 80640
rect 10905 80640 11595 80760
rect 13305 80640 13860 80760
rect 13740 80460 13860 80640
rect 14205 80655 14595 80775
rect 15405 80640 16095 80760
rect 17940 80640 19095 80760
rect 13740 80340 14460 80460
rect 8805 80025 9195 80145
rect 10005 80025 11295 80145
rect 14340 80160 14460 80340
rect 17940 80190 18060 80640
rect 19905 80640 20895 80760
rect 23505 80640 24495 80760
rect 24705 80640 26295 80760
rect 27705 80640 28095 80760
rect 28305 80655 28695 80775
rect 30405 80655 30795 80775
rect 37605 80640 38160 80760
rect 14340 80040 14895 80160
rect 2505 79740 2895 79860
rect 9240 79860 9360 79980
rect 9240 79740 12195 79860
rect 27105 79740 28095 79860
rect 34140 79860 34260 80595
rect 34740 80460 34860 80610
rect 34440 80400 34860 80460
rect 34395 80340 34860 80400
rect 34395 80205 34605 80340
rect 36405 80040 36795 80160
rect 38040 80160 38160 80640
rect 40140 80190 40260 80895
rect 40905 80655 41295 80775
rect 43440 80205 43560 80610
rect 45705 80640 47760 80760
rect 47640 80460 47760 80640
rect 51540 80760 51660 80895
rect 51540 80640 51960 80760
rect 47640 80400 48960 80460
rect 47640 80340 49005 80400
rect 48795 80205 49005 80340
rect 38040 80040 39495 80160
rect 42405 80025 42795 80145
rect 43305 80040 43560 80205
rect 43305 79995 43500 80040
rect 44505 80040 45495 80160
rect 47505 80040 47895 80160
rect 50040 80160 50160 80595
rect 49905 80040 50160 80160
rect 50805 80025 51195 80145
rect 51840 79905 51960 80640
rect 52440 80190 52560 80895
rect 53205 80640 53760 80760
rect 53640 80190 53760 80640
rect 54105 80640 55695 80760
rect 56505 80640 57180 80760
rect 57705 80640 58860 80760
rect 58740 80460 58860 80640
rect 59205 80640 62160 80760
rect 58740 80400 61845 80460
rect 58740 80340 61905 80400
rect 61695 80205 61905 80340
rect 54405 80040 58680 80160
rect 59205 80025 60195 80145
rect 61890 80100 61905 80205
rect 62040 80190 62160 80640
rect 63105 80640 66495 80760
rect 66705 80640 67395 80760
rect 68505 80640 68760 80760
rect 68640 80460 68760 80640
rect 69105 80655 71895 80775
rect 73305 80655 74295 80775
rect 75540 80640 76995 80760
rect 68640 80340 69960 80460
rect 62805 80040 63795 80160
rect 64905 80040 65595 80160
rect 69840 80190 69960 80340
rect 74940 80205 75060 80595
rect 67605 80025 67995 80145
rect 75540 79905 75660 80640
rect 80505 80640 81060 80760
rect 77640 80160 77760 80595
rect 76605 80040 77760 80160
rect 78240 80160 78360 80595
rect 80940 80460 81060 80640
rect 83400 80760 83595 80805
rect 81705 80640 82860 80760
rect 80940 80340 81360 80460
rect 78240 80040 78795 80160
rect 81240 80190 81360 80340
rect 82740 80190 82860 80640
rect 83340 80595 83595 80760
rect 83340 80190 83460 80595
rect 80205 80040 80595 80160
rect 84840 80160 84960 80610
rect 91500 80760 91695 80805
rect 91440 80595 91695 80760
rect 84840 80040 85995 80160
rect 87540 80160 87660 80595
rect 91440 80205 91560 80595
rect 87405 80040 87660 80160
rect 88005 80040 88995 80160
rect 91440 80040 91695 80205
rect 91500 79995 91695 80040
rect 34140 79740 34695 79860
rect 41805 79740 43695 79860
rect 51705 79740 51960 79905
rect 51705 79695 51900 79740
rect 64605 79740 70695 79860
rect 70905 79740 71295 79860
rect 72105 79740 74595 79860
rect 75405 79740 75660 79905
rect 75405 79695 75600 79740
rect 2940 79560 3060 79695
rect 2940 79440 5895 79560
rect 10605 79440 12795 79560
rect 14805 79440 15495 79560
rect 16305 79440 19395 79560
rect 27405 79440 28995 79560
rect 31305 79440 32295 79560
rect 32505 79440 34995 79560
rect 36705 79440 38595 79560
rect 41640 79560 41760 79695
rect 40005 79440 41760 79560
rect 51540 79560 51660 79695
rect 51540 79440 54195 79560
rect 57405 79440 59895 79560
rect 61305 79440 63195 79560
rect 65505 79440 66795 79560
rect 71340 79440 73095 79560
rect 1605 79140 4680 79260
rect 5205 79140 7995 79260
rect 17505 79140 18795 79260
rect 34305 79140 37095 79260
rect 43305 79140 46395 79260
rect 46605 79140 48195 79260
rect 48405 79140 59595 79260
rect 71340 79260 71460 79440
rect 73305 79440 75495 79560
rect 82605 79440 85095 79560
rect 87405 79440 88395 79560
rect 66405 79140 71460 79260
rect 76305 79140 78195 79260
rect 81405 79140 85695 79260
rect 87105 79140 90195 79260
rect 91005 79140 93165 79260
rect 6705 78840 22095 78960
rect 23805 78840 26595 78960
rect 26805 78840 30195 78960
rect 31005 78840 31695 78960
rect 33705 78840 38280 78960
rect 38805 78840 39195 78960
rect 39405 78840 42060 78960
rect 6540 78660 6660 78795
rect 405 78540 6660 78660
rect 8505 78540 13995 78660
rect 17205 78540 18495 78660
rect 22605 78540 24795 78660
rect 25005 78540 28680 78660
rect 29205 78540 32895 78660
rect 34605 78540 34995 78660
rect 41940 78660 42060 78840
rect 43605 78840 43995 78960
rect 52005 78840 55995 78960
rect 58905 78840 63495 78960
rect 67305 78840 73395 78960
rect 74805 78840 75795 78960
rect 76740 78840 86295 78960
rect 41940 78540 45195 78660
rect 47805 78540 48195 78660
rect 50205 78540 52395 78660
rect 52605 78540 55695 78660
rect 58305 78540 58995 78660
rect 59805 78540 64995 78660
rect 76740 78660 76860 78840
rect 67605 78540 76860 78660
rect 77205 78540 81195 78660
rect 86805 78540 88095 78660
rect 3105 78240 5295 78360
rect 30405 78240 31095 78360
rect 41805 78240 45795 78360
rect 50505 78240 56595 78360
rect 60705 78240 62295 78360
rect 65805 78240 66795 78360
rect 70005 78240 70995 78360
rect 71205 78240 74595 78360
rect 76005 78240 79695 78360
rect 80805 78240 90795 78360
rect 7905 77940 10395 78060
rect 16605 77940 17595 78060
rect 23205 77940 28095 78060
rect 28905 77940 32295 78060
rect 39405 77940 40695 78060
rect 43905 77940 48795 78060
rect 51105 77940 52695 78060
rect 62805 77940 64395 78060
rect 65205 77940 67695 78060
rect 73905 77940 76095 78060
rect 79005 77940 82695 78060
rect 82905 77940 85995 78060
rect 86205 77940 90495 78060
rect 21105 77640 31095 77760
rect 32205 77640 32895 77760
rect 39105 77640 41295 77760
rect 44805 77640 45195 77760
rect 53205 77640 54495 77760
rect 59505 77640 60495 77760
rect 64005 77640 68295 77760
rect 71805 77640 75060 77760
rect 74940 77505 75060 77640
rect 75705 77640 80580 77760
rect 81105 77640 85095 77760
rect 92250 77640 93165 77760
rect 11805 77340 14595 77460
rect 16605 77340 20595 77460
rect 22005 77340 24195 77460
rect 37905 77340 40095 77460
rect 44805 77340 46695 77460
rect 47505 77340 51495 77460
rect 55905 77340 57195 77460
rect 60405 77340 61995 77460
rect 63105 77340 68595 77460
rect 69705 77340 73995 77460
rect 75105 77340 76695 77460
rect 82005 77340 83895 77460
rect 1605 77040 4995 77160
rect 7005 77040 8295 77160
rect 49305 77040 53295 77160
rect 54105 77040 58395 77160
rect 61905 77040 62295 77160
rect 62505 77040 66195 77160
rect 85305 77040 87795 77160
rect 17505 76740 20295 76860
rect 26505 76740 31695 76860
rect 31905 76740 33060 76860
rect 5505 76440 10095 76560
rect 19605 76440 19995 76560
rect 22305 76440 22995 76560
rect 32940 76560 33060 76740
rect 37905 76740 38595 76860
rect 39705 76740 40395 76860
rect 55605 76740 56595 76860
rect 57705 76740 59295 76860
rect 60000 76860 60195 76905
rect 59940 76695 60195 76860
rect 60990 76695 61005 76800
rect 61305 76740 63360 76860
rect 32940 76440 35295 76560
rect 36105 76440 39195 76560
rect 1005 76155 1995 76275
rect 2205 76140 3795 76260
rect 4605 76155 7695 76275
rect 10905 76155 11295 76275
rect 12405 76140 13095 76260
rect 13440 76140 16395 76260
rect 13440 75960 13560 76140
rect 21405 76155 21795 76275
rect 24405 76155 24795 76275
rect 25005 76140 26295 76260
rect 27390 76095 27405 76200
rect 28905 76155 29295 76275
rect 32505 76140 34560 76260
rect 27195 75960 27405 76095
rect 12540 75840 13560 75960
rect 26340 75900 27405 75960
rect 26340 75840 27345 75900
rect 12540 75690 12660 75840
rect 705 75525 2295 75645
rect 2505 75540 3495 75660
rect 20505 75540 23895 75660
rect 26340 75660 26460 75840
rect 26205 75540 26460 75660
rect 27540 75660 27660 76110
rect 34440 75705 34560 76140
rect 38340 75960 38460 76110
rect 35205 75840 38460 75960
rect 26805 75540 27660 75660
rect 28605 75540 30795 75660
rect 38640 75690 38760 76440
rect 41940 76440 42495 76560
rect 39405 76140 40395 76260
rect 41940 75960 42060 76440
rect 59940 76560 60060 76695
rect 53505 76440 60060 76560
rect 60795 76560 61005 76695
rect 60795 76500 61395 76560
rect 60825 76440 61395 76500
rect 62205 76440 63060 76560
rect 42405 76140 44595 76260
rect 49605 76140 50895 76260
rect 45240 75960 45360 76110
rect 52305 76140 53895 76260
rect 56940 76140 58095 76260
rect 56040 75960 56160 76110
rect 41940 75840 42360 75960
rect 45240 75840 46260 75960
rect 37005 75525 37395 75645
rect 38805 75540 40695 75660
rect 42240 75405 42360 75840
rect 43905 75540 44895 75660
rect 46140 75660 46260 75840
rect 55440 75840 56160 75960
rect 46140 75540 46395 75660
rect 47805 75525 49095 75645
rect 50505 75525 52395 75645
rect 52605 75540 52995 75660
rect 55440 75660 55560 75840
rect 54405 75540 55560 75660
rect 56940 75660 57060 76140
rect 59205 76260 59400 76305
rect 59205 76095 59460 76260
rect 55905 75540 57060 75660
rect 59340 75660 59460 76095
rect 61740 75705 61860 76110
rect 59340 75540 60195 75660
rect 61740 75540 61995 75705
rect 61800 75495 61995 75540
rect 62940 75660 63060 76440
rect 63240 76260 63360 76740
rect 68505 76740 72495 76860
rect 75105 76740 77595 76860
rect 82305 76740 84195 76860
rect 84405 76740 89895 76860
rect 90105 76740 91395 76860
rect 63705 76440 65160 76560
rect 65040 76260 65160 76440
rect 66405 76440 68805 76560
rect 68595 76320 68805 76440
rect 72405 76440 73695 76560
rect 77505 76440 77895 76560
rect 87540 76440 88395 76560
rect 63240 76140 63660 76260
rect 65040 76140 67380 76260
rect 63540 75960 63660 76140
rect 65340 75960 65460 76140
rect 67905 76140 68160 76260
rect 63540 75840 65160 75960
rect 65340 75840 65760 75960
rect 65040 75705 65160 75840
rect 62940 75540 63495 75660
rect 63705 75540 64695 75660
rect 65040 75540 65295 75705
rect 65100 75495 65295 75540
rect 65640 75660 65760 75840
rect 68040 75705 68160 76140
rect 68805 76140 70395 76260
rect 65640 75540 67395 75660
rect 70905 75540 72195 75660
rect 73140 75660 73260 76110
rect 77640 76140 78795 76260
rect 76440 75705 76560 76095
rect 73140 75540 74895 75660
rect 77640 75690 77760 76140
rect 79605 76155 80280 76275
rect 80805 76155 81195 76275
rect 81600 76260 81795 76305
rect 81540 76095 81795 76260
rect 83940 76140 85695 76260
rect 81540 75690 81660 76095
rect 82440 75660 82560 76095
rect 83940 75960 84060 76140
rect 87540 76260 87660 76440
rect 88605 76440 89595 76560
rect 85905 76140 87660 76260
rect 88005 76140 89760 76260
rect 83640 75840 84060 75960
rect 83640 75690 83760 75840
rect 89640 75690 89760 76140
rect 90705 76155 91095 76275
rect 82440 75540 82995 75660
rect 84405 75525 85395 75645
rect 1905 75240 5295 75360
rect 10605 75240 11595 75360
rect 13305 75240 14895 75360
rect 18405 75240 18795 75360
rect 19605 75240 19995 75360
rect 20205 75240 22095 75360
rect 27105 75240 27795 75360
rect 28905 75240 29295 75360
rect 35505 75240 36195 75360
rect 46005 75240 49695 75360
rect 54705 75240 55095 75360
rect 58005 75240 58380 75360
rect 58905 75240 61095 75360
rect 66705 75240 69495 75360
rect 71205 75240 71595 75360
rect 76005 75240 77295 75360
rect 89205 75240 91395 75360
rect 7605 74940 9495 75060
rect 23805 74940 25095 75060
rect 25305 74940 26295 75060
rect 30705 74940 32895 75060
rect 52605 74940 55695 75060
rect 58740 75060 58860 75195
rect 57105 74940 58860 75060
rect 61905 74940 63195 75060
rect 73005 74940 79560 75060
rect 4305 74640 6495 74760
rect 13905 74640 15960 74760
rect 6405 74340 7695 74460
rect 8805 74340 11295 74460
rect 11505 74340 11880 74460
rect 12405 74340 14295 74460
rect 15840 74460 15960 74640
rect 16305 74640 17595 74760
rect 24105 74640 26595 74760
rect 29805 74640 31995 74760
rect 32205 74640 33795 74760
rect 36405 74640 43995 74760
rect 49605 74640 52095 74760
rect 53505 74640 53895 74760
rect 55005 74640 56295 74760
rect 57405 74640 60195 74760
rect 60405 74640 61395 74760
rect 61605 74640 64095 74760
rect 65805 74640 66795 74760
rect 67005 74640 70095 74760
rect 71205 74640 72495 74760
rect 74505 74640 78195 74760
rect 79440 74760 79560 74940
rect 79905 74940 81195 75060
rect 86205 74940 87495 75060
rect 88305 74940 88695 75060
rect 88905 74940 91095 75060
rect 79440 74640 79995 74760
rect 80805 74640 81495 74760
rect 85005 74640 85695 74760
rect 15840 74340 25995 74460
rect 34605 74340 42495 74460
rect 42705 74340 44295 74460
rect 44505 74340 45795 74460
rect 48405 74340 50895 74460
rect 63105 74340 63495 74460
rect 64905 74340 68295 74460
rect 70140 74460 70260 74595
rect 70140 74340 70695 74460
rect 77205 74340 80295 74460
rect 85605 74340 86295 74460
rect 87405 74340 88095 74460
rect 15405 74040 19095 74160
rect 22005 74040 25695 74160
rect 47805 74040 49395 74160
rect 52305 74040 56595 74160
rect 56805 74040 57195 74160
rect 62205 74040 64395 74160
rect 69405 74040 70995 74160
rect 71805 74040 74895 74160
rect 80805 74040 83895 74160
rect 87105 74040 88395 74160
rect 19905 73740 24795 73860
rect 36105 73740 37095 73860
rect 37305 73740 37680 73860
rect 38205 73740 38895 73860
rect 47205 73740 50895 73860
rect 52005 73740 56895 73860
rect 59205 73740 59895 73860
rect 61005 73740 61695 73860
rect 63105 73740 69495 73860
rect 75705 73740 76695 73860
rect 90405 73740 91860 73860
rect 91740 73605 91860 73740
rect 6105 73440 7395 73560
rect 23505 73440 25395 73560
rect 25605 73440 27195 73560
rect 31305 73440 32295 73560
rect 35505 73440 36495 73560
rect 39405 73440 41895 73560
rect 42705 73440 44895 73560
rect 45105 73440 45795 73560
rect 48105 73440 49695 73560
rect 51705 73440 58695 73560
rect 62805 73440 65895 73560
rect 68505 73440 69795 73560
rect 74205 73440 79995 73560
rect 84705 73440 85695 73560
rect 91740 73440 91995 73605
rect 91800 73395 91995 73440
rect 2805 73140 3495 73260
rect 3705 73140 8295 73260
rect 8505 73140 10395 73260
rect 14640 73140 15195 73260
rect 1905 72840 2460 72960
rect 2340 72405 2460 72840
rect 4305 72840 4695 72960
rect 5805 72855 7095 72975
rect 8640 72840 8895 72960
rect 8640 72660 8760 72840
rect 11205 72840 12795 72960
rect 14640 72660 14760 73140
rect 39105 73140 40260 73260
rect 16605 72855 16695 72975
rect 16905 72855 16995 72975
rect 18105 72840 19695 72960
rect 20505 72855 21195 72975
rect 24105 72840 24795 72960
rect 33405 72840 34095 72960
rect 7740 72540 8760 72660
rect 13140 72540 14760 72660
rect 27240 72660 27360 72810
rect 27240 72540 29460 72660
rect 4905 72225 5895 72345
rect 7740 72360 7860 72540
rect 6705 72300 8460 72360
rect 6705 72240 8505 72300
rect 8295 72105 8505 72240
rect 10005 72240 12195 72360
rect 13140 72390 13260 72540
rect 14640 72390 14760 72540
rect 15405 72240 17295 72360
rect 23205 72240 25695 72360
rect 25905 72240 27795 72360
rect 28005 72225 28695 72345
rect 29340 72360 29460 72540
rect 29340 72240 29595 72360
rect 31305 72240 32895 72360
rect 33705 72225 34395 72345
rect 35040 72360 35160 73095
rect 35040 72240 36195 72360
rect 40140 72390 40260 73140
rect 55605 73140 57360 73260
rect 41505 72840 42495 72960
rect 45705 72840 46860 72960
rect 43140 72660 43260 72810
rect 43140 72540 45060 72660
rect 40905 72225 41295 72345
rect 42105 72225 42795 72345
rect 44940 72360 45060 72540
rect 44940 72240 45360 72360
rect 2205 71940 2595 72060
rect 20205 71940 21795 72060
rect 22005 71940 28995 72060
rect 35805 71940 39195 72060
rect 42795 72060 43005 72180
rect 45240 72105 45360 72240
rect 42795 71940 44595 72060
rect 45240 71940 45495 72105
rect 45300 71895 45495 71940
rect 46740 72060 46860 72840
rect 47505 72840 48495 72960
rect 49905 72840 52860 72960
rect 52740 72660 52860 72840
rect 53505 72840 54195 72960
rect 55005 72840 55695 72960
rect 52740 72540 53160 72660
rect 53040 72390 53160 72540
rect 48105 72225 49395 72345
rect 53205 72240 55995 72360
rect 46740 71940 47595 72060
rect 56340 72060 56460 72795
rect 57240 72390 57360 73140
rect 60705 73140 62895 73260
rect 57705 72840 58260 72960
rect 58140 72405 58260 72840
rect 59640 72390 59760 73095
rect 60105 72840 60960 72960
rect 60840 72660 60960 72840
rect 61305 72855 61995 72975
rect 60840 72540 62460 72660
rect 60405 72240 61095 72360
rect 62340 72390 62460 72540
rect 62640 72105 62760 73140
rect 67305 73140 67695 73260
rect 71205 73140 72795 73260
rect 77805 73140 78495 73260
rect 78705 73140 79095 73260
rect 83805 73140 84195 73260
rect 86505 73140 87060 73260
rect 62940 72405 63060 72780
rect 66540 72660 66660 72810
rect 69105 72840 70695 72960
rect 71040 72840 71295 72960
rect 63405 72540 66660 72660
rect 64905 72240 66195 72360
rect 66405 72240 66795 72360
rect 56340 71940 56895 72060
rect 61905 71940 62595 72060
rect 67440 72060 67560 72795
rect 68340 72660 68460 72810
rect 68040 72600 68460 72660
rect 67995 72540 68460 72600
rect 67995 72405 68205 72540
rect 71040 72660 71160 72840
rect 74205 72840 74895 72960
rect 75240 72840 75495 72960
rect 75240 72660 75360 72840
rect 77205 72840 77895 72960
rect 81795 72960 82005 73095
rect 81795 72900 82695 72960
rect 81840 72840 82695 72900
rect 70305 72540 71160 72660
rect 74940 72540 75360 72660
rect 71805 72240 73395 72360
rect 74940 72105 75060 72540
rect 76140 72405 76260 72795
rect 76905 72225 77595 72345
rect 78840 72360 78960 72795
rect 83340 72405 83460 72795
rect 83895 72660 84105 72795
rect 83895 72600 84660 72660
rect 83940 72540 84660 72600
rect 78540 72300 78960 72360
rect 78495 72240 78960 72300
rect 78495 72105 78705 72240
rect 79305 72225 79695 72345
rect 81405 72225 82395 72345
rect 84540 72390 84660 72540
rect 85440 72405 85560 72795
rect 86640 72660 86760 72810
rect 86340 72600 86760 72660
rect 86295 72540 86760 72600
rect 86940 72660 87060 73140
rect 87405 72840 91395 72960
rect 86940 72540 87660 72660
rect 86295 72405 86505 72540
rect 87540 72390 87660 72540
rect 67440 71940 68295 72060
rect 4005 71640 4995 71760
rect 10905 71640 13095 71760
rect 19005 71640 20895 71760
rect 24705 71640 28095 71760
rect 30105 71640 31695 71760
rect 48405 71640 51195 71760
rect 52005 71640 54195 71760
rect 55005 71640 57795 71760
rect 61305 71640 64995 71760
rect 67005 71640 68595 71760
rect 70305 71640 73095 71760
rect 77205 71640 80295 71760
rect 84705 71640 86895 71760
rect 16605 71340 23295 71460
rect 23505 71340 23895 71460
rect 32205 71340 37995 71460
rect 49605 71340 50295 71460
rect 59505 71340 65595 71460
rect 65805 71340 66195 71460
rect 67800 71460 67995 71505
rect 67740 71295 67995 71460
rect 70005 71340 72660 71460
rect 1605 71040 2895 71160
rect 3105 71040 3195 71160
rect 3405 71040 7995 71160
rect 8205 71040 10995 71160
rect 20505 71040 29895 71160
rect 30105 71040 33795 71160
rect 34140 71040 35895 71160
rect 5205 70740 8595 70860
rect 11505 70740 15795 70860
rect 18840 70740 20295 70860
rect 11805 70440 17895 70560
rect 18840 70560 18960 70740
rect 21105 70740 26895 70860
rect 34140 70860 34260 71040
rect 43605 71040 53595 71160
rect 58740 71040 63495 71160
rect 31905 70740 34260 70860
rect 36705 70740 45195 70860
rect 45405 70740 49995 70860
rect 58740 70860 58860 71040
rect 67740 71160 67860 71295
rect 64305 71040 67860 71160
rect 72540 71160 72660 71340
rect 73605 71340 90795 71460
rect 72540 71040 77595 71160
rect 78405 71040 78795 71160
rect 79005 71040 80595 71160
rect 56805 70740 58860 70860
rect 59205 70740 60795 70860
rect 63105 70740 67380 70860
rect 67905 70740 69495 70860
rect 70605 70740 75195 70860
rect 18105 70440 18960 70560
rect 19605 70440 27195 70560
rect 27405 70440 31395 70560
rect 32640 70440 35295 70560
rect 7305 70140 9195 70260
rect 22605 70140 24195 70260
rect 24405 70140 25095 70260
rect 32640 70260 32760 70440
rect 36405 70440 43695 70560
rect 45705 70440 49095 70560
rect 54405 70440 55395 70560
rect 60105 70440 63195 70560
rect 65505 70440 70680 70560
rect 71205 70440 78195 70560
rect 79005 70440 82095 70560
rect 82305 70440 83295 70560
rect 29205 70140 32760 70260
rect 33105 70140 44160 70260
rect 405 69840 11595 69960
rect 18405 69840 19395 69960
rect 26205 69840 34995 69960
rect 36105 69840 40395 69960
rect 44040 69960 44160 70140
rect 53505 70140 54795 70260
rect 55005 70140 55395 70260
rect 58905 70140 64995 70260
rect 69405 70140 72195 70260
rect 73305 70140 84795 70260
rect 44040 69840 46095 69960
rect 49305 69840 59895 69960
rect 61605 69840 62895 69960
rect 67605 69840 69195 69960
rect 80505 69840 84495 69960
rect 88605 69840 91395 69960
rect 13305 69540 17295 69660
rect 21105 69540 23895 69660
rect 24105 69540 40995 69660
rect 43305 69540 43995 69660
rect 49005 69540 53280 69660
rect 53805 69540 62760 69660
rect 7605 69240 14595 69360
rect 25905 69240 28380 69360
rect 28905 69240 32760 69360
rect 1305 68940 3495 69060
rect 15705 68940 16095 69060
rect 32640 69060 32760 69240
rect 34605 69240 36495 69360
rect 57405 69240 62295 69360
rect 62640 69360 62760 69540
rect 65205 69540 69795 69660
rect 76305 69540 77295 69660
rect 78405 69540 82995 69660
rect 85905 69540 87495 69660
rect 62640 69240 64095 69360
rect 68205 69240 69495 69360
rect 76605 69240 77895 69360
rect 82905 69240 83595 69360
rect 85005 69240 88695 69360
rect 32640 68940 35595 69060
rect 38205 68940 39195 69060
rect 40005 68940 43995 69060
rect 46605 68940 52395 69060
rect 58305 68940 66780 69060
rect 67305 68940 68595 69060
rect 71205 68940 72195 69060
rect 74805 68940 80295 69060
rect 81405 68940 83295 69060
rect 11205 68640 16260 68760
rect 705 68355 1095 68475
rect 1905 68355 2280 68475
rect 4605 68340 5895 68460
rect 6705 68340 7695 68460
rect 8505 68340 10095 68460
rect 2640 67860 2760 68295
rect 7740 68160 7860 68310
rect 10740 68160 10860 68310
rect 11805 68340 12195 68460
rect 15705 68460 15900 68505
rect 16140 68460 16260 68640
rect 17205 68640 18195 68760
rect 32505 68640 33195 68760
rect 44505 68640 45195 68760
rect 65940 68640 67695 68760
rect 15705 68295 15960 68460
rect 16140 68340 18360 68460
rect 7740 68040 10860 68160
rect 15840 68160 15960 68295
rect 15840 68040 18060 68160
rect 2640 67740 3195 67860
rect 4905 67740 5595 67860
rect 8205 67740 10395 67860
rect 9105 67440 9495 67560
rect 10740 67560 10860 68040
rect 12105 67740 15495 67860
rect 17940 67890 18060 68040
rect 16605 67725 17580 67845
rect 18240 67860 18360 68340
rect 19005 68355 19695 68475
rect 23505 68340 25095 68460
rect 25440 68340 25695 68460
rect 22740 68160 22860 68310
rect 25440 68160 25560 68340
rect 22140 68100 22860 68160
rect 22095 68040 22860 68100
rect 23040 68040 25560 68160
rect 22095 67905 22305 68040
rect 18240 67740 18495 67860
rect 19905 67740 20595 67860
rect 23040 67890 23160 68040
rect 26805 67740 27195 67860
rect 10740 67440 13395 67560
rect 27540 67560 27660 68310
rect 28305 68340 29295 68460
rect 29505 68355 30795 68475
rect 35505 68355 42195 68475
rect 42405 68340 43395 68460
rect 28605 67740 31695 67860
rect 32040 67860 32160 68310
rect 45840 68340 46395 68460
rect 45840 68160 45960 68340
rect 47505 68340 48495 68460
rect 49905 68340 54195 68460
rect 56205 68355 57195 68475
rect 60405 68340 61695 68460
rect 62400 68460 62595 68505
rect 62340 68295 62595 68460
rect 64005 68355 64395 68475
rect 37005 68040 40560 68160
rect 32040 67740 32595 67860
rect 40440 67860 40560 68040
rect 44940 68040 45960 68160
rect 40440 67740 42495 67860
rect 42705 67740 43695 67860
rect 44940 67860 45060 68040
rect 44505 67740 45060 67860
rect 45405 67725 46095 67845
rect 56805 67740 57495 67860
rect 62340 67605 62460 68295
rect 65940 68160 66060 68640
rect 69705 68640 70695 68760
rect 73605 68640 74295 68760
rect 76695 68640 79695 68760
rect 76695 68520 76905 68640
rect 92205 68760 92400 68805
rect 92205 68595 92460 68760
rect 67005 68340 68460 68460
rect 65640 68040 66060 68160
rect 68340 68160 68460 68340
rect 68805 68340 75360 68460
rect 75240 68205 75360 68340
rect 76005 68355 76695 68475
rect 80400 68460 80595 68505
rect 68340 68100 68760 68160
rect 68340 68040 68805 68100
rect 75240 68040 75495 68205
rect 65640 67890 65760 68040
rect 68595 67905 68805 68040
rect 75300 67995 75495 68040
rect 63105 67725 63495 67845
rect 77340 67905 77460 68310
rect 79140 67905 79260 68310
rect 80340 68295 80595 68460
rect 80340 67905 80460 68295
rect 70605 67725 74295 67845
rect 77340 67740 77595 67905
rect 77400 67695 77595 67740
rect 79005 67740 79260 67905
rect 79005 67695 79200 67740
rect 81540 67860 81660 68595
rect 82005 68340 82395 68460
rect 84405 68340 84660 68460
rect 84540 67905 84660 68340
rect 81540 67740 82095 67860
rect 85740 67605 85860 68595
rect 89205 68340 90960 68460
rect 88395 68160 88605 68295
rect 88395 68100 88860 68160
rect 88440 68040 88860 68100
rect 88740 67890 88860 68040
rect 90840 67890 90960 68340
rect 91305 68355 91995 68475
rect 92340 68160 92460 68595
rect 91740 68100 92460 68160
rect 91695 68040 92460 68100
rect 91695 67905 91905 68040
rect 26205 67440 27660 67560
rect 28605 67440 32895 67560
rect 35505 67440 42195 67560
rect 47205 67440 47595 67560
rect 60105 67440 61980 67560
rect 69105 67440 69795 67560
rect 75105 67440 75795 67560
rect 81105 67440 82995 67560
rect 87705 67440 88095 67560
rect 2805 67140 4395 67260
rect 12405 67140 12795 67260
rect 16005 67140 18495 67260
rect 22305 67140 25395 67260
rect 26505 67140 27795 67260
rect 28005 67140 28695 67260
rect 31305 67140 32580 67260
rect 33105 67140 34395 67260
rect 43905 67140 49695 67260
rect 49905 67140 53295 67260
rect 54405 67140 57795 67260
rect 58605 67140 60195 67260
rect 63405 67140 64380 67260
rect 64905 67140 68595 67260
rect 69405 67140 70095 67260
rect 71805 67140 76395 67260
rect 76605 67140 78795 67260
rect 80805 67140 82095 67260
rect 88605 67140 91395 67260
rect 1605 66840 6195 66960
rect 6405 66840 7995 66960
rect 8805 66840 11595 66960
rect 17505 66840 21795 66960
rect 32505 66840 36795 66960
rect 43305 66840 58995 66960
rect 67605 66840 71295 66960
rect 72405 66840 79995 66960
rect 80205 66840 82695 66960
rect 82905 66840 83595 66960
rect 90105 66840 91395 66960
rect 17805 66540 19680 66660
rect 20205 66540 21195 66660
rect 37305 66540 39795 66660
rect 40605 66540 41895 66660
rect 44205 66540 45495 66660
rect 53805 66540 55695 66660
rect 60405 66540 65595 66660
rect 67905 66540 68895 66660
rect 69705 66540 73695 66660
rect 76605 66540 76995 66660
rect 78405 66540 80895 66660
rect 85905 66540 87195 66660
rect 14805 66240 16680 66360
rect 17205 66240 24795 66360
rect 28005 66240 29595 66360
rect 34605 66240 36495 66360
rect 37605 66240 37995 66360
rect 41205 66240 45795 66360
rect 46005 66240 48195 66360
rect 49605 66240 59595 66360
rect 61005 66240 63495 66360
rect 67305 66240 69195 66360
rect 70005 66240 70995 66360
rect 84105 66240 84495 66360
rect 89505 66240 90195 66360
rect 90405 66240 91695 66360
rect 9405 65940 9795 66060
rect 10005 65940 13095 66060
rect 14505 65940 14895 66060
rect 15105 65940 25095 66060
rect 28305 65940 31995 66060
rect 36405 65940 39495 66060
rect 40305 65940 40695 66060
rect 40905 65940 41595 66060
rect 51405 65940 53895 66060
rect 55905 65940 59295 66060
rect 67005 65940 69495 66060
rect 71205 65940 71595 66060
rect 73905 65940 76995 66060
rect 77205 65940 77895 66060
rect 85905 65940 86595 66060
rect 3705 65640 5595 65760
rect 13005 65640 22395 65760
rect 23805 65640 27195 65760
rect 37005 65640 40995 65760
rect 42105 65640 43695 65760
rect 49605 65640 49995 65760
rect 52005 65640 52995 65760
rect 64605 65640 67680 65760
rect 68205 65640 72195 65760
rect 76005 65640 76695 65760
rect 79305 65640 84495 65760
rect 89205 65640 91095 65760
rect 4605 65340 6795 65460
rect 11205 65340 11895 65460
rect 16605 65340 17295 65460
rect 18105 65340 19995 65460
rect 30105 65460 30300 65505
rect 30105 65295 30360 65460
rect 36705 65340 40395 65460
rect 59505 65340 61095 65460
rect 66105 65340 68295 65460
rect 69105 65340 70395 65460
rect 75105 65340 75495 65460
rect 85005 65340 85860 65460
rect 1005 65055 1395 65175
rect 2505 65040 3360 65160
rect 1905 64440 2595 64560
rect 3240 64590 3360 65040
rect 3840 64860 3960 65295
rect 4305 65055 4680 65175
rect 4995 64860 5205 64995
rect 7140 65040 7995 65160
rect 3840 64740 4860 64860
rect 4995 64800 5760 64860
rect 5040 64740 5760 64800
rect 4740 64560 4860 64740
rect 4740 64440 5295 64560
rect 5640 64560 5760 64740
rect 7140 64605 7260 65040
rect 17805 65040 18060 65160
rect 10140 64605 10260 65010
rect 17940 64605 18060 65040
rect 27540 65040 28095 65160
rect 19305 64740 20880 64860
rect 5640 64440 6495 64560
rect 10140 64440 10395 64605
rect 10200 64395 10395 64440
rect 12405 64425 15195 64545
rect 16005 64425 16395 64545
rect 17940 64440 18195 64605
rect 18000 64395 18195 64440
rect 21195 64560 21405 64695
rect 21195 64500 24495 64560
rect 21240 64440 24495 64500
rect 26640 64560 26760 65010
rect 27540 64590 27660 65040
rect 30240 65160 30360 65295
rect 30240 65040 35295 65160
rect 40440 65040 41295 65160
rect 36240 64605 36360 64995
rect 40440 64605 40560 65040
rect 42105 65160 42300 65205
rect 42105 64995 42360 65160
rect 43605 65040 43995 65160
rect 44640 65040 50595 65160
rect 42240 64605 42360 64995
rect 44640 64605 44760 65040
rect 51405 65040 52395 65160
rect 53400 65160 53595 65205
rect 53340 64995 53595 65160
rect 25905 64440 26760 64560
rect 53340 64590 53460 64995
rect 54540 64605 54660 65295
rect 55440 64605 55560 65010
rect 54540 64440 54795 64605
rect 54600 64395 54795 64440
rect 55440 64440 55695 64605
rect 55500 64395 55695 64440
rect 6105 64140 8295 64260
rect 8505 64140 9195 64260
rect 11805 64140 13995 64260
rect 14205 64140 15060 64260
rect 7005 63840 7695 63960
rect 14940 63960 15060 64140
rect 19905 64140 23295 64260
rect 29805 64140 31095 64260
rect 40005 64140 41895 64260
rect 56040 64260 56160 65040
rect 70440 65040 71895 65160
rect 57540 64605 57660 64995
rect 60840 64860 60960 65010
rect 59640 64740 60960 64860
rect 59640 64560 59760 64740
rect 58305 64440 59760 64560
rect 60105 64425 60495 64545
rect 61440 64560 61560 65010
rect 61440 64440 61995 64560
rect 63105 64440 68280 64560
rect 68805 64440 69195 64560
rect 69540 64305 69660 65010
rect 70140 64305 70260 65010
rect 70440 64590 70560 65040
rect 72705 65055 73395 65175
rect 73605 65040 74595 65160
rect 76140 64860 76260 65295
rect 75240 64800 76260 64860
rect 75195 64740 76260 64800
rect 75195 64605 75405 64740
rect 72405 64440 73995 64560
rect 76440 64305 76560 65010
rect 77505 65040 78195 65160
rect 80205 65040 81195 65160
rect 79305 64440 79695 64560
rect 53805 64140 56160 64260
rect 77040 64140 78795 64260
rect 14940 63840 17295 63960
rect 25305 63840 25995 63960
rect 37605 63840 40995 63960
rect 45405 63840 49095 63960
rect 54405 63840 55080 63960
rect 55605 63840 58695 63960
rect 59805 63840 61395 63960
rect 73005 63840 73395 63960
rect 73605 63840 74295 63960
rect 77040 63960 77160 64140
rect 81840 64275 81960 65010
rect 82440 64560 82560 64995
rect 85140 64605 85260 64995
rect 85740 64605 85860 65340
rect 86205 65340 88695 65460
rect 86805 65040 88095 65160
rect 88440 64605 88560 65340
rect 89640 64605 89760 64995
rect 82305 64440 82560 64560
rect 83205 64425 83595 64545
rect 81840 64140 82095 64275
rect 81900 64095 82095 64140
rect 84405 64140 84495 64260
rect 84705 64140 86295 64260
rect 88305 64140 88695 64260
rect 76005 63840 77160 63960
rect 87405 63840 87795 63960
rect 9105 63540 10695 63660
rect 11505 63540 16095 63660
rect 18705 63540 22095 63660
rect 25605 63540 25995 63660
rect 26205 63540 28395 63660
rect 31605 63540 32895 63660
rect 48105 63540 51795 63660
rect 64005 63540 67095 63660
rect 75705 63540 77295 63660
rect 79905 63540 83295 63660
rect 84105 63540 85095 63660
rect 89505 63540 90495 63660
rect 17205 63240 23880 63360
rect 24405 63240 29895 63360
rect 35805 63240 39795 63360
rect 40605 63240 41760 63360
rect 10005 62940 11595 63060
rect 18105 62940 19395 63060
rect 24105 62940 29595 63060
rect 41640 63060 41760 63240
rect 67905 63240 71895 63360
rect 72705 63240 74895 63360
rect 77805 63240 84795 63360
rect 41640 62940 44295 63060
rect 49005 62940 53595 63060
rect 55005 62940 56595 63060
rect 62205 62940 80595 63060
rect 12105 62640 13695 62760
rect 16905 62640 19995 62760
rect 23805 62640 37995 62760
rect 40740 62640 43095 62760
rect 40740 62505 40860 62640
rect 54705 62640 62895 62760
rect 72105 62640 75795 62760
rect 82905 62640 83595 62760
rect 23205 62340 33960 62460
rect 33840 62205 33960 62340
rect 38805 62340 40695 62460
rect 43605 62340 45195 62460
rect 46740 62340 55695 62460
rect 10605 62040 13395 62160
rect 13605 62040 16395 62160
rect 16605 62040 18195 62160
rect 34005 62040 36495 62160
rect 46740 62160 46860 62340
rect 57105 62340 60195 62460
rect 63705 62340 70995 62460
rect 72105 62340 73995 62460
rect 85440 62340 88395 62460
rect 36705 62040 46860 62160
rect 54105 62040 54795 62160
rect 69705 62040 76095 62160
rect 81105 62040 81495 62160
rect 85440 62160 85560 62340
rect 83205 62040 85560 62160
rect 25005 61740 30795 61860
rect 31005 61740 31695 61860
rect 32805 61740 33795 61860
rect 34005 61740 35460 61860
rect 16305 61440 18795 61560
rect 19005 61440 20595 61560
rect 21705 61440 25695 61560
rect 35340 61560 35460 61740
rect 39705 61740 48795 61860
rect 52905 61740 55095 61860
rect 55305 61740 57195 61860
rect 57405 61740 61095 61860
rect 62805 61740 63495 61860
rect 64905 61740 66795 61860
rect 67005 61740 68295 61860
rect 69705 61740 70095 61860
rect 74205 61740 75195 61860
rect 78405 61740 80295 61860
rect 86505 61740 86895 61860
rect 87105 61740 89295 61860
rect 89505 61740 90495 61860
rect 35340 61440 37095 61560
rect 40605 61440 42495 61560
rect 49905 61440 52395 61560
rect 65505 61440 69795 61560
rect 73305 61440 76995 61560
rect 77205 61440 77595 61560
rect 82305 61440 86895 61560
rect 1905 61140 4695 61260
rect 4905 61140 5895 61260
rect 7605 61140 11295 61260
rect 27105 61140 34395 61260
rect 3240 60840 3795 60960
rect 2505 60555 2895 60675
rect 3240 60105 3360 60840
rect 20205 60840 21495 60960
rect 24240 60840 25995 60960
rect 3705 60540 4995 60660
rect 5205 60540 7395 60660
rect 7605 60555 7995 60675
rect 8805 60540 10095 60660
rect 18105 60555 19095 60675
rect 21405 60540 22095 60660
rect 11805 60240 14295 60360
rect 1005 59940 1395 60060
rect 7740 60000 8295 60060
rect 7695 59940 8295 60000
rect 7695 59805 7905 59940
rect 19605 59940 22395 60060
rect 24240 60060 24360 60840
rect 28305 60840 28695 60960
rect 24705 60540 27195 60660
rect 27540 60540 28695 60660
rect 27540 60360 27660 60540
rect 29040 60360 29160 61140
rect 35205 61140 40095 61260
rect 43005 61140 49395 61260
rect 49605 61140 49995 61260
rect 56505 61140 58695 61260
rect 58905 61140 59595 61260
rect 60405 61140 61695 61260
rect 65805 61140 66195 61260
rect 74805 61140 76095 61260
rect 84405 61140 86295 61260
rect 86940 61260 87060 61380
rect 86940 61140 91395 61260
rect 32205 60840 33195 60960
rect 37305 60840 39195 60960
rect 39405 60840 39795 60960
rect 41040 60840 42195 60960
rect 29805 60555 30795 60675
rect 32505 60540 33195 60660
rect 33405 60540 34995 60660
rect 39495 60360 39705 60495
rect 26940 60240 27660 60360
rect 28440 60240 29160 60360
rect 38040 60300 39705 60360
rect 41040 60360 41160 60840
rect 61005 60840 63105 60960
rect 41505 60540 42795 60660
rect 43005 60540 43995 60660
rect 38040 60240 39660 60300
rect 41040 60240 42660 60360
rect 26940 60090 27060 60240
rect 28440 60090 28560 60240
rect 23505 59940 24360 60060
rect 31605 59940 35295 60060
rect 38040 60060 38160 60240
rect 42540 60090 42660 60240
rect 47640 60105 47760 60540
rect 48540 60360 48660 60540
rect 48540 60240 49395 60360
rect 35505 59940 38160 60060
rect 38805 59925 40395 60045
rect 41205 60000 41760 60060
rect 41205 59940 41805 60000
rect 41595 59805 41805 59940
rect 43305 59940 43695 60060
rect 43905 59940 44595 60060
rect 47505 59940 47760 60105
rect 50340 60090 50460 60795
rect 50640 60105 50760 60510
rect 52905 60540 53295 60660
rect 62895 60720 63105 60840
rect 63405 60840 64260 60960
rect 54405 60540 55395 60660
rect 54240 60105 54360 60540
rect 57705 60555 58095 60675
rect 63105 60555 63795 60675
rect 47505 59895 47700 59940
rect 50640 59940 50895 60105
rect 50700 59895 50895 59940
rect 51705 59895 52395 60015
rect 54240 59940 54495 60105
rect 54300 59895 54495 59940
rect 56205 59940 57495 60060
rect 2205 59640 3795 59760
rect 10905 59640 15195 59760
rect 25740 59640 26595 59760
rect 7305 59340 10095 59460
rect 19005 59340 20895 59460
rect 22005 59340 23595 59460
rect 25740 59460 25860 59640
rect 59340 59760 59460 60495
rect 61140 60060 61260 60495
rect 62040 60105 62160 60495
rect 60705 59940 61260 60060
rect 64140 60060 64260 60840
rect 76905 60840 77295 60960
rect 80805 60840 82995 60960
rect 89340 60840 91260 60960
rect 69105 60540 70395 60660
rect 71505 60540 72495 60660
rect 72840 60540 73395 60660
rect 65940 60105 66060 60495
rect 72840 60360 72960 60540
rect 78540 60540 78795 60660
rect 72540 60240 72960 60360
rect 63405 59940 64260 60060
rect 64905 59925 65295 60045
rect 68805 59940 69195 60060
rect 70905 59925 71295 60045
rect 72540 59805 72660 60240
rect 78540 60105 78660 60540
rect 80940 60600 84195 60660
rect 80895 60540 84195 60600
rect 80895 60390 81105 60540
rect 87105 60540 87360 60660
rect 86040 60105 86160 60495
rect 87240 60105 87360 60540
rect 89340 60660 89460 60840
rect 91140 60705 91260 60840
rect 88905 60540 89460 60660
rect 89805 60660 90000 60705
rect 89805 60495 90060 60660
rect 76605 59925 76995 60045
rect 84105 59940 85395 60060
rect 88740 60060 88860 60495
rect 88305 59940 88860 60060
rect 89940 60060 90060 60495
rect 90195 60360 90405 60495
rect 90195 60300 90960 60360
rect 90240 60240 90960 60300
rect 90840 60090 90960 60240
rect 89940 60000 90660 60060
rect 89940 59940 90705 60000
rect 90495 59805 90705 59940
rect 92040 60060 92160 60795
rect 92040 59940 92460 60060
rect 58005 59640 59460 59760
rect 60105 59640 61395 59760
rect 69705 59640 70095 59760
rect 24405 59340 25860 59460
rect 27105 59340 27495 59460
rect 29805 59340 31395 59460
rect 32205 59340 43095 59460
rect 49605 59340 51195 59460
rect 51405 59340 54495 59460
rect 54705 59340 68295 59460
rect 69105 59340 72795 59460
rect 76905 59340 79095 59460
rect 86805 59340 88095 59460
rect 89205 59340 91995 59460
rect 405 59040 6195 59160
rect 7605 59040 10395 59160
rect 12405 59040 13095 59160
rect 15105 59040 17895 59160
rect 18705 59040 21195 59160
rect 24105 59040 26595 59160
rect 28005 59040 30495 59160
rect 51540 59100 52395 59160
rect 51495 59040 52395 59100
rect 51495 58905 51705 59040
rect 57705 59040 66195 59160
rect 70005 59040 71895 59160
rect 73305 59040 76395 59160
rect 87705 59040 89595 59160
rect 92340 58905 92460 59940
rect 1905 58740 4995 58860
rect 10305 58740 12795 58860
rect 13440 58740 26295 58860
rect 2505 58440 4095 58560
rect 4305 58440 11295 58560
rect 13440 58560 13560 58740
rect 33705 58740 39960 58860
rect 39840 58605 39960 58740
rect 49605 58740 50895 58860
rect 52905 58740 58395 58860
rect 59205 58740 63195 58860
rect 73905 58740 75195 58860
rect 78405 58740 78795 58860
rect 91005 58740 91395 58860
rect 92205 58740 92460 58905
rect 92205 58695 92400 58740
rect 11505 58440 13560 58560
rect 15705 58440 16695 58560
rect 17805 58440 19095 58560
rect 24105 58440 24495 58560
rect 24705 58440 25395 58560
rect 38205 58440 39195 58560
rect 40005 58440 43995 58560
rect 46905 58440 47895 58560
rect 51405 58440 51795 58560
rect 54405 58440 55095 58560
rect 62805 58440 63195 58560
rect 73740 58560 73860 58695
rect 66705 58440 73860 58560
rect 76605 58440 79095 58560
rect 5805 58140 7695 58260
rect 7905 58140 12495 58260
rect 21705 58140 22995 58260
rect 26505 58140 28395 58260
rect 32805 58140 34095 58260
rect 41505 58140 43695 58260
rect 48405 58140 52095 58260
rect 69405 58140 73395 58260
rect 76305 58140 79395 58260
rect 84705 58140 86895 58260
rect 90405 58140 91095 58260
rect 13605 57840 17295 57960
rect 19305 57840 22695 57960
rect 24705 57840 25395 57960
rect 26205 57840 27795 57960
rect 28905 57840 30195 57960
rect 38505 57840 39195 57960
rect 40605 57840 41895 57960
rect 42105 57840 45495 57960
rect 46305 57840 46995 57960
rect 48105 57840 53160 57960
rect 1005 57540 3795 57660
rect 4005 57540 6195 57660
rect 9105 57540 9495 57660
rect 9705 57540 12195 57660
rect 33405 57540 33795 57660
rect 37305 57540 37695 57660
rect 40905 57540 41895 57660
rect 4605 57240 5295 57360
rect 8805 57240 9060 57360
rect 1005 56625 1395 56745
rect 2940 56760 3060 57195
rect 8940 56805 9060 57240
rect 10800 57360 10995 57405
rect 10740 57195 10995 57360
rect 12840 57240 13695 57360
rect 2940 56640 3795 56760
rect 6105 56640 7695 56760
rect 7905 56625 8295 56745
rect 8940 56640 9195 56805
rect 9000 56595 9195 56640
rect 9840 56760 9960 57195
rect 10740 56790 10860 57195
rect 12840 56805 12960 57240
rect 14505 57240 16395 57360
rect 17205 57240 19560 57360
rect 9840 56640 10095 56760
rect 11505 56625 11895 56745
rect 13605 56625 13995 56745
rect 14205 56640 15795 56760
rect 19440 56790 19560 57240
rect 19740 56805 19860 57210
rect 22605 57240 23295 57360
rect 23640 57240 24495 57360
rect 23640 57060 23760 57240
rect 25305 57360 25500 57405
rect 25305 57195 25560 57360
rect 20505 56940 23760 57060
rect 18405 56625 18795 56745
rect 19740 56640 19995 56805
rect 19800 56595 19995 56640
rect 21705 56625 22695 56745
rect 23805 56625 25095 56745
rect 10695 56460 10905 56580
rect 5805 56340 10905 56460
rect 16905 56340 17595 56460
rect 25440 56475 25560 57195
rect 25740 57060 25860 57495
rect 42105 57540 43395 57660
rect 45105 57540 45795 57660
rect 49905 57540 52395 57660
rect 26595 57060 26805 57195
rect 25740 56940 26160 57060
rect 26595 57000 27060 57060
rect 26640 56940 27060 57000
rect 26040 56760 26160 56940
rect 26040 56640 26595 56760
rect 26940 56760 27060 56940
rect 26940 56640 27495 56760
rect 28440 56760 28560 57195
rect 29205 57255 29595 57375
rect 29805 57240 32895 57360
rect 35505 57240 36660 57360
rect 33495 57060 33705 57195
rect 33240 57000 33705 57060
rect 33240 56940 33660 57000
rect 33240 56790 33360 56940
rect 35025 56805 35145 57195
rect 28440 56640 29895 56760
rect 30105 56625 32880 56745
rect 34305 56640 34680 56760
rect 25740 56460 25860 56580
rect 36540 56505 36660 57240
rect 39105 57240 39495 57360
rect 36840 56760 36960 57195
rect 40440 56805 40560 57195
rect 36840 56640 37395 56760
rect 42105 56625 42495 56745
rect 42840 56505 42960 57210
rect 44505 57240 46395 57360
rect 48195 57060 48405 57195
rect 43740 57000 48405 57060
rect 50640 57240 51495 57360
rect 43740 56940 48360 57000
rect 43740 56505 43860 56940
rect 50640 56805 50760 57240
rect 53040 57360 53160 57840
rect 58305 57840 61095 57960
rect 75405 57840 78495 57960
rect 81405 57840 82095 57960
rect 83205 57840 83895 57960
rect 86805 57840 87495 57960
rect 88605 57840 88995 57960
rect 55005 57540 55995 57660
rect 79305 57540 82395 57660
rect 84240 57540 84795 57660
rect 52905 57240 53160 57360
rect 55305 57240 56280 57360
rect 58440 57240 58995 57360
rect 44205 56625 44595 56745
rect 45405 56640 47595 56760
rect 49905 56640 50280 56760
rect 51405 56595 51795 56715
rect 56640 56760 56760 57195
rect 52605 56640 56760 56760
rect 57240 56760 57360 57195
rect 57840 56805 57960 57195
rect 58440 56805 58560 57240
rect 61695 57405 61905 57495
rect 60405 57285 62295 57405
rect 61740 57240 61860 57285
rect 66405 57255 67395 57375
rect 63795 57060 64005 57195
rect 57105 56640 57360 56760
rect 59895 56760 60105 56895
rect 59505 56700 60105 56760
rect 62940 57000 64005 57060
rect 62940 56940 63960 57000
rect 59505 56640 60060 56700
rect 62940 56505 63060 56940
rect 68340 56760 68460 57195
rect 76440 57060 76560 57210
rect 80805 57240 81660 57360
rect 75540 56940 76560 57060
rect 81540 57060 81660 57240
rect 82005 57255 82695 57375
rect 81540 57000 83760 57060
rect 81540 56940 83805 57000
rect 63405 56595 64095 56715
rect 68340 56640 68595 56760
rect 70905 56625 73395 56745
rect 75540 56760 75660 56940
rect 83595 56805 83805 56940
rect 74205 56640 75660 56760
rect 76005 56640 78795 56760
rect 84240 56790 84360 57540
rect 85905 57540 87795 57660
rect 90705 57540 91395 57660
rect 86205 57240 86760 57360
rect 86640 56505 86760 57240
rect 86940 57240 88395 57360
rect 86940 56790 87060 57240
rect 89505 57240 89895 57360
rect 90840 56805 90960 57195
rect 25740 56340 28695 56460
rect 30705 56340 31395 56460
rect 31605 56340 32295 56460
rect 33405 56340 35595 56460
rect 36540 56340 36795 56505
rect 36600 56295 36795 56340
rect 38505 56340 39795 56460
rect 43605 56340 43860 56505
rect 43605 56295 43800 56340
rect 46605 56340 48195 56460
rect 52305 56340 54795 56460
rect 62940 56490 63300 56505
rect 62940 56340 63195 56490
rect 63000 56295 63195 56340
rect 66105 56340 66795 56460
rect 74205 56340 79695 56460
rect 2805 56040 4695 56160
rect 4905 56040 12495 56160
rect 12705 56040 20295 56160
rect 21105 56040 22995 56160
rect 25305 56040 26295 56160
rect 27105 56040 27495 56160
rect 34605 56040 34995 56160
rect 36105 56040 38595 56160
rect 47805 56040 49695 56160
rect 53805 56040 56295 56160
rect 67605 56040 69795 56160
rect 75405 56040 76995 56160
rect 79305 56040 80295 56160
rect 81405 56040 82695 56160
rect 82905 56040 84795 56160
rect 88005 56040 88695 56160
rect 9105 55740 10095 55860
rect 10305 55740 13395 55860
rect 15705 55740 17295 55860
rect 26805 55740 31380 55860
rect 31905 55740 34695 55860
rect 61605 55740 63495 55860
rect 66405 55740 66795 55860
rect 68505 55740 69495 55860
rect 77505 55740 82095 55860
rect 24405 55440 26895 55560
rect 27705 55440 29295 55560
rect 29505 55440 30360 55560
rect 15105 55140 22995 55260
rect 23205 55140 27195 55260
rect 30240 55260 30360 55440
rect 32205 55440 34995 55560
rect 38205 55440 41895 55560
rect 45105 55440 47895 55560
rect 55605 55440 60195 55560
rect 70005 55440 76095 55560
rect 30240 55140 36195 55260
rect 36405 55140 43395 55260
rect 45705 55140 50295 55260
rect 58605 55140 60795 55260
rect 75705 55140 77295 55260
rect 90405 55140 91695 55260
rect 10605 54840 13095 54960
rect 25005 54840 25695 54960
rect 28305 54840 32160 54960
rect 19005 54540 24660 54660
rect 405 54240 4995 54360
rect 5205 54240 6495 54360
rect 24540 54360 24660 54540
rect 25005 54540 29595 54660
rect 32040 54660 32160 54840
rect 32505 54840 36495 54960
rect 43905 54840 49095 54960
rect 49905 54840 53460 54960
rect 32040 54540 35280 54660
rect 35805 54540 39495 54660
rect 41205 54540 45795 54660
rect 47805 54540 48795 54660
rect 53340 54660 53460 54840
rect 62505 54840 65295 54960
rect 65505 54840 75195 54960
rect 79005 54840 83895 54960
rect 88305 54840 91395 54960
rect 53340 54540 58395 54660
rect 65205 54540 67395 54660
rect 68205 54540 71595 54660
rect 90705 54540 91695 54660
rect 24540 54240 25995 54360
rect 29505 54240 37095 54360
rect 43305 54240 49995 54360
rect 50805 54240 52395 54360
rect 53205 54240 54195 54360
rect 54405 54240 63795 54360
rect 75405 54240 78195 54360
rect 78405 54240 78795 54360
rect 86205 54240 87795 54360
rect 3105 53940 11295 54060
rect 14505 53940 16095 54060
rect 17805 53940 18495 54060
rect 23505 53940 24195 54060
rect 26505 53940 28395 54060
rect 36705 53940 37395 54060
rect 40005 53940 47580 54060
rect 48105 53940 48495 54060
rect 55005 53940 67695 54060
rect 69705 53940 71895 54060
rect 73605 53940 79095 54060
rect 83505 53940 85695 54060
rect 89205 53940 91395 54060
rect 4305 53640 5295 53760
rect 20805 53640 23295 53760
rect 26205 53640 28695 53760
rect 33105 53640 34095 53760
rect 34305 53640 35595 53760
rect 43005 53640 45195 53760
rect 62805 53640 65595 53760
rect 83805 53640 86895 53760
rect 9240 53340 10095 53460
rect 9240 53205 9360 53340
rect 11805 53340 14295 53460
rect 15405 53340 16695 53460
rect 18105 53340 18795 53460
rect 19605 53340 19995 53460
rect 20205 53340 23595 53460
rect 26340 53340 27795 53460
rect 8205 53040 9195 53160
rect 26340 53160 26460 53340
rect 46305 53340 47295 53460
rect 48405 53340 53595 53460
rect 67305 53340 67995 53460
rect 70605 53340 73395 53460
rect 76905 53340 79395 53460
rect 88605 53340 91095 53460
rect 25905 53040 26460 53160
rect 38805 53040 41295 53160
rect 41505 53040 43095 53160
rect 55605 53040 55995 53160
rect 58305 53040 61095 53160
rect 77805 53040 79395 53160
rect 79605 53040 81495 53160
rect 81705 53040 83295 53160
rect 90300 53160 90495 53205
rect 90240 52995 90495 53160
rect 2205 52740 3495 52860
rect 6705 52755 7395 52875
rect 8040 52740 9495 52860
rect 8040 52560 8160 52740
rect 12705 52755 13695 52875
rect 7740 52440 8160 52560
rect 1005 52110 1095 52230
rect 1305 52110 1395 52230
rect 5505 52140 6495 52260
rect 7740 52290 7860 52440
rect 10140 52305 10260 52695
rect 11040 52560 11160 52710
rect 19005 52740 20895 52860
rect 23805 52740 25095 52860
rect 11040 52440 13260 52560
rect 13140 52305 13260 52440
rect 12105 52140 12495 52260
rect 13140 52140 13395 52305
rect 13200 52095 13395 52140
rect 14940 52260 15060 52695
rect 14205 52140 15060 52260
rect 21540 52305 21660 52710
rect 23340 52440 25995 52560
rect 21540 52140 21795 52305
rect 21600 52095 21795 52140
rect 23340 52290 23460 52440
rect 26640 52260 26760 52710
rect 30705 52740 33495 52860
rect 35505 52740 36060 52860
rect 28395 52560 28605 52695
rect 28395 52500 29760 52560
rect 28440 52440 29760 52500
rect 25005 52140 26760 52260
rect 27705 52140 29295 52260
rect 29640 52260 29760 52440
rect 34440 52305 34560 52695
rect 29640 52140 31995 52260
rect 35940 52290 36060 52740
rect 44505 52755 44895 52875
rect 36195 52560 36405 52695
rect 36195 52500 37260 52560
rect 36240 52440 37305 52500
rect 37095 52305 37305 52440
rect 38340 52260 38460 52695
rect 38805 52440 42495 52560
rect 42795 52560 43005 52695
rect 42795 52500 43560 52560
rect 42840 52440 43560 52500
rect 38340 52140 38895 52260
rect 43440 52290 43560 52440
rect 46740 52260 46860 52710
rect 47295 52560 47505 52695
rect 47295 52500 47760 52560
rect 47340 52440 47805 52500
rect 47595 52305 47805 52440
rect 46740 52140 47280 52260
rect 47940 52005 48060 52710
rect 51705 52755 52395 52875
rect 53205 52740 54495 52860
rect 56505 52740 56895 52860
rect 48840 52305 48960 52695
rect 50040 52560 50160 52710
rect 49440 52500 50160 52560
rect 49395 52440 50160 52500
rect 49395 52305 49605 52440
rect 50640 52005 50760 52710
rect 63705 52740 65595 52860
rect 65805 52740 67395 52860
rect 71505 52740 74895 52860
rect 78105 52740 78960 52860
rect 58995 52560 59205 52695
rect 51840 52440 59460 52560
rect 51840 52260 51960 52440
rect 51105 52140 51960 52260
rect 52305 52125 53595 52245
rect 55005 52125 55395 52245
rect 55605 52140 56595 52260
rect 59340 52260 59460 52440
rect 60405 52440 65460 52560
rect 65340 52260 65460 52440
rect 65340 52140 65895 52260
rect 68340 52260 68460 52695
rect 67305 52140 68460 52260
rect 70140 52260 70260 52695
rect 75495 52560 75705 52695
rect 75495 52500 75960 52560
rect 75540 52440 75960 52500
rect 70140 52140 75180 52260
rect 75840 52260 75960 52440
rect 77340 52305 77460 52695
rect 78840 52305 78960 52740
rect 83205 52740 83760 52860
rect 80895 52560 81105 52695
rect 80895 52500 83160 52560
rect 80940 52440 83205 52500
rect 82995 52305 83205 52440
rect 79605 52125 80595 52245
rect 83640 52290 83760 52740
rect 86805 52740 87195 52860
rect 85440 52305 85560 52695
rect 2505 51840 3495 51960
rect 3705 51840 9795 51960
rect 13005 51840 14595 51960
rect 14805 51840 15495 51960
rect 25905 51840 26595 51960
rect 31005 51840 31695 51960
rect 37905 51840 44595 51960
rect 49305 51840 49695 51960
rect 60705 51840 61095 51960
rect 66405 51840 67995 51960
rect 69705 51840 70395 51960
rect 82605 51840 83895 51960
rect 705 51540 8895 51660
rect 13305 51540 13695 51660
rect 16605 51540 19095 51660
rect 19305 51540 21195 51660
rect 22005 51540 24795 51660
rect 26205 51540 26895 51660
rect 27705 51540 28095 51660
rect 32205 51540 33795 51660
rect 34005 51540 38595 51660
rect 42405 51540 44895 51660
rect 47505 51540 48195 51660
rect 53805 51540 55995 51660
rect 66705 51540 71895 51660
rect 81405 51540 84795 51660
rect 86040 51660 86160 52710
rect 89505 52740 89895 52860
rect 88140 52305 88260 52695
rect 90240 52560 90360 52995
rect 89640 52440 90360 52560
rect 91140 52740 91695 52860
rect 86505 52125 86895 52245
rect 89640 52260 89760 52440
rect 91140 52290 91260 52740
rect 89040 52200 89760 52260
rect 88995 52140 89760 52200
rect 88995 52005 89205 52140
rect 86040 51540 88695 51660
rect 9705 51240 10380 51360
rect 10905 51240 13395 51360
rect 29205 51240 30495 51360
rect 34305 51240 39495 51360
rect 41805 51240 46995 51360
rect 49005 51240 51495 51360
rect 57705 51240 60795 51360
rect 79305 51240 80895 51360
rect 82005 51240 85695 51360
rect 86805 51240 87495 51360
rect 1905 50940 11295 51060
rect 13005 50940 15195 51060
rect 17505 50940 20595 51060
rect 22305 50940 30195 51060
rect 31305 50940 33195 51060
rect 34005 50940 37695 51060
rect 44205 50940 46695 51060
rect 46905 50940 47895 51060
rect 48105 50940 52095 51060
rect 58905 50940 66195 51060
rect 67905 50940 72195 51060
rect 76305 50940 76995 51060
rect 79005 50940 81495 51060
rect 82905 50940 83295 51060
rect 23205 50640 24195 50760
rect 28605 50640 29895 50760
rect 34905 50640 35580 50760
rect 36105 50640 36495 50760
rect 38505 50640 40995 50760
rect 43605 50640 45195 50760
rect 49005 50640 49395 50760
rect 63405 50640 68595 50760
rect 79005 50640 79995 50760
rect 80205 50640 81795 50760
rect 85905 50640 86295 50760
rect 88005 50640 90195 50760
rect 5805 50340 7995 50460
rect 11505 50340 14895 50460
rect 15705 50340 16695 50460
rect 17505 50340 18495 50460
rect 18705 50340 28095 50460
rect 30405 50340 33795 50460
rect 37005 50340 37995 50460
rect 40905 50340 41595 50460
rect 42705 50340 49260 50460
rect 6405 50040 7095 50160
rect 9405 50040 10695 50160
rect 19005 50040 23295 50160
rect 24405 50040 26295 50160
rect 30405 50040 32895 50160
rect 33105 50040 34095 50160
rect 35205 50040 37395 50160
rect 38505 50040 38895 50160
rect 39105 50040 40095 50160
rect 43905 50040 44595 50160
rect 44805 50040 46095 50160
rect 47205 50040 48195 50160
rect 49140 50160 49260 50340
rect 58140 50340 59895 50460
rect 58140 50205 58260 50340
rect 71805 50340 73395 50460
rect 75705 50340 76995 50460
rect 83805 50340 84495 50460
rect 49140 50040 50895 50160
rect 57105 50040 58095 50160
rect 66405 50040 67095 50160
rect 67305 50040 70995 50160
rect 78405 50040 79695 50160
rect 84405 50040 85695 50160
rect 87705 50040 88095 50160
rect 91005 50040 91695 50160
rect 3105 49740 3495 49860
rect 16905 49740 17295 49860
rect 25005 49740 25695 49860
rect 27105 49740 28560 49860
rect 705 49440 1095 49560
rect 1440 49440 2295 49560
rect 1440 48990 1560 49440
rect 4305 49440 5595 49560
rect 8805 49440 10695 49560
rect 10905 49440 11460 49560
rect 5340 49140 6795 49260
rect 5340 48990 5460 49140
rect 11340 49260 11460 49440
rect 11805 49455 12195 49575
rect 13605 49440 15360 49560
rect 11340 49140 11760 49260
rect 4605 48840 5295 48960
rect 6105 48840 8295 48960
rect 9405 48825 10395 48945
rect 11640 48960 11760 49140
rect 11640 48840 13095 48960
rect 13305 48840 14595 48960
rect 15240 48960 15360 49440
rect 19605 49440 20295 49560
rect 20640 49440 21495 49560
rect 17595 49260 17805 49395
rect 20640 49260 20760 49440
rect 17595 49200 18360 49260
rect 17640 49140 18405 49200
rect 18195 49005 18405 49140
rect 15240 48840 16995 48960
rect 19740 49140 20760 49260
rect 22140 49260 22260 49410
rect 22905 49440 24795 49560
rect 28440 49560 28560 49740
rect 31005 49860 31200 49905
rect 31005 49695 31260 49860
rect 32505 49740 33660 49860
rect 28440 49440 28695 49560
rect 29505 49455 30195 49575
rect 22140 49140 24060 49260
rect 19740 48990 19860 49140
rect 22605 48840 23595 48960
rect 23940 48960 24060 49140
rect 26640 49005 26760 49395
rect 27540 49005 27660 49395
rect 31140 49005 31260 49695
rect 32205 49440 32760 49560
rect 32640 49005 32760 49440
rect 33540 49005 33660 49740
rect 41505 49740 42195 49860
rect 46605 49740 47895 49860
rect 51705 49740 52395 49860
rect 52605 49740 53295 49860
rect 54405 49740 55395 49860
rect 56205 49740 58995 49860
rect 61605 49740 62595 49860
rect 65805 49740 66795 49860
rect 67005 49740 68295 49860
rect 69405 49740 72495 49860
rect 73305 49740 73695 49860
rect 82605 49860 82800 49905
rect 82605 49710 82860 49860
rect 82500 49695 82860 49710
rect 86505 49740 88395 49860
rect 90705 49860 90900 49905
rect 90705 49695 90960 49860
rect 35805 49440 36495 49560
rect 39105 49440 40260 49560
rect 37140 49005 37260 49395
rect 38295 49260 38505 49395
rect 38295 49200 38760 49260
rect 38340 49140 38760 49200
rect 23940 48840 25095 48960
rect 28605 48840 29895 48960
rect 38640 48990 38760 49140
rect 40140 49005 40260 49440
rect 40440 48960 40560 49695
rect 41205 49440 42060 49560
rect 41940 49260 42060 49440
rect 43095 49560 43305 49695
rect 42705 49500 43305 49560
rect 42705 49440 43260 49500
rect 44805 49440 47160 49560
rect 41940 49140 42360 49260
rect 40440 48840 40995 48960
rect 42240 48990 42360 49140
rect 47040 48990 47160 49440
rect 49605 49440 51195 49560
rect 43005 48840 44295 48960
rect 48405 48825 49095 48945
rect 19695 48705 19905 48780
rect 10905 48540 12495 48660
rect 19605 48495 19905 48705
rect 30405 48540 30795 48660
rect 32205 48540 32895 48660
rect 38805 48540 39195 48660
rect 42795 48660 43005 48780
rect 49440 48705 49560 49410
rect 52305 49440 55260 49560
rect 51705 48825 52395 48945
rect 53805 48840 54195 48960
rect 55140 48990 55260 49440
rect 56040 49440 57495 49560
rect 41805 48540 43005 48660
rect 43605 48540 48495 48660
rect 56040 48660 56160 49440
rect 60705 49440 62295 49560
rect 63105 49440 63480 49560
rect 64005 49455 64395 49575
rect 67305 49440 67560 49560
rect 65340 49005 65460 49395
rect 56805 48825 57795 48945
rect 58605 48825 58995 48945
rect 59205 48840 60195 48960
rect 61905 48825 62595 48945
rect 64005 48840 64695 48960
rect 67440 48960 67560 49440
rect 67440 48840 68295 48960
rect 55005 48540 56160 48660
rect 57795 48660 58005 48780
rect 57795 48540 59595 48660
rect 65205 48540 65895 48660
rect 68640 48660 68760 49410
rect 72405 49440 74595 49560
rect 75705 49440 77295 49560
rect 77640 49440 79695 49560
rect 77640 49260 77760 49440
rect 81705 49440 82395 49560
rect 74640 49140 77760 49260
rect 69105 48840 71295 48960
rect 71505 48840 73995 48960
rect 74640 48705 74760 49140
rect 82740 48990 82860 49695
rect 85005 49455 85995 49575
rect 83640 49005 83760 49395
rect 86940 49005 87060 49395
rect 75405 48840 80295 48960
rect 80505 48840 82095 48960
rect 89040 48705 89160 49695
rect 89340 49005 89460 49695
rect 90240 49005 90360 49395
rect 90840 48705 90960 49695
rect 66705 48540 68760 48660
rect 85605 48540 86595 48660
rect 87405 48540 88095 48660
rect 90705 48660 90960 48705
rect 90705 48540 91395 48660
rect 90705 48495 90900 48540
rect 2205 48240 2895 48360
rect 3105 48240 3795 48360
rect 9105 48240 14160 48360
rect 12705 47940 13695 48060
rect 14040 48060 14160 48240
rect 16005 48240 17895 48360
rect 25905 48240 31095 48360
rect 36105 48240 36495 48360
rect 40905 48240 43095 48360
rect 44205 48240 45195 48360
rect 45405 48240 46395 48360
rect 52905 48240 57495 48360
rect 60105 48240 61695 48360
rect 62505 48240 65595 48360
rect 68505 48240 69495 48360
rect 70605 48240 71595 48360
rect 75105 48240 75495 48360
rect 78705 48240 79095 48360
rect 80805 48240 84495 48360
rect 88605 48240 89895 48360
rect 14040 47940 18795 48060
rect 22605 47940 24795 48060
rect 26205 47940 26895 48060
rect 27105 47940 30795 48060
rect 31905 47940 33495 48060
rect 34305 47940 34695 48060
rect 40605 47940 42795 48060
rect 45705 47940 49095 48060
rect 50805 47940 51495 48060
rect 70305 47940 71295 48060
rect 77205 47940 83895 48060
rect 88905 47940 91695 48060
rect 7305 47640 10695 47760
rect 25305 47640 32595 47760
rect 34905 47640 35295 47760
rect 37905 47640 43395 47760
rect 47205 47640 48795 47760
rect 57705 47640 61095 47760
rect 63405 47640 73095 47760
rect 74505 47640 77895 47760
rect 79905 47640 80895 47760
rect 81705 47640 83295 47760
rect 85005 47640 86895 47760
rect 87105 47640 88095 47760
rect 4905 47340 6495 47460
rect 6705 47340 11595 47460
rect 11805 47340 20295 47460
rect 30405 47340 32295 47460
rect 32505 47340 33795 47460
rect 39105 47340 41595 47460
rect 41805 47340 42195 47460
rect 44205 47340 49695 47460
rect 49905 47340 50895 47460
rect 61905 47340 73395 47460
rect 74205 47340 76395 47460
rect 80205 47340 86295 47460
rect 90105 47340 91095 47460
rect 91305 47340 91695 47460
rect 21405 47040 24495 47160
rect 25605 47040 27795 47160
rect 28005 47040 35595 47160
rect 37005 47040 45495 47160
rect 46305 47040 57495 47160
rect 65505 47040 67695 47160
rect 80505 47040 83595 47160
rect 2805 46740 5895 46860
rect 14505 46740 15195 46860
rect 22005 46740 25695 46860
rect 29505 46740 33195 46860
rect 38805 46740 39495 46860
rect 40305 46740 42495 46860
rect 43305 46740 45795 46860
rect 49005 46740 55695 46860
rect 61005 46740 66195 46860
rect 67605 46740 71895 46860
rect 73905 46740 75795 46860
rect 88005 46740 88395 46860
rect 25305 46440 27660 46560
rect 12105 46140 15195 46260
rect 24405 46140 26295 46260
rect 27540 46260 27660 46440
rect 28005 46440 28695 46560
rect 32205 46440 34695 46560
rect 36405 46440 37095 46560
rect 41505 46440 46995 46560
rect 47805 46440 53895 46560
rect 57105 46440 60195 46560
rect 60405 46440 63195 46560
rect 73005 46440 76095 46560
rect 76905 46440 83295 46560
rect 86505 46440 88395 46560
rect 27540 46140 32895 46260
rect 42705 46140 44895 46260
rect 57405 46140 61995 46260
rect 64905 46140 69795 46260
rect 70005 46140 74595 46260
rect 77505 46140 81195 46260
rect 81405 46140 83595 46260
rect 7605 45840 11295 45960
rect 20805 45840 25080 45960
rect 25605 45840 26595 45960
rect 31305 45840 34095 45960
rect 36105 45840 39495 45960
rect 43905 45840 45495 45960
rect 48705 45840 52995 45960
rect 60105 45840 62595 45960
rect 64605 45840 65895 45960
rect 76005 45840 82695 45960
rect 83505 45840 86895 45960
rect 89205 45840 90495 45960
rect 92205 45960 92400 46005
rect 92205 45795 92460 45960
rect 11340 45660 11460 45795
rect 11340 45540 13695 45660
rect 20040 45540 24195 45660
rect 5505 45240 8895 45360
rect 9105 45240 10695 45360
rect 20040 45360 20160 45540
rect 28605 45540 28995 45660
rect 29205 45540 29895 45660
rect 30705 45540 32595 45660
rect 32805 45540 34395 45660
rect 37305 45540 40395 45660
rect 43605 45540 47580 45660
rect 48105 45540 51795 45660
rect 58305 45540 61995 45660
rect 63705 45540 64095 45660
rect 69705 45540 73095 45660
rect 74805 45540 75195 45660
rect 81105 45540 81795 45660
rect 88305 45540 90795 45660
rect 16605 45240 20160 45360
rect 26115 45240 27195 45360
rect 34500 45360 34695 45405
rect 34440 45195 34695 45360
rect 44805 45240 46605 45360
rect 2205 44955 2595 45075
rect 3405 44955 4095 45075
rect 7905 44955 8295 45075
rect 9300 45060 9495 45105
rect 9240 44895 9495 45060
rect 10305 44940 11880 45060
rect 12405 44955 13095 45075
rect 14100 45060 14295 45105
rect 14040 44895 14295 45060
rect 17805 44940 19695 45060
rect 21240 44940 21795 45060
rect 9240 44760 9360 44895
rect 8640 44640 9360 44760
rect 705 44325 1095 44445
rect 1905 44340 4395 44460
rect 4605 44340 6195 44460
rect 7005 44340 7395 44460
rect 8640 44490 8760 44640
rect 14040 44490 14160 44895
rect 15705 44340 16395 44460
rect 9705 44040 12195 44160
rect 13995 44160 14205 44280
rect 13005 44040 14205 44160
rect 17040 44160 17160 44910
rect 21240 44760 21360 44940
rect 22605 44940 22860 45060
rect 20340 44640 21360 44760
rect 20340 44460 20460 44640
rect 22740 44505 22860 44940
rect 25395 44760 25605 44895
rect 25140 44700 25605 44760
rect 28440 44940 28995 45060
rect 25140 44640 25560 44700
rect 18105 44340 20460 44460
rect 20805 44340 21495 44460
rect 25140 44460 25260 44640
rect 23805 44340 25260 44460
rect 28440 44460 28560 44940
rect 31500 45060 31695 45105
rect 31440 44895 31695 45060
rect 34440 45060 34560 45195
rect 33840 44940 34560 45060
rect 25605 44340 28560 44460
rect 30240 44460 30360 44895
rect 31440 44505 31560 44895
rect 33540 44760 33660 44910
rect 32040 44700 33660 44760
rect 31995 44640 33660 44700
rect 31995 44505 32205 44640
rect 28905 44340 31080 44460
rect 33840 44460 33960 44940
rect 39795 45060 40005 45195
rect 46395 45120 46605 45240
rect 49905 45240 50295 45360
rect 66405 45240 66960 45360
rect 38640 45000 40005 45060
rect 38640 44940 39960 45000
rect 35040 44760 35160 44910
rect 38640 44760 38760 44940
rect 40995 44760 41205 44895
rect 34740 44640 35160 44760
rect 35640 44700 38760 44760
rect 35595 44640 38760 44700
rect 39240 44700 41205 44760
rect 39240 44640 41160 44700
rect 33240 44340 33960 44460
rect 33240 44205 33360 44340
rect 34740 44460 34860 44640
rect 34305 44340 34860 44460
rect 35595 44505 35805 44640
rect 39240 44460 39360 44640
rect 37905 44340 39360 44460
rect 39540 44340 40395 44460
rect 39540 44205 39660 44340
rect 41640 44460 41760 44910
rect 42405 44940 42960 45060
rect 42840 44760 42960 44940
rect 43740 44940 44895 45060
rect 42840 44700 43260 44760
rect 42840 44640 43305 44700
rect 43095 44505 43305 44640
rect 41640 44340 42495 44460
rect 43740 44490 43860 44940
rect 46605 44940 47160 45060
rect 47040 44760 47160 44940
rect 47505 44955 47895 45075
rect 48705 44940 50595 45060
rect 52605 44940 55395 45060
rect 55605 44955 57195 45075
rect 59205 44985 59595 45105
rect 63705 44940 65295 45060
rect 60540 44760 60660 44910
rect 47040 44640 48360 44760
rect 48240 44490 48360 44640
rect 59640 44640 60660 44760
rect 45705 44325 46095 44445
rect 49005 44340 49395 44460
rect 52005 44325 52695 44445
rect 54105 44325 54495 44445
rect 59640 44460 59760 44640
rect 61140 44505 61260 44910
rect 62205 44640 62760 44760
rect 56505 44340 59760 44460
rect 60105 44340 60795 44460
rect 61140 44340 61395 44505
rect 61200 44295 61395 44340
rect 62640 44460 62760 44640
rect 62640 44340 63195 44460
rect 63540 44460 63660 44910
rect 65940 44505 66060 44910
rect 63540 44340 64095 44460
rect 65940 44340 66195 44505
rect 66000 44295 66195 44340
rect 16605 44040 17160 44160
rect 23505 44040 24495 44160
rect 25905 44040 27195 44160
rect 29505 44040 30495 44160
rect 33105 44040 33360 44205
rect 33105 43995 33300 44040
rect 35505 44040 35895 44160
rect 36105 44040 36795 44160
rect 39405 44040 39660 44205
rect 39405 43995 39600 44040
rect 47505 44040 48495 44160
rect 53805 44040 62295 44160
rect 66540 44160 66660 44895
rect 66840 44460 66960 45240
rect 73605 45240 76695 45360
rect 78105 45240 79095 45360
rect 88500 45360 88695 45405
rect 88440 45195 88695 45360
rect 91605 45240 91995 45360
rect 68640 44505 68760 44940
rect 73305 44940 74295 45060
rect 74505 44940 74880 45060
rect 75405 44940 76860 45060
rect 69840 44505 69960 44895
rect 68505 44340 68760 44505
rect 68505 44295 68700 44340
rect 71940 44460 72060 44895
rect 76740 44760 76860 44940
rect 77205 44955 79695 45075
rect 82305 44940 82995 45060
rect 84405 44940 85395 45060
rect 80595 44760 80805 44895
rect 76740 44640 80460 44760
rect 80595 44700 81360 44760
rect 80640 44640 81405 44700
rect 80340 44490 80460 44640
rect 81195 44505 81405 44640
rect 86640 44505 86760 44895
rect 87540 44505 87660 44895
rect 70605 44340 72060 44460
rect 73605 44325 78495 44445
rect 83505 44400 84060 44460
rect 83505 44340 84105 44400
rect 83895 44205 84105 44340
rect 84705 44340 85695 44460
rect 88440 44205 88560 45195
rect 89340 44505 89460 44895
rect 90240 44505 90360 44895
rect 91305 44325 91995 44445
rect 64005 44040 66660 44160
rect 75705 44040 76995 44160
rect 90105 44040 91395 44160
rect 9405 43740 10095 43860
rect 16305 43740 19395 43860
rect 21105 43740 22095 43860
rect 24540 43860 24660 43995
rect 24540 43740 25995 43860
rect 32805 43740 33495 43860
rect 36705 43740 37095 43860
rect 40905 43740 41895 43860
rect 45405 43740 46095 43860
rect 46305 43740 46695 43860
rect 64605 43740 64995 43860
rect 65805 43740 68295 43860
rect 76305 43740 76695 43860
rect 88005 43740 88995 43860
rect 92340 43860 92460 45795
rect 91905 43740 92460 43860
rect 2205 43440 4095 43560
rect 4305 43440 8595 43560
rect 25305 43440 27495 43560
rect 36405 43440 37395 43560
rect 42105 43440 42795 43560
rect 47805 43440 49395 43560
rect 49605 43440 55995 43560
rect 60105 43440 61695 43560
rect 68205 43440 73395 43560
rect 77505 43440 81195 43560
rect 86505 43440 90495 43560
rect 6105 43140 12195 43260
rect 13605 43140 16995 43260
rect 17205 43140 17295 43260
rect 18705 43140 19995 43260
rect 23505 43140 24495 43260
rect 28305 43140 30195 43260
rect 32505 43140 33495 43260
rect 38205 43140 44295 43260
rect 56805 43140 57195 43260
rect 61605 43140 64095 43260
rect 65205 43140 66495 43260
rect 78105 43140 78495 43260
rect 78705 43140 80295 43260
rect 83205 43140 84195 43260
rect 3405 42840 3795 42960
rect 4005 42840 7695 42960
rect 28140 42960 28260 43095
rect 24405 42840 28260 42960
rect 31005 42840 32595 42960
rect 35205 42840 35895 42960
rect 40005 42840 43095 42960
rect 45540 42840 50295 42960
rect 8505 42540 10995 42660
rect 16005 42540 18795 42660
rect 25005 42540 31395 42660
rect 33405 42540 33795 42660
rect 34140 42540 34695 42660
rect 2805 42240 4995 42360
rect 7605 42240 14595 42360
rect 20205 42240 23295 42360
rect 24105 42240 30795 42360
rect 31740 42240 31995 42360
rect 11805 41940 12795 42060
rect 17805 41940 19605 42060
rect 19395 41820 19605 41940
rect 22605 42000 23160 42060
rect 22605 41940 23205 42000
rect 1005 41640 1395 41760
rect 3405 41760 3600 41805
rect 3405 41595 3660 41760
rect 4605 41640 6360 41760
rect 3540 41190 3660 41595
rect 6240 41190 6360 41640
rect 6705 41640 8295 41760
rect 9105 41640 9360 41760
rect 2505 41040 3495 41160
rect 7605 41025 8595 41145
rect 9240 41160 9360 41640
rect 10305 41640 10995 41760
rect 14505 41640 14895 41760
rect 15105 41640 16395 41760
rect 12540 41205 12660 41595
rect 15540 41460 15660 41640
rect 19605 41640 21495 41760
rect 22995 41805 23205 41940
rect 31740 42060 31860 42240
rect 34140 42360 34260 42540
rect 45540 42660 45660 42840
rect 51105 42840 51795 42960
rect 55305 42840 55995 42960
rect 62805 42840 63795 42960
rect 68040 42840 68895 42960
rect 68040 42705 68160 42840
rect 70305 42840 71295 42960
rect 72705 42840 76995 42960
rect 79905 42840 80895 42960
rect 88305 42840 88695 42960
rect 89505 42840 91995 42960
rect 41205 42540 45660 42660
rect 47805 42540 60495 42660
rect 63540 42540 67995 42660
rect 32205 42240 34260 42360
rect 34605 42240 37560 42360
rect 27105 41940 31860 42060
rect 32805 41940 34095 42060
rect 37440 42060 37560 42240
rect 37905 42240 38295 42360
rect 43605 42240 44595 42360
rect 56505 42240 58995 42360
rect 63540 42360 63660 42540
rect 71205 42540 71595 42660
rect 71940 42540 77595 42660
rect 62640 42240 63660 42360
rect 37440 41940 40995 42060
rect 49905 41940 51195 42060
rect 62640 42060 62760 42240
rect 64005 42240 64695 42360
rect 67905 42240 68295 42360
rect 70005 42240 70695 42360
rect 71940 42360 72060 42540
rect 82305 42540 83295 42660
rect 84405 42540 85695 42660
rect 71040 42240 72060 42360
rect 71040 42060 71160 42240
rect 72405 42240 73695 42360
rect 75240 42240 77595 42360
rect 75240 42060 75360 42240
rect 79005 42240 81495 42360
rect 87105 42240 87495 42360
rect 90405 42240 90795 42360
rect 61905 41940 62760 42060
rect 69840 41940 71160 42060
rect 74040 41940 75360 42060
rect 26805 41655 27495 41775
rect 31605 41655 31995 41775
rect 36405 41640 39060 41760
rect 15540 41340 15960 41460
rect 9240 41040 11295 41160
rect 14640 41100 15195 41160
rect 14595 41040 15195 41100
rect 14595 40905 14805 41040
rect 15840 41160 15960 41340
rect 23640 41205 23760 41595
rect 24840 41340 27060 41460
rect 15840 41040 16695 41160
rect 22605 41025 22995 41145
rect 24840 41160 24960 41340
rect 24405 41040 24960 41160
rect 26940 41190 27060 41340
rect 29595 41460 29805 41595
rect 35295 41460 35505 41595
rect 28005 41400 29805 41460
rect 34740 41400 35505 41460
rect 38940 41460 39060 41640
rect 39405 41640 40395 41760
rect 40740 41640 42495 41760
rect 28005 41340 29760 41400
rect 34740 41340 35460 41400
rect 38940 41340 39360 41460
rect 25605 41040 26295 41160
rect 30105 41100 30360 41160
rect 30105 41040 30405 41100
rect 1905 40740 4695 40860
rect 4905 40740 5295 40860
rect 25305 40740 25980 40860
rect 26295 40860 26505 40980
rect 30195 40905 30405 41040
rect 34740 41160 34860 41340
rect 31905 41040 34860 41160
rect 35205 41040 36495 41160
rect 39240 41160 39360 41340
rect 40740 41460 40860 41640
rect 43905 41640 45195 41760
rect 50505 41640 50895 41760
rect 39705 41340 40860 41460
rect 50340 41205 50460 41610
rect 52605 41640 54195 41760
rect 55005 41640 55695 41760
rect 57405 41655 58095 41775
rect 39240 41040 40095 41160
rect 26295 40740 28095 40860
rect 32505 40740 36195 40860
rect 39240 40860 39360 41040
rect 40905 41025 41595 41145
rect 43005 41040 43395 41160
rect 45105 41025 48495 41145
rect 50205 41040 50460 41205
rect 50205 40995 50400 41040
rect 51540 41160 51660 41595
rect 51105 41040 52695 41160
rect 52905 41025 55395 41145
rect 56640 41160 56760 41595
rect 59640 41205 59760 41895
rect 62505 41640 62895 41760
rect 63705 41640 63960 41760
rect 56640 41040 56895 41160
rect 57705 41025 58095 41145
rect 58305 41025 58695 41145
rect 59640 41040 59895 41205
rect 59700 40995 59895 41040
rect 61440 41160 61560 41595
rect 61305 41040 61560 41160
rect 63840 41205 63960 41640
rect 64305 41640 65760 41760
rect 63840 41040 64095 41205
rect 63900 40995 64095 41040
rect 65640 41190 65760 41640
rect 67005 41640 67695 41760
rect 68040 41640 69495 41760
rect 68040 41190 68160 41640
rect 69840 41760 69960 41940
rect 69705 41640 69960 41760
rect 71340 41640 71595 41760
rect 70440 41205 70560 41595
rect 71340 41205 71460 41640
rect 72540 41205 72660 41595
rect 66705 41040 67995 41160
rect 68805 41040 69795 41160
rect 74040 41160 74160 41940
rect 76140 42000 77295 42060
rect 75495 41760 75705 41895
rect 76095 41940 77295 42000
rect 76095 41805 76305 41940
rect 82005 41940 83295 42060
rect 83505 41940 84195 42060
rect 89505 41940 89895 42060
rect 75495 41700 75960 41760
rect 75540 41640 75960 41700
rect 75840 41205 75960 41640
rect 76440 41640 78795 41760
rect 73905 41040 74160 41160
rect 37905 40740 39360 40860
rect 49905 40740 52095 40860
rect 72405 40740 72795 40860
rect 73005 40740 74295 40860
rect 76440 40890 76560 41640
rect 79605 41640 80295 41760
rect 81240 41640 82095 41760
rect 81240 41205 81360 41640
rect 86595 41760 86805 41895
rect 86595 41700 87795 41760
rect 86640 41640 87795 41700
rect 86640 41460 86760 41640
rect 84540 41400 86760 41460
rect 84495 41340 86760 41400
rect 84495 41205 84705 41340
rect 77505 41040 79695 41160
rect 82605 41025 83295 41145
rect 87405 41040 88095 41160
rect 88440 41160 88560 41595
rect 88440 41040 90195 41160
rect 79740 40860 79860 40980
rect 82395 40860 82605 40980
rect 79740 40740 82605 40860
rect 84105 40740 85395 40860
rect 7905 40440 13695 40560
rect 22005 40440 24795 40560
rect 27705 40440 28395 40560
rect 34005 40440 36495 40560
rect 38205 40440 41295 40560
rect 42405 40440 43695 40560
rect 43905 40440 44295 40560
rect 58005 40440 58995 40560
rect 60705 40440 63195 40560
rect 66405 40440 68595 40560
rect 68940 40440 71895 40560
rect 405 40140 2295 40260
rect 4605 40140 4995 40260
rect 15105 40140 16095 40260
rect 16305 40140 17295 40260
rect 17505 40140 21195 40260
rect 30405 40140 36795 40260
rect 37005 40140 37395 40260
rect 38505 40140 39495 40260
rect 44805 40140 49095 40260
rect 54405 40140 56295 40260
rect 68940 40260 69060 40440
rect 78105 40440 80295 40560
rect 64005 40140 69060 40260
rect 70440 40140 72195 40260
rect 10305 39840 26760 39960
rect 3405 39540 24495 39660
rect 26640 39660 26760 39840
rect 28005 39840 28395 39960
rect 32505 39840 38595 39960
rect 38940 39900 40395 39960
rect 38895 39840 40395 39900
rect 38895 39705 39105 39840
rect 42105 39840 43395 39960
rect 44505 39840 46395 39960
rect 58005 39840 59895 39960
rect 70440 39960 70560 40140
rect 73905 40140 74295 40260
rect 60105 39840 70560 39960
rect 84105 39840 84795 39960
rect 85005 39840 90195 39960
rect 90405 39840 91095 39960
rect 26640 39540 34095 39660
rect 34305 39540 35595 39660
rect 40905 39540 49695 39660
rect 50805 39540 54495 39660
rect 55605 39540 66495 39660
rect 70905 39540 74295 39660
rect 82005 39540 87195 39660
rect 10005 39240 10995 39360
rect 12405 39240 19095 39360
rect 30705 39240 33195 39360
rect 38505 39240 40395 39360
rect 62805 39240 66795 39360
rect 69705 39240 76995 39360
rect 77205 39240 78495 39360
rect 88905 39240 90195 39360
rect 1005 38940 7695 39060
rect 13305 38940 19695 39060
rect 25605 38940 27195 39060
rect 28005 38940 28695 39060
rect 31305 38940 34695 39060
rect 36405 38940 42795 39060
rect 46905 38940 49395 39060
rect 50805 38940 53595 39060
rect 56505 38940 69195 39060
rect 74205 38940 76095 39060
rect 88305 38940 91995 39060
rect 405 38640 10695 38760
rect 21105 38640 23295 38760
rect 25005 38640 26895 38760
rect 32205 38640 36195 38760
rect 40605 38640 41895 38760
rect 44205 38640 45795 38760
rect 48405 38640 49695 38760
rect 61305 38640 64995 38760
rect 65205 38640 65895 38760
rect 68205 38640 70395 38760
rect 86505 38640 88695 38760
rect 90105 38640 90795 38760
rect 4305 38340 7095 38460
rect 7305 38340 9495 38460
rect 10905 38340 12495 38460
rect 14805 38340 20595 38460
rect 20805 38340 23595 38460
rect 27405 38340 33495 38460
rect 36705 38340 40095 38460
rect 43005 38340 49995 38460
rect 56805 38340 59295 38460
rect 59505 38340 65895 38460
rect 66105 38340 67395 38460
rect 67605 38340 71295 38460
rect 71505 38340 74895 38460
rect 78405 38340 79995 38460
rect 80805 38340 82995 38460
rect 86640 38340 87495 38460
rect 86640 38205 86760 38340
rect 4005 38040 13395 38160
rect 15705 38040 16695 38160
rect 17805 38040 21360 38160
rect 21240 37905 21360 38040
rect 24105 38040 26295 38160
rect 27705 38040 31995 38160
rect 34605 38040 37695 38160
rect 49305 38040 50295 38160
rect 51405 38040 56295 38160
rect 60405 38040 61395 38160
rect 64905 38040 66795 38160
rect 69405 38040 74595 38160
rect 79005 38040 81495 38160
rect 84540 38040 86595 38160
rect 705 37740 3195 37860
rect 6105 37740 11295 37860
rect 11505 37740 12195 37860
rect 14205 37740 16995 37860
rect 21405 37740 27195 37860
rect 37905 37740 40695 37860
rect 42705 37740 46095 37860
rect 67605 37740 69495 37860
rect 84540 37860 84660 38040
rect 91005 38040 91995 38160
rect 77805 37740 84660 37860
rect 18105 37440 18795 37560
rect 22605 37440 25695 37560
rect 26805 37440 29295 37560
rect 30540 37440 31395 37560
rect 1305 37140 1860 37260
rect 1740 36705 1860 37140
rect 2205 37140 3795 37260
rect 5505 37140 6795 37260
rect 7005 37140 7695 37260
rect 15405 37155 15795 37275
rect 9540 36960 9660 37110
rect 8805 36840 9660 36960
rect 10140 36705 10260 37110
rect 18705 37155 19695 37275
rect 24405 37155 25395 37275
rect 27405 37140 28380 37260
rect 10140 36540 10395 36705
rect 10200 36495 10395 36540
rect 15705 36540 19995 36660
rect 20805 36540 25395 36660
rect 26340 36690 26460 37095
rect 27240 36960 27360 37110
rect 27240 36840 28260 36960
rect 26505 36525 27495 36645
rect 1005 36240 2580 36360
rect 3105 36240 6195 36360
rect 10305 36240 10695 36360
rect 15405 36240 15795 36360
rect 22905 36240 24495 36360
rect 25905 36240 26895 36360
rect 28140 36360 28260 36840
rect 28740 36705 28860 37110
rect 30540 36960 30660 37440
rect 32205 37440 32895 37560
rect 33105 37440 35295 37560
rect 38040 37440 39495 37560
rect 34005 37260 34200 37305
rect 34005 37095 34260 37260
rect 36705 37140 37095 37260
rect 32295 36960 32505 37095
rect 30105 36840 30660 36960
rect 31440 36900 32505 36960
rect 31440 36840 32460 36900
rect 28605 36540 28860 36705
rect 28605 36495 28800 36540
rect 29805 36540 30195 36660
rect 31440 36690 31560 36840
rect 33240 36660 33360 37095
rect 33240 36540 33795 36660
rect 28140 36240 28695 36360
rect 34140 36360 34260 37095
rect 35040 36705 35160 37095
rect 38040 36690 38160 37440
rect 41505 37440 45495 37560
rect 47340 37440 49395 37560
rect 39405 37155 40095 37275
rect 43605 37140 44595 37260
rect 40695 36960 40905 37095
rect 40695 36900 43995 36960
rect 40740 36840 43995 36900
rect 45240 36705 45360 37110
rect 36105 36525 36495 36645
rect 41505 36510 41880 36630
rect 42405 36600 43860 36660
rect 42405 36540 43905 36600
rect 33405 36240 34260 36360
rect 43695 36405 43905 36540
rect 45105 36540 45360 36705
rect 45105 36495 45300 36540
rect 47340 36660 47460 37440
rect 52605 37440 53295 37560
rect 60705 37440 61695 37560
rect 61905 37440 62295 37560
rect 68505 37440 68895 37560
rect 71340 37440 72495 37560
rect 47805 37140 49260 37260
rect 49140 36690 49260 37140
rect 50205 37155 50895 37275
rect 52005 37140 52260 37260
rect 52140 36705 52260 37140
rect 53640 36960 53760 37110
rect 56205 37140 57495 37260
rect 57840 37140 58395 37260
rect 57840 36960 57960 37140
rect 63405 37155 64095 37275
rect 65040 37140 65895 37260
rect 52905 36840 53760 36960
rect 56940 36840 57960 36960
rect 46305 36540 47460 36660
rect 56940 36690 57060 36840
rect 61140 36690 61260 37095
rect 55305 36540 56295 36660
rect 60405 36525 61095 36645
rect 65040 36690 65160 37140
rect 67005 37140 67860 37260
rect 67740 37005 67860 37140
rect 71340 37260 71460 37440
rect 72705 37440 73095 37560
rect 82605 37440 83295 37560
rect 84705 37440 85395 37560
rect 85605 37440 85995 37560
rect 87105 37560 87300 37605
rect 87105 37395 87360 37560
rect 88005 37440 88995 37560
rect 70140 37140 71460 37260
rect 67740 36840 67995 37005
rect 67800 36795 67995 36840
rect 61905 36540 64260 36660
rect 45705 36240 46095 36360
rect 11505 35940 12795 36060
rect 13605 35940 16395 36060
rect 17205 35940 20595 36060
rect 25140 35940 25995 36060
rect 25140 35805 25260 35940
rect 28305 35940 28995 36060
rect 33240 36060 33360 36195
rect 49905 36240 52695 36360
rect 61005 36240 62295 36360
rect 64140 36360 64260 36540
rect 65805 36525 66195 36645
rect 68940 36660 69060 37095
rect 67305 36540 69060 36660
rect 70140 36660 70260 37140
rect 71805 37140 72360 37260
rect 72240 37005 72360 37140
rect 72240 36840 72495 37005
rect 72300 36795 72495 36840
rect 74940 36705 75060 37095
rect 70005 36540 70260 36660
rect 70605 36525 71895 36645
rect 75840 36690 75960 37395
rect 76140 36705 76260 37110
rect 77205 37260 77400 37305
rect 77205 37095 77460 37260
rect 76140 36540 76395 36705
rect 76200 36495 76395 36540
rect 77340 36690 77460 37095
rect 79140 37140 79395 37260
rect 79140 36705 79260 37140
rect 80040 36405 80160 37110
rect 81405 37140 81960 37260
rect 80595 36960 80805 37095
rect 80340 36900 80805 36960
rect 80340 36840 80760 36900
rect 80340 36690 80460 36840
rect 81840 36690 81960 37140
rect 82695 36960 82905 37095
rect 82140 36900 82905 36960
rect 82095 36840 82860 36900
rect 82095 36705 82305 36840
rect 83205 36540 84195 36660
rect 85740 36660 85860 37095
rect 87240 36960 87360 37395
rect 87240 36900 88260 36960
rect 87240 36840 88305 36900
rect 88095 36705 88305 36840
rect 89940 36705 90060 37095
rect 91140 36705 91260 37095
rect 85305 36540 85860 36660
rect 87105 36525 87495 36645
rect 89205 36540 89595 36660
rect 64140 36240 65295 36360
rect 70905 36240 71295 36360
rect 79005 36240 79680 36360
rect 83505 36240 83895 36360
rect 85605 36240 85995 36360
rect 31005 35940 33360 36060
rect 35205 35940 40695 36060
rect 44805 35940 53295 36060
rect 58905 35940 74295 36060
rect 74505 35940 76095 36060
rect 85005 35940 85695 36060
rect 85905 35940 87495 36060
rect 88605 35940 90195 36060
rect 91005 35940 91395 36060
rect 705 35640 1395 35760
rect 4005 35640 4395 35760
rect 7305 35640 7995 35760
rect 8205 35640 9195 35760
rect 9405 35640 10695 35760
rect 10905 35640 16695 35760
rect 17505 35640 18495 35760
rect 24105 35640 25095 35760
rect 26205 35640 27795 35760
rect 29505 35640 34695 35760
rect 37605 35640 42795 35760
rect 43005 35640 46995 35760
rect 59505 35640 60195 35760
rect 65505 35640 69795 35760
rect 73905 35640 76695 35760
rect 79005 35640 90495 35760
rect 11205 35340 11895 35460
rect 12105 35340 16080 35460
rect 16605 35340 22095 35460
rect 23505 35340 29595 35460
rect 30405 35340 31380 35460
rect 31905 35340 37395 35460
rect 37605 35340 38895 35460
rect 40005 35340 42495 35460
rect 44805 35340 46695 35460
rect 63105 35340 64995 35460
rect 74805 35340 79395 35460
rect 82605 35340 89595 35460
rect 91605 35340 91995 35460
rect 1305 35040 1695 35160
rect 3105 35040 4395 35160
rect 4605 35040 5295 35160
rect 6105 35040 8595 35160
rect 8805 35040 13695 35160
rect 13905 35040 14295 35160
rect 20205 35040 20895 35160
rect 22005 35040 24795 35160
rect 25605 35040 27360 35160
rect 27240 34905 27360 35040
rect 28305 35040 28695 35160
rect 28905 35040 35295 35160
rect 40305 35040 54195 35160
rect 55005 35040 55995 35160
rect 61005 35040 64095 35160
rect 67305 35040 67995 35160
rect 70905 35040 72195 35160
rect 75105 35040 75795 35160
rect 76905 35040 78795 35160
rect 80505 35040 82095 35160
rect 84105 35040 84795 35160
rect 14505 34740 15495 34860
rect 17805 34740 19095 34860
rect 19305 34740 21195 34860
rect 21405 34740 25395 34860
rect 27405 34740 31695 34860
rect 37305 34740 38895 34860
rect 42705 34740 44895 34860
rect 45105 34740 45495 34860
rect 45840 34740 50595 34860
rect 1905 34440 3795 34560
rect 5805 34440 6960 34560
rect 6840 34305 6960 34440
rect 12705 34440 17295 34560
rect 18105 34440 21660 34560
rect 21540 34305 21660 34440
rect 25005 34440 26295 34560
rect 27105 34440 30195 34560
rect 33105 34440 36180 34560
rect 36705 34440 40695 34560
rect 45840 34560 45960 34740
rect 50805 34740 52695 34860
rect 57495 34860 57705 34995
rect 57495 34800 61695 34860
rect 57540 34740 61695 34800
rect 62505 34740 62895 34860
rect 63105 34740 64395 34860
rect 72405 34740 76395 34860
rect 76605 34740 77295 34860
rect 77505 34740 79095 34860
rect 79305 34740 83595 34860
rect 88005 34740 88695 34860
rect 89505 34740 90195 34860
rect 91005 34740 91695 34860
rect 42405 34440 45960 34560
rect 53205 34440 58095 34560
rect 4905 34140 5295 34260
rect 7005 34140 7695 34260
rect 10305 34140 11295 34260
rect -360 33840 495 33960
rect 2505 33855 3495 33975
rect 1605 33225 3495 33345
rect 4140 33105 4260 34095
rect 12705 34140 13095 34260
rect 21705 34140 22395 34260
rect 22605 34140 24495 34260
rect 29205 34140 30195 34260
rect 6105 33960 6300 34005
rect 6105 33795 6360 33960
rect 6705 33840 6960 33960
rect 6240 33390 6360 33795
rect 4905 33225 5595 33345
rect 6840 33105 6960 33840
rect 9405 33840 9795 33960
rect 10605 33840 15195 33960
rect 16005 33840 17595 33960
rect 18405 33840 19995 33960
rect 20205 33840 22560 33960
rect 10440 33405 10560 33795
rect 7905 33225 8295 33345
rect 11805 33240 13395 33360
rect 14205 33240 14595 33360
rect 18705 33225 19095 33345
rect 19905 33240 22095 33360
rect 22440 33360 22560 33840
rect 25905 33855 26595 33975
rect 27825 33405 27945 34095
rect 34605 34140 35595 34260
rect 51405 34140 52395 34260
rect 53505 34140 53895 34260
rect 59205 34140 60960 34260
rect 31605 33840 32280 33960
rect 28395 33660 28605 33795
rect 28140 33600 28605 33660
rect 28140 33540 28560 33600
rect 28140 33405 28260 33540
rect 29340 33405 29460 33795
rect 33795 33960 34005 34095
rect 32805 33900 34005 33960
rect 32805 33840 33960 33900
rect 43605 33855 43995 33975
rect 45105 33855 46095 33975
rect 47805 33840 49095 33960
rect 50505 33855 50895 33975
rect 54405 33840 54795 33960
rect 57600 33960 57795 34005
rect 29940 33600 36495 33660
rect 29895 33540 36495 33600
rect 29895 33405 30105 33540
rect 52095 33660 52305 33795
rect 57540 33795 57795 33960
rect 59805 33855 60495 33975
rect 52095 33600 52860 33660
rect 52140 33540 52905 33600
rect 22440 33240 22680 33360
rect 23205 33240 24795 33360
rect 28305 33240 28695 33360
rect 31305 33300 33045 33360
rect 33240 33300 39495 33360
rect 31305 33240 33105 33300
rect 32895 33105 33105 33240
rect -360 32940 1095 33060
rect 4140 32940 4395 33105
rect 4200 32895 4395 32940
rect 6705 32940 6960 33105
rect 6705 32895 6900 32940
rect 20805 32940 21495 33060
rect 26505 32940 26895 33060
rect 33090 33000 33105 33105
rect 33195 33240 39495 33300
rect 33195 33105 33405 33240
rect 40695 33360 40905 33495
rect 52695 33405 52905 33540
rect 40695 33300 41295 33360
rect 40740 33240 41295 33300
rect 43905 33240 44895 33360
rect 57540 33360 57660 33795
rect 60840 33660 60960 34140
rect 61605 34140 63195 34260
rect 63795 34140 73095 34260
rect 63795 34020 64005 34140
rect 74805 34140 75195 34260
rect 76305 34140 78195 34260
rect 90105 34140 90795 34260
rect 63840 33660 63960 33810
rect 65505 33840 66360 33960
rect 64695 33660 64905 33795
rect 58305 33540 60060 33660
rect 60840 33540 63960 33660
rect 64140 33600 64905 33660
rect 66240 33660 66360 33840
rect 66705 33855 68595 33975
rect 69300 33960 69495 34005
rect 69240 33795 69495 33960
rect 71805 33855 72495 33975
rect 81705 33840 82695 33960
rect 82905 33855 83295 33975
rect 66240 33600 67260 33660
rect 64140 33540 64860 33600
rect 66240 33540 67305 33600
rect 59940 33390 60060 33540
rect 58605 33240 59295 33360
rect 63540 33360 63660 33540
rect 64140 33390 64260 33540
rect 67095 33405 67305 33540
rect 62205 33240 63660 33360
rect 69240 33360 69360 33795
rect 75540 33540 76395 33660
rect 75540 33390 75660 33540
rect 80040 33405 80160 33795
rect 78240 33240 79560 33360
rect 35505 32940 38295 33060
rect 41205 32940 41595 33060
rect 46005 32940 47295 33060
rect 49305 32940 52995 33060
rect 53805 32940 61395 33060
rect 78240 33060 78360 33240
rect 77205 32940 78360 33060
rect 79440 33060 79560 33240
rect 83640 33390 83760 34095
rect 84105 33840 84360 33960
rect 80340 33240 81795 33360
rect 80340 33060 80460 33240
rect 84240 33105 84360 33840
rect 86805 33840 87360 33960
rect 87240 33405 87360 33840
rect 88740 33405 88860 33795
rect 90240 33405 90360 33795
rect 79440 32940 80460 33060
rect 84105 32940 84360 33105
rect 84105 32895 84300 32940
rect 3705 32640 4995 32760
rect 9105 32640 10395 32760
rect 11205 32640 12795 32760
rect 16305 32640 17295 32760
rect 17505 32640 19695 32760
rect 25005 32640 25695 32760
rect 28605 32640 34095 32760
rect 35205 32640 39495 32760
rect 47805 32640 48495 32760
rect 54105 32640 58695 32760
rect 59505 32640 60195 32760
rect 73005 32640 75495 32760
rect 79305 32640 80595 32760
rect 82905 32640 85995 32760
rect 11040 32460 11160 32595
rect 7005 32340 11160 32460
rect 16905 32340 17895 32460
rect 19305 32340 20895 32460
rect 24105 32340 25995 32460
rect 30705 32340 33495 32460
rect 34605 32340 35295 32460
rect 36405 32340 39195 32460
rect 44805 32340 48795 32460
rect 55905 32340 58095 32460
rect 59205 32340 65595 32460
rect 69105 32340 71895 32460
rect 81705 32340 84795 32460
rect 3405 32040 11595 32160
rect 21240 32040 22995 32160
rect 2205 31740 2895 31860
rect 4305 31740 8895 31860
rect 21240 31860 21360 32040
rect 24405 32040 25095 32160
rect 29805 32040 34860 32160
rect 19905 31740 21360 31860
rect 21540 31740 24195 31860
rect 21540 31560 21660 31740
rect 28605 31740 33195 31860
rect 34740 31860 34860 32040
rect 36705 32040 44295 32160
rect 56805 32040 57795 32160
rect 69405 32040 72495 32160
rect 34740 31740 36195 31860
rect 36405 31740 37095 31860
rect 37905 31740 49695 31860
rect 58905 31740 61095 31860
rect 67005 31740 67395 31860
rect 81405 31740 86595 31860
rect 705 31440 21660 31560
rect 24540 31440 25560 31560
rect 1305 31140 20895 31260
rect 24540 31260 24660 31440
rect 24105 31140 24660 31260
rect 25440 31260 25560 31440
rect 25905 31440 27495 31560
rect 27705 31440 29880 31560
rect 30405 31440 35595 31560
rect 38505 31440 40095 31560
rect 48405 31440 53595 31560
rect 65205 31440 69195 31560
rect 70905 31440 73995 31560
rect 76905 31440 80595 31560
rect 83805 31440 87795 31560
rect 25440 31140 29595 31260
rect 30705 31140 31380 31260
rect 31905 31140 32295 31260
rect 38205 31140 41295 31260
rect 41505 31140 51795 31260
rect 54105 31140 59895 31260
rect 60105 31140 63195 31260
rect 66405 31140 68895 31260
rect 79005 31140 80295 31260
rect 4605 30840 8895 30960
rect 15705 30840 21195 30960
rect 23205 30840 23595 30960
rect 25005 30840 33495 30960
rect 37005 30840 37695 30960
rect 51105 30840 71295 30960
rect 76305 30840 79395 30960
rect 81105 30840 83595 30960
rect 85305 30840 88995 30960
rect 13605 30540 20295 30660
rect 22005 30540 23880 30660
rect 24405 30540 30495 30660
rect 31605 30540 32295 30660
rect 33405 30540 36495 30660
rect 53505 30540 54795 30660
rect 68040 30540 70695 30660
rect 1605 30240 4395 30360
rect 8205 30240 9195 30360
rect 10605 30240 11595 30360
rect 31305 30240 34995 30360
rect 12105 29940 13695 30060
rect 15105 29940 17460 30060
rect 17340 29805 17460 29940
rect 22305 29940 25695 30060
rect 32295 30090 32505 30240
rect 37005 30240 40695 30360
rect 40905 30240 48195 30360
rect 48405 30240 50760 30360
rect 50640 30105 50760 30240
rect 68040 30360 68160 30540
rect 62505 30240 65760 30360
rect 33705 29940 34260 30060
rect 6105 29640 7395 29760
rect 7605 29640 11595 29760
rect 17505 29640 19695 29760
rect 31305 29640 31695 29760
rect 34140 29760 34260 29940
rect 34605 29940 35895 30060
rect 38205 29940 50280 30060
rect 50805 29940 52695 30060
rect 64005 29940 64695 30060
rect 65640 30060 65760 30240
rect 67740 30240 68160 30360
rect 65640 29940 67095 30060
rect 36495 29760 36705 29895
rect 34140 29700 36705 29760
rect 34140 29640 36660 29700
rect 39105 29640 42795 29760
rect 53505 29640 54495 29760
rect 55140 29640 58695 29760
rect 1740 28605 1860 29310
rect 4605 29340 4860 29460
rect 2640 28905 2760 29295
rect 3840 28860 3960 29310
rect 4740 28905 4860 29340
rect 6705 29340 7995 29460
rect 9690 29295 9705 29400
rect 10005 29340 11295 29460
rect 5340 28905 5460 29295
rect 9495 29160 9705 29295
rect 12240 29160 12360 29310
rect 9495 29100 9960 29160
rect 11940 29100 12360 29160
rect 9540 29040 9960 29100
rect 9840 28905 9960 29040
rect 3405 28740 3960 28860
rect 6405 28740 7695 28860
rect 7905 28725 8895 28845
rect 9705 28860 9960 28905
rect 11895 29040 12360 29100
rect 11895 28905 12105 29040
rect 9705 28740 10095 28860
rect 9705 28695 9900 28740
rect 12840 28605 12960 29310
rect 14505 29355 15495 29475
rect 18705 29355 19095 29475
rect 20100 29460 20295 29505
rect 13395 29160 13605 29295
rect 13140 29100 13605 29160
rect 13140 29040 13560 29100
rect 13140 28890 13260 29040
rect 13905 28740 14595 28860
rect 16740 28860 16860 29310
rect 20040 29295 20295 29460
rect 22605 29340 22995 29460
rect 24405 29355 25395 29475
rect 28005 29340 28860 29460
rect 20040 28890 20160 29295
rect 20895 29160 21105 29295
rect 20895 29100 28395 29160
rect 20940 29040 28395 29100
rect 28740 29160 28860 29340
rect 29205 29340 31395 29460
rect 32205 29355 33495 29475
rect 33705 29340 37080 29460
rect 37905 29355 38595 29475
rect 43905 29355 44295 29475
rect 45405 29355 46095 29475
rect 49005 29355 49395 29475
rect 50505 29355 51195 29475
rect 55140 29460 55260 29640
rect 62595 29760 62805 29895
rect 67740 29805 67860 30240
rect 68505 30240 69195 30360
rect 73305 30240 81795 30360
rect 86805 30240 89295 30360
rect 89505 30240 90495 30360
rect 77805 29940 80895 30060
rect 84705 29940 85095 30060
rect 61605 29700 62805 29760
rect 61605 29640 62760 29700
rect 63915 29640 64995 29760
rect 67740 29640 67995 29805
rect 67800 29595 67995 29640
rect 69705 29640 70995 29760
rect 73605 29640 74595 29760
rect 75405 29640 76395 29760
rect 83205 29640 83895 29760
rect 87105 29640 87795 29760
rect 51405 29340 55260 29460
rect 55605 29340 56895 29460
rect 57705 29355 58395 29475
rect 28740 29040 34695 29160
rect 40140 28905 40260 29310
rect 59340 29160 59460 29310
rect 41505 29040 44760 29160
rect 15405 28740 16860 28860
rect 17805 28740 19995 28860
rect 24705 28740 29295 28860
rect 36705 28725 37395 28845
rect 40005 28740 40260 28905
rect 44640 28890 44760 29040
rect 54240 29040 59460 29160
rect 40005 28695 40200 28740
rect 47505 28740 47895 28860
rect 48105 28725 48495 28845
rect 54240 28860 54360 29040
rect 53205 28740 54360 28860
rect 54705 28725 55695 28845
rect 60705 28740 61395 28860
rect 63240 28860 63360 29295
rect 64140 29160 64260 29310
rect 64140 29040 64560 29160
rect 64440 28905 64560 29040
rect 65205 29160 65400 29205
rect 65205 29100 65460 29160
rect 65205 28995 65505 29100
rect 65295 28905 65505 28995
rect 63240 28740 63795 28860
rect 64440 28740 64695 28905
rect 64500 28695 64695 28740
rect 3105 28440 5595 28560
rect 26505 28440 30795 28560
rect 33705 28440 35895 28560
rect 43305 28440 43695 28560
rect 43905 28440 44580 28560
rect 45105 28440 49395 28560
rect 65205 28440 65595 28560
rect 65940 28560 66060 29310
rect 66540 28860 66660 29310
rect 69105 29340 69795 29460
rect 72105 29340 73260 29460
rect 66540 28740 68295 28860
rect 70440 28860 70560 29310
rect 73140 29160 73260 29340
rect 74040 29160 74160 29310
rect 76095 29160 76305 29295
rect 73140 29040 74160 29160
rect 70440 28740 70995 28860
rect 72405 28800 72660 28860
rect 72405 28740 72705 28800
rect 72495 28605 72705 28740
rect 74040 28605 74160 29040
rect 75540 29100 76305 29160
rect 77340 29340 77895 29460
rect 75540 29040 76260 29100
rect 75540 28860 75660 29040
rect 74505 28740 75660 28860
rect 77340 28860 77460 29340
rect 76905 28740 77460 28860
rect 79125 28860 79245 29295
rect 78405 28740 79245 28860
rect 79440 28605 79560 29310
rect 65940 28440 66495 28560
rect 76005 28440 76395 28560
rect 79305 28440 79560 28605
rect 80040 28560 80160 29310
rect 82605 29340 83295 29460
rect 85005 29355 85995 29475
rect 88305 29340 88695 29460
rect 81495 29160 81705 29295
rect 81495 29100 83895 29160
rect 81540 29040 83895 29100
rect 80505 28740 81180 28860
rect 81705 28725 82095 28845
rect 82905 28725 83595 28845
rect 84405 28740 85095 28860
rect 86505 28740 88995 28860
rect 89205 28725 91095 28845
rect 80040 28440 81795 28560
rect 79305 28395 79500 28440
rect 87105 28440 88095 28560
rect 5940 28140 8295 28260
rect 705 27840 1395 27960
rect 2205 27840 4995 27960
rect 5940 27960 6060 28140
rect 11805 28140 12495 28260
rect 16305 28140 16995 28260
rect 19905 28140 20595 28260
rect 23205 28140 25395 28260
rect 29805 28140 30495 28260
rect 38340 28140 46695 28260
rect 38340 28005 38460 28140
rect 47505 28140 52995 28260
rect 53205 28140 56595 28260
rect 58605 28140 59595 28260
rect 59805 28140 63195 28260
rect 63405 28140 64395 28260
rect 64605 28140 67695 28260
rect 68505 28140 69495 28260
rect 82305 28140 83880 28260
rect 84405 28140 85695 28260
rect 88005 28140 89595 28260
rect 5205 27840 6060 27960
rect 25905 27840 26580 27960
rect 27105 27840 31395 27960
rect 33405 27840 34995 27960
rect 37005 27840 38295 27960
rect 42705 27840 45495 27960
rect 49605 27840 53595 27960
rect 57405 27840 59595 27960
rect 61005 27840 64095 27960
rect 66405 27840 67095 27960
rect 69405 27840 77595 27960
rect 82005 27840 85995 27960
rect 1905 27540 4095 27660
rect 4305 27540 6495 27660
rect 6705 27540 10695 27660
rect 31905 27540 32895 27660
rect 33105 27540 35595 27660
rect 35805 27540 40695 27660
rect 43905 27540 45195 27660
rect 55905 27540 60795 27660
rect 71805 27540 76095 27660
rect 78105 27540 80595 27660
rect 84705 27540 85395 27660
rect 88905 27540 89295 27660
rect 13005 27240 16095 27360
rect 16305 27240 18795 27360
rect 19005 27240 23295 27360
rect 24105 27240 24795 27360
rect 25605 27240 27195 27360
rect 29205 27240 29895 27360
rect 30105 27240 35880 27360
rect 36405 27240 41295 27360
rect 51105 27240 64695 27360
rect 64905 27240 67095 27360
rect 67305 27240 69495 27360
rect 73305 27240 74595 27360
rect 75405 27240 76560 27360
rect 76440 27105 76560 27240
rect 88605 27240 89595 27360
rect 1005 26940 3495 27060
rect 10905 26940 13695 27060
rect 13905 26940 14295 27060
rect 21105 26940 23595 27060
rect 23805 26940 25095 27060
rect 37605 26940 39495 27060
rect 40605 26940 41895 27060
rect 42105 26940 46095 27060
rect 46305 26940 49995 27060
rect 55005 26940 56895 27060
rect 60105 26940 61095 27060
rect 76440 26940 76695 27105
rect 76500 26895 76695 26940
rect 79905 26940 84495 27060
rect 4005 26640 6060 26760
rect 5940 26460 6060 26640
rect 17505 26640 18195 26760
rect 22005 26640 22395 26760
rect 31905 26640 32595 26760
rect 34905 26640 36195 26760
rect 40905 26640 42795 26760
rect 43005 26640 44895 26760
rect 46905 26640 48795 26760
rect 54405 26640 57795 26760
rect 58005 26640 61995 26760
rect 65505 26640 66195 26760
rect 70605 26640 74595 26760
rect 78300 26760 78495 26805
rect 78240 26595 78495 26760
rect 82605 26640 84195 26760
rect 4905 26340 5760 26460
rect 5940 26340 6660 26460
rect 1005 26040 1695 26160
rect 2505 26040 3195 26160
rect 3405 26040 4395 26160
rect 5640 26160 5760 26340
rect 5640 26040 6360 26160
rect 2205 25425 2895 25545
rect 3105 25440 4095 25560
rect 4440 25560 4560 26010
rect 4440 25440 5595 25560
rect 6240 25590 6360 26040
rect 6540 25305 6660 26340
rect 7605 26340 8295 26460
rect 12105 26340 13095 26460
rect 13305 26340 19995 26460
rect 20205 26340 21495 26460
rect 24405 26340 25395 26460
rect 25605 26340 27495 26460
rect 29505 26340 30195 26460
rect 36105 26340 39495 26460
rect 46605 26340 47460 26460
rect 8640 25605 8760 26010
rect 9705 26160 9900 26205
rect 9705 25995 9960 26160
rect 10305 26055 11295 26175
rect 12405 26040 13995 26160
rect 17940 26040 19395 26160
rect 7005 25425 7395 25545
rect 8640 25440 8895 25605
rect 8700 25395 8895 25440
rect 9840 25590 9960 25995
rect 11205 25440 13095 25560
rect 13305 25425 14595 25545
rect 14940 25560 15060 26010
rect 17940 25605 18060 26040
rect 21840 26040 22395 26160
rect 21840 25905 21960 26040
rect 23400 26160 23595 26205
rect 18540 25740 19995 25860
rect 14940 25440 16395 25560
rect 18540 25590 18660 25740
rect 21705 25740 21960 25905
rect 23340 25995 23595 26160
rect 24705 26040 25260 26160
rect 26340 26100 30195 26160
rect 21705 25695 21900 25740
rect 23340 25590 23460 25995
rect 25140 25590 25260 26040
rect 26295 26040 30195 26100
rect 26295 25890 26505 26040
rect 31605 26055 31995 26175
rect 32640 26040 33195 26160
rect 29205 25425 29895 25545
rect 30840 25560 30960 26010
rect 32640 25860 32760 26040
rect 33540 26040 34395 26160
rect 33540 25860 33660 26040
rect 38340 25860 38460 26010
rect 40005 26040 40395 26160
rect 40605 26040 43995 26160
rect 32340 25740 32760 25860
rect 32940 25740 33660 25860
rect 37440 25740 38460 25860
rect 30840 25440 31695 25560
rect 32340 25590 32460 25740
rect 32940 25590 33060 25740
rect 37440 25605 37560 25740
rect 34905 25425 35595 25545
rect 37305 25440 37560 25605
rect 37305 25395 37500 25440
rect 38205 25425 39180 25545
rect 39705 25440 40095 25560
rect 41205 25440 42195 25560
rect 43605 25425 46395 25545
rect 47340 25560 47460 26340
rect 63105 26340 64395 26460
rect 69105 26460 69300 26505
rect 69105 26295 69360 26460
rect 70005 26460 70200 26505
rect 70005 26295 70260 26460
rect 70905 26340 71295 26460
rect 71505 26340 72795 26460
rect 49005 26040 50895 26160
rect 51600 26160 51795 26205
rect 51540 25995 51795 26160
rect 52605 26055 52995 26175
rect 53205 26040 53595 26160
rect 57705 26055 58395 26175
rect 51540 25860 51660 25995
rect 59040 25860 59160 26010
rect 51240 25800 51660 25860
rect 58740 25800 59160 25860
rect 51195 25740 51660 25800
rect 58695 25740 59160 25800
rect 51195 25605 51405 25740
rect 47340 25440 49260 25560
rect 11505 25140 11895 25260
rect 15405 25140 16995 25260
rect 25905 25140 27195 25260
rect 27405 25140 31095 25260
rect 49140 25260 49260 25440
rect 49605 25440 49995 25560
rect 50205 25425 50595 25545
rect 58695 25605 58905 25740
rect 59640 25605 59760 25995
rect 52305 25425 52695 25545
rect 54105 25425 57795 25545
rect 60540 25305 60660 26010
rect 60840 25590 60960 26295
rect 61140 26040 65295 26160
rect 49140 25140 49995 25260
rect 17040 24960 17160 25095
rect 61140 25260 61260 26040
rect 62205 25425 62595 25545
rect 67740 25560 67860 26010
rect 69240 25605 69360 26295
rect 70140 25605 70260 26295
rect 71940 26040 72495 26160
rect 67740 25440 68880 25560
rect 71940 25590 72060 26040
rect 74295 25860 74505 25995
rect 73740 25800 74505 25860
rect 73740 25740 74460 25800
rect 73740 25560 73860 25740
rect 75840 25605 75960 25995
rect 78240 25605 78360 26595
rect 79905 26340 80895 26460
rect 81105 26340 83505 26460
rect 83295 26220 83505 26340
rect 87240 26460 87360 27195
rect 85905 26340 87360 26460
rect 82440 26040 82695 26160
rect 78795 25860 79005 25995
rect 78795 25800 80760 25860
rect 78840 25740 80805 25800
rect 80595 25605 80805 25740
rect 72705 25440 73860 25560
rect 60705 25140 61260 25260
rect 61605 25140 63495 25260
rect 66405 25140 67395 25260
rect 74205 25140 75495 25260
rect 81540 25260 81660 25995
rect 82440 25305 82560 26040
rect 83505 26055 83895 26175
rect 87840 25890 87960 27195
rect 84840 25560 84960 25710
rect 88140 25740 89295 25860
rect 88140 25560 88260 25740
rect 84240 25440 84960 25560
rect 85140 25500 88260 25560
rect 85095 25440 88260 25500
rect 80505 25140 81660 25260
rect 82305 25140 82560 25305
rect 82305 25095 82500 25140
rect 84240 25260 84360 25440
rect 85095 25305 85305 25440
rect 83805 25140 84360 25260
rect 85275 25200 85305 25305
rect 17040 24840 19095 24960
rect 20805 24840 24195 24960
rect 34305 24840 37395 24960
rect 38640 24840 40095 24960
rect 38640 24705 38760 24840
rect 40305 24840 47295 24960
rect 62505 24840 65295 24960
rect 67905 24840 69795 24960
rect 77505 24840 79395 24960
rect 5805 24540 10395 24660
rect 22905 24540 26295 24660
rect 28905 24540 33495 24660
rect 34605 24540 38595 24660
rect 39405 24540 42195 24660
rect 44205 24540 53295 24660
rect 74805 24540 76095 24660
rect 83205 24540 85395 24660
rect 16140 24240 25995 24360
rect 6105 23940 8895 24060
rect 9105 23940 14895 24060
rect 16140 24060 16260 24240
rect 32505 24240 37860 24360
rect 15705 23940 16260 24060
rect 21405 23940 29295 24060
rect 31605 23940 34695 24060
rect 37740 24060 37860 24240
rect 46305 24240 48495 24360
rect 58905 24240 64995 24360
rect 79305 24240 82095 24360
rect 37740 23940 43695 24060
rect 49005 23940 54795 24060
rect 55005 23940 57195 24060
rect 57405 23940 57795 24060
rect 58005 23940 65595 24060
rect 65805 23940 68295 24060
rect 77340 23940 78495 24060
rect 1605 23640 6195 23760
rect 24105 23640 26580 23760
rect 27105 23640 31260 23760
rect 2505 23340 4995 23460
rect 7305 23340 12495 23460
rect 15105 23340 27795 23460
rect 31140 23460 31260 23640
rect 65505 23640 69795 23760
rect 77340 23760 77460 23940
rect 85740 23805 85860 25095
rect 89640 25005 89760 25995
rect 90105 25740 90660 25860
rect 90540 25305 90660 25740
rect 70005 23640 77460 23760
rect 31140 23340 34395 23460
rect 35205 23340 44595 23460
rect 51405 23340 54195 23460
rect 64605 23340 72495 23460
rect 72705 23340 77595 23460
rect 19905 23040 22395 23160
rect 24240 23040 28695 23160
rect 24240 22905 24360 23040
rect 35040 23160 35160 23295
rect 32505 23040 35160 23160
rect 36405 23040 43095 23160
rect 78105 23040 79095 23160
rect 79905 23040 81495 23160
rect 1905 22740 3195 22860
rect 3405 22740 6495 22860
rect 16305 22740 17595 22860
rect 23505 22740 24180 22860
rect 24705 22740 26895 22860
rect 28005 22740 28995 22860
rect 29205 22740 31980 22860
rect 36240 22860 36360 22995
rect 32505 22740 36360 22860
rect 36705 22740 42960 22860
rect 4005 22440 4695 22560
rect 22905 22440 23895 22560
rect 31005 22440 33195 22560
rect 33405 22440 33795 22560
rect 42840 22560 42960 22740
rect 49305 22740 51495 22860
rect 57105 22740 62595 22860
rect 71505 22740 74295 22860
rect 74505 22740 75495 22860
rect 75705 22740 76995 22860
rect 89505 22740 91095 22860
rect 42840 22440 48795 22560
rect 52905 22440 55995 22560
rect 64905 22440 66195 22560
rect 73605 22440 74295 22560
rect 74505 22440 80595 22560
rect 80805 22440 81195 22560
rect 10905 22140 12195 22260
rect 13905 22140 15795 22260
rect 16605 22140 17295 22260
rect 18705 22140 19995 22260
rect 20805 22140 21495 22260
rect 22305 22140 36495 22260
rect 49440 22140 54495 22260
rect 49440 22005 49560 22140
rect 63105 22140 64095 22260
rect 69705 22140 70395 22260
rect 76905 22140 77895 22260
rect 82005 22140 84360 22260
rect 8505 21840 9795 21960
rect 10605 21840 13095 21960
rect 13305 21840 14295 21960
rect 14505 21840 20460 21960
rect 6705 21540 7695 21660
rect 7905 21555 9495 21675
rect 18105 21555 19095 21675
rect 20340 21660 20460 21840
rect 22605 21840 27780 21960
rect 28305 21840 28395 21960
rect 28605 21840 32295 21960
rect 33840 21840 37080 21960
rect 20340 21540 25695 21660
rect 28905 21555 30195 21675
rect 33840 21660 33960 21840
rect 37605 21840 38595 21960
rect 38805 21840 39495 21960
rect 42705 21840 44595 21960
rect 44805 21840 46095 21960
rect 48105 21840 49395 21960
rect 65205 21840 65895 21960
rect 66105 21840 68595 21960
rect 73905 21840 74595 21960
rect 76005 21960 76200 22005
rect 76005 21795 76260 21960
rect 82605 21840 83895 21960
rect 32805 21540 33960 21660
rect 34305 21540 35460 21660
rect 16440 21105 16560 21495
rect 26895 21360 27105 21495
rect 26640 21300 27105 21360
rect 26640 21240 27060 21300
rect 3705 20925 4995 21045
rect 12705 20925 13095 21045
rect 21705 20925 22695 21045
rect 24405 20940 25095 21060
rect 26640 21060 26760 21240
rect 26205 20940 26760 21060
rect 27405 20940 28995 21060
rect 30705 20925 31395 21045
rect 10605 20640 14295 20760
rect 16005 20640 17295 20760
rect 17505 20640 18795 20760
rect 20205 20640 21795 20760
rect 23505 20595 23595 20805
rect 28005 20640 28695 20760
rect 32640 20760 32760 21510
rect 35340 21360 35460 21540
rect 35805 21540 37095 21660
rect 37305 21540 37695 21660
rect 38340 21540 40095 21660
rect 35340 21240 36360 21360
rect 33405 20940 33795 21060
rect 36240 20805 36360 21240
rect 38340 21060 38460 21540
rect 41505 21555 41895 21675
rect 44340 21540 45495 21660
rect 44340 21360 44460 21540
rect 46905 21555 47280 21675
rect 49005 21555 49680 21675
rect 50205 21660 50400 21705
rect 50205 21495 50460 21660
rect 51195 21660 51405 21795
rect 50805 21600 51405 21660
rect 50805 21540 51360 21600
rect 52305 21555 53295 21675
rect 55605 21555 56595 21675
rect 57405 21540 58995 21660
rect 47595 21360 47805 21495
rect 50340 21360 50460 21495
rect 44040 21240 44460 21360
rect 44640 21240 47460 21360
rect 47595 21300 48060 21360
rect 47640 21240 48060 21300
rect 50340 21300 52560 21360
rect 50340 21240 52605 21300
rect 38205 20940 38460 21060
rect 44040 21060 44160 21240
rect 43305 20940 44160 21060
rect 44640 21060 44760 21240
rect 47340 21105 47460 21240
rect 47940 21105 48060 21240
rect 52395 21105 52605 21240
rect 44505 20940 44760 21060
rect 45105 20940 45795 21060
rect 47340 20940 47595 21105
rect 47400 20895 47595 20940
rect 47940 20940 48180 21105
rect 48000 20895 48180 20940
rect 48705 20925 49080 21045
rect 49605 20940 50295 21060
rect 51105 20940 51495 21060
rect 54405 20940 55695 21060
rect 32640 20640 33195 20760
rect 41505 20640 41895 20760
rect 44895 20760 45105 20880
rect 43605 20640 45105 20760
rect 52440 20760 52560 20895
rect 59340 21060 59460 21795
rect 59805 21540 61095 21660
rect 62205 21540 63795 21660
rect 58905 20940 59460 21060
rect 60705 20925 61395 21045
rect 66705 20940 67095 21060
rect 52440 20640 56595 20760
rect 68040 20760 68160 21510
rect 71805 21540 72795 21660
rect 68940 21060 69060 21495
rect 74040 21105 74160 21495
rect 76140 21105 76260 21795
rect 77805 21540 78480 21660
rect 68505 20940 69060 21060
rect 69705 20925 70095 21045
rect 72105 20940 73095 21060
rect 78840 21060 78960 21495
rect 76905 20940 78960 21060
rect 80340 21060 80460 21495
rect 80940 21360 81060 21795
rect 81405 21540 81960 21660
rect 81840 21360 81960 21540
rect 80940 21240 81660 21360
rect 81840 21240 82095 21360
rect 80340 20940 80895 21060
rect 81540 21060 81660 21240
rect 83205 21225 83595 21345
rect 81540 20940 82395 21060
rect 67605 20640 68160 20760
rect 74505 20640 75195 20760
rect 83205 20640 83895 20760
rect 2205 20340 4695 20460
rect 4905 20340 10095 20460
rect 10905 20340 11895 20460
rect 12105 20340 13995 20460
rect 14205 20340 27195 20460
rect 30105 20340 31695 20460
rect 32505 20340 34095 20460
rect 34905 20340 37695 20460
rect 39405 20340 40995 20460
rect 46605 20340 46995 20460
rect 49905 20340 52095 20460
rect 53805 20340 54495 20460
rect 54705 20340 55095 20460
rect 57105 20340 57795 20460
rect 59505 20340 64095 20460
rect 64305 20340 65895 20460
rect 69405 20340 73560 20460
rect 4905 20040 7095 20160
rect 7305 20040 10095 20160
rect 15405 20040 16695 20160
rect 41505 20040 42195 20160
rect 43005 20040 44295 20160
rect 44505 20040 47295 20160
rect 47505 20040 47895 20160
rect 48105 20040 58095 20160
rect 70305 20040 71895 20160
rect 73440 20160 73560 20340
rect 73905 20340 75795 20460
rect 76005 20340 79395 20460
rect 79605 20340 82095 20460
rect 84240 20460 84360 22140
rect 85740 21360 85860 22695
rect 89205 22140 90795 22260
rect 88740 21540 90195 21660
rect 85740 21240 85995 21360
rect 88740 21360 88860 21540
rect 88005 21240 88860 21360
rect 90705 20940 93165 21060
rect 83505 20340 84360 20460
rect 73440 20040 74295 20160
rect 89505 20040 90195 20160
rect 1905 19740 5295 19860
rect 16305 19740 18795 19860
rect 27405 19740 29595 19860
rect 31905 19740 40095 19860
rect 40305 19740 58695 19860
rect 83805 19740 85095 19860
rect 85905 19740 89595 19860
rect 7605 19440 12795 19560
rect 13005 19440 15495 19560
rect 20505 19440 23295 19560
rect 23505 19440 26595 19560
rect 32505 19440 34695 19560
rect 40005 19440 41295 19560
rect 42105 19440 46395 19560
rect 46605 19440 50160 19560
rect 50040 19305 50160 19440
rect 53205 19440 54195 19560
rect 70905 19440 72195 19560
rect 83205 19440 85395 19560
rect 88005 19440 89460 19560
rect 8205 19140 10695 19260
rect 10905 19140 11295 19260
rect 16605 19140 16995 19260
rect 17205 19140 17895 19260
rect 37140 19140 41595 19260
rect 37140 19005 37260 19140
rect 50205 19140 51795 19260
rect 62805 19140 64995 19260
rect 82305 19140 83295 19260
rect 89340 19260 89460 19440
rect 89340 19140 91395 19260
rect 3105 18840 4095 18960
rect 9705 18840 12195 18960
rect 12405 18840 14595 18960
rect 19605 18840 19995 18960
rect 22905 18840 27795 18960
rect 32505 18840 37095 18960
rect 43005 18840 45495 18960
rect 45705 18840 48495 18960
rect 53805 18840 58395 18960
rect 58605 18840 59295 18960
rect 60405 18840 61695 18960
rect 77505 18840 81195 18960
rect 8505 18540 9795 18660
rect 24405 18540 25395 18660
rect 31005 18540 31695 18660
rect 33390 18495 33405 18600
rect 33705 18540 34995 18660
rect 37905 18540 40695 18660
rect 47340 18540 48195 18660
rect 1440 17790 1560 18495
rect 2505 18240 3795 18360
rect 4005 18240 4995 18360
rect 5340 18240 5595 18360
rect 5340 18060 5460 18240
rect 3540 17940 5460 18060
rect 3540 17790 3660 17940
rect -360 17640 495 17760
rect 2205 17625 2895 17745
rect 6240 17760 6360 18210
rect 11205 18240 11595 18360
rect 12600 18360 12795 18405
rect 12540 18195 12795 18360
rect 6240 17640 7095 17760
rect 12540 17790 12660 18195
rect 13740 18060 13860 18210
rect 15705 18240 16395 18360
rect 17040 18240 19395 18360
rect 17040 18060 17160 18240
rect 19740 18240 21495 18360
rect 13740 17940 14460 18060
rect 16140 18000 17160 18060
rect 7905 17640 9195 17760
rect 10005 17625 10695 17745
rect 10905 17640 11895 17760
rect 14340 17760 14460 17940
rect 16095 17940 17160 18000
rect 16095 17805 16305 17940
rect 19740 17805 19860 18240
rect 26205 18240 26895 18360
rect 28005 18240 28695 18360
rect 30405 18360 30600 18405
rect 30405 18195 30660 18360
rect 32790 18195 32805 18300
rect 33195 18360 33405 18495
rect 33105 18300 33405 18360
rect 33105 18240 33345 18300
rect 34605 18240 35595 18360
rect 22140 18000 24195 18060
rect 22095 17940 24195 18000
rect 22095 17805 22305 17940
rect 30540 17805 30660 18195
rect 32595 18060 32805 18195
rect 32595 18000 33360 18060
rect 32640 17940 33360 18000
rect 14340 17640 14895 17760
rect 20805 17625 21195 17745
rect 27105 17625 27495 17745
rect 33240 17790 33360 17940
rect 35940 17790 36060 18495
rect 36540 18240 38295 18360
rect 36540 17790 36660 18240
rect 39705 18240 40995 18360
rect 43905 18255 46095 18375
rect 42240 17805 42360 18210
rect 31905 17625 32295 17745
rect 34005 17625 34395 17745
rect 42105 17640 42360 17805
rect 46440 17790 46560 18495
rect 46905 18240 47160 18360
rect 47040 17805 47160 18240
rect 47340 18060 47460 18540
rect 51405 18540 52395 18660
rect 52605 18540 52995 18660
rect 63705 18540 67695 18660
rect 50505 18240 50895 18360
rect 47340 17940 47760 18060
rect 42105 17595 42300 17640
rect 43305 17625 43695 17745
rect 43905 17640 44595 17760
rect 47640 17505 47760 17940
rect 47940 17760 48060 18195
rect 48840 17940 49995 18060
rect 48840 17790 48960 17940
rect 52095 18060 52305 18195
rect 56040 18240 57195 18360
rect 52095 18000 52860 18060
rect 52140 17940 52860 18000
rect 47940 17640 48195 17760
rect 51405 17625 52395 17745
rect 52740 17760 52860 17940
rect 52740 17640 53295 17760
rect 54105 17625 54495 17745
rect 56040 17760 56160 18240
rect 58005 18240 59160 18360
rect 59040 17790 59160 18240
rect 60105 18240 60795 18360
rect 62505 18240 63195 18360
rect 64305 18240 66060 18360
rect 65940 17790 66060 18240
rect 66540 17790 66660 18540
rect 70305 18240 70695 18360
rect 70905 18285 71595 18405
rect 76005 18240 79680 18360
rect 80205 18240 80595 18360
rect 82905 18255 83295 18375
rect 85605 18240 86160 18360
rect 55605 17640 56160 17760
rect 59805 17625 60495 17745
rect 67440 17760 67560 18195
rect 72240 17805 72360 18195
rect 81795 18060 82005 18195
rect 81795 18000 84195 18060
rect 81840 17940 84195 18000
rect 85305 17955 85695 18075
rect 86040 18060 86160 18240
rect 89040 18240 89895 18360
rect 86040 17940 88095 18060
rect 67440 17640 67995 17760
rect 14205 17340 15195 17460
rect 16005 17340 17295 17460
rect 20505 17340 21795 17460
rect 31305 17340 34695 17460
rect 34905 17340 37995 17460
rect 38805 17340 41295 17460
rect 42705 17340 45195 17460
rect 47640 17340 47895 17505
rect 47700 17295 47895 17340
rect 56205 17340 57495 17460
rect 58995 17460 59205 17580
rect 73605 17640 75195 17760
rect 77205 17640 80595 17760
rect 81705 17640 82095 17760
rect 84240 17760 84360 17910
rect 83205 17640 84360 17760
rect 58995 17340 61995 17460
rect 74505 17340 78795 17460
rect 79815 17340 82695 17460
rect 85800 17460 85995 17505
rect 85740 17400 85995 17460
rect 85695 17295 85995 17400
rect 85695 17205 85905 17295
rect 6105 17040 8295 17160
rect 10005 17040 13095 17160
rect 52005 17040 55395 17160
rect 59505 17040 61395 17160
rect 63105 17040 66495 17160
rect 72105 17040 79095 17160
rect 19305 16740 22095 16860
rect 65205 16740 66780 16860
rect 67305 16740 70080 16860
rect 70605 16740 79395 16860
rect 80505 16740 82695 16860
rect 705 16440 12795 16560
rect 21405 16440 22695 16560
rect 28005 16440 34995 16560
rect 35805 16440 69495 16560
rect 76440 16440 83895 16560
rect 6705 16140 12495 16260
rect 16905 16140 19095 16260
rect 24405 16140 28695 16260
rect 30705 16140 34995 16260
rect 59505 16140 64395 16260
rect 65505 16140 70395 16260
rect 76440 16260 76560 16440
rect 89040 16305 89160 18240
rect 91005 18240 91860 18360
rect 90405 17940 91560 18060
rect 89640 17160 89760 17895
rect 91440 17505 91560 17940
rect 89640 17040 90135 17160
rect 91740 17160 91860 18240
rect 90345 17040 90360 17160
rect 91740 17040 92460 17160
rect 91005 16740 91995 16860
rect 92340 16305 92460 17040
rect 71505 16140 76560 16260
rect 76905 16140 77295 16260
rect 77505 16140 87795 16260
rect 92205 16140 92460 16305
rect 92205 16095 92400 16140
rect 1605 15840 5895 15960
rect 13005 15840 35595 15960
rect 37905 15840 39495 15960
rect 39705 15840 40095 15960
rect 65205 15840 68295 15960
rect 74505 15840 74895 15960
rect 14805 15540 19995 15660
rect 28905 15540 31395 15660
rect 35505 15540 43395 15660
rect 47505 15540 53895 15660
rect 54105 15540 56295 15660
rect 69105 15540 78195 15660
rect 78405 15540 81795 15660
rect 82605 15540 90495 15660
rect 705 15240 6195 15360
rect 24705 15240 25395 15360
rect 32640 15240 36795 15360
rect 1005 14940 2295 15060
rect 2505 14940 4695 15060
rect 15105 14940 15795 15060
rect 16005 14940 17895 15060
rect 25905 14940 31095 15060
rect 32640 15060 32760 15240
rect 38040 15240 41895 15360
rect 31305 14940 32760 15060
rect 38040 15060 38160 15240
rect 64605 15240 67395 15360
rect 33105 14940 38160 15060
rect 47205 14940 53295 15060
rect 53505 14940 55095 15060
rect 69405 14940 72495 15060
rect 74505 14940 76260 15060
rect 16305 14640 18495 14760
rect 20805 14640 23595 14760
rect 26340 14640 28395 14760
rect 26340 14505 26460 14640
rect 32505 14640 38295 14760
rect 40605 14640 42495 14760
rect 42705 14640 45795 14760
rect 46005 14640 57495 14760
rect 63405 14640 65595 14760
rect 71805 14640 73995 14760
rect 76140 14760 76260 14940
rect 76605 14940 80895 15060
rect 81705 14940 82395 15060
rect 85905 14940 87195 15060
rect 88005 14940 89895 15060
rect 76140 14640 77295 14760
rect 4005 14340 11595 14460
rect 19605 14340 19995 14460
rect 24705 14340 26295 14460
rect 30105 14340 31995 14460
rect 32805 14340 36795 14460
rect 37005 14340 37995 14460
rect 43605 14340 44895 14460
rect 46905 14340 60495 14460
rect 64005 14340 64995 14460
rect 70305 14340 70695 14460
rect 74505 14340 77895 14460
rect 79605 14340 79995 14460
rect 85905 14340 87795 14460
rect 1305 14040 3195 14160
rect 6105 14040 9495 14160
rect 13005 14040 15495 14160
rect 15705 14040 16395 14160
rect 16605 14040 17295 14160
rect 23805 14040 24795 14160
rect 25005 14040 28995 14160
rect 49005 14040 50295 14160
rect 55005 14040 55695 14160
rect 57840 14040 62295 14160
rect 2700 13860 2895 13905
rect 2640 13695 2895 13860
rect 13605 13740 15195 13860
rect 20205 13755 20595 13875
rect 23205 13740 24495 13860
rect 25905 13755 26295 13875
rect 30705 13755 33495 13875
rect 2640 13305 2760 13695
rect 5640 13305 5760 13710
rect 3705 13125 4695 13245
rect 5505 13140 5760 13305
rect 5505 13095 5700 13140
rect 7305 13125 7995 13245
rect 10440 13260 10560 13710
rect 36105 13740 36495 13860
rect 38505 13740 39960 13860
rect 8805 13140 10560 13260
rect 11805 13140 12495 13260
rect 14205 13125 16995 13245
rect 18705 13125 19695 13245
rect 22905 13125 23595 13245
rect 25005 13140 25395 13260
rect 25605 13125 25995 13245
rect 27705 13125 28695 13245
rect 29505 13125 29895 13245
rect 31605 13125 32295 13245
rect 34440 13260 34560 13695
rect 34440 13140 35595 13260
rect 39840 13290 39960 13740
rect 44505 13740 46695 13860
rect 49905 13755 50895 13875
rect 55440 13740 56295 13860
rect 53640 13440 54495 13560
rect 53640 13290 53760 13440
rect 55440 13290 55560 13740
rect 57840 13290 57960 14040
rect 74805 14040 75780 14160
rect 76305 14040 76680 14160
rect 80505 14040 83295 14160
rect 58305 13740 59895 13860
rect 61005 13755 61695 13875
rect 63105 13740 64395 13860
rect 65805 13860 66000 13905
rect 65805 13695 66060 13860
rect 67605 13740 68160 13860
rect 37005 13140 37995 13260
rect 41505 13125 43995 13245
rect 46005 13125 46395 13245
rect 47805 13125 49095 13245
rect 50205 13125 50595 13245
rect 52005 13125 52995 13245
rect 58605 13140 59295 13260
rect 60405 13125 60780 13245
rect 61605 13140 62895 13260
rect 64305 13140 64995 13260
rect 65940 13290 66060 13695
rect 68040 13290 68160 13740
rect 69705 13755 70095 13875
rect 75105 13740 75495 13860
rect 68805 13140 69495 13260
rect 70605 13140 71295 13260
rect 73140 13260 73260 13710
rect 76995 13860 77205 13995
rect 76305 13800 77205 13860
rect 76305 13740 77160 13800
rect 79440 13560 79560 13710
rect 80205 13740 85395 13860
rect 90105 13740 92760 13860
rect 79440 13440 82095 13560
rect 73140 13140 74595 13260
rect 75705 13125 77595 13245
rect 78405 13125 79095 13245
rect 80505 13140 81195 13260
rect 1005 12840 1995 12960
rect 14505 12840 15495 12960
rect 25995 12960 26205 13080
rect 25995 12840 30795 12960
rect 39105 12840 39495 12960
rect 60840 12960 60960 13080
rect 60840 12840 63495 12960
rect 77595 12960 77805 13080
rect 77595 12840 81795 12960
rect 82005 12840 84195 12960
rect 84405 12840 85995 12960
rect 6705 12540 9195 12660
rect 12405 12540 13095 12660
rect 13305 12540 20895 12660
rect 47205 12540 52695 12660
rect 69705 12540 71595 12660
rect 72405 12540 75495 12660
rect 26205 12240 29295 12360
rect 34005 12240 37095 12360
rect 44805 12240 53295 12360
rect 54105 12240 55995 12360
rect 61005 12240 69195 12360
rect 16605 11940 17295 12060
rect 22905 11940 31095 12060
rect 31305 11940 32295 12060
rect 32505 11940 35895 12060
rect 40005 11940 46995 12060
rect 67005 11940 70995 12060
rect 76605 11940 78495 12060
rect 82905 11940 88695 12060
rect 4305 11640 5295 11760
rect 5505 11640 8595 11760
rect 12105 11640 13995 11760
rect 25005 11640 26595 11760
rect 27405 11640 28980 11760
rect 29505 11640 32895 11760
rect 47805 11640 48495 11760
rect 48705 11640 54495 11760
rect 57105 11640 61395 11760
rect 64905 11640 68595 11760
rect 72405 11640 79095 11760
rect 1005 11340 5895 11460
rect 6105 11340 7995 11460
rect 8205 11340 10695 11460
rect 28905 11340 35595 11460
rect 35805 11340 38295 11460
rect 38505 11340 40395 11460
rect 60405 11340 63795 11460
rect 84705 11340 85695 11460
rect 1905 11040 2895 11160
rect 8505 11040 9195 11160
rect 11505 11040 12480 11160
rect 13005 11040 16395 11160
rect 17805 11040 18495 11160
rect 19605 11040 27195 11160
rect 30105 11040 32895 11160
rect 33105 11040 33795 11160
rect 34605 11040 35295 11160
rect 36705 11040 40395 11160
rect 45405 11040 48195 11160
rect 49005 11040 50295 11160
rect 50505 11040 51195 11160
rect 53505 11040 54195 11160
rect 58005 11040 61095 11160
rect 61305 11040 61995 11160
rect 67305 11040 68595 11160
rect 76305 11040 76995 11160
rect 79305 11040 83280 11160
rect 83805 11040 84195 11160
rect 705 10740 1395 10860
rect 27705 10740 33195 10860
rect 33405 10740 36195 10860
rect 36405 10740 36960 10860
rect 2805 10455 5895 10575
rect 6705 10440 7395 10560
rect 8205 10560 8400 10605
rect 8205 10395 8460 10560
rect 9705 10440 10095 10560
rect 11040 10440 12195 10560
rect 8340 9990 8460 10395
rect 11040 9990 11160 10440
rect 13140 10440 13395 10560
rect 13140 10005 13260 10440
rect 14205 10455 14895 10575
rect 1005 9825 1395 9945
rect 4905 9825 5295 9945
rect 15840 9960 15960 10410
rect 17205 10440 17895 10560
rect 19095 10560 19305 10695
rect 18705 10500 19305 10560
rect 18705 10440 19260 10500
rect 19440 10440 20295 10560
rect 19440 10260 19560 10440
rect 21105 10440 21360 10560
rect 18840 10140 19560 10260
rect 18840 9990 18960 10140
rect 21240 10005 21360 10440
rect 22305 10440 23295 10560
rect 13905 9840 15960 9960
rect 19605 9825 20595 9945
rect 24840 9960 24960 10410
rect 26505 10440 26895 10560
rect 28905 10560 29100 10605
rect 28905 10395 29160 10560
rect 31005 10440 31695 10560
rect 23805 9840 24960 9960
rect 25305 9840 25995 9960
rect 29040 9990 29160 10395
rect 26805 9840 27795 9960
rect 33405 9825 34095 9945
rect 35640 9960 35760 10395
rect 36840 9990 36960 10740
rect 40905 10740 44895 10860
rect 55305 10740 55995 10860
rect 64605 10740 65295 10860
rect 70605 10740 71595 10860
rect 74805 10740 76395 10860
rect 82140 10740 84795 10860
rect 39105 10440 44595 10560
rect 37095 10260 37305 10395
rect 37095 10200 38160 10260
rect 37140 10140 38160 10200
rect 38040 9990 38160 10140
rect 40440 9990 40560 10440
rect 51105 10440 51495 10560
rect 46440 10260 46560 10410
rect 50940 10260 51060 10410
rect 54405 10440 55260 10560
rect 46440 10140 48960 10260
rect 34905 9840 35760 9960
rect 42405 9840 42795 9960
rect 45105 9825 45495 9945
rect 48105 9825 48495 9945
rect 48840 9960 48960 10140
rect 50640 10140 51060 10260
rect 55140 10260 55260 10440
rect 56505 10440 57195 10560
rect 82140 10620 82260 10740
rect 85005 10740 86295 10860
rect 55140 10140 55560 10260
rect 50640 9960 50760 10140
rect 48840 9840 50760 9960
rect 53205 9840 53895 9960
rect 55440 9990 55560 10140
rect 62940 10260 63060 10425
rect 66105 10440 66795 10560
rect 72600 10560 72780 10605
rect 61905 10140 63060 10260
rect 63540 10200 64860 10260
rect 63495 10140 64860 10200
rect 63495 10005 63705 10140
rect 54105 9840 54795 9960
rect 56205 9825 57495 9945
rect 60105 9825 61095 9945
rect 64740 9990 64860 10140
rect 67440 10005 67560 10410
rect 64905 9825 66195 9945
rect 67305 9840 67560 10005
rect 72540 10395 72780 10560
rect 73305 10455 73995 10575
rect 75705 10440 79095 10560
rect 79905 10455 80895 10575
rect 81705 10455 82095 10575
rect 83040 10440 84195 10560
rect 72540 9990 72660 10395
rect 83040 9990 83160 10440
rect 85140 10440 89595 10560
rect 85140 10005 85260 10440
rect 67305 9795 67500 9840
rect 76905 9840 78795 9960
rect 5040 9540 6195 9660
rect 705 9240 1995 9360
rect 5040 9360 5160 9540
rect 9105 9540 10095 9660
rect 19440 9660 19560 9780
rect 18405 9540 19560 9660
rect 22605 9540 26295 9660
rect 31605 9540 32895 9660
rect 51705 9540 52260 9660
rect 2205 9240 5160 9360
rect 5505 9240 6795 9360
rect 11805 9240 17295 9360
rect 22305 9240 24495 9360
rect 36405 9240 37395 9360
rect 43905 9240 49095 9360
rect 49305 9240 49995 9360
rect 52140 9360 52260 9540
rect 67905 9540 69795 9660
rect 72405 9540 73095 9660
rect 76005 9540 80595 9660
rect 86805 9540 89895 9660
rect 52140 9240 58095 9360
rect 58305 9240 58695 9360
rect 67005 9240 69195 9360
rect 74805 9240 78195 9360
rect 13905 8940 22395 9060
rect 29805 8940 31995 9060
rect 36240 9060 36360 9195
rect 32205 8940 36360 9060
rect 44805 8940 46995 9060
rect 50805 8940 51795 9060
rect 52005 8940 52395 9060
rect 61605 8940 68895 9060
rect 79005 8940 83595 9060
rect 83805 8940 84795 9060
rect 4305 8640 8895 8760
rect 12705 8640 14295 8760
rect 14505 8640 16095 8760
rect 25005 8640 28395 8760
rect 41205 8640 44295 8760
rect 62505 8640 67095 8760
rect 71205 8640 74895 8760
rect 82005 8640 88095 8760
rect 24405 8340 30495 8460
rect 34305 8340 39795 8460
rect 46905 8340 50595 8460
rect 69105 8340 75195 8460
rect 82605 8340 85695 8460
rect 13305 8040 18195 8160
rect 27405 8040 30195 8160
rect 35505 8040 38595 8160
rect 68805 8040 85395 8160
rect 86805 8040 88995 8160
rect 15105 7740 16395 7860
rect 16605 7740 16995 7860
rect 30705 7740 39795 7860
rect 40005 7740 50595 7860
rect 55605 7740 61695 7860
rect 61905 7740 65595 7860
rect 6405 7440 8295 7560
rect 8505 7440 14295 7560
rect 15705 7440 17595 7560
rect 20805 7440 25395 7560
rect 67605 7440 77295 7560
rect 80805 7440 81195 7560
rect 86805 7440 90195 7560
rect 90405 7440 91695 7560
rect 1905 7140 3795 7260
rect 4005 7140 11895 7260
rect 28005 7140 35295 7260
rect 52305 7140 55395 7260
rect 64905 7140 74595 7260
rect 84105 7140 86895 7260
rect 13005 6840 13395 6960
rect 13605 6840 13995 6960
rect 17805 6840 19095 6960
rect 19305 6840 21195 6960
rect 25905 6840 27195 6960
rect 41505 6840 47895 6960
rect 49305 6840 53595 6960
rect 56805 6840 65295 6960
rect 83505 6840 85995 6960
rect 7605 6540 9195 6660
rect 23805 6540 29595 6660
rect 35805 6540 36795 6660
rect 39405 6540 42495 6660
rect 42705 6540 42795 6660
rect 43005 6540 45195 6660
rect 46305 6540 48195 6660
rect 57405 6540 59595 6660
rect 59805 6540 62295 6660
rect 76005 6540 77295 6660
rect 89205 6540 91095 6660
rect 2505 6240 3195 6360
rect 3405 6240 4695 6360
rect 17640 6240 20895 6360
rect 2340 5940 2895 6060
rect 2340 5460 2460 5940
rect 6540 5940 7695 6060
rect 6540 5490 6660 5940
rect 9705 5955 10395 6075
rect 2205 5340 2460 5460
rect 8805 5340 9495 5460
rect 11040 5460 11160 5910
rect 16740 5505 16860 5895
rect 17640 5760 17760 6240
rect 36840 6360 36960 6495
rect 36840 6240 45795 6360
rect 46005 6240 47295 6360
rect 49005 6240 49395 6360
rect 53205 6240 54495 6360
rect 54705 6240 55695 6360
rect 66105 6240 70695 6360
rect 81705 6240 82395 6360
rect 82605 6240 84195 6360
rect 87405 6240 88095 6360
rect 18000 6060 18195 6105
rect 17340 5640 17760 5760
rect 17940 5895 18195 6060
rect 19905 5955 22095 6075
rect 23340 5940 24795 6060
rect 10305 5340 11160 5460
rect 12105 5340 12495 5460
rect 14505 5340 15195 5460
rect 17340 5490 17460 5640
rect 17940 5490 18060 5895
rect 23340 5760 23460 5940
rect 26205 5955 26595 6075
rect 28005 5940 28995 6060
rect 33195 6075 33405 6195
rect 31005 5955 33495 6075
rect 33240 5940 33360 5955
rect 38805 5940 41295 6060
rect 48705 5955 51195 6075
rect 56505 5955 57795 6075
rect 58005 5940 58995 6060
rect 21405 5640 23460 5760
rect 29040 5760 29160 5910
rect 36240 5760 36360 5910
rect 60705 5940 61695 6060
rect 61905 5940 63195 6060
rect 64005 5955 64395 6075
rect 66705 5940 67995 6060
rect 71805 5985 72795 6105
rect 29040 5640 41160 5760
rect 18105 5340 18795 5460
rect 27705 5340 29295 5460
rect 29640 5460 29760 5640
rect 29640 5340 31395 5460
rect 32205 5325 32580 5445
rect 33105 5325 33795 5445
rect 34605 5340 35595 5460
rect 37305 5340 38295 5460
rect 38505 5340 39195 5460
rect 41040 5490 41160 5640
rect 42105 5640 44595 5760
rect 40005 5340 40395 5460
rect 41205 5340 42795 5460
rect 45705 5340 48495 5460
rect 51105 5325 52095 5445
rect 54705 5325 55095 5445
rect 60105 5340 62895 5460
rect 63705 5340 64695 5460
rect 75540 5490 75660 6195
rect 76605 5940 77895 6060
rect 85200 6060 85395 6105
rect 85140 5895 85395 6060
rect 89805 5955 91395 6075
rect 78840 5640 83895 5760
rect 68505 5340 68895 5460
rect 10005 5040 10695 5160
rect 21105 5040 25995 5160
rect 29295 5160 29505 5280
rect 78840 5460 78960 5640
rect 85140 5460 85260 5895
rect 86805 5325 88095 5445
rect 88905 5325 90495 5445
rect 29295 5040 30495 5160
rect 41505 5040 41895 5160
rect 46305 5040 46995 5160
rect 47205 5040 48195 5160
rect 55605 5040 57495 5160
rect 57705 5040 59295 5160
rect 66405 5040 72195 5160
rect 72405 5040 76095 5160
rect 76305 5040 76995 5160
rect 3705 4740 4695 4860
rect 6105 4740 10095 4860
rect 10305 4740 12195 4860
rect 14205 4740 16695 4860
rect 19305 4740 20595 4860
rect 31305 4740 42495 4860
rect 47805 4740 48495 4860
rect 49905 4740 50295 4860
rect 50505 4740 51495 4860
rect 51705 4740 54795 4860
rect 55005 4740 56295 4860
rect 59205 4740 60795 4860
rect 65805 4740 70095 4860
rect 89505 4740 90195 4860
rect 8205 4440 9195 4560
rect 22605 4440 25995 4560
rect 26805 4440 40695 4560
rect 45705 4440 48795 4560
rect 52905 4440 53595 4560
rect 85905 4440 86595 4560
rect 87405 4440 91995 4560
rect 1605 4140 1995 4260
rect 2205 4140 7395 4260
rect 7605 4140 9795 4260
rect 13905 4140 18495 4260
rect 23205 4140 25695 4260
rect 25905 4140 29895 4260
rect 39105 4140 42195 4260
rect 43605 4140 48495 4260
rect 49305 4140 53295 4260
rect 89805 4140 90795 4260
rect 8205 3840 10995 3960
rect 12705 3840 13395 3960
rect 15105 3840 15795 3960
rect 16005 3840 22095 3960
rect 22740 3840 30195 3960
rect 22740 3705 22860 3840
rect 30405 3840 31695 3960
rect 38505 3840 48195 3960
rect 49005 3840 56895 3960
rect 57105 3840 61395 3960
rect 61605 3840 65295 3960
rect 73905 3840 75195 3960
rect 77505 3840 77895 3960
rect 405 3540 1395 3660
rect 4305 3540 6195 3660
rect 16605 3540 17595 3660
rect 19605 3540 22695 3660
rect 34005 3540 36495 3660
rect 39240 3540 51195 3660
rect 4005 3240 8895 3360
rect 9105 3240 11295 3360
rect 11505 3240 13095 3360
rect 13305 3240 24495 3360
rect 25605 3240 26895 3360
rect 30105 3240 31395 3360
rect 33405 3240 36195 3360
rect 39240 3360 39360 3540
rect 51405 3540 52995 3660
rect 37005 3240 39360 3360
rect 40305 3240 50595 3360
rect 53505 3240 55995 3360
rect 56205 3240 57495 3360
rect 60705 3240 63660 3360
rect 25005 2940 29295 3060
rect 29505 2940 32595 3060
rect 36705 2940 39495 3060
rect 43800 3060 43995 3105
rect 43740 2940 43995 3060
rect 43800 2895 43995 2940
rect 44205 2940 45960 3060
rect 1740 2640 4095 2760
rect 1740 2190 1860 2640
rect 4905 2640 5595 2760
rect 5940 2190 6060 2895
rect 6405 2640 11895 2760
rect 12240 2190 12360 2895
rect 12900 2760 13095 2805
rect 12840 2595 13095 2760
rect 15105 2640 16260 2760
rect 12840 2190 12960 2595
rect 16140 2460 16260 2640
rect 16905 2640 17295 2760
rect 20205 2655 20895 2775
rect 21705 2640 24195 2760
rect 26205 2640 27795 2760
rect 28605 2640 28995 2760
rect 29340 2640 30795 2760
rect 29340 2460 29460 2640
rect 34605 2655 35295 2775
rect 37305 2655 37995 2775
rect 41340 2640 43395 2760
rect 41340 2460 41460 2640
rect 44805 2640 45495 2760
rect 13905 2340 15960 2460
rect 16140 2340 16560 2460
rect 2505 2040 3495 2160
rect 3705 2040 5295 2160
rect 9105 2025 9495 2145
rect 15840 2190 15960 2340
rect 14205 2040 14595 2160
rect 16440 2160 16560 2340
rect 28140 2340 45360 2460
rect 28140 2190 28260 2340
rect 45240 2190 45360 2340
rect 45840 2190 45960 2940
rect 46305 2640 46995 2760
rect 50805 2640 53295 2760
rect 54600 2760 54795 2805
rect 47505 2340 48660 2460
rect 48540 2190 48660 2340
rect 16440 2040 18195 2160
rect 21405 2025 22095 2145
rect 22905 2025 23295 2145
rect 25905 2040 27495 2160
rect 29505 2025 29895 2145
rect 30705 2025 31095 2145
rect 31905 2025 32295 2145
rect 33105 2025 33795 2145
rect 34905 2040 39195 2160
rect 40305 2025 40995 2145
rect 42705 2025 43095 2145
rect 43905 2025 44595 2145
rect 47205 2025 47895 2145
rect 51105 2040 52695 2160
rect 5295 1860 5505 1980
rect 5295 1740 7095 1860
rect 7905 1740 8385 1860
rect 19305 1740 20595 1860
rect 28095 1860 28305 1980
rect 26505 1740 28305 1860
rect 36405 1740 37995 1860
rect 38205 1740 38595 1860
rect 39195 1860 39405 1980
rect 39195 1740 41595 1860
rect 53205 1740 53895 1860
rect 54240 1860 54360 2610
rect 54540 2595 54795 2760
rect 61995 2760 62205 2895
rect 61605 2700 62205 2760
rect 61605 2640 62160 2700
rect 62505 2655 63195 2775
rect 54540 2190 54660 2595
rect 56640 2460 56760 2610
rect 55605 2340 56760 2460
rect 63540 2190 63660 3240
rect 72705 3240 74295 3360
rect 78405 3240 80595 3360
rect 64005 2640 64695 2760
rect 66105 2655 66495 2775
rect 68505 2655 69495 2775
rect 73905 2640 75195 2760
rect 79605 2640 80595 2760
rect 82905 2655 83895 2775
rect 71040 2340 72960 2460
rect 57105 2025 60495 2145
rect 61305 2040 62895 2160
rect 65805 2040 67395 2160
rect 71040 2160 71160 2340
rect 72840 2160 72960 2340
rect 72105 1995 72480 2115
rect 73005 1995 76695 2115
rect 77805 1995 78195 2115
rect 88005 2025 88995 2145
rect 54240 1740 55260 1860
rect 13605 1440 18195 1560
rect 19005 1440 23895 1560
rect 24105 1440 24795 1560
rect 29205 1440 35295 1560
rect 35505 1440 36795 1560
rect 45105 1440 47295 1560
rect 55140 1560 55260 1740
rect 64905 1740 66195 1860
rect 55140 1440 55395 1560
rect 55605 1440 61695 1560
rect 61905 1440 62295 1560
rect 63405 1440 66495 1560
rect 11205 1140 22395 1260
rect 27105 1140 35160 1260
rect 4905 840 25695 960
rect 35040 960 35160 1140
rect 48105 1140 61095 1260
rect 35040 840 36195 960
rect 42405 840 60195 960
rect 64605 840 67995 960
rect 11505 540 19995 660
rect 32205 540 41595 660
rect 43005 540 50895 660
rect 52005 540 56295 660
use INVX1  _889_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 80850 0 -1 27450
box -180 -120 1080 4080
use NOR2X1  _890_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 76050 0 1 19650
box -180 -120 1380 4080
use NAND2X1  _891_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 77850 0 1 19650
box -180 -120 1380 4080
use INVX1  _892_
timestamp 1727136778
transform 1 0 81150 0 -1 19650
box -180 -120 1080 4080
use INVX1  _893_
timestamp 1727136778
transform -1 0 79650 0 1 19650
box -180 -120 1080 4080
use INVX2  _894_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 82950 0 -1 19650
box -180 -120 1080 4080
use NOR2X1  _895_
timestamp 1727136778
transform -1 0 79950 0 -1 27450
box -180 -120 1380 4080
use NAND2X1  _896_
timestamp 1727136778
transform -1 0 78150 0 -1 27450
box -180 -120 1380 4080
use INVX1  _897_
timestamp 1727136778
transform 1 0 77250 0 1 35250
box -180 -120 1080 4080
use NOR2X1  _898_
timestamp 1727136778
transform -1 0 83550 0 -1 27450
box -180 -120 1380 4080
use AOI21X1  _899_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 79350 0 1 27450
box -180 -120 1680 4080
use NOR2X1  _900_
timestamp 1727136778
transform -1 0 89250 0 1 35250
box -180 -120 1380 4080
use OAI21X1  _901_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 87150 0 1 35250
box -180 -120 1680 4080
use INVX1  _902_
timestamp 1727136778
transform 1 0 87450 0 -1 35250
box -180 -120 1080 4080
use INVX4  _903_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 73950 0 1 27450
box -180 -120 1380 4080
use OAI21X1  _904_
timestamp 1727136778
transform -1 0 81750 0 1 19650
box -180 -120 1680 4080
use INVX1  _905_
timestamp 1727136778
transform -1 0 86550 0 -1 35250
box -180 -120 1080 4080
use NOR2X1  _906_
timestamp 1727136778
transform -1 0 64650 0 -1 35250
box -180 -120 1380 4080
use INVX1  _907_
timestamp 1727136778
transform 1 0 75150 0 -1 35250
box -180 -120 1080 4080
use INVX1  _908_
timestamp 1727136778
transform 1 0 89850 0 -1 43050
box -180 -120 1080 4080
use OAI21X1  _909_
timestamp 1727136778
transform 1 0 84450 0 1 27450
box -180 -120 1680 4080
use OAI21X1  _910_
timestamp 1727136778
transform 1 0 83250 0 -1 35250
box -180 -120 1680 4080
use AOI22X1  _911_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 81750 0 1 27450
box -210 -120 1980 4080
use NAND2X1  _912_
timestamp 1727136778
transform 1 0 86850 0 1 27450
box -180 -120 1380 4080
use OAI21X1  _913_
timestamp 1727136778
transform -1 0 85050 0 1 35250
box -180 -120 1680 4080
use OAI21X1  _914_
timestamp 1727136778
transform -1 0 80550 0 1 35250
box -180 -120 1680 4080
use NAND2X1  _915_
timestamp 1727136778
transform 1 0 79050 0 -1 35250
box -180 -120 1380 4080
use NOR2X1  _916_
timestamp 1727136778
transform -1 0 85950 0 1 43050
box -180 -120 1380 4080
use NOR2X1  _917_
timestamp 1727136778
transform 1 0 87750 0 -1 43050
box -180 -120 1380 4080
use OAI22X1  _918_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 82950 0 -1 43050
box -180 -120 1980 4080
use OR2X2  _919_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 81450 0 1 35250
box -180 -120 1680 4080
use INVX1  _920_
timestamp 1727136778
transform -1 0 84450 0 -1 43050
box -180 -120 1080 4080
use AOI22X1  _921_
timestamp 1727136778
transform 1 0 85350 0 -1 43050
box -210 -120 1980 4080
use NAND3X1  _922_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 81150 0 -1 35250
box -180 -120 1680 4080
use AND2X2  _923_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 88950 0 -1 35250
box -180 -120 1680 4095
use OAI21X1  _924_
timestamp 1727136778
transform 1 0 88950 0 1 27450
box -180 -120 1680 4080
use INVX1  _925_
timestamp 1727136778
transform -1 0 90750 0 1 19650
box -180 -120 1080 4080
use INVX1  _926_
timestamp 1727136778
transform -1 0 65850 0 1 66450
box -180 -120 1080 4080
use NAND2X1  _927_
timestamp 1727136778
transform 1 0 73350 0 -1 50850
box -180 -120 1380 4080
use OAI21X1  _928_
timestamp 1727136778
transform 1 0 70950 0 -1 50850
box -180 -120 1680 4080
use INVX1  _929_
timestamp 1727136778
transform 1 0 63450 0 1 66450
box -180 -120 1080 4080
use NAND2X1  _930_
timestamp 1727136778
transform 1 0 55650 0 1 58650
box -180 -120 1380 4080
use OAI21X1  _931_
timestamp 1727136778
transform -1 0 59250 0 1 58650
box -180 -120 1680 4080
use INVX1  _932_
timestamp 1727136778
transform 1 0 62250 0 -1 66450
box -180 -120 1080 4080
use NAND2X1  _933_
timestamp 1727136778
transform -1 0 67650 0 -1 50850
box -180 -120 1380 4080
use OAI21X1  _934_
timestamp 1727136778
transform 1 0 68550 0 -1 50850
box -180 -120 1680 4080
use INVX1  _935_
timestamp 1727136778
transform -1 0 81750 0 1 74250
box -180 -120 1080 4080
use NAND2X1  _936_
timestamp 1727136778
transform 1 0 61650 0 1 66450
box -180 -120 1380 4080
use OAI21X1  _937_
timestamp 1727136778
transform -1 0 61650 0 -1 66450
box -180 -120 1680 4080
use INVX1  _938_
timestamp 1727136778
transform -1 0 60750 0 -1 82050
box -180 -120 1080 4080
use NAND2X1  _939_
timestamp 1727136778
transform 1 0 55350 0 1 66450
box -180 -120 1380 4080
use OAI21X1  _940_
timestamp 1727136778
transform 1 0 52350 0 -1 66450
box -180 -120 1680 4080
use INVX1  _941_
timestamp 1727136778
transform -1 0 49950 0 -1 74250
box -180 -120 1080 4080
use NAND2X1  _942_
timestamp 1727136778
transform 1 0 54750 0 -1 58650
box -180 -120 1380 4080
use OAI21X1  _943_
timestamp 1727136778
transform 1 0 52650 0 -1 58650
box -180 -120 1680 4080
use INVX1  _944_
timestamp 1727136778
transform -1 0 80850 0 1 50850
box -180 -120 1080 4080
use NAND2X1  _945_
timestamp 1727136778
transform 1 0 83850 0 -1 50850
box -180 -120 1380 4080
use OAI21X1  _946_
timestamp 1727136778
transform 1 0 81750 0 -1 50850
box -180 -120 1680 4080
use INVX4  _947_
timestamp 1727136778
transform 1 0 85350 0 1 11850
box -180 -120 1380 4080
use NAND2X1  _948_
timestamp 1727136778
transform 1 0 79050 0 -1 43050
box -180 -120 1380 4080
use OAI21X1  _949_
timestamp 1727136778
transform 1 0 76950 0 -1 43050
box -180 -120 1680 4080
use INVX1  _950_
timestamp 1727136778
transform -1 0 70950 0 1 27450
box -180 -120 1080 4080
use INVX1  _951_
timestamp 1727136778
transform 1 0 58950 0 -1 27450
box -180 -120 1080 4080
use INVX2  _952_
timestamp 1727136778
transform 1 0 35550 0 1 50850
box -180 -120 1080 4080
use NOR2X1  _953_
timestamp 1727136778
transform 1 0 40050 0 -1 19650
box -180 -120 1380 4080
use AND2X2  _954_
timestamp 1727136778
transform -1 0 38850 0 1 19650
box -180 -120 1680 4095
use NAND2X1  _955_
timestamp 1727136778
transform 1 0 41850 0 1 11850
box -180 -120 1380 4080
use NAND2X1  _956_
timestamp 1727136778
transform 1 0 48150 0 1 27450
box -180 -120 1380 4080
use NAND2X1  _957_
timestamp 1727136778
transform 1 0 52650 0 -1 27450
box -180 -120 1380 4080
use OR2X2  _958_
timestamp 1727136778
transform 1 0 54750 0 -1 27450
box -180 -120 1680 4080
use NAND2X1  _959_
timestamp 1727136778
transform 1 0 54750 0 1 19650
box -180 -120 1380 4080
use AND2X2  _960_
timestamp 1727136778
transform 1 0 47850 0 1 19650
box -180 -120 1680 4095
use OAI21X1  _961_
timestamp 1727136778
transform -1 0 53850 0 1 19650
box -180 -120 1680 4080
use NAND2X1  _962_
timestamp 1727136778
transform 1 0 57150 0 -1 27450
box -180 -120 1380 4080
use INVX1  _963_
timestamp 1727136778
transform 1 0 44250 0 -1 19650
box -180 -120 1080 4080
use NAND2X1  _964_
timestamp 1727136778
transform -1 0 40950 0 1 27450
box -180 -120 1380 4080
use NAND2X1  _965_
timestamp 1727136778
transform 1 0 37950 0 1 27450
box -180 -120 1380 4080
use OR2X2  _966_
timestamp 1727136778
transform 1 0 50550 0 -1 27450
box -180 -120 1680 4080
use INVX1  _967_
timestamp 1727136778
transform -1 0 44850 0 1 27450
box -180 -120 1080 4080
use INVX1  _968_
timestamp 1727136778
transform 1 0 39150 0 1 50850
box -180 -120 1080 4080
use OAI21X1  _969_
timestamp 1727136778
transform -1 0 43350 0 1 27450
box -180 -120 1680 4080
use NAND3X1  _970_
timestamp 1727136778
transform 1 0 45750 0 -1 19650
box -180 -120 1680 4080
use NOR2X1  _971_
timestamp 1727136778
transform 1 0 46050 0 -1 27450
box -180 -120 1380 4080
use AND2X2  _972_
timestamp 1727136778
transform -1 0 49650 0 -1 27450
box -180 -120 1680 4095
use OAI21X1  _973_
timestamp 1727136778
transform 1 0 45750 0 1 19650
box -180 -120 1680 4080
use NAND3X1  _974_
timestamp 1727136778
transform -1 0 54150 0 1 11850
box -180 -120 1680 4080
use INVX1  _975_
timestamp 1727136778
transform 1 0 46350 0 1 11850
box -180 -120 1080 4080
use NAND2X1  _976_
timestamp 1727136778
transform 1 0 39450 0 1 19650
box -180 -120 1380 4080
use INVX2  _977_
timestamp 1727136778
transform 1 0 32250 0 1 58650
box -180 -120 1080 4080
use NAND2X1  _978_
timestamp 1727136778
transform 1 0 37950 0 -1 27450
box -180 -120 1380 4080
use OAI21X1  _979_
timestamp 1727136778
transform 1 0 31650 0 1 19650
box -180 -120 1680 4080
use OAI21X1  _980_
timestamp 1727136778
transform 1 0 43950 0 1 11850
box -180 -120 1680 4080
use AOI21X1  _981_
timestamp 1727136778
transform 1 0 55050 0 1 11850
box -180 -120 1680 4080
use OAI21X1  _982_
timestamp 1727136778
transform -1 0 53550 0 -1 11850
box -180 -120 1680 4080
use OAI21X1  _983_
timestamp 1727136778
transform -1 0 43050 0 1 19650
box -180 -120 1680 4080
use AND2X2  _984_
timestamp 1727136778
transform -1 0 38250 0 -1 35250
box -180 -120 1680 4095
use NAND3X1  _985_
timestamp 1727136778
transform -1 0 37050 0 1 27450
box -180 -120 1680 4080
use AOI22X1  _986_
timestamp 1727136778
transform -1 0 27750 0 -1 35250
box -210 -120 1980 4080
use INVX1  _987_
timestamp 1727136778
transform -1 0 25050 0 1 11850
box -180 -120 1080 4080
use NAND2X1  _988_
timestamp 1727136778
transform -1 0 22050 0 1 19650
box -180 -120 1380 4080
use INVX1  _989_
timestamp 1727136778
transform -1 0 28050 0 -1 19650
box -180 -120 1080 4080
use NAND3X1  _990_
timestamp 1727136778
transform 1 0 28350 0 1 11850
box -180 -120 1680 4080
use NAND2X1  _991_
timestamp 1727136778
transform 1 0 36450 0 1 58650
box -180 -120 1380 4080
use NOR2X1  _992_
timestamp 1727136778
transform -1 0 37050 0 -1 27450
box -180 -120 1380 4080
use OAI21X1  _993_
timestamp 1727136778
transform 1 0 30750 0 1 11850
box -180 -120 1680 4080
use NAND3X1  _994_
timestamp 1727136778
transform 1 0 39450 0 1 11850
box -180 -120 1680 4080
use AOI21X1  _995_
timestamp 1727136778
transform -1 0 43350 0 -1 19650
box -180 -120 1680 4080
use OAI21X1  _996_
timestamp 1727136778
transform 1 0 25950 0 1 11850
box -180 -120 1680 4080
use NAND3X1  _997_
timestamp 1727136778
transform -1 0 23250 0 1 11850
box -180 -120 1680 4080
use NAND3X1  _998_
timestamp 1727136778
transform 1 0 24450 0 -1 11850
box -180 -120 1680 4080
use NAND2X1  _999_
timestamp 1727136778
transform 1 0 33450 0 1 27450
box -180 -120 1380 4080
use INVX1  _1000_
timestamp 1727136778
transform 1 0 33750 0 1 19650
box -180 -120 1080 4080
use AND2X2  _1001_
timestamp 1727136778
transform 1 0 42150 0 -1 27450
box -180 -120 1680 4095
use NAND2X1  _1002_
timestamp 1727136778
transform 1 0 35550 0 1 19650
box -180 -120 1380 4080
use INVX1  _1003_
timestamp 1727136778
transform -1 0 45150 0 -1 27450
box -180 -120 1080 4080
use OAI21X1  _1004_
timestamp 1727136778
transform 1 0 37650 0 -1 19650
box -180 -120 1680 4080
use NAND3X1  _1005_
timestamp 1727136778
transform -1 0 36750 0 -1 19650
box -180 -120 1680 4080
use OAI21X1  _1006_
timestamp 1727136778
transform 1 0 30750 0 -1 19650
box -180 -120 1680 4080
use INVX1  _1007_
timestamp 1727136778
transform -1 0 26250 0 1 19650
box -180 -120 1080 4080
use OAI21X1  _1008_
timestamp 1727136778
transform 1 0 27150 0 1 19650
box -180 -120 1680 4080
use NAND3X1  _1009_
timestamp 1727136778
transform -1 0 31050 0 1 19650
box -180 -120 1680 4080
use AND2X2  _1010_
timestamp 1727136778
transform 1 0 34950 0 1 11850
box -180 -120 1680 4095
use NAND3X1  _1011_
timestamp 1727136778
transform -1 0 34950 0 -1 11850
box -180 -120 1680 4080
use AOI21X1  _1012_
timestamp 1727136778
transform -1 0 23850 0 -1 11850
box -180 -120 1680 4080
use AOI21X1  _1013_
timestamp 1727136778
transform -1 0 38550 0 1 11850
box -180 -120 1680 4080
use NAND2X1  _1014_
timestamp 1727136778
transform -1 0 34350 0 1 11850
box -180 -120 1380 4080
use OAI21X1  _1015_
timestamp 1727136778
transform -1 0 32550 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1016_
timestamp 1727136778
transform -1 0 32550 0 1 4050
box -180 -120 1680 4080
use AOI21X1  _1017_
timestamp 1727136778
transform 1 0 33450 0 1 4050
box -180 -120 1680 4080
use OAI21X1  _1018_
timestamp 1727136778
transform -1 0 37350 0 1 4050
box -180 -120 1680 4080
use AOI21X1  _1019_
timestamp 1727136778
transform -1 0 28050 0 -1 11850
box -180 -120 1680 4080
use OAI21X1  _1020_
timestamp 1727136778
transform -1 0 24450 0 1 19650
box -180 -120 1680 4080
use AND2X2  _1021_
timestamp 1727136778
transform -1 0 23250 0 1 58650
box -180 -120 1680 4095
use NAND2X1  _1022_
timestamp 1727136778
transform -1 0 22050 0 1 27450
box -180 -120 1380 4080
use INVX1  _1023_
timestamp 1727136778
transform 1 0 17550 0 1 35250
box -180 -120 1080 4080
use INVX2  _1024_
timestamp 1727136778
transform 1 0 22950 0 -1 74250
box -180 -120 1080 4080
use NAND2X1  _1025_
timestamp 1727136778
transform 1 0 22050 0 -1 35250
box -180 -120 1380 4080
use OAI21X1  _1026_
timestamp 1727136778
transform 1 0 19350 0 1 35250
box -180 -120 1680 4080
use NAND2X1  _1027_
timestamp 1727136778
transform 1 0 22950 0 1 27450
box -180 -120 1380 4080
use INVX1  _1028_
timestamp 1727136778
transform 1 0 16050 0 -1 27450
box -180 -120 1080 4080
use NAND3X1  _1029_
timestamp 1727136778
transform -1 0 15450 0 -1 27450
box -180 -120 1680 4080
use NOR2X1  _1030_
timestamp 1727136778
transform -1 0 25350 0 -1 35250
box -180 -120 1380 4080
use AOI22X1  _1031_
timestamp 1727136778
transform 1 0 19650 0 -1 35250
box -210 -120 1980 4080
use OAI21X1  _1032_
timestamp 1727136778
transform -1 0 20250 0 1 27450
box -180 -120 1680 4080
use AOI21X1  _1033_
timestamp 1727136778
transform -1 0 17850 0 1 19650
box -180 -120 1680 4080
use AOI21X1  _1034_
timestamp 1727136778
transform -1 0 26550 0 -1 19650
box -180 -120 1680 4080
use OAI21X1  _1035_
timestamp 1727136778
transform -1 0 17850 0 1 27450
box -180 -120 1680 4080
use NAND3X1  _1036_
timestamp 1727136778
transform -1 0 19350 0 -1 27450
box -180 -120 1680 4080
use AOI21X1  _1037_
timestamp 1727136778
transform -1 0 17550 0 -1 19650
box -180 -120 1680 4080
use NAND2X1  _1038_
timestamp 1727136778
transform 1 0 24750 0 1 27450
box -180 -120 1380 4080
use INVX1  _1039_
timestamp 1727136778
transform -1 0 21150 0 -1 27450
box -180 -120 1080 4080
use AND2X2  _1040_
timestamp 1727136778
transform -1 0 32550 0 1 27450
box -180 -120 1680 4095
use AND2X2  _1041_
timestamp 1727136778
transform -1 0 41250 0 -1 27450
box -180 -120 1680 4095
use NAND2X1  _1042_
timestamp 1727136778
transform 1 0 28950 0 1 27450
box -180 -120 1380 4080
use INVX2  _1043_
timestamp 1727136778
transform 1 0 34950 0 -1 35250
box -180 -120 1080 4080
use NAND2X1  _1044_
timestamp 1727136778
transform 1 0 34050 0 -1 27450
box -180 -120 1380 4080
use OAI21X1  _1045_
timestamp 1727136778
transform 1 0 31950 0 -1 27450
box -180 -120 1680 4080
use NAND3X1  _1046_
timestamp 1727136778
transform -1 0 25950 0 -1 27450
box -180 -120 1680 4080
use OAI21X1  _1047_
timestamp 1727136778
transform 1 0 26550 0 1 27450
box -180 -120 1680 4080
use OAI21X1  _1048_
timestamp 1727136778
transform -1 0 31050 0 -1 27450
box -180 -120 1680 4080
use NAND3X1  _1049_
timestamp 1727136778
transform -1 0 23550 0 -1 27450
box -180 -120 1680 4080
use AND2X2  _1050_
timestamp 1727136778
transform 1 0 22650 0 -1 19650
box -180 -120 1680 4095
use OAI21X1  _1051_
timestamp 1727136778
transform -1 0 12150 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1052_
timestamp 1727136778
transform 1 0 18450 0 -1 19650
box -180 -120 1680 4080
use NAND3X1  _1053_
timestamp 1727136778
transform 1 0 18450 0 1 19650
box -180 -120 1680 4080
use NAND2X1  _1054_
timestamp 1727136778
transform -1 0 22050 0 -1 19650
box -180 -120 1380 4080
use NAND3X1  _1055_
timestamp 1727136778
transform -1 0 16050 0 1 11850
box -180 -120 1680 4080
use NAND3X1  _1056_
timestamp 1727136778
transform 1 0 15450 0 -1 11850
box -180 -120 1680 4080
use OAI21X1  _1057_
timestamp 1727136778
transform -1 0 30150 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1058_
timestamp 1727136778
transform 1 0 19350 0 1 11850
box -180 -120 1680 4080
use OAI21X1  _1059_
timestamp 1727136778
transform 1 0 16950 0 1 11850
box -180 -120 1680 4080
use NAND3X1  _1060_
timestamp 1727136778
transform -1 0 19050 0 -1 11850
box -180 -120 1680 4080
use INVX4  _1061_
timestamp 1727136778
transform -1 0 45450 0 1 58650
box -180 -120 1380 4080
use NOR2X1  _1062_
timestamp 1727136778
transform -1 0 30150 0 -1 19650
box -180 -120 1380 4080
use OAI21X1  _1063_
timestamp 1727136778
transform 1 0 32850 0 -1 19650
box -180 -120 1680 4080
use XNOR2X1  _1064_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727153789
transform 1 0 21150 0 1 4050
box -180 -120 2280 4080
use INVX1  _1065_
timestamp 1727136778
transform -1 0 15150 0 -1 4050
box -180 -120 1080 4080
use NAND3X1  _1066_
timestamp 1727136778
transform 1 0 15750 0 -1 4050
box -180 -120 1680 4080
use AOI21X1  _1067_
timestamp 1727136778
transform 1 0 19950 0 -1 11850
box -180 -120 1680 4080
use AOI21X1  _1068_
timestamp 1727136778
transform -1 0 14550 0 -1 11850
box -180 -120 1680 4080
use OAI21X1  _1069_
timestamp 1727136778
transform 1 0 18750 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1070_
timestamp 1727136778
transform 1 0 29850 0 -1 4050
box -180 -120 1680 4080
use NAND2X1  _1071_
timestamp 1727136778
transform 1 0 24150 0 1 4050
box -180 -120 1380 4080
use INVX1  _1072_
timestamp 1727136778
transform -1 0 4050 0 -1 4050
box -180 -120 1080 4080
use OAI21X1  _1073_
timestamp 1727136778
transform -1 0 16050 0 1 4050
box -180 -120 1680 4080
use AOI21X1  _1074_
timestamp 1727136778
transform -1 0 13650 0 1 11850
box -180 -120 1680 4080
use OAI21X1  _1075_
timestamp 1727136778
transform -1 0 13350 0 1 27450
box -180 -120 1680 4080
use NAND3X1  _1076_
timestamp 1727136778
transform -1 0 16350 0 -1 35250
box -180 -120 1680 4080
use AOI22X1  _1077_
timestamp 1727136778
transform 1 0 17250 0 -1 35250
box -210 -120 1980 4080
use INVX1  _1078_
timestamp 1727136778
transform -1 0 8250 0 1 35250
box -180 -120 1080 4080
use NAND2X1  _1079_
timestamp 1727136778
transform -1 0 14850 0 1 35250
box -180 -120 1380 4080
use INVX1  _1080_
timestamp 1727136778
transform -1 0 13950 0 -1 35250
box -180 -120 1080 4080
use NAND3X1  _1081_
timestamp 1727136778
transform -1 0 4950 0 -1 35250
box -180 -120 1680 4080
use NAND2X1  _1082_
timestamp 1727136778
transform -1 0 16650 0 1 35250
box -180 -120 1380 4080
use NOR2X1  _1083_
timestamp 1727136778
transform -1 0 12750 0 1 35250
box -180 -120 1380 4080
use OAI21X1  _1084_
timestamp 1727136778
transform -1 0 7350 0 -1 35250
box -180 -120 1680 4080
use AOI21X1  _1085_
timestamp 1727136778
transform -1 0 6750 0 1 27450
box -180 -120 1680 4080
use OAI21X1  _1086_
timestamp 1727136778
transform 1 0 10650 0 -1 35250
box -180 -120 1680 4080
use NAND3X1  _1087_
timestamp 1727136778
transform 1 0 8250 0 -1 35250
box -180 -120 1680 4080
use AOI22X1  _1088_
timestamp 1727136778
transform -1 0 11250 0 -1 27450
box -210 -120 1980 4080
use NAND2X1  _1089_
timestamp 1727136778
transform 1 0 29850 0 -1 43050
box -180 -120 1380 4080
use INVX1  _1090_
timestamp 1727136778
transform 1 0 23850 0 -1 43050
box -180 -120 1080 4080
use AND2X2  _1091_
timestamp 1727136778
transform -1 0 29850 0 -1 35250
box -180 -120 1680 4095
use AND2X2  _1092_
timestamp 1727136778
transform -1 0 32250 0 1 35250
box -180 -120 1680 4095
use NAND2X1  _1093_
timestamp 1727136778
transform 1 0 28650 0 1 35250
box -180 -120 1380 4080
use AOI22X1  _1094_
timestamp 1727136778
transform 1 0 32850 0 1 50850
box -210 -120 1980 4080
use INVX1  _1095_
timestamp 1727136778
transform -1 0 28950 0 -1 43050
box -180 -120 1080 4080
use NAND3X1  _1096_
timestamp 1727136778
transform -1 0 27150 0 -1 43050
box -180 -120 1680 4080
use OAI21X1  _1097_
timestamp 1727136778
transform -1 0 25350 0 1 35250
box -180 -120 1680 4080
use OAI21X1  _1098_
timestamp 1727136778
transform -1 0 27750 0 1 35250
box -180 -120 1680 4080
use NAND3X1  _1099_
timestamp 1727136778
transform -1 0 23250 0 1 35250
box -180 -120 1680 4080
use AND2X2  _1100_
timestamp 1727136778
transform -1 0 2250 0 1 35250
box -180 -120 1680 4095
use OAI21X1  _1101_
timestamp 1727136778
transform -1 0 2550 0 -1 27450
box -180 -120 1680 4080
use AOI21X1  _1102_
timestamp 1727136778
transform -1 0 15750 0 1 27450
box -180 -120 1680 4080
use NAND3X1  _1103_
timestamp 1727136778
transform 1 0 9750 0 1 27450
box -180 -120 1680 4080
use NAND3X1  _1104_
timestamp 1727136778
transform 1 0 7350 0 1 27450
box -180 -120 1680 4080
use NAND2X1  _1105_
timestamp 1727136778
transform 1 0 3150 0 1 35250
box -180 -120 1380 4080
use NAND3X1  _1106_
timestamp 1727136778
transform -1 0 2550 0 1 27450
box -180 -120 1680 4080
use NAND3X1  _1107_
timestamp 1727136778
transform 1 0 3150 0 1 11850
box -180 -120 1680 4080
use OAI21X1  _1108_
timestamp 1727136778
transform 1 0 13650 0 -1 19650
box -180 -120 1680 4080
use NAND3X1  _1109_
timestamp 1727136778
transform -1 0 7050 0 -1 27450
box -180 -120 1680 4080
use OAI21X1  _1110_
timestamp 1727136778
transform -1 0 4650 0 -1 27450
box -180 -120 1680 4080
use NAND3X1  _1111_
timestamp 1727136778
transform -1 0 2550 0 1 19650
box -180 -120 1680 4080
use NAND2X1  _1112_
timestamp 1727136778
transform -1 0 31950 0 -1 35250
box -180 -120 1380 4080
use INVX1  _1113_
timestamp 1727136778
transform 1 0 7350 0 -1 19650
box -180 -120 1080 4080
use AOI22X1  _1114_
timestamp 1727136778
transform -1 0 28650 0 -1 27450
box -210 -120 1980 4080
use INVX1  _1115_
timestamp 1727136778
transform -1 0 8850 0 -1 27450
box -180 -120 1080 4080
use OAI21X1  _1116_
timestamp 1727136778
transform -1 0 10950 0 1 19650
box -180 -120 1680 4080
use NOR2X1  _1117_
timestamp 1727136778
transform 1 0 11850 0 1 19650
box -180 -120 1380 4080
use NAND2X1  _1118_
timestamp 1727136778
transform -1 0 6750 0 1 19650
box -180 -120 1380 4080
use NAND3X1  _1119_
timestamp 1727136778
transform 1 0 7650 0 1 11850
box -180 -120 1680 4080
use NAND2X1  _1120_
timestamp 1727136778
transform 1 0 7650 0 1 19650
box -180 -120 1380 4080
use OAI21X1  _1121_
timestamp 1727136778
transform 1 0 13950 0 1 19650
box -180 -120 1680 4080
use NAND3X1  _1122_
timestamp 1727136778
transform -1 0 12750 0 -1 19650
box -180 -120 1680 4080
use NAND2X1  _1123_
timestamp 1727136778
transform -1 0 11250 0 1 11850
box -180 -120 1380 4080
use NAND3X1  _1124_
timestamp 1727136778
transform 1 0 8250 0 -1 11850
box -180 -120 1680 4080
use AOI21X1  _1125_
timestamp 1727136778
transform 1 0 3150 0 1 19650
box -180 -120 1680 4080
use AOI21X1  _1126_
timestamp 1727136778
transform -1 0 2550 0 1 11850
box -180 -120 1680 4080
use NAND3X1  _1127_
timestamp 1727136778
transform 1 0 9150 0 -1 19650
box -180 -120 1680 4080
use NAND3X1  _1128_
timestamp 1727136778
transform -1 0 6750 0 -1 19650
box -180 -120 1680 4080
use NAND2X1  _1129_
timestamp 1727136778
transform -1 0 4350 0 -1 19650
box -180 -120 1380 4080
use OAI21X1  _1130_
timestamp 1727136778
transform 1 0 5850 0 -1 11850
box -180 -120 1680 4080
use AOI21X1  _1131_
timestamp 1727136778
transform -1 0 7050 0 1 4050
box -180 -120 1680 4080
use AOI21X1  _1132_
timestamp 1727136778
transform -1 0 13650 0 1 4050
box -180 -120 1680 4080
use OAI21X1  _1133_
timestamp 1727136778
transform -1 0 2550 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1134_
timestamp 1727136778
transform -1 0 4950 0 -1 11850
box -180 -120 1680 4080
use AOI21X1  _1135_
timestamp 1727136778
transform 1 0 3150 0 1 4050
box -180 -120 1680 4080
use OAI21X1  _1136_
timestamp 1727136778
transform -1 0 6450 0 -1 4050
box -180 -120 1680 4080
use NAND3X1  _1137_
timestamp 1727136778
transform -1 0 2550 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1138_
timestamp 1727136778
transform 1 0 7650 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1139_
timestamp 1727136778
transform 1 0 9450 0 -1 4050
box -180 -120 1680 4080
use AOI21X1  _1140_
timestamp 1727136778
transform 1 0 27450 0 -1 4050
box -180 -120 1680 4080
use INVX1  _1141_
timestamp 1727136778
transform 1 0 34350 0 -1 4050
box -180 -120 1080 4080
use INVX1  _1142_
timestamp 1727136778
transform 1 0 38250 0 1 4050
box -180 -120 1080 4080
use NOR2X1  _1143_
timestamp 1727136778
transform 1 0 50250 0 1 19650
box -180 -120 1380 4080
use INVX1  _1144_
timestamp 1727136778
transform 1 0 55050 0 -1 19650
box -180 -120 1080 4080
use OAI21X1  _1145_
timestamp 1727136778
transform 1 0 45750 0 1 27450
box -180 -120 1680 4080
use AOI21X1  _1146_
timestamp 1727136778
transform -1 0 52050 0 -1 19650
box -180 -120 1680 4080
use OAI21X1  _1147_
timestamp 1727136778
transform -1 0 45150 0 1 19650
box -180 -120 1680 4080
use NAND3X1  _1148_
timestamp 1727136778
transform 1 0 48150 0 -1 19650
box -180 -120 1680 4080
use AOI21X1  _1149_
timestamp 1727136778
transform -1 0 49650 0 1 11850
box -180 -120 1680 4080
use AND2X2  _1150_
timestamp 1727136778
transform 1 0 42750 0 -1 11850
box -180 -120 1680 4095
use NAND3X1  _1151_
timestamp 1727136778
transform 1 0 50250 0 1 11850
box -180 -120 1680 4080
use AOI21X1  _1152_
timestamp 1727136778
transform -1 0 49350 0 -1 11850
box -180 -120 1680 4080
use OAI21X1  _1153_
timestamp 1727136778
transform 1 0 35850 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1154_
timestamp 1727136778
transform 1 0 37950 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1155_
timestamp 1727136778
transform 1 0 40350 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1156_
timestamp 1727136778
transform -1 0 41550 0 1 4050
box -180 -120 1680 4080
use OAI21X1  _1157_
timestamp 1727136778
transform -1 0 18150 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1158_
timestamp 1727136778
transform 1 0 18150 0 -1 4050
box -180 -120 1680 4080
use AOI22X1  _1159_
timestamp 1727136778
transform -1 0 28050 0 1 4050
box -210 -120 1980 4080
use NAND3X1  _1160_
timestamp 1727136778
transform 1 0 7050 0 -1 4050
box -180 -120 1680 4080
use OAI21X1  _1161_
timestamp 1727136778
transform 1 0 11850 0 -1 4050
box -180 -120 1680 4080
use AOI21X1  _1162_
timestamp 1727136778
transform 1 0 20550 0 -1 4050
box -180 -120 1680 4080
use NAND3X1  _1163_
timestamp 1727136778
transform 1 0 49950 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1164_
timestamp 1727136778
transform 1 0 56850 0 -1 19650
box -180 -120 1680 4080
use NAND2X1  _1165_
timestamp 1727136778
transform -1 0 60150 0 1 27450
box -180 -120 1380 4080
use OR2X2  _1166_
timestamp 1727136778
transform 1 0 62550 0 -1 27450
box -180 -120 1680 4080
use NAND2X1  _1167_
timestamp 1727136778
transform 1 0 64950 0 -1 27450
box -180 -120 1380 4080
use AOI22X1  _1168_
timestamp 1727136778
transform -1 0 54150 0 1 27450
box -210 -120 1980 4080
use OAI21X1  _1169_
timestamp 1727136778
transform 1 0 60450 0 -1 27450
box -180 -120 1680 4080
use OAI21X1  _1170_
timestamp 1727136778
transform 1 0 52950 0 -1 19650
box -180 -120 1680 4080
use NAND3X1  _1171_
timestamp 1727136778
transform 1 0 61350 0 -1 19650
box -180 -120 1680 4080
use AOI21X1  _1172_
timestamp 1727136778
transform 1 0 58950 0 -1 19650
box -180 -120 1680 4080
use OAI21X1  _1173_
timestamp 1727136778
transform 1 0 61350 0 1 11850
box -180 -120 1680 4080
use OAI21X1  _1174_
timestamp 1727136778
transform 1 0 54450 0 -1 11850
box -180 -120 1680 4080
use NAND3X1  _1175_
timestamp 1727136778
transform -1 0 58350 0 -1 11850
box -180 -120 1680 4080
use INVX1  _1176_
timestamp 1727136778
transform 1 0 55050 0 1 4050
box -180 -120 1080 4080
use AOI22X1  _1177_
timestamp 1727136778
transform -1 0 46950 0 -1 11850
box -210 -120 1980 4080
use OAI21X1  _1178_
timestamp 1727136778
transform -1 0 46350 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1179_
timestamp 1727136778
transform 1 0 50550 0 1 4050
box -180 -120 1680 4080
use AOI21X1  _1180_
timestamp 1727136778
transform 1 0 32250 0 -1 4050
box -180 -120 1680 4080
use NOR3X1  _1181_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 49950 0 -1 4050
box -180 -120 2880 4095
use INVX1  _1182_
timestamp 1727136778
transform -1 0 60450 0 1 11850
box -180 -120 1080 4080
use NAND3X1  _1183_
timestamp 1727136778
transform 1 0 57450 0 1 11850
box -180 -120 1680 4080
use INVX1  _1184_
timestamp 1727136778
transform -1 0 55950 0 1 27450
box -180 -120 1080 4080
use OAI21X1  _1185_
timestamp 1727136778
transform -1 0 58050 0 1 27450
box -180 -120 1680 4080
use OR2X2  _1186_
timestamp 1727136778
transform 1 0 61050 0 1 19650
box -180 -120 1680 4080
use NAND2X1  _1187_
timestamp 1727136778
transform -1 0 51450 0 1 27450
box -180 -120 1380 4080
use NOR2X1  _1188_
timestamp 1727136778
transform -1 0 67950 0 -1 27450
box -180 -120 1380 4080
use INVX1  _1189_
timestamp 1727136778
transform 1 0 56850 0 1 19650
box -180 -120 1080 4080
use OAI21X1  _1190_
timestamp 1727136778
transform 1 0 58650 0 1 19650
box -180 -120 1680 4080
use NAND3X1  _1191_
timestamp 1727136778
transform -1 0 64650 0 1 19650
box -180 -120 1680 4080
use INVX1  _1192_
timestamp 1727136778
transform 1 0 67650 0 -1 19650
box -180 -120 1080 4080
use INVX1  _1193_
timestamp 1727136778
transform 1 0 65850 0 1 11850
box -180 -120 1080 4080
use OAI21X1  _1194_
timestamp 1727136778
transform 1 0 63450 0 1 11850
box -180 -120 1680 4080
use NAND3X1  _1195_
timestamp 1727136778
transform 1 0 67650 0 1 11850
box -180 -120 1680 4080
use AOI21X1  _1196_
timestamp 1727136778
transform 1 0 59250 0 -1 11850
box -180 -120 1680 4080
use NOR3X1  _1197_
timestamp 1727136778
transform -1 0 64350 0 -1 11850
box -180 -120 2880 4095
use OAI21X1  _1198_
timestamp 1727136778
transform 1 0 46950 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1199_
timestamp 1727136778
transform 1 0 42450 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1200_
timestamp 1727136778
transform 1 0 52950 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1201_
timestamp 1727136778
transform -1 0 58050 0 1 4050
box -180 -120 1680 4080
use INVX1  _1202_
timestamp 1727136778
transform 1 0 61350 0 1 4050
box -180 -120 1080 4080
use OAI21X1  _1203_
timestamp 1727136778
transform 1 0 53550 0 -1 4050
box -180 -120 1680 4080
use AOI21X1  _1204_
timestamp 1727136778
transform -1 0 57150 0 -1 4050
box -180 -120 1680 4080
use OAI21X1  _1205_
timestamp 1727136778
transform 1 0 40650 0 -1 4050
box -180 -120 1680 4080
use AOI21X1  _1206_
timestamp 1727136778
transform -1 0 2550 0 -1 4050
box -180 -120 1680 4080
use NAND2X1  _1207_
timestamp 1727136778
transform 1 0 11850 0 -1 27450
box -180 -120 1380 4080
use OAI21X1  _1208_
timestamp 1727136778
transform -1 0 2550 0 -1 19650
box -180 -120 1680 4080
use NAND2X1  _1209_
timestamp 1727136778
transform 1 0 36150 0 -1 50850
box -180 -120 1380 4080
use INVX1  _1210_
timestamp 1727136778
transform -1 0 24150 0 -1 50850
box -180 -120 1080 4080
use NOR2X1  _1211_
timestamp 1727136778
transform -1 0 34050 0 -1 35250
box -180 -120 1380 4080
use OAI21X1  _1212_
timestamp 1727136778
transform 1 0 28050 0 1 43050
box -180 -120 1680 4080
use NAND2X1  _1213_
timestamp 1727136778
transform 1 0 31650 0 -1 50850
box -180 -120 1380 4080
use OR2X2  _1214_
timestamp 1727136778
transform 1 0 33750 0 -1 50850
box -180 -120 1680 4080
use NAND3X1  _1215_
timestamp 1727136778
transform -1 0 22650 0 -1 50850
box -180 -120 1680 4080
use AND2X2  _1216_
timestamp 1727136778
transform -1 0 31050 0 -1 50850
box -180 -120 1680 4095
use NOR2X1  _1217_
timestamp 1727136778
transform 1 0 30450 0 1 43050
box -180 -120 1380 4080
use OAI21X1  _1218_
timestamp 1727136778
transform -1 0 28950 0 -1 50850
box -180 -120 1680 4080
use NAND2X1  _1219_
timestamp 1727136778
transform 1 0 19050 0 -1 50850
box -180 -120 1380 4080
use AOI21X1  _1220_
timestamp 1727136778
transform -1 0 4650 0 1 27450
box -180 -120 1680 4080
use NAND2X1  _1221_
timestamp 1727136778
transform -1 0 24450 0 -1 58650
box -180 -120 1380 4080
use AND2X2  _1222_
timestamp 1727136778
transform -1 0 30450 0 -1 66450
box -180 -120 1680 4095
use OAI21X1  _1223_
timestamp 1727136778
transform 1 0 27150 0 -1 58650
box -180 -120 1680 4080
use AND2X2  _1224_
timestamp 1727136778
transform -1 0 33450 0 -1 58650
box -180 -120 1680 4095
use OAI21X1  _1225_
timestamp 1727136778
transform 1 0 29550 0 -1 58650
box -180 -120 1680 4080
use NAND3X1  _1226_
timestamp 1727136778
transform -1 0 26550 0 -1 58650
box -180 -120 1680 4080
use INVX1  _1227_
timestamp 1727136778
transform 1 0 24150 0 1 58650
box -180 -120 1080 4080
use NAND2X1  _1228_
timestamp 1727136778
transform 1 0 30150 0 1 58650
box -180 -120 1380 4080
use AOI22X1  _1229_
timestamp 1727136778
transform 1 0 33750 0 1 58650
box -210 -120 1980 4080
use INVX1  _1230_
timestamp 1727136778
transform 1 0 28350 0 1 58650
box -180 -120 1080 4080
use NAND3X1  _1231_
timestamp 1727136778
transform -1 0 27450 0 1 58650
box -180 -120 1680 4080
use NAND2X1  _1232_
timestamp 1727136778
transform 1 0 11850 0 -1 58650
box -180 -120 1380 4080
use AOI21X1  _1233_
timestamp 1727136778
transform 1 0 5250 0 1 35250
box -180 -120 1680 4080
use NAND2X1  _1234_
timestamp 1727136778
transform 1 0 17250 0 -1 66450
box -180 -120 1380 4080
use XOR2X1  _1235_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727152697
transform 1 0 14250 0 1 58650
box -180 -120 2265 4080
use NAND2X1  _1236_
timestamp 1727136778
transform -1 0 5850 0 1 50850
box -180 -120 1380 4080
use OAI21X1  _1237_
timestamp 1727136778
transform 1 0 9150 0 1 35250
box -180 -120 1680 4080
use XNOR2X1  _1238_
timestamp 1727153789
transform 1 0 11550 0 1 58650
box -180 -120 2280 4080
use NAND2X1  _1239_
timestamp 1727136778
transform -1 0 9150 0 -1 58650
box -180 -120 1380 4080
use NAND3X1  _1240_
timestamp 1727136778
transform -1 0 8250 0 1 50850
box -180 -120 1680 4080
use AND2X2  _1241_
timestamp 1727136778
transform -1 0 4950 0 -1 58650
box -180 -120 1680 4095
use NAND2X1  _1242_
timestamp 1727136778
transform 1 0 10050 0 -1 58650
box -180 -120 1380 4080
use NAND2X1  _1243_
timestamp 1727136778
transform 1 0 5850 0 -1 58650
box -180 -120 1380 4080
use NAND3X1  _1244_
timestamp 1727136778
transform 1 0 3450 0 1 58650
box -180 -120 1680 4080
use NAND3X1  _1245_
timestamp 1727136778
transform -1 0 4650 0 -1 50850
box -180 -120 1680 4080
use OAI21X1  _1246_
timestamp 1727136778
transform -1 0 2550 0 -1 35250
box -180 -120 1680 4080
use AOI22X1  _1247_
timestamp 1727136778
transform -1 0 2850 0 -1 58650
box -210 -120 1980 4080
use AOI21X1  _1248_
timestamp 1727136778
transform 1 0 8850 0 1 50850
box -180 -120 1680 4080
use OAI21X1  _1249_
timestamp 1727136778
transform 1 0 1050 0 1 43050
box -180 -120 1680 4080
use NAND3X1  _1250_
timestamp 1727136778
transform -1 0 4950 0 1 43050
box -180 -120 1680 4080
use AND2X2  _1251_
timestamp 1727136778
transform -1 0 18150 0 -1 50850
box -180 -120 1680 4095
use NAND3X1  _1252_
timestamp 1727136778
transform 1 0 7650 0 -1 50850
box -180 -120 1680 4080
use OAI21X1  _1253_
timestamp 1727136778
transform 1 0 1050 0 -1 50850
box -180 -120 1680 4080
use NAND3X1  _1254_
timestamp 1727136778
transform -1 0 11250 0 -1 50850
box -180 -120 1680 4080
use NAND3X1  _1255_
timestamp 1727136778
transform -1 0 2550 0 -1 43050
box -180 -120 1680 4080
use AOI21X1  _1256_
timestamp 1727136778
transform 1 0 5550 0 1 11850
box -180 -120 1680 4080
use AOI22X1  _1257_
timestamp 1727136778
transform -1 0 16050 0 -1 50850
box -210 -120 1980 4080
use AOI21X1  _1258_
timestamp 1727136778
transform 1 0 5850 0 1 43050
box -180 -120 1680 4080
use OAI21X1  _1259_
timestamp 1727136778
transform -1 0 14250 0 1 43050
box -180 -120 1680 4080
use AOI21X1  _1260_
timestamp 1727136778
transform -1 0 13950 0 -1 43050
box -180 -120 1680 4080
use INVX1  _1261_
timestamp 1727136778
transform 1 0 14850 0 -1 43050
box -180 -120 1080 4080
use NAND3X1  _1262_
timestamp 1727136778
transform 1 0 3450 0 -1 43050
box -180 -120 1680 4080
use OAI21X1  _1263_
timestamp 1727136778
transform -1 0 11850 0 1 43050
box -180 -120 1680 4080
use AOI21X1  _1264_
timestamp 1727136778
transform 1 0 7950 0 -1 43050
box -180 -120 1680 4080
use OAI21X1  _1265_
timestamp 1727136778
transform -1 0 11850 0 -1 43050
box -180 -120 1680 4080
use OAI21X1  _1266_
timestamp 1727136778
transform -1 0 11550 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1267_
timestamp 1727136778
transform -1 0 7050 0 -1 43050
box -180 -120 1680 4080
use NAND3X1  _1268_
timestamp 1727136778
transform 1 0 16650 0 -1 43050
box -180 -120 1680 4080
use NAND3X1  _1269_
timestamp 1727136778
transform 1 0 19050 0 -1 43050
box -180 -120 1680 4080
use AND2X2  _1270_
timestamp 1727136778
transform 1 0 35550 0 -1 43050
box -180 -120 1680 4095
use XOR2X1  _1271_
timestamp 1727152697
transform -1 0 48750 0 -1 43050
box -180 -120 2265 4080
use NOR2X1  _1272_
timestamp 1727136778
transform 1 0 75450 0 -1 50850
box -180 -120 1380 4080
use NOR2X1  _1273_
timestamp 1727136778
transform -1 0 72450 0 -1 43050
box -180 -120 1380 4080
use OAI21X1  _1274_
timestamp 1727136778
transform 1 0 62850 0 -1 43050
box -180 -120 1680 4080
use AOI21X1  _1275_
timestamp 1727136778
transform 1 0 59850 0 1 35250
box -180 -120 1680 4080
use OAI21X1  _1276_
timestamp 1727136778
transform -1 0 68550 0 -1 43050
box -180 -120 1680 4080
use OAI21X1  _1277_
timestamp 1727136778
transform 1 0 62250 0 1 35250
box -180 -120 1680 4080
use NAND2X1  _1278_
timestamp 1727136778
transform 1 0 71850 0 1 27450
box -180 -120 1380 4080
use OAI21X1  _1279_
timestamp 1727136778
transform 1 0 70950 0 -1 27450
box -180 -120 1680 4080
use INVX1  _1280_
timestamp 1727136778
transform -1 0 54450 0 -1 35250
box -180 -120 1080 4080
use INVX1  _1281_
timestamp 1727136778
transform -1 0 58950 0 1 35250
box -180 -120 1080 4080
use OAI21X1  _1282_
timestamp 1727136778
transform -1 0 62550 0 -1 35250
box -180 -120 1680 4080
use OAI21X1  _1283_
timestamp 1727136778
transform -1 0 57150 0 1 35250
box -180 -120 1680 4080
use NAND3X1  _1284_
timestamp 1727136778
transform -1 0 26550 0 -1 4050
box -180 -120 1680 4080
use INVX1  _1285_
timestamp 1727136778
transform -1 0 49950 0 1 4050
box -180 -120 1080 4080
use NAND2X1  _1286_
timestamp 1727136778
transform -1 0 24150 0 -1 4050
box -180 -120 1380 4080
use NAND3X1  _1287_
timestamp 1727136778
transform 1 0 28950 0 1 4050
box -180 -120 1680 4080
use NAND3X1  _1288_
timestamp 1727136778
transform 1 0 45150 0 -1 4050
box -180 -120 1680 4080
use AOI21X1  _1289_
timestamp 1727136778
transform 1 0 43050 0 -1 4050
box -180 -120 1680 4080
use OAI21X1  _1290_
timestamp 1727136778
transform -1 0 49050 0 -1 4050
box -180 -120 1680 4080
use AOI21X1  _1291_
timestamp 1727136778
transform -1 0 37650 0 -1 4050
box -180 -120 1680 4080
use NAND2X1  _1292_
timestamp 1727136778
transform -1 0 34950 0 -1 43050
box -180 -120 1380 4080
use OAI21X1  _1293_
timestamp 1727136778
transform -1 0 41250 0 -1 43050
box -180 -120 1680 4080
use INVX1  _1294_
timestamp 1727136778
transform 1 0 19350 0 1 43050
box -180 -120 1080 4080
use AOI21X1  _1295_
timestamp 1727136778
transform 1 0 16950 0 1 43050
box -180 -120 1680 4080
use OAI21X1  _1296_
timestamp 1727136778
transform -1 0 26550 0 -1 50850
box -180 -120 1680 4080
use INVX1  _1297_
timestamp 1727136778
transform 1 0 24750 0 1 50850
box -180 -120 1080 4080
use AOI21X1  _1298_
timestamp 1727136778
transform 1 0 5250 0 -1 50850
box -180 -120 1680 4080
use OAI21X1  _1299_
timestamp 1727136778
transform 1 0 12150 0 -1 50850
box -180 -120 1680 4080
use NAND2X1  _1300_
timestamp 1727136778
transform -1 0 25650 0 -1 66450
box -180 -120 1380 4080
use NOR2X1  _1301_
timestamp 1727136778
transform 1 0 31050 0 1 50850
box -180 -120 1380 4080
use NAND2X1  _1302_
timestamp 1727136778
transform -1 0 30150 0 1 66450
box -180 -120 1380 4080
use NAND2X1  _1303_
timestamp 1727136778
transform -1 0 32550 0 -1 66450
box -180 -120 1380 4080
use OAI22X1  _1304_
timestamp 1727136778
transform -1 0 28050 0 -1 66450
box -180 -120 1980 4080
use XNOR2X1  _1305_
timestamp 1727153789
transform -1 0 23550 0 -1 66450
box -180 -120 2280 4080
use XNOR2X1  _1306_
timestamp 1727153789
transform 1 0 12150 0 -1 66450
box -180 -120 2280 4080
use NOR2X1  _1307_
timestamp 1727136778
transform 1 0 5550 0 1 58650
box -180 -120 1380 4080
use AOI21X1  _1308_
timestamp 1727136778
transform -1 0 2550 0 1 58650
box -180 -120 1680 4080
use NAND2X1  _1309_
timestamp 1727136778
transform 1 0 20250 0 1 66450
box -180 -120 1380 4080
use NAND2X1  _1310_
timestamp 1727136778
transform 1 0 24450 0 -1 74250
box -180 -120 1380 4080
use INVX1  _1311_
timestamp 1727136778
transform 1 0 16950 0 -1 74250
box -180 -120 1080 4080
use AND2X2  _1312_
timestamp 1727136778
transform -1 0 28050 0 -1 74250
box -180 -120 1680 4095
use AND2X2  _1313_
timestamp 1727136778
transform -1 0 22050 0 -1 74250
box -180 -120 1680 4095
use NAND2X1  _1314_
timestamp 1727136778
transform -1 0 19650 0 -1 74250
box -180 -120 1380 4080
use AOI22X1  _1315_
timestamp 1727136778
transform 1 0 19950 0 1 74250
box -210 -120 1980 4080
use INVX1  _1316_
timestamp 1727136778
transform -1 0 12750 0 1 74250
box -180 -120 1080 4080
use AOI21X1  _1317_
timestamp 1727136778
transform 1 0 14550 0 -1 74250
box -180 -120 1680 4080
use INVX2  _1318_
timestamp 1727136778
transform 1 0 42150 0 1 66450
box -180 -120 1080 4080
use OAI21X1  _1319_
timestamp 1727136778
transform -1 0 32550 0 1 66450
box -180 -120 1680 4080
use OAI21X1  _1320_
timestamp 1727136778
transform -1 0 28050 0 1 66450
box -180 -120 1680 4080
use AOI21X1  _1321_
timestamp 1727136778
transform -1 0 25950 0 1 66450
box -180 -120 1680 4080
use OAI22X1  _1322_
timestamp 1727136778
transform -1 0 19350 0 1 66450
box -180 -120 1980 4080
use NAND3X1  _1323_
timestamp 1727136778
transform -1 0 23550 0 1 66450
box -180 -120 1680 4080
use NAND3X1  _1324_
timestamp 1727136778
transform -1 0 13950 0 -1 74250
box -180 -120 1680 4080
use NOR2X1  _1325_
timestamp 1727136778
transform -1 0 16650 0 1 66450
box -180 -120 1380 4080
use NAND3X1  _1326_
timestamp 1727136778
transform -1 0 11550 0 -1 74250
box -180 -120 1680 4080
use NAND2X1  _1327_
timestamp 1727136778
transform -1 0 2250 0 -1 74250
box -180 -120 1380 4080
use NOR2X1  _1328_
timestamp 1727136778
transform -1 0 2250 0 -1 66450
box -180 -120 1380 4080
use NOR2X1  _1329_
timestamp 1727136778
transform 1 0 9750 0 1 58650
box -180 -120 1380 4080
use OAI21X1  _1330_
timestamp 1727136778
transform -1 0 9150 0 1 58650
box -180 -120 1680 4080
use AOI21X1  _1331_
timestamp 1727136778
transform 1 0 3150 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1332_
timestamp 1727136778
transform 1 0 7350 0 -1 66450
box -180 -120 1680 4080
use XOR2X1  _1333_
timestamp 1727152697
transform 1 0 12450 0 1 66450
box -180 -120 2265 4080
use NAND3X1  _1334_
timestamp 1727136778
transform 1 0 7950 0 -1 74250
box -180 -120 1680 4080
use NAND2X1  _1335_
timestamp 1727136778
transform -1 0 1950 0 1 66450
box -180 -120 1380 4080
use NAND3X1  _1336_
timestamp 1727136778
transform 1 0 7650 0 1 66450
box -180 -120 1680 4080
use NAND3X1  _1337_
timestamp 1727136778
transform 1 0 17250 0 1 58650
box -180 -120 1680 4080
use NOR3X1  _1338_
timestamp 1727136778
transform 1 0 1050 0 1 50850
box -180 -120 2880 4095
use AOI21X1  _1339_
timestamp 1727136778
transform 1 0 10950 0 1 50850
box -180 -120 1680 4080
use AOI21X1  _1340_
timestamp 1727136778
transform 1 0 10050 0 1 66450
box -180 -120 1680 4080
use NAND3X1  _1341_
timestamp 1727136778
transform 1 0 2850 0 1 66450
box -180 -120 1680 4080
use OAI21X1  _1342_
timestamp 1727136778
transform -1 0 4350 0 -1 66450
box -180 -120 1680 4080
use AOI21X1  _1343_
timestamp 1727136778
transform 1 0 5250 0 -1 66450
box -180 -120 1680 4080
use OAI21X1  _1344_
timestamp 1727136778
transform -1 0 14850 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1345_
timestamp 1727136778
transform -1 0 23850 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1346_
timestamp 1727136778
transform 1 0 13950 0 -1 58650
box -180 -120 1680 4080
use OAI21X1  _1347_
timestamp 1727136778
transform 1 0 15750 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1348_
timestamp 1727136778
transform -1 0 21750 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1349_
timestamp 1727136778
transform -1 0 22650 0 1 43050
box -180 -120 1680 4080
use AOI21X1  _1350_
timestamp 1727136778
transform 1 0 8250 0 1 43050
box -180 -120 1680 4080
use OAI21X1  _1351_
timestamp 1727136778
transform 1 0 14850 0 1 43050
box -180 -120 1680 4080
use NAND3X1  _1352_
timestamp 1727136778
transform 1 0 26550 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1353_
timestamp 1727136778
transform -1 0 19650 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1354_
timestamp 1727136778
transform 1 0 25650 0 1 43050
box -180 -120 1680 4080
use NAND2X1  _1355_
timestamp 1727136778
transform -1 0 33750 0 1 43050
box -180 -120 1380 4080
use AND2X2  _1356_
timestamp 1727136778
transform 1 0 49650 0 -1 43050
box -180 -120 1680 4095
use OAI21X1  _1357_
timestamp 1727136778
transform 1 0 51750 0 -1 43050
box -180 -120 1680 4080
use OAI21X1  _1358_
timestamp 1727136778
transform 1 0 54150 0 -1 43050
box -180 -120 1680 4080
use AND2X2  _1359_
timestamp 1727136778
transform 1 0 68850 0 -1 27450
box -180 -120 1680 4095
use NAND2X1  _1360_
timestamp 1727136778
transform 1 0 67950 0 1 27450
box -180 -120 1380 4080
use OAI21X1  _1361_
timestamp 1727136778
transform -1 0 64650 0 1 27450
box -180 -120 1680 4080
use OAI21X1  _1362_
timestamp 1727136778
transform 1 0 65550 0 1 27450
box -180 -120 1680 4080
use AOI21X1  _1363_
timestamp 1727136778
transform -1 0 62550 0 1 27450
box -180 -120 1680 4080
use AOI22X1  _1364_
timestamp 1727136778
transform 1 0 58650 0 -1 35250
box -210 -120 1980 4080
use OAI21X1  _1365_
timestamp 1727136778
transform -1 0 73950 0 1 19650
box -180 -120 1680 4080
use AOI21X1  _1366_
timestamp 1727136778
transform -1 0 25050 0 1 43050
box -180 -120 1680 4080
use AOI22X1  _1367_
timestamp 1727136778
transform 1 0 21150 0 -1 43050
box -210 -120 1980 4080
use NOR2X1  _1368_
timestamp 1727136778
transform 1 0 31950 0 -1 43050
box -180 -120 1380 4080
use NAND3X1  _1369_
timestamp 1727136778
transform 1 0 44250 0 -1 43050
box -180 -120 1680 4080
use AOI21X1  _1370_
timestamp 1727136778
transform 1 0 34350 0 1 43050
box -180 -120 1680 4080
use INVX1  _1371_
timestamp 1727136778
transform 1 0 37950 0 -1 43050
box -180 -120 1080 4080
use NAND2X1  _1372_
timestamp 1727136778
transform -1 0 20550 0 -1 66450
box -180 -120 1380 4080
use OAI21X1  _1373_
timestamp 1727136778
transform 1 0 14850 0 -1 66450
box -180 -120 1680 4080
use INVX1  _1374_
timestamp 1727136778
transform -1 0 8850 0 1 74250
box -180 -120 1080 4080
use AOI21X1  _1375_
timestamp 1727136778
transform -1 0 6750 0 1 66450
box -180 -120 1680 4080
use NAND2X1  _1376_
timestamp 1727136778
transform -1 0 20550 0 1 82050
box -180 -120 1380 4080
use INVX1  _1377_
timestamp 1727136778
transform -1 0 14250 0 1 82050
box -180 -120 1080 4080
use NOR2X1  _1378_
timestamp 1727136778
transform -1 0 19050 0 1 74250
box -180 -120 1380 4080
use OAI21X1  _1379_
timestamp 1727136778
transform -1 0 16950 0 1 74250
box -180 -120 1680 4080
use NAND2X1  _1380_
timestamp 1727136778
transform -1 0 18750 0 1 82050
box -180 -120 1380 4080
use OR2X2  _1381_
timestamp 1727136778
transform -1 0 16650 0 1 82050
box -180 -120 1680 4080
use NAND3X1  _1382_
timestamp 1727136778
transform -1 0 12450 0 1 82050
box -180 -120 1680 4080
use AND2X2  _1383_
timestamp 1727136778
transform -1 0 16650 0 -1 89850
box -180 -120 1680 4095
use NOR2X1  _1384_
timestamp 1727136778
transform -1 0 18750 0 -1 89850
box -180 -120 1380 4080
use OAI21X1  _1385_
timestamp 1727136778
transform -1 0 14250 0 -1 89850
box -180 -120 1680 4080
use NAND2X1  _1386_
timestamp 1727136778
transform -1 0 4650 0 -1 89850
box -180 -120 1380 4080
use OR2X2  _1387_
timestamp 1727136778
transform 1 0 9750 0 -1 66450
box -180 -120 1680 4080
use NAND2X1  _1388_
timestamp 1727136778
transform 1 0 24150 0 -1 82050
box -180 -120 1380 4080
use NAND2X1  _1389_
timestamp 1727136778
transform -1 0 28350 0 1 74250
box -180 -120 1380 4080
use NAND2X1  _1390_
timestamp 1727136778
transform -1 0 26550 0 1 74250
box -180 -120 1380 4080
use AOI22X1  _1391_
timestamp 1727136778
transform -1 0 24450 0 1 74250
box -210 -120 1980 4080
use INVX1  _1392_
timestamp 1727136778
transform 1 0 30750 0 -1 82050
box -180 -120 1080 4080
use OAI21X1  _1393_
timestamp 1727136778
transform 1 0 28650 0 -1 82050
box -180 -120 1680 4080
use XNOR2X1  _1394_
timestamp 1727153789
transform 1 0 21150 0 -1 82050
box -180 -120 2280 4080
use AOI21X1  _1395_
timestamp 1727136778
transform 1 0 6450 0 1 82050
box -180 -120 1680 4080
use NAND3X1  _1396_
timestamp 1727136778
transform -1 0 10350 0 1 82050
box -180 -120 1680 4080
use INVX1  _1397_
timestamp 1727136778
transform -1 0 1950 0 1 89850
box -180 -120 1080 4080
use OAI21X1  _1398_
timestamp 1727136778
transform -1 0 6450 0 1 89850
box -180 -120 1680 4080
use AND2X2  _1399_
timestamp 1727136778
transform -1 0 11850 0 -1 89850
box -180 -120 1680 4095
use NAND2X1  _1400_
timestamp 1727136778
transform -1 0 5850 0 1 82050
box -180 -120 1380 4080
use INVX1  _1401_
timestamp 1727136778
transform -1 0 1650 0 1 82050
box -180 -120 1080 4080
use NAND2X1  _1402_
timestamp 1727136778
transform -1 0 3750 0 1 82050
box -180 -120 1380 4080
use NAND3X1  _1403_
timestamp 1727136778
transform 1 0 5550 0 -1 89850
box -180 -120 1680 4080
use NAND3X1  _1404_
timestamp 1727136778
transform -1 0 8850 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1405_
timestamp 1727136778
transform 1 0 5550 0 -1 74250
box -180 -120 1680 4080
use AOI22X1  _1406_
timestamp 1727136778
transform -1 0 2850 0 -1 89850
box -210 -120 1980 4080
use OR2X2  _1407_
timestamp 1727136778
transform -1 0 2550 0 -1 82050
box -180 -120 1680 4080
use NAND2X1  _1408_
timestamp 1727136778
transform -1 0 6750 0 -1 82050
box -180 -120 1380 4080
use AOI21X1  _1409_
timestamp 1727136778
transform -1 0 4950 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1410_
timestamp 1727136778
transform 1 0 3450 0 1 74250
box -180 -120 1680 4080
use NAND3X1  _1411_
timestamp 1727136778
transform -1 0 7050 0 1 74250
box -180 -120 1680 4080
use NAND3X1  _1412_
timestamp 1727136778
transform 1 0 9750 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1413_
timestamp 1727136778
transform -1 0 2550 0 1 74250
box -180 -120 1680 4080
use NAND3X1  _1414_
timestamp 1727136778
transform -1 0 10950 0 1 74250
box -180 -120 1680 4080
use NAND2X1  _1415_
timestamp 1727136778
transform -1 0 20850 0 1 58650
box -180 -120 1380 4080
use NAND3X1  _1416_
timestamp 1727136778
transform 1 0 28950 0 1 50850
box -180 -120 1680 4080
use AOI21X1  _1417_
timestamp 1727136778
transform 1 0 16050 0 -1 58650
box -180 -120 1680 4080
use OAI21X1  _1418_
timestamp 1727136778
transform -1 0 19950 0 -1 58650
box -180 -120 1680 4080
use NAND3X1  _1419_
timestamp 1727136778
transform 1 0 20850 0 -1 58650
box -180 -120 1680 4080
use NAND2X1  _1420_
timestamp 1727136778
transform -1 0 38250 0 1 50850
box -180 -120 1380 4080
use AOI21X1  _1421_
timestamp 1727136778
transform -1 0 38550 0 1 35250
box -180 -120 1680 4080
use NAND2X1  _1422_
timestamp 1727136778
transform 1 0 42150 0 -1 43050
box -180 -120 1380 4080
use OAI21X1  _1423_
timestamp 1727136778
transform -1 0 40650 0 1 35250
box -180 -120 1680 4080
use INVX1  _1424_
timestamp 1727136778
transform 1 0 43350 0 -1 35250
box -180 -120 1080 4080
use NOR2X1  _1425_
timestamp 1727136778
transform -1 0 46350 0 -1 35250
box -180 -120 1380 4080
use OAI21X1  _1426_
timestamp 1727136778
transform 1 0 46950 0 -1 35250
box -180 -120 1680 4080
use NOR2X1  _1427_
timestamp 1727136778
transform 1 0 69450 0 -1 43050
box -180 -120 1380 4080
use NOR2X1  _1428_
timestamp 1727136778
transform -1 0 65850 0 1 35250
box -180 -120 1380 4080
use AOI21X1  _1429_
timestamp 1727136778
transform 1 0 65550 0 1 19650
box -180 -120 1680 4080
use OAI21X1  _1430_
timestamp 1727136778
transform 1 0 67650 0 1 19650
box -180 -120 1680 4080
use NOR2X1  _1431_
timestamp 1727136778
transform -1 0 72150 0 1 35250
box -180 -120 1380 4080
use NOR2X1  _1432_
timestamp 1727136778
transform 1 0 71550 0 -1 35250
box -180 -120 1380 4080
use AOI22X1  _1433_
timestamp 1727136778
transform -1 0 67050 0 -1 35250
box -210 -120 1980 4080
use OAI21X1  _1434_
timestamp 1727136778
transform 1 0 70050 0 1 19650
box -180 -120 1680 4080
use INVX1  _1435_
timestamp 1727136778
transform 1 0 89550 0 -1 11850
box -180 -120 1080 4080
use INVX1  _1436_
timestamp 1727136778
transform -1 0 87450 0 1 43050
box -180 -120 1080 4080
use OAI21X1  _1437_
timestamp 1727136778
transform -1 0 59850 0 -1 43050
box -180 -120 1680 4080
use INVX1  _1438_
timestamp 1727136778
transform 1 0 40350 0 -1 50850
box -180 -120 1080 4080
use OAI21X1  _1439_
timestamp 1727136778
transform 1 0 19350 0 -1 89850
box -180 -120 1680 4080
use INVX1  _1440_
timestamp 1727136778
transform -1 0 19050 0 1 89850
box -180 -120 1080 4080
use AOI21X1  _1441_
timestamp 1727136778
transform 1 0 7950 0 -1 89850
box -180 -120 1680 4080
use NAND2X1  _1442_
timestamp 1727136778
transform 1 0 27450 0 1 82050
box -180 -120 1380 4080
use INVX1  _1443_
timestamp 1727136778
transform -1 0 32250 0 -1 89850
box -180 -120 1080 4080
use NOR2X1  _1444_
timestamp 1727136778
transform -1 0 22650 0 1 82050
box -180 -120 1380 4080
use OAI22X1  _1445_
timestamp 1727136778
transform -1 0 27750 0 -1 82050
box -180 -120 1980 4080
use NAND2X1  _1446_
timestamp 1727136778
transform 1 0 23550 0 1 82050
box -180 -120 1380 4080
use NOR2X1  _1447_
timestamp 1727136778
transform 1 0 25650 0 1 82050
box -180 -120 1380 4080
use INVX1  _1448_
timestamp 1727136778
transform 1 0 27150 0 -1 89850
box -180 -120 1080 4080
use NAND3X1  _1449_
timestamp 1727136778
transform -1 0 30450 0 -1 89850
box -180 -120 1680 4080
use INVX1  _1450_
timestamp 1727136778
transform -1 0 24450 0 -1 89850
box -180 -120 1080 4080
use OAI21X1  _1451_
timestamp 1727136778
transform 1 0 25050 0 -1 89850
box -180 -120 1680 4080
use NAND2X1  _1452_
timestamp 1727136778
transform 1 0 28950 0 -1 74250
box -180 -120 1380 4080
use NAND2X1  _1453_
timestamp 1727136778
transform 1 0 31650 0 1 74250
box -180 -120 1380 4080
use OR2X2  _1454_
timestamp 1727136778
transform 1 0 29250 0 1 74250
box -180 -120 1680 4080
use INVX1  _1455_
timestamp 1727136778
transform 1 0 43350 0 -1 82050
box -180 -120 1080 4080
use OAI21X1  _1456_
timestamp 1727136778
transform -1 0 34050 0 -1 82050
box -180 -120 1680 4080
use AND2X2  _1457_
timestamp 1727136778
transform -1 0 31050 0 1 82050
box -180 -120 1680 4095
use AOI21X1  _1458_
timestamp 1727136778
transform -1 0 25650 0 1 89850
box -180 -120 1680 4080
use INVX1  _1459_
timestamp 1727136778
transform -1 0 8250 0 1 89850
box -180 -120 1080 4080
use NAND3X1  _1460_
timestamp 1727136778
transform 1 0 26550 0 1 89850
box -180 -120 1680 4080
use NAND3X1  _1461_
timestamp 1727136778
transform 1 0 11250 0 1 89850
box -180 -120 1680 4080
use OAI21X1  _1462_
timestamp 1727136778
transform -1 0 4350 0 1 89850
box -180 -120 1680 4080
use INVX1  _1463_
timestamp 1727136778
transform -1 0 22650 0 -1 89850
box -180 -120 1080 4080
use OAI21X1  _1464_
timestamp 1727136778
transform -1 0 14850 0 1 89850
box -180 -120 1680 4080
use NAND3X1  _1465_
timestamp 1727136778
transform -1 0 17250 0 1 89850
box -180 -120 1680 4080
use NAND3X1  _1466_
timestamp 1727136778
transform -1 0 10650 0 1 89850
box -180 -120 1680 4080
use OAI21X1  _1467_
timestamp 1727136778
transform -1 0 21150 0 1 89850
box -180 -120 1680 4080
use NAND3X1  _1468_
timestamp 1727136778
transform 1 0 22050 0 1 89850
box -180 -120 1680 4080
use NAND2X1  _1469_
timestamp 1727136778
transform -1 0 18150 0 -1 82050
box -180 -120 1380 4080
use NAND3X1  _1470_
timestamp 1727136778
transform -1 0 14850 0 1 74250
box -180 -120 1680 4080
use AOI21X1  _1471_
timestamp 1727136778
transform 1 0 12150 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1472_
timestamp 1727136778
transform 1 0 14550 0 -1 82050
box -180 -120 1680 4080
use NAND3X1  _1473_
timestamp 1727136778
transform 1 0 18750 0 -1 82050
box -180 -120 1680 4080
use NAND2X1  _1474_
timestamp 1727136778
transform 1 0 42150 0 -1 50850
box -180 -120 1380 4080
use NOR3X1  _1475_
timestamp 1727136778
transform 1 0 41550 0 1 35250
box -180 -120 2880 4095
use AOI21X1  _1476_
timestamp 1727136778
transform 1 0 45150 0 1 35250
box -180 -120 1680 4080
use INVX1  _1477_
timestamp 1727136778
transform 1 0 47250 0 1 35250
box -180 -120 1080 4080
use OAI21X1  _1478_
timestamp 1727136778
transform 1 0 49050 0 1 35250
box -180 -120 1680 4080
use OAI21X1  _1479_
timestamp 1727136778
transform 1 0 53250 0 1 35250
box -180 -120 1680 4080
use NAND2X1  _1480_
timestamp 1727136778
transform -1 0 64650 0 -1 19650
box -180 -120 1380 4080
use NAND2X1  _1481_
timestamp 1727136778
transform -1 0 66750 0 -1 19650
box -180 -120 1380 4080
use NAND2X1  _1482_
timestamp 1727136778
transform 1 0 70050 0 1 11850
box -180 -120 1380 4080
use NAND2X1  _1483_
timestamp 1727136778
transform 1 0 80850 0 1 11850
box -180 -120 1380 4080
use OAI21X1  _1484_
timestamp 1727136778
transform -1 0 84450 0 1 11850
box -180 -120 1680 4080
use AOI21X1  _1485_
timestamp 1727136778
transform 1 0 82950 0 -1 11850
box -180 -120 1680 4080
use AOI22X1  _1486_
timestamp 1727136778
transform -1 0 86850 0 -1 11850
box -210 -120 1980 4080
use INVX1  _1487_
timestamp 1727136778
transform 1 0 87750 0 -1 11850
box -180 -120 1080 4080
use OAI21X1  _1488_
timestamp 1727136778
transform 1 0 33150 0 -1 89850
box -180 -120 1680 4080
use INVX1  _1489_
timestamp 1727136778
transform 1 0 35250 0 -1 89850
box -180 -120 1080 4080
use INVX1  _1490_
timestamp 1727136778
transform -1 0 36450 0 1 74250
box -180 -120 1080 4080
use NAND2X1  _1491_
timestamp 1727136778
transform -1 0 44550 0 1 82050
box -180 -120 1380 4080
use OAI21X1  _1492_
timestamp 1727136778
transform -1 0 33150 0 1 82050
box -180 -120 1680 4080
use OAI21X1  _1493_
timestamp 1727136778
transform -1 0 35550 0 1 82050
box -180 -120 1680 4080
use OR2X2  _1494_
timestamp 1727136778
transform 1 0 38850 0 1 82050
box -180 -120 1680 4080
use INVX1  _1495_
timestamp 1727136778
transform 1 0 44850 0 -1 82050
box -180 -120 1080 4080
use OAI21X1  _1496_
timestamp 1727136778
transform 1 0 36450 0 1 82050
box -180 -120 1680 4080
use NAND2X1  _1497_
timestamp 1727136778
transform 1 0 39450 0 -1 82050
box -180 -120 1380 4080
use OAI21X1  _1498_
timestamp 1727136778
transform 1 0 41250 0 -1 82050
box -180 -120 1680 4080
use INVX1  _1499_
timestamp 1727136778
transform 1 0 33750 0 1 74250
box -180 -120 1080 4080
use NAND3X1  _1500_
timestamp 1727136778
transform 1 0 37050 0 -1 82050
box -180 -120 1680 4080
use NAND2X1  _1501_
timestamp 1727136778
transform 1 0 41250 0 1 82050
box -180 -120 1380 4080
use NOR2X1  _1502_
timestamp 1727136778
transform 1 0 41250 0 -1 89850
box -180 -120 1380 4080
use NAND2X1  _1503_
timestamp 1727136778
transform 1 0 42150 0 1 89850
box -180 -120 1380 4080
use INVX1  _1504_
timestamp 1727136778
transform 1 0 43350 0 -1 89850
box -180 -120 1080 4080
use OAI21X1  _1505_
timestamp 1727136778
transform -1 0 38250 0 -1 89850
box -180 -120 1680 4080
use OR2X2  _1506_
timestamp 1727136778
transform -1 0 41250 0 1 89850
box -180 -120 1680 4080
use NAND3X1  _1507_
timestamp 1727136778
transform -1 0 38850 0 1 89850
box -180 -120 1680 4080
use NAND2X1  _1508_
timestamp 1727136778
transform -1 0 34350 0 1 89850
box -180 -120 1380 4080
use NAND3X1  _1509_
timestamp 1727136778
transform 1 0 31050 0 1 89850
box -180 -120 1680 4080
use NAND2X1  _1510_
timestamp 1727136778
transform -1 0 30150 0 1 89850
box -180 -120 1380 4080
use NAND3X1  _1511_
timestamp 1727136778
transform 1 0 34950 0 1 89850
box -180 -120 1680 4080
use NAND2X1  _1512_
timestamp 1727136778
transform -1 0 42150 0 1 50850
box -180 -120 1380 4080
use NOR2X1  _1513_
timestamp 1727136778
transform 1 0 50250 0 1 43050
box -180 -120 1380 4080
use NOR2X1  _1514_
timestamp 1727136778
transform -1 0 46950 0 1 43050
box -180 -120 1380 4080
use NAND3X1  _1515_
timestamp 1727136778
transform 1 0 47850 0 1 43050
box -180 -120 1680 4080
use NAND2X1  _1516_
timestamp 1727136778
transform -1 0 39450 0 -1 50850
box -180 -120 1380 4080
use AOI22X1  _1517_
timestamp 1727136778
transform 1 0 43350 0 1 43050
box -210 -120 1980 4080
use AOI21X1  _1518_
timestamp 1727136778
transform -1 0 49950 0 -1 50850
box -180 -120 1680 4080
use NAND2X1  _1519_
timestamp 1727136778
transform 1 0 44250 0 -1 50850
box -180 -120 1380 4080
use OAI21X1  _1520_
timestamp 1727136778
transform 1 0 46050 0 -1 50850
box -180 -120 1680 4080
use AOI21X1  _1521_
timestamp 1727136778
transform 1 0 38850 0 1 43050
box -180 -120 1680 4080
use OAI21X1  _1522_
timestamp 1727136778
transform 1 0 41250 0 1 43050
box -180 -120 1680 4080
use AOI22X1  _1523_
timestamp 1727136778
transform 1 0 43050 0 1 50850
box -210 -120 1980 4080
use OAI21X1  _1524_
timestamp 1727136778
transform 1 0 49650 0 1 50850
box -180 -120 1680 4080
use OR2X2  _1525_
timestamp 1727136778
transform -1 0 83850 0 1 43050
box -180 -120 1680 4080
use NAND3X1  _1526_
timestamp 1727136778
transform -1 0 76350 0 1 35250
box -180 -120 1680 4080
use INVX1  _1527_
timestamp 1727136778
transform 1 0 67350 0 -1 11850
box -180 -120 1080 4080
use OAI21X1  _1528_
timestamp 1727136778
transform 1 0 65250 0 -1 11850
box -180 -120 1680 4080
use NAND2X1  _1529_
timestamp 1727136778
transform 1 0 69150 0 -1 11850
box -180 -120 1380 4080
use NAND2X1  _1530_
timestamp 1727136778
transform -1 0 73950 0 1 35250
box -180 -120 1380 4080
use OAI21X1  _1531_
timestamp 1727136778
transform -1 0 77850 0 1 11850
box -180 -120 1680 4080
use AOI21X1  _1532_
timestamp 1727136778
transform 1 0 78750 0 1 11850
box -180 -120 1680 4080
use AOI22X1  _1533_
timestamp 1727136778
transform -1 0 82050 0 -1 11850
box -210 -120 1980 4080
use INVX1  _1534_
timestamp 1727136778
transform -1 0 78450 0 1 4050
box -180 -120 1080 4080
use INVX1  _1535_
timestamp 1727136778
transform -1 0 57450 0 -1 43050
box -180 -120 1080 4080
use NAND2X1  _1536_
timestamp 1727136778
transform 1 0 47850 0 1 50850
box -180 -120 1380 4080
use INVX1  _1537_
timestamp 1727136778
transform 1 0 42450 0 1 58650
box -180 -120 1080 4080
use AOI21X1  _1538_
timestamp 1727136778
transform 1 0 39150 0 -1 89850
box -180 -120 1680 4080
use OAI21X1  _1539_
timestamp 1727136778
transform 1 0 34650 0 -1 82050
box -180 -120 1680 4080
use NOR2X1  _1540_
timestamp 1727136778
transform -1 0 40950 0 1 74250
box -180 -120 1380 4080
use NAND3X1  _1541_
timestamp 1727136778
transform -1 0 43650 0 -1 74250
box -180 -120 1680 4080
use OAI22X1  _1542_
timestamp 1727136778
transform -1 0 38850 0 1 74250
box -180 -120 1980 4080
use NAND2X1  _1543_
timestamp 1727136778
transform 1 0 40050 0 -1 74250
box -180 -120 1380 4080
use XNOR2X1  _1544_
timestamp 1727153789
transform 1 0 37050 0 -1 74250
box -180 -120 2280 4080
use XOR2X1  _1545_
timestamp 1727152697
transform -1 0 39150 0 1 66450
box -180 -120 2265 4080
use XOR2X1  _1546_
timestamp 1727152697
transform -1 0 39750 0 -1 66450
box -180 -120 2265 4080
use NOR2X1  _1547_
timestamp 1727136778
transform -1 0 41550 0 -1 58650
box -180 -120 1380 4080
use OAI21X1  _1548_
timestamp 1727136778
transform -1 0 47250 0 1 50850
box -180 -120 1680 4080
use OAI21X1  _1549_
timestamp 1727136778
transform -1 0 43650 0 -1 58650
box -180 -120 1680 4080
use NAND3X1  _1550_
timestamp 1727136778
transform 1 0 52350 0 1 43050
box -180 -120 1680 4080
use AOI21X1  _1551_
timestamp 1727136778
transform 1 0 58950 0 1 4050
box -180 -120 1680 4080
use OAI21X1  _1552_
timestamp 1727136778
transform 1 0 62850 0 1 4050
box -180 -120 1680 4080
use INVX1  _1553_
timestamp 1727136778
transform -1 0 76950 0 1 27450
box -180 -120 1080 4080
use AOI21X1  _1554_
timestamp 1727136778
transform 1 0 78750 0 -1 19650
box -180 -120 1680 4080
use AOI21X1  _1555_
timestamp 1727136778
transform 1 0 78150 0 -1 11850
box -180 -120 1680 4080
use AOI22X1  _1556_
timestamp 1727136778
transform -1 0 76650 0 1 4050
box -210 -120 1980 4080
use INVX1  _1557_
timestamp 1727136778
transform -1 0 73950 0 1 4050
box -180 -120 1080 4080
use NAND3X1  _1558_
timestamp 1727136778
transform 1 0 37950 0 -1 58650
box -180 -120 1680 4080
use INVX1  _1559_
timestamp 1727136778
transform 1 0 53250 0 -1 50850
box -180 -120 1080 4080
use NAND3X1  _1560_
timestamp 1727136778
transform 1 0 55050 0 -1 50850
box -180 -120 1680 4080
use NAND2X1  _1561_
timestamp 1727136778
transform -1 0 41550 0 1 58650
box -180 -120 1380 4080
use OAI21X1  _1562_
timestamp 1727136778
transform 1 0 40650 0 -1 66450
box -180 -120 1680 4080
use INVX1  _1563_
timestamp 1727136778
transform 1 0 55950 0 1 50850
box -180 -120 1080 4080
use INVX1  _1564_
timestamp 1727136778
transform -1 0 31650 0 -1 74250
box -180 -120 1080 4080
use NAND2X1  _1565_
timestamp 1727136778
transform -1 0 33750 0 -1 74250
box -180 -120 1380 4080
use OAI21X1  _1566_
timestamp 1727136778
transform -1 0 36150 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1567_
timestamp 1727136778
transform 1 0 43650 0 1 66450
box -180 -120 1680 4080
use XOR2X1  _1568_
timestamp 1727152697
transform 1 0 50250 0 1 66450
box -180 -120 2265 4080
use NAND3X1  _1569_
timestamp 1727136778
transform 1 0 59550 0 -1 50850
box -180 -120 1680 4080
use AOI21X1  _1570_
timestamp 1727136778
transform 1 0 50850 0 -1 50850
box -180 -120 1680 4080
use INVX1  _1571_
timestamp 1727136778
transform -1 0 55050 0 1 50850
box -180 -120 1080 4080
use OAI21X1  _1572_
timestamp 1727136778
transform 1 0 52050 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1573_
timestamp 1727136778
transform 1 0 61950 0 -1 50850
box -180 -120 1680 4080
use NAND2X1  _1574_
timestamp 1727136778
transform -1 0 61950 0 -1 4050
box -180 -120 1380 4080
use NOR2X1  _1575_
timestamp 1727136778
transform 1 0 65250 0 -1 4050
box -180 -120 1380 4080
use AOI21X1  _1576_
timestamp 1727136778
transform 1 0 62850 0 -1 4050
box -180 -120 1680 4080
use OAI21X1  _1577_
timestamp 1727136778
transform 1 0 67050 0 -1 4050
box -180 -120 1680 4080
use NOR2X1  _1578_
timestamp 1727136778
transform 1 0 85950 0 -1 50850
box -180 -120 1380 4080
use NOR2X1  _1579_
timestamp 1727136778
transform -1 0 78150 0 -1 35250
box -180 -120 1380 4080
use AOI21X1  _1580_
timestamp 1727136778
transform -1 0 77550 0 -1 11850
box -180 -120 1680 4080
use AOI22X1  _1581_
timestamp 1727136778
transform 1 0 73650 0 -1 11850
box -210 -120 1980 4080
use INVX1  _1582_
timestamp 1727136778
transform -1 0 68550 0 1 4050
box -180 -120 1080 4080
use AOI21X1  _1583_
timestamp 1727136778
transform -1 0 58650 0 -1 50850
box -180 -120 1680 4080
use NAND3X1  _1584_
timestamp 1727136778
transform 1 0 44550 0 -1 74250
box -180 -120 1680 4080
use NAND2X1  _1585_
timestamp 1727136778
transform 1 0 46950 0 -1 74250
box -180 -120 1380 4080
use OAI21X1  _1586_
timestamp 1727136778
transform 1 0 54450 0 1 43050
box -180 -120 1680 4080
use NAND2X1  _1587_
timestamp 1727136778
transform 1 0 38550 0 -1 4050
box -180 -120 1380 4080
use XNOR2X1  _1588_
timestamp 1727153789
transform -1 0 60150 0 -1 4050
box -180 -120 2280 4080
use NAND2X1  _1589_
timestamp 1727136778
transform 1 0 74250 0 1 11850
box -180 -120 1380 4080
use OAI21X1  _1590_
timestamp 1727136778
transform 1 0 72150 0 1 11850
box -180 -120 1680 4080
use AOI21X1  _1591_
timestamp 1727136778
transform -1 0 72750 0 -1 11850
box -180 -120 1680 4080
use AOI22X1  _1592_
timestamp 1727136778
transform -1 0 66750 0 1 4050
box -210 -120 1980 4080
use NAND2X1  _1593_
timestamp 1727136778
transform -1 0 66450 0 -1 43050
box -180 -120 1380 4080
use OAI21X1  _1594_
timestamp 1727136778
transform 1 0 64950 0 1 43050
box -180 -120 1680 4080
use NAND2X1  _1595_
timestamp 1727136778
transform 1 0 60150 0 1 58650
box -180 -120 1380 4080
use OAI21X1  _1596_
timestamp 1727136778
transform -1 0 63450 0 1 58650
box -180 -120 1680 4080
use NAND2X1  _1597_
timestamp 1727136778
transform 1 0 60450 0 1 43050
box -180 -120 1380 4080
use OAI21X1  _1598_
timestamp 1727136778
transform -1 0 64050 0 1 43050
box -180 -120 1680 4080
use NAND2X1  _1599_
timestamp 1727136778
transform -1 0 59550 0 -1 58650
box -180 -120 1380 4080
use OAI21X1  _1600_
timestamp 1727136778
transform -1 0 61950 0 -1 58650
box -180 -120 1680 4080
use NAND2X1  _1601_
timestamp 1727136778
transform 1 0 49950 0 1 58650
box -180 -120 1380 4080
use OAI21X1  _1602_
timestamp 1727136778
transform -1 0 51450 0 -1 66450
box -180 -120 1680 4080
use NAND2X1  _1603_
timestamp 1727136778
transform 1 0 44550 0 -1 58650
box -180 -120 1380 4080
use OAI21X1  _1604_
timestamp 1727136778
transform -1 0 48150 0 -1 58650
box -180 -120 1680 4080
use NAND2X1  _1605_
timestamp 1727136778
transform -1 0 68250 0 1 50850
box -180 -120 1380 4080
use OAI21X1  _1606_
timestamp 1727136778
transform -1 0 79050 0 -1 50850
box -180 -120 1680 4080
use NAND2X1  _1607_
timestamp 1727136778
transform 1 0 66750 0 1 35250
box -180 -120 1380 4080
use OAI21X1  _1608_
timestamp 1727136778
transform -1 0 70050 0 1 35250
box -180 -120 1680 4080
use DFFPOSX1  _1609_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726828622
transform -1 0 71850 0 1 50850
box -195 -120 3795 4080
use DFFPOSX1  _1610_
timestamp 1726828622
transform -1 0 54750 0 1 58650
box -195 -120 3795 4080
use DFFPOSX1  _1611_
timestamp 1726828622
transform -1 0 73650 0 1 43050
box -195 -120 3795 4080
use DFFPOSX1  _1612_
timestamp 1726828622
transform -1 0 59250 0 -1 66450
box -195 -120 3795 4080
use DFFPOSX1  _1613_
timestamp 1726828622
transform -1 0 49350 0 -1 66450
box -195 -120 3795 4080
use DFFPOSX1  _1614_
timestamp 1726828622
transform -1 0 51750 0 -1 58650
box -195 -120 3795 4080
use DFFPOSX1  _1615_
timestamp 1726828622
transform -1 0 79050 0 1 50850
box -195 -120 3795 4080
use DFFPOSX1  _1616_
timestamp 1726828622
transform 1 0 72450 0 -1 43050
box -195 -120 3795 4080
use DFFPOSX1  _1617_
timestamp 1726828622
transform -1 0 76050 0 -1 27450
box -195 -120 3795 4080
use DFFPOSX1  _1618_
timestamp 1726828622
transform -1 0 58050 0 -1 35250
box -195 -120 3795 4080
use DFFPOSX1  _1619_
timestamp 1726828622
transform -1 0 73950 0 -1 19650
box -195 -120 3795 4080
use DFFPOSX1  _1620_
timestamp 1726828622
transform 1 0 82050 0 1 4050
box -195 -120 3795 4080
use DFFPOSX1  _1621_
timestamp 1726828622
transform -1 0 82050 0 1 4050
box -195 -120 3795 4080
use DFFPOSX1  _1622_
timestamp 1726828622
transform 1 0 76350 0 -1 4050
box -195 -120 3795 4080
use DFFPOSX1  _1623_
timestamp 1726828622
transform 1 0 70650 0 -1 4050
box -195 -120 3795 4080
use DFFPOSX1  _1624_
timestamp 1726828622
transform -1 0 72150 0 1 4050
box -195 -120 3795 4080
use DFFPOSX1  _1625_
timestamp 1726828622
transform -1 0 70050 0 1 43050
box -195 -120 3795 4080
use DFFPOSX1  _1626_
timestamp 1726828622
transform -1 0 65550 0 -1 58650
box -195 -120 3795 4080
use DFFPOSX1  _1627_
timestamp 1726828622
transform -1 0 59550 0 1 43050
box -195 -120 3795 4080
use DFFPOSX1  _1628_
timestamp 1726828622
transform -1 0 62550 0 1 50850
box -195 -120 3795 4080
use DFFPOSX1  _1629_
timestamp 1726828622
transform -1 0 45750 0 -1 66450
box -195 -120 3795 4080
use DFFPOSX1  _1630_
timestamp 1726828622
transform -1 0 49050 0 1 58650
box -195 -120 3795 4080
use DFFPOSX1  _1631_
timestamp 1726828622
transform -1 0 75450 0 1 50850
box -195 -120 3795 4080
use DFFPOSX1  _1632_
timestamp 1726828622
transform -1 0 70650 0 -1 35250
box -195 -120 3795 4080
use DFFSR  _1633_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727133863
transform -1 0 88950 0 1 19650
box -180 -120 7380 4095
use DFFSR  _1634_
timestamp 1727133863
transform -1 0 91050 0 -1 19650
box -180 -120 7380 4095
use DFFSR  _1635_
timestamp 1727133863
transform -1 0 90750 0 -1 27450
box -180 -120 7380 4095
use INVX1  _1636_
timestamp 1727136778
transform -1 0 89550 0 -1 82050
box -180 -120 1080 4080
use INVX4  _1637_
timestamp 1727136778
transform 1 0 88950 0 1 89850
box -180 -120 1380 4080
use OAI21X1  _1638_
timestamp 1727136778
transform -1 0 81750 0 -1 82050
box -180 -120 1680 4080
use NOR2X1  _1639_
timestamp 1727136778
transform 1 0 78450 0 -1 82050
box -180 -120 1380 4080
use INVX1  _1640_
timestamp 1727136778
transform 1 0 78450 0 1 82050
box -180 -120 1080 4080
use INVX2  _1641_
timestamp 1727136778
transform -1 0 57150 0 1 82050
box -180 -120 1080 4080
use NAND2X1  _1642_
timestamp 1727136778
transform -1 0 48750 0 1 82050
box -180 -120 1380 4080
use INVX2  _1643_
timestamp 1727136778
transform -1 0 46050 0 -1 89850
box -180 -120 1080 4080
use NAND2X1  _1644_
timestamp 1727136778
transform -1 0 59250 0 1 82050
box -180 -120 1380 4080
use NAND2X1  _1645_
timestamp 1727136778
transform -1 0 67050 0 -1 82050
box -180 -120 1380 4080
use AOI22X1  _1646_
timestamp 1727136778
transform -1 0 63450 0 -1 82050
box -210 -120 1980 4080
use INVX2  _1647_
timestamp 1727136778
transform 1 0 47850 0 1 89850
box -180 -120 1080 4080
use INVX1  _1648_
timestamp 1727136778
transform 1 0 86850 0 -1 82050
box -180 -120 1080 4080
use INVX1  _1649_
timestamp 1727136778
transform -1 0 65250 0 -1 82050
box -180 -120 1080 4080
use OAI21X1  _1650_
timestamp 1727136778
transform -1 0 68250 0 1 82050
box -180 -120 1680 4080
use NAND2X1  _1651_
timestamp 1727136778
transform 1 0 64650 0 1 82050
box -180 -120 1380 4080
use NAND2X1  _1652_
timestamp 1727136778
transform -1 0 55650 0 1 82050
box -180 -120 1380 4080
use OAI21X1  _1653_
timestamp 1727136778
transform 1 0 62550 0 1 82050
box -180 -120 1680 4080
use OAI21X1  _1654_
timestamp 1727136778
transform 1 0 87150 0 1 82050
box -180 -120 1680 4080
use AOI21X1  _1655_
timestamp 1727136778
transform -1 0 86550 0 1 82050
box -180 -120 1680 4080
use NOR2X1  _1656_
timestamp 1727136778
transform 1 0 89250 0 -1 89850
box -180 -120 1380 4080
use OAI21X1  _1657_
timestamp 1727136778
transform 1 0 86850 0 -1 89850
box -180 -120 1680 4080
use OAI21X1  _1658_
timestamp 1727136778
transform 1 0 84750 0 -1 89850
box -180 -120 1680 4080
use XOR2X1  _1659_
timestamp 1727152697
transform -1 0 82350 0 1 82050
box -180 -120 2265 4080
use NOR2X1  _1660_
timestamp 1727136778
transform -1 0 83850 0 -1 89850
box -180 -120 1380 4080
use OAI21X1  _1661_
timestamp 1727136778
transform 1 0 80550 0 -1 89850
box -180 -120 1680 4080
use NAND2X1  _1662_
timestamp 1727136778
transform -1 0 53250 0 1 89850
box -180 -120 1380 4080
use NAND3X1  _1663_
timestamp 1727136778
transform -1 0 50850 0 1 82050
box -180 -120 1680 4080
use AOI22X1  _1664_
timestamp 1727136778
transform -1 0 53550 0 1 82050
box -210 -120 1980 4080
use INVX1  _1665_
timestamp 1727136778
transform -1 0 55650 0 -1 66450
box -180 -120 1080 4080
use NOR2X1  _1666_
timestamp 1727136778
transform -1 0 58650 0 1 66450
box -180 -120 1380 4080
use OAI21X1  _1667_
timestamp 1727136778
transform 1 0 57750 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1668_
timestamp 1727136778
transform 1 0 55950 0 -1 89850
box -180 -120 1680 4080
use OAI21X1  _1669_
timestamp 1727136778
transform -1 0 62250 0 -1 89850
box -180 -120 1680 4080
use AOI21X1  _1670_
timestamp 1727136778
transform 1 0 62850 0 -1 89850
box -180 -120 1680 4080
use INVX1  _1671_
timestamp 1727136778
transform 1 0 78750 0 1 89850
box -180 -120 1080 4080
use OAI21X1  _1672_
timestamp 1727136778
transform -1 0 86550 0 1 89850
box -180 -120 1680 4080
use MUX2X1  _1673_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 82350 0 1 89850
box -180 -120 1965 4080
use NAND2X1  _1674_
timestamp 1727136778
transform -1 0 81750 0 1 89850
box -180 -120 1380 4080
use INVX1  _1675_
timestamp 1727136778
transform -1 0 84150 0 1 82050
box -180 -120 1080 4080
use OAI21X1  _1676_
timestamp 1727136778
transform 1 0 82350 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1677_
timestamp 1727136778
transform -1 0 74850 0 1 82050
box -180 -120 1680 4080
use MUX2X1  _1678_
timestamp 1727136778
transform -1 0 75750 0 -1 82050
box -180 -120 1965 4080
use NAND2X1  _1679_
timestamp 1727136778
transform -1 0 68850 0 -1 82050
box -180 -120 1380 4080
use NAND2X1  _1680_
timestamp 1727136778
transform 1 0 69750 0 -1 82050
box -180 -120 1380 4080
use AOI21X1  _1681_
timestamp 1727136778
transform -1 0 61650 0 1 82050
box -180 -120 1680 4080
use NAND2X1  _1682_
timestamp 1727136778
transform 1 0 68850 0 1 82050
box -180 -120 1380 4080
use NAND3X1  _1683_
timestamp 1727136778
transform 1 0 70950 0 1 82050
box -180 -120 1680 4080
use AOI22X1  _1684_
timestamp 1727136778
transform 1 0 75750 0 1 82050
box -210 -120 1980 4080
use OAI21X1  _1685_
timestamp 1727136778
transform -1 0 64050 0 1 89850
box -180 -120 1680 4080
use OAI21X1  _1686_
timestamp 1727136778
transform 1 0 64950 0 1 89850
box -180 -120 1680 4080
use NAND2X1  _1687_
timestamp 1727136778
transform -1 0 77850 0 -1 89850
box -180 -120 1380 4080
use NAND2X1  _1688_
timestamp 1727136778
transform 1 0 78450 0 -1 89850
box -180 -120 1380 4080
use INVX1  _1689_
timestamp 1727136778
transform 1 0 73650 0 -1 35250
box -180 -120 1080 4080
use NOR2X1  _1690_
timestamp 1727136778
transform 1 0 76650 0 1 89850
box -180 -120 1380 4080
use OAI21X1  _1691_
timestamp 1727136778
transform -1 0 75750 0 1 89850
box -180 -120 1680 4080
use NAND2X1  _1692_
timestamp 1727136778
transform 1 0 53850 0 -1 89850
box -180 -120 1380 4080
use NAND3X1  _1693_
timestamp 1727136778
transform 1 0 46950 0 -1 89850
box -180 -120 1680 4080
use AOI22X1  _1694_
timestamp 1727136778
transform -1 0 51150 0 -1 89850
box -210 -120 1980 4080
use INVX1  _1695_
timestamp 1727136778
transform -1 0 44850 0 1 89850
box -180 -120 1080 4080
use NOR2X1  _1696_
timestamp 1727136778
transform -1 0 46950 0 1 89850
box -180 -120 1380 4080
use OAI21X1  _1697_
timestamp 1727136778
transform -1 0 51150 0 1 89850
box -180 -120 1680 4080
use OAI21X1  _1698_
timestamp 1727136778
transform 1 0 51750 0 -1 89850
box -180 -120 1680 4080
use OAI21X1  _1699_
timestamp 1727136778
transform -1 0 59850 0 -1 89850
box -180 -120 1680 4080
use AOI21X1  _1700_
timestamp 1727136778
transform -1 0 60150 0 1 89850
box -180 -120 1680 4080
use OAI21X1  _1701_
timestamp 1727136778
transform -1 0 55350 0 1 89850
box -180 -120 1680 4080
use OAI21X1  _1702_
timestamp 1727136778
transform 1 0 56250 0 1 89850
box -180 -120 1680 4080
use XOR2X1  _1703_
timestamp 1727152697
transform -1 0 70950 0 1 89850
box -180 -120 2265 4080
use INVX1  _1704_
timestamp 1727136778
transform -1 0 72750 0 -1 58650
box -180 -120 1080 4080
use INVX1  _1705_
timestamp 1727136778
transform 1 0 61050 0 1 89850
box -180 -120 1080 4080
use OAI21X1  _1706_
timestamp 1727136778
transform -1 0 66750 0 -1 89850
box -180 -120 1680 4080
use INVX1  _1707_
timestamp 1727136778
transform -1 0 67950 0 1 89850
box -180 -120 1080 4080
use AOI22X1  _1708_
timestamp 1727136778
transform 1 0 67650 0 -1 89850
box -210 -120 1980 4080
use NAND2X1  _1709_
timestamp 1727136778
transform -1 0 56250 0 -1 74250
box -180 -120 1380 4080
use AND2X2  _1710_
timestamp 1727136778
transform -1 0 59550 0 1 74250
box -180 -120 1680 4095
use NAND2X1  _1711_
timestamp 1727136778
transform -1 0 54750 0 1 74250
box -180 -120 1380 4080
use AOI22X1  _1712_
timestamp 1727136778
transform -1 0 57450 0 1 74250
box -210 -120 1980 4080
use OAI21X1  _1713_
timestamp 1727136778
transform -1 0 52650 0 1 74250
box -180 -120 1680 4080
use OAI21X1  _1714_
timestamp 1727136778
transform 1 0 56850 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1715_
timestamp 1727136778
transform -1 0 60750 0 -1 74250
box -180 -120 1680 4080
use AOI21X1  _1716_
timestamp 1727136778
transform 1 0 61650 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1717_
timestamp 1727136778
transform -1 0 67950 0 1 66450
box -180 -120 1680 4080
use OAI21X1  _1718_
timestamp 1727136778
transform 1 0 68850 0 1 66450
box -180 -120 1680 4080
use XOR2X1  _1719_
timestamp 1727152697
transform 1 0 71250 0 1 66450
box -180 -120 2265 4080
use XNOR2X1  _1720_
timestamp 1727153789
transform 1 0 63750 0 -1 66450
box -180 -120 2280 4080
use NAND2X1  _1721_
timestamp 1727136778
transform 1 0 70350 0 -1 89850
box -180 -120 1380 4080
use NAND3X1  _1722_
timestamp 1727136778
transform 1 0 71850 0 1 89850
box -180 -120 1680 4080
use NAND3X1  _1723_
timestamp 1727136778
transform 1 0 72150 0 -1 89850
box -180 -120 1680 4080
use NAND2X1  _1724_
timestamp 1727136778
transform -1 0 73350 0 1 58650
box -180 -120 1380 4080
use OAI21X1  _1725_
timestamp 1727136778
transform 1 0 66750 0 -1 66450
box -180 -120 1680 4080
use INVX1  _1726_
timestamp 1727136778
transform -1 0 64950 0 1 58650
box -180 -120 1080 4080
use OAI21X1  _1727_
timestamp 1727136778
transform -1 0 67350 0 1 58650
box -180 -120 1680 4080
use NAND2X1  _1728_
timestamp 1727136778
transform -1 0 46650 0 1 82050
box -180 -120 1380 4080
use AND2X2  _1729_
timestamp 1727136778
transform 1 0 46350 0 -1 82050
box -180 -120 1680 4095
use NAND2X1  _1730_
timestamp 1727136778
transform -1 0 49950 0 -1 82050
box -180 -120 1380 4080
use AOI22X1  _1731_
timestamp 1727136778
transform -1 0 52650 0 -1 82050
box -210 -120 1980 4080
use OAI21X1  _1732_
timestamp 1727136778
transform 1 0 53250 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1733_
timestamp 1727136778
transform 1 0 55650 0 -1 82050
box -180 -120 1680 4080
use OAI21X1  _1734_
timestamp 1727136778
transform 1 0 74850 0 -1 74250
box -180 -120 1680 4080
use AOI21X1  _1735_
timestamp 1727136778
transform 1 0 73950 0 1 66450
box -180 -120 1680 4080
use OAI21X1  _1736_
timestamp 1727136778
transform -1 0 80250 0 1 66450
box -180 -120 1680 4080
use OAI21X1  _1737_
timestamp 1727136778
transform 1 0 76350 0 1 66450
box -180 -120 1680 4080
use INVX1  _1738_
timestamp 1727136778
transform 1 0 76950 0 1 58650
box -180 -120 1080 4080
use XOR2X1  _1739_
timestamp 1727152697
transform 1 0 73950 0 1 58650
box -180 -120 2265 4080
use INVX1  _1740_
timestamp 1727136778
transform -1 0 78450 0 -1 66450
box -180 -120 1080 4080
use AOI21X1  _1741_
timestamp 1727136778
transform 1 0 78750 0 1 58650
box -180 -120 1680 4080
use NAND2X1  _1742_
timestamp 1727136778
transform 1 0 52950 0 -1 74250
box -180 -120 1380 4080
use AND2X2  _1743_
timestamp 1727136778
transform -1 0 43350 0 1 74250
box -180 -120 1680 4095
use NAND2X1  _1744_
timestamp 1727136778
transform -1 0 45450 0 1 74250
box -180 -120 1380 4080
use AOI22X1  _1745_
timestamp 1727136778
transform -1 0 50250 0 1 74250
box -210 -120 1980 4080
use OAI21X1  _1746_
timestamp 1727136778
transform 1 0 46350 0 1 74250
box -180 -120 1680 4080
use OAI21X1  _1747_
timestamp 1727136778
transform 1 0 50850 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1748_
timestamp 1727136778
transform -1 0 77850 0 1 74250
box -180 -120 1680 4080
use AOI21X1  _1749_
timestamp 1727136778
transform 1 0 78750 0 1 74250
box -180 -120 1680 4080
use OAI21X1  _1750_
timestamp 1727136778
transform 1 0 82050 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1751_
timestamp 1727136778
transform 1 0 80850 0 1 66450
box -180 -120 1680 4080
use INVX1  _1752_
timestamp 1727136778
transform -1 0 80250 0 -1 66450
box -180 -120 1080 4080
use XOR2X1  _1753_
timestamp 1727152697
transform 1 0 81150 0 1 58650
box -180 -120 2265 4080
use INVX1  _1754_
timestamp 1727136778
transform 1 0 77550 0 1 27450
box -180 -120 1080 4080
use OAI21X1  _1755_
timestamp 1727136778
transform 1 0 81150 0 -1 66450
box -180 -120 1680 4080
use INVX1  _1756_
timestamp 1727136778
transform 1 0 73050 0 -1 74250
box -180 -120 1080 4080
use AND2X2  _1757_
timestamp 1727136778
transform -1 0 67350 0 -1 74250
box -180 -120 1680 4095
use NAND2X1  _1758_
timestamp 1727136778
transform 1 0 64050 0 -1 74250
box -180 -120 1380 4080
use AOI22X1  _1759_
timestamp 1727136778
transform 1 0 60450 0 1 74250
box -210 -120 1980 4080
use OAI21X1  _1760_
timestamp 1727136778
transform 1 0 68250 0 -1 74250
box -180 -120 1680 4080
use OAI22X1  _1761_
timestamp 1727136778
transform -1 0 72150 0 -1 74250
box -180 -120 1980 4080
use OAI21X1  _1762_
timestamp 1727136778
transform -1 0 78750 0 -1 74250
box -180 -120 1680 4080
use AOI21X1  _1763_
timestamp 1727136778
transform 1 0 79650 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1764_
timestamp 1727136778
transform 1 0 84150 0 -1 74250
box -180 -120 1680 4080
use OAI21X1  _1765_
timestamp 1727136778
transform 1 0 86550 0 -1 74250
box -180 -120 1680 4080
use NAND2X1  _1766_
timestamp 1727136778
transform 1 0 88050 0 -1 58650
box -180 -120 1380 4080
use INVX1  _1767_
timestamp 1727136778
transform 1 0 73650 0 -1 66450
box -180 -120 1080 4080
use AOI21X1  _1768_
timestamp 1727136778
transform -1 0 73050 0 -1 66450
box -180 -120 1680 4080
use AOI21X1  _1769_
timestamp 1727136778
transform -1 0 70650 0 -1 66450
box -180 -120 1680 4080
use OAI21X1  _1770_
timestamp 1727136778
transform -1 0 76650 0 -1 66450
box -180 -120 1680 4080
use OR2X2  _1771_
timestamp 1727136778
transform 1 0 83250 0 1 66450
box -180 -120 1680 4080
use AOI22X1  _1772_
timestamp 1727136778
transform 1 0 83550 0 -1 66450
box -210 -120 1980 4080
use INVX1  _1773_
timestamp 1727136778
transform -1 0 88050 0 1 89850
box -180 -120 1080 4080
use NAND2X1  _1774_
timestamp 1727136778
transform -1 0 85350 0 1 58650
box -180 -120 1380 4080
use NAND2X1  _1775_
timestamp 1727136778
transform -1 0 87150 0 -1 58650
box -180 -120 1380 4080
use OAI21X1  _1776_
timestamp 1727136778
transform 1 0 85950 0 -1 66450
box -180 -120 1680 4080
use NAND2X1  _1777_
timestamp 1727136778
transform 1 0 74550 0 1 74250
box -180 -120 1380 4080
use AND2X2  _1778_
timestamp 1727136778
transform 1 0 67650 0 1 74250
box -180 -120 1680 4095
use NAND2X1  _1779_
timestamp 1727136778
transform 1 0 65550 0 1 74250
box -180 -120 1380 4080
use AOI22X1  _1780_
timestamp 1727136778
transform 1 0 63150 0 1 74250
box -210 -120 1980 4080
use OAI21X1  _1781_
timestamp 1727136778
transform 1 0 70050 0 1 74250
box -180 -120 1680 4080
use OAI21X1  _1782_
timestamp 1727136778
transform 1 0 72150 0 1 74250
box -180 -120 1680 4080
use OAI21X1  _1783_
timestamp 1727136778
transform 1 0 84750 0 -1 82050
box -180 -120 1680 4080
use AOI21X1  _1784_
timestamp 1727136778
transform 1 0 82650 0 1 74250
box -180 -120 1680 4080
use OAI21X1  _1785_
timestamp 1727136778
transform -1 0 88950 0 1 74250
box -180 -120 1680 4080
use OAI21X1  _1786_
timestamp 1727136778
transform 1 0 89550 0 1 74250
box -180 -120 1680 4080
use NAND2X1  _1787_
timestamp 1727136778
transform -1 0 89850 0 -1 4050
box -180 -120 1380 4080
use NAND2X1  _1788_
timestamp 1727136778
transform 1 0 86250 0 1 58650
box -180 -120 1380 4080
use INVX1  _1789_
timestamp 1727136778
transform 1 0 90150 0 -1 66450
box -180 -120 1080 4080
use NAND3X1  _1790_
timestamp 1727136778
transform 1 0 90450 0 1 58650
box -180 -120 1680 4080
use NAND2X1  _1791_
timestamp 1727136778
transform 1 0 90150 0 1 35250
box -180 -120 1380 4080
use NOR2X1  _1792_
timestamp 1727136778
transform 1 0 70050 0 1 58650
box -180 -120 1380 4080
use NAND2X1  _1793_
timestamp 1727136778
transform 1 0 68250 0 1 58650
box -180 -120 1380 4080
use NOR2X1  _1794_
timestamp 1727136778
transform 1 0 73650 0 -1 58650
box -180 -120 1380 4080
use NAND3X1  _1795_
timestamp 1727136778
transform -1 0 85050 0 -1 58650
box -180 -120 1680 4080
use NOR2X1  _1796_
timestamp 1727136778
transform 1 0 81750 0 -1 58650
box -180 -120 1380 4080
use AND2X2  _1797_
timestamp 1727136778
transform -1 0 77250 0 -1 58650
box -180 -120 1680 4095
use NAND3X1  _1798_
timestamp 1727136778
transform -1 0 89550 0 1 58650
box -180 -120 1680 4080
use NAND2X1  _1799_
timestamp 1727136778
transform -1 0 89550 0 -1 66450
box -180 -120 1380 4080
use NAND2X1  _1800_
timestamp 1727136778
transform -1 0 89250 0 1 50850
box -180 -120 1380 4080
use NAND2X1  _1801_
timestamp 1727136778
transform 1 0 81450 0 1 50850
box -180 -120 1380 4080
use NOR2X1  _1802_
timestamp 1727136778
transform 1 0 71850 0 -1 82050
box -180 -120 1380 4080
use OAI21X1  _1803_
timestamp 1727136778
transform 1 0 88650 0 1 4050
box -180 -120 1680 4080
use NOR2X1  _1804_
timestamp 1727136778
transform -1 0 89550 0 1 66450
box -180 -120 1380 4080
use AOI21X1  _1805_
timestamp 1727136778
transform 1 0 90450 0 1 66450
box -180 -120 1680 4080
use XOR2X1  _1806_
timestamp 1727152697
transform -1 0 87750 0 1 66450
box -180 -120 2265 4080
use OAI21X1  _1807_
timestamp 1727136778
transform 1 0 85650 0 1 50850
box -180 -120 1680 4080
use NAND3X1  _1808_
timestamp 1727136778
transform 1 0 83250 0 1 50850
box -180 -120 1680 4080
use AOI21X1  _1809_
timestamp 1727136778
transform 1 0 85050 0 1 74250
box -180 -120 1680 4080
use XOR2X1  _1810_
timestamp 1727152697
transform 1 0 88950 0 -1 74250
box -180 -120 2265 4080
use NAND3X1  _1811_
timestamp 1727136778
transform 1 0 86250 0 1 4050
box -180 -120 1680 4080
use INVX1  _1812_
timestamp 1727136778
transform 1 0 90150 0 -1 58650
box -180 -120 1080 4080
use NAND3X1  _1813_
timestamp 1727136778
transform -1 0 91650 0 1 50850
box -180 -120 1680 4080
use NAND2X1  _1814_
timestamp 1727136778
transform -1 0 91350 0 -1 50850
box -180 -120 1380 4080
use NAND3X1  _1815_
timestamp 1727136778
transform 1 0 88050 0 -1 50850
box -180 -120 1680 4080
use NAND3X1  _1816_
timestamp 1727136778
transform -1 0 91650 0 1 43050
box -180 -120 1680 4080
use NAND2X1  _1817_
timestamp 1727136778
transform -1 0 89250 0 1 43050
box -180 -120 1380 4080
use BUFX2  _1818_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 50550 0 -1 35250
box -180 -120 1380 4080
use BUFX2  _1819_
timestamp 1727136778
transform -1 0 40350 0 -1 35250
box -180 -120 1380 4080
use BUFX2  _1820_
timestamp 1727136778
transform -1 0 70350 0 -1 19650
box -180 -120 1380 4080
use BUFX2  _1821_
timestamp 1727136778
transform -1 0 85950 0 -1 4050
box -180 -120 1380 4080
use BUFX2  _1822_
timestamp 1727136778
transform 1 0 82650 0 -1 4050
box -180 -120 1380 4080
use BUFX2  _1823_
timestamp 1727136778
transform 1 0 80550 0 -1 4050
box -180 -120 1380 4080
use BUFX2  _1824_
timestamp 1727136778
transform 1 0 75150 0 -1 4050
box -180 -120 1380 4080
use BUFX2  _1825_
timestamp 1727136778
transform 1 0 69450 0 -1 4050
box -180 -120 1380 4080
use BUFX2  _1826_
timestamp 1727136778
transform 1 0 86550 0 -1 4050
box -180 -120 1380 4080
use BUFX2  BUFX2_insert0
timestamp 1727136778
transform 1 0 59550 0 1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert1
timestamp 1727136778
transform -1 0 34650 0 1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert2
timestamp 1727136778
transform -1 0 36150 0 1 35250
box -180 -120 1380 4080
use BUFX2  BUFX2_insert3
timestamp 1727136778
transform -1 0 35550 0 -1 58650
box -180 -120 1380 4080
use BUFX2  BUFX2_insert4
timestamp 1727136778
transform -1 0 67650 0 -1 58650
box -180 -120 1380 4080
use BUFX2  BUFX2_insert5
timestamp 1727136778
transform -1 0 57750 0 -1 58650
box -180 -120 1380 4080
use BUFX2  BUFX2_insert6
timestamp 1727136778
transform -1 0 42450 0 -1 35250
box -180 -120 1380 4080
use BUFX2  BUFX2_insert7
timestamp 1727136778
transform -1 0 52650 0 -1 35250
box -180 -120 1380 4080
use BUFX2  BUFX2_insert13
timestamp 1727136778
transform 1 0 78450 0 1 43050
box -180 -120 1380 4080
use BUFX2  BUFX2_insert14
timestamp 1727136778
transform -1 0 58950 0 1 50850
box -180 -120 1380 4080
use BUFX2  BUFX2_insert15
timestamp 1727136778
transform -1 0 66450 0 1 50850
box -180 -120 1380 4080
use BUFX2  BUFX2_insert16
timestamp 1727136778
transform -1 0 61950 0 -1 43050
box -180 -120 1380 4080
use BUFX2  BUFX2_insert17
timestamp 1727136778
transform 1 0 38550 0 1 58650
box -180 -120 1380 4080
use BUFX2  BUFX2_insert18
timestamp 1727136778
transform -1 0 36450 0 1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert19
timestamp 1727136778
transform 1 0 46050 0 1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert20
timestamp 1727136778
transform -1 0 37950 0 1 43050
box -180 -120 1380 4080
use BUFX2  BUFX2_insert21
timestamp 1727136778
transform 1 0 80250 0 1 43050
box -180 -120 1380 4080
use BUFX2  BUFX2_insert22
timestamp 1727136778
transform -1 0 64650 0 1 50850
box -180 -120 1380 4080
use BUFX2  BUFX2_insert23
timestamp 1727136778
transform 1 0 64350 0 -1 50850
box -180 -120 1380 4080
use BUFX2  BUFX2_insert24
timestamp 1727136778
transform 1 0 79650 0 -1 50850
box -180 -120 1380 4080
use BUFX2  BUFX2_insert25
timestamp 1727136778
transform -1 0 36750 0 -1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert26
timestamp 1727136778
transform -1 0 41250 0 1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert27
timestamp 1727136778
transform -1 0 37350 0 -1 58650
box -180 -120 1380 4080
use BUFX2  BUFX2_insert28
timestamp 1727136778
transform 1 0 48150 0 1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert29
timestamp 1727136778
transform -1 0 34350 0 1 35250
box -180 -120 1380 4080
use BUFX2  BUFX2_insert30
timestamp 1727136778
transform 1 0 51150 0 1 35250
box -180 -120 1380 4080
use BUFX2  BUFX2_insert31
timestamp 1727136778
transform -1 0 34650 0 -1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert32
timestamp 1727136778
transform 1 0 53250 0 1 66450
box -180 -120 1380 4080
use BUFX2  BUFX2_insert33
timestamp 1727136778
transform -1 0 77550 0 -1 82050
box -180 -120 1380 4080
use BUFX2  BUFX2_insert34
timestamp 1727136778
transform -1 0 91650 0 -1 82050
box -180 -120 1380 4080
use BUFX2  BUFX2_insert35
timestamp 1727136778
transform -1 0 75750 0 -1 89850
box -180 -120 1380 4080
use BUFX2  BUFX2_insert36
timestamp 1727136778
transform -1 0 90750 0 1 82050
box -180 -120 1380 4080
use CLKBUF1  CLKBUF1_insert8 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 71250 0 -1 58650
box -180 -120 3180 4080
use CLKBUF1  CLKBUF1_insert9
timestamp 1727136778
transform -1 0 77550 0 1 43050
box -180 -120 3180 4080
use CLKBUF1  CLKBUF1_insert10
timestamp 1727136778
transform -1 0 90450 0 1 11850
box -180 -120 3180 4080
use CLKBUF1  CLKBUF1_insert11
timestamp 1727136778
transform -1 0 80850 0 -1 58650
box -180 -120 3180 4080
use CLKBUF1  CLKBUF1_insert12
timestamp 1727136778
transform -1 0 77850 0 -1 19650
box -180 -120 3180 4080
use FILL  FILL89850x150 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1700315010
transform -1 0 90150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL90150x150
timestamp 1700315010
transform -1 0 90450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL90150x4050
timestamp 1700315010
transform 1 0 90150 0 1 4050
box -180 -120 480 4080
use FILL  FILL90150x89850
timestamp 1700315010
transform 1 0 90150 0 1 89850
box -180 -120 480 4080
use FILL  FILL90450x150
timestamp 1700315010
transform -1 0 90750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL90450x4050
timestamp 1700315010
transform 1 0 90450 0 1 4050
box -180 -120 480 4080
use FILL  FILL90450x7950
timestamp 1700315010
transform -1 0 90750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL90450x11850
timestamp 1700315010
transform 1 0 90450 0 1 11850
box -180 -120 480 4080
use FILL  FILL90450x27450
timestamp 1700315010
transform 1 0 90450 0 1 27450
box -180 -120 480 4080
use FILL  FILL90450x31350
timestamp 1700315010
transform -1 0 90750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL90450x85950
timestamp 1700315010
transform -1 0 90750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL90450x89850
timestamp 1700315010
transform 1 0 90450 0 1 89850
box -180 -120 480 4080
use FILL  FILL90750x150
timestamp 1700315010
transform -1 0 91050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL90750x4050
timestamp 1700315010
transform 1 0 90750 0 1 4050
box -180 -120 480 4080
use FILL  FILL90750x7950
timestamp 1700315010
transform -1 0 91050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL90750x11850
timestamp 1700315010
transform 1 0 90750 0 1 11850
box -180 -120 480 4080
use FILL  FILL90750x19650
timestamp 1700315010
transform 1 0 90750 0 1 19650
box -180 -120 480 4080
use FILL  FILL90750x23550
timestamp 1700315010
transform -1 0 91050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL90750x27450
timestamp 1700315010
transform 1 0 90750 0 1 27450
box -180 -120 480 4080
use FILL  FILL90750x31350
timestamp 1700315010
transform -1 0 91050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL90750x39150
timestamp 1700315010
transform -1 0 91050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL90750x82050
timestamp 1700315010
transform 1 0 90750 0 1 82050
box -180 -120 480 4080
use FILL  FILL90750x85950
timestamp 1700315010
transform -1 0 91050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL90750x89850
timestamp 1700315010
transform 1 0 90750 0 1 89850
box -180 -120 480 4080
use FILL  FILL91050x150
timestamp 1700315010
transform -1 0 91350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL91050x4050
timestamp 1700315010
transform 1 0 91050 0 1 4050
box -180 -120 480 4080
use FILL  FILL91050x7950
timestamp 1700315010
transform -1 0 91350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL91050x11850
timestamp 1700315010
transform 1 0 91050 0 1 11850
box -180 -120 480 4080
use FILL  FILL91050x15750
timestamp 1700315010
transform -1 0 91350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL91050x19650
timestamp 1700315010
transform 1 0 91050 0 1 19650
box -180 -120 480 4080
use FILL  FILL91050x23550
timestamp 1700315010
transform -1 0 91350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL91050x27450
timestamp 1700315010
transform 1 0 91050 0 1 27450
box -180 -120 480 4080
use FILL  FILL91050x31350
timestamp 1700315010
transform -1 0 91350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL91050x39150
timestamp 1700315010
transform -1 0 91350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL91050x54750
timestamp 1700315010
transform -1 0 91350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL91050x62550
timestamp 1700315010
transform -1 0 91350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL91050x70350
timestamp 1700315010
transform -1 0 91350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL91050x74250
timestamp 1700315010
transform 1 0 91050 0 1 74250
box -180 -120 480 4080
use FILL  FILL91050x82050
timestamp 1700315010
transform 1 0 91050 0 1 82050
box -180 -120 480 4080
use FILL  FILL91050x85950
timestamp 1700315010
transform -1 0 91350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL91050x89850
timestamp 1700315010
transform 1 0 91050 0 1 89850
box -180 -120 480 4080
use FILL  FILL91350x150
timestamp 1700315010
transform -1 0 91650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL91350x4050
timestamp 1700315010
transform 1 0 91350 0 1 4050
box -180 -120 480 4080
use FILL  FILL91350x7950
timestamp 1700315010
transform -1 0 91650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL91350x11850
timestamp 1700315010
transform 1 0 91350 0 1 11850
box -180 -120 480 4080
use FILL  FILL91350x15750
timestamp 1700315010
transform -1 0 91650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL91350x19650
timestamp 1700315010
transform 1 0 91350 0 1 19650
box -180 -120 480 4080
use FILL  FILL91350x23550
timestamp 1700315010
transform -1 0 91650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL91350x27450
timestamp 1700315010
transform 1 0 91350 0 1 27450
box -180 -120 480 4080
use FILL  FILL91350x31350
timestamp 1700315010
transform -1 0 91650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL91350x35250
timestamp 1700315010
transform 1 0 91350 0 1 35250
box -180 -120 480 4080
use FILL  FILL91350x39150
timestamp 1700315010
transform -1 0 91650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL91350x46950
timestamp 1700315010
transform -1 0 91650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL91350x54750
timestamp 1700315010
transform -1 0 91650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL91350x62550
timestamp 1700315010
transform -1 0 91650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL91350x70350
timestamp 1700315010
transform -1 0 91650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL91350x74250
timestamp 1700315010
transform 1 0 91350 0 1 74250
box -180 -120 480 4080
use FILL  FILL91350x82050
timestamp 1700315010
transform 1 0 91350 0 1 82050
box -180 -120 480 4080
use FILL  FILL91350x85950
timestamp 1700315010
transform -1 0 91650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL91350x89850
timestamp 1700315010
transform 1 0 91350 0 1 89850
box -180 -120 480 4080
use FILL  FILL91650x150
timestamp 1700315010
transform -1 0 91950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL91650x4050
timestamp 1700315010
transform 1 0 91650 0 1 4050
box -180 -120 480 4080
use FILL  FILL91650x7950
timestamp 1700315010
transform -1 0 91950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL91650x11850
timestamp 1700315010
transform 1 0 91650 0 1 11850
box -180 -120 480 4080
use FILL  FILL91650x15750
timestamp 1700315010
transform -1 0 91950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL91650x19650
timestamp 1700315010
transform 1 0 91650 0 1 19650
box -180 -120 480 4080
use FILL  FILL91650x23550
timestamp 1700315010
transform -1 0 91950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL91650x27450
timestamp 1700315010
transform 1 0 91650 0 1 27450
box -180 -120 480 4080
use FILL  FILL91650x31350
timestamp 1700315010
transform -1 0 91950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL91650x35250
timestamp 1700315010
transform 1 0 91650 0 1 35250
box -180 -120 480 4080
use FILL  FILL91650x39150
timestamp 1700315010
transform -1 0 91950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL91650x43050
timestamp 1700315010
transform 1 0 91650 0 1 43050
box -180 -120 480 4080
use FILL  FILL91650x46950
timestamp 1700315010
transform -1 0 91950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL91650x50850
timestamp 1700315010
transform 1 0 91650 0 1 50850
box -180 -120 480 4080
use FILL  FILL91650x54750
timestamp 1700315010
transform -1 0 91950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL91650x62550
timestamp 1700315010
transform -1 0 91950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL91650x70350
timestamp 1700315010
transform -1 0 91950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL91650x74250
timestamp 1700315010
transform 1 0 91650 0 1 74250
box -180 -120 480 4080
use FILL  FILL91650x78150
timestamp 1700315010
transform -1 0 91950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL91650x82050
timestamp 1700315010
transform 1 0 91650 0 1 82050
box -180 -120 480 4080
use FILL  FILL91650x85950
timestamp 1700315010
transform -1 0 91950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL91650x89850
timestamp 1700315010
transform 1 0 91650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__889_
timestamp 1700315010
transform 1 0 79950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__890_
timestamp 1700315010
transform -1 0 74250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__891_
timestamp 1700315010
transform -1 0 76350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__892_
timestamp 1700315010
transform 1 0 80250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__893_
timestamp 1700315010
transform -1 0 78150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__894_
timestamp 1700315010
transform 1 0 82050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__895_
timestamp 1700315010
transform -1 0 78450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__896_
timestamp 1700315010
transform -1 0 76350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__897_
timestamp 1700315010
transform 1 0 76350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__898_
timestamp 1700315010
transform -1 0 82050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__899_
timestamp 1700315010
transform 1 0 78450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__900_
timestamp 1700315010
transform -1 0 87450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__901_
timestamp 1700315010
transform -1 0 85350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__902_
timestamp 1700315010
transform 1 0 86550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__903_
timestamp 1700315010
transform 1 0 73050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__904_
timestamp 1700315010
transform -1 0 79950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__905_
timestamp 1700315010
transform -1 0 85050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__906_
timestamp 1700315010
transform -1 0 62850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__907_
timestamp 1700315010
transform 1 0 74550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__908_
timestamp 1700315010
transform 1 0 88950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__909_
timestamp 1700315010
transform 1 0 83550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__910_
timestamp 1700315010
transform 1 0 82650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__911_
timestamp 1700315010
transform 1 0 80850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__912_
timestamp 1700315010
transform 1 0 85950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__913_
timestamp 1700315010
transform -1 0 83250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__914_
timestamp 1700315010
transform -1 0 78450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__915_
timestamp 1700315010
transform 1 0 78150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__916_
timestamp 1700315010
transform -1 0 84150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__917_
timestamp 1700315010
transform 1 0 87150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__918_
timestamp 1700315010
transform -1 0 80550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__919_
timestamp 1700315010
transform 1 0 80550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__920_
timestamp 1700315010
transform -1 0 83250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__921_
timestamp 1700315010
transform 1 0 84450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__922_
timestamp 1700315010
transform 1 0 80250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__923_
timestamp 1700315010
transform 1 0 88350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__924_
timestamp 1700315010
transform 1 0 88050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__925_
timestamp 1700315010
transform -1 0 89250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__926_
timestamp 1700315010
transform -1 0 64650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__927_
timestamp 1700315010
transform 1 0 72450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__928_
timestamp 1700315010
transform 1 0 70050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__929_
timestamp 1700315010
transform 1 0 62850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__930_
timestamp 1700315010
transform 1 0 54750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__931_
timestamp 1700315010
transform -1 0 57150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__932_
timestamp 1700315010
transform 1 0 61650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__933_
timestamp 1700315010
transform -1 0 65850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__934_
timestamp 1700315010
transform 1 0 67650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__935_
timestamp 1700315010
transform -1 0 80550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__936_
timestamp 1700315010
transform 1 0 60750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__937_
timestamp 1700315010
transform -1 0 59550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__938_
timestamp 1700315010
transform -1 0 59550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__939_
timestamp 1700315010
transform 1 0 54450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__940_
timestamp 1700315010
transform 1 0 51450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__941_
timestamp 1700315010
transform -1 0 48450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__942_
timestamp 1700315010
transform 1 0 54150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__943_
timestamp 1700315010
transform 1 0 51750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__944_
timestamp 1700315010
transform -1 0 79350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__945_
timestamp 1700315010
transform 1 0 83250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__946_
timestamp 1700315010
transform 1 0 80850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__947_
timestamp 1700315010
transform 1 0 84450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__948_
timestamp 1700315010
transform 1 0 78450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__949_
timestamp 1700315010
transform 1 0 76050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__950_
timestamp 1700315010
transform -1 0 69450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__951_
timestamp 1700315010
transform 1 0 58350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__952_
timestamp 1700315010
transform 1 0 34650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__953_
timestamp 1700315010
transform 1 0 39150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__954_
timestamp 1700315010
transform -1 0 37050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__955_
timestamp 1700315010
transform 1 0 40950 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__956_
timestamp 1700315010
transform 1 0 47250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__957_
timestamp 1700315010
transform 1 0 52050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__958_
timestamp 1700315010
transform 1 0 53850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__959_
timestamp 1700315010
transform 1 0 53850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__960_
timestamp 1700315010
transform 1 0 47250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__961_
timestamp 1700315010
transform -1 0 51750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__962_
timestamp 1700315010
transform 1 0 56250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__963_
timestamp 1700315010
transform 1 0 43350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__964_
timestamp 1700315010
transform -1 0 39450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__965_
timestamp 1700315010
transform 1 0 37050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__966_
timestamp 1700315010
transform 1 0 49650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__967_
timestamp 1700315010
transform -1 0 43650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__968_
timestamp 1700315010
transform 1 0 38250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__969_
timestamp 1700315010
transform -1 0 41250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__970_
timestamp 1700315010
transform 1 0 45150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__971_
timestamp 1700315010
transform 1 0 45150 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__972_
timestamp 1700315010
transform -1 0 47550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__973_
timestamp 1700315010
transform 1 0 45150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__974_
timestamp 1700315010
transform -1 0 52050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__975_
timestamp 1700315010
transform 1 0 45450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__976_
timestamp 1700315010
transform 1 0 38850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__977_
timestamp 1700315010
transform 1 0 31350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__978_
timestamp 1700315010
transform 1 0 37050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__979_
timestamp 1700315010
transform 1 0 31050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__980_
timestamp 1700315010
transform 1 0 43050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__981_
timestamp 1700315010
transform 1 0 54150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__982_
timestamp 1700315010
transform -1 0 51750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__983_
timestamp 1700315010
transform -1 0 40950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__984_
timestamp 1700315010
transform -1 0 36150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__985_
timestamp 1700315010
transform -1 0 34950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__986_
timestamp 1700315010
transform -1 0 25650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__987_
timestamp 1700315010
transform -1 0 23550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__988_
timestamp 1700315010
transform -1 0 20250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__989_
timestamp 1700315010
transform -1 0 26850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__990_
timestamp 1700315010
transform 1 0 27450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__991_
timestamp 1700315010
transform 1 0 35550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__992_
timestamp 1700315010
transform -1 0 35550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__993_
timestamp 1700315010
transform 1 0 29850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__994_
timestamp 1700315010
transform 1 0 38550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__995_
timestamp 1700315010
transform -1 0 41550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__996_
timestamp 1700315010
transform 1 0 25050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__997_
timestamp 1700315010
transform -1 0 21150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__998_
timestamp 1700315010
transform 1 0 23850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__999_
timestamp 1700315010
transform 1 0 32550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1000_
timestamp 1700315010
transform 1 0 33150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1001_
timestamp 1700315010
transform 1 0 41250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1002_
timestamp 1700315010
transform 1 0 34650 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1003_
timestamp 1700315010
transform -1 0 43950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1004_
timestamp 1700315010
transform 1 0 36750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1005_
timestamp 1700315010
transform -1 0 34650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1006_
timestamp 1700315010
transform 1 0 30150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1007_
timestamp 1700315010
transform -1 0 24750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1008_
timestamp 1700315010
transform 1 0 26250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1009_
timestamp 1700315010
transform -1 0 28950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1010_
timestamp 1700315010
transform 1 0 34350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1011_
timestamp 1700315010
transform -1 0 32850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1012_
timestamp 1700315010
transform -1 0 21750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1013_
timestamp 1700315010
transform -1 0 36750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1014_
timestamp 1700315010
transform -1 0 32550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1015_
timestamp 1700315010
transform -1 0 30450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1016_
timestamp 1700315010
transform -1 0 30750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1017_
timestamp 1700315010
transform 1 0 32550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1018_
timestamp 1700315010
transform -1 0 35250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1019_
timestamp 1700315010
transform -1 0 26250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1020_
timestamp 1700315010
transform -1 0 22350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1021_
timestamp 1700315010
transform -1 0 21150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1022_
timestamp 1700315010
transform -1 0 20550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1023_
timestamp 1700315010
transform 1 0 16650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1024_
timestamp 1700315010
transform 1 0 22050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1025_
timestamp 1700315010
transform 1 0 21450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1026_
timestamp 1700315010
transform 1 0 18450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1027_
timestamp 1700315010
transform 1 0 22050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1028_
timestamp 1700315010
transform 1 0 15450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1029_
timestamp 1700315010
transform -1 0 13350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1030_
timestamp 1700315010
transform -1 0 23550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1031_
timestamp 1700315010
transform 1 0 19050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1032_
timestamp 1700315010
transform -1 0 18150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1033_
timestamp 1700315010
transform -1 0 15750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1034_
timestamp 1700315010
transform -1 0 24450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1035_
timestamp 1700315010
transform -1 0 16050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1036_
timestamp 1700315010
transform -1 0 17250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1037_
timestamp 1700315010
transform -1 0 15450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1038_
timestamp 1700315010
transform 1 0 24150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1039_
timestamp 1700315010
transform -1 0 19650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1040_
timestamp 1700315010
transform -1 0 30450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1041_
timestamp 1700315010
transform -1 0 39450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1042_
timestamp 1700315010
transform 1 0 28050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1043_
timestamp 1700315010
transform 1 0 34050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1044_
timestamp 1700315010
transform 1 0 33450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1045_
timestamp 1700315010
transform 1 0 31050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1046_
timestamp 1700315010
transform -1 0 23850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1047_
timestamp 1700315010
transform 1 0 25950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1048_
timestamp 1700315010
transform -1 0 28950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1049_
timestamp 1700315010
transform -1 0 21450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1050_
timestamp 1700315010
transform 1 0 22050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1051_
timestamp 1700315010
transform -1 0 10050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1052_
timestamp 1700315010
transform 1 0 17550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1053_
timestamp 1700315010
transform 1 0 17850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1054_
timestamp 1700315010
transform -1 0 20250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1055_
timestamp 1700315010
transform -1 0 13950 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1056_
timestamp 1700315010
transform 1 0 14550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1057_
timestamp 1700315010
transform -1 0 28350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1058_
timestamp 1700315010
transform 1 0 18450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1059_
timestamp 1700315010
transform 1 0 16050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1060_
timestamp 1700315010
transform -1 0 17250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1061_
timestamp 1700315010
transform -1 0 43650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1062_
timestamp 1700315010
transform -1 0 28350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1063_
timestamp 1700315010
transform 1 0 32250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1064_
timestamp 1700315010
transform 1 0 20250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1065_
timestamp 1700315010
transform -1 0 13650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1066_
timestamp 1700315010
transform 1 0 15150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1067_
timestamp 1700315010
transform 1 0 19050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1068_
timestamp 1700315010
transform -1 0 12450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1069_
timestamp 1700315010
transform 1 0 18150 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1070_
timestamp 1700315010
transform 1 0 28950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1071_
timestamp 1700315010
transform 1 0 23250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1072_
timestamp 1700315010
transform -1 0 2850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1073_
timestamp 1700315010
transform -1 0 13950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1074_
timestamp 1700315010
transform -1 0 11550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1075_
timestamp 1700315010
transform -1 0 11550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1076_
timestamp 1700315010
transform -1 0 14250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1077_
timestamp 1700315010
transform 1 0 16350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1078_
timestamp 1700315010
transform -1 0 7050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1079_
timestamp 1700315010
transform -1 0 13050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1080_
timestamp 1700315010
transform -1 0 12450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1081_
timestamp 1700315010
transform -1 0 2850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1082_
timestamp 1700315010
transform -1 0 15150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1083_
timestamp 1700315010
transform -1 0 10950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1084_
timestamp 1700315010
transform -1 0 5250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1085_
timestamp 1700315010
transform -1 0 4950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1086_
timestamp 1700315010
transform 1 0 9750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1087_
timestamp 1700315010
transform 1 0 7350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1088_
timestamp 1700315010
transform -1 0 9150 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1089_
timestamp 1700315010
transform 1 0 28950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1090_
timestamp 1700315010
transform 1 0 22950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1091_
timestamp 1700315010
transform -1 0 28050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1092_
timestamp 1700315010
transform -1 0 30150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1093_
timestamp 1700315010
transform 1 0 27750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1094_
timestamp 1700315010
transform 1 0 32250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1095_
timestamp 1700315010
transform -1 0 27450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1096_
timestamp 1700315010
transform -1 0 25050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1097_
timestamp 1700315010
transform -1 0 23550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1098_
timestamp 1700315010
transform -1 0 25650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1099_
timestamp 1700315010
transform -1 0 21150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1100_
timestamp 1700315010
transform -1 0 450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1101_
timestamp 1700315010
transform -1 0 450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1102_
timestamp 1700315010
transform -1 0 13650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1103_
timestamp 1700315010
transform 1 0 8850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1104_
timestamp 1700315010
transform 1 0 6750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1105_
timestamp 1700315010
transform 1 0 2250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1106_
timestamp 1700315010
transform -1 0 450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1107_
timestamp 1700315010
transform 1 0 2550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1108_
timestamp 1700315010
transform 1 0 12750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1109_
timestamp 1700315010
transform -1 0 4950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1110_
timestamp 1700315010
transform -1 0 2850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1111_
timestamp 1700315010
transform -1 0 450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1112_
timestamp 1700315010
transform -1 0 30150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1113_
timestamp 1700315010
transform 1 0 6750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1114_
timestamp 1700315010
transform -1 0 26250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1115_
timestamp 1700315010
transform -1 0 7350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1116_
timestamp 1700315010
transform -1 0 9150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1117_
timestamp 1700315010
transform 1 0 10950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1118_
timestamp 1700315010
transform -1 0 4950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1119_
timestamp 1700315010
transform 1 0 7050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1120_
timestamp 1700315010
transform 1 0 6750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1121_
timestamp 1700315010
transform 1 0 13050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1122_
timestamp 1700315010
transform -1 0 10950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1123_
timestamp 1700315010
transform -1 0 9450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1124_
timestamp 1700315010
transform 1 0 7350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1125_
timestamp 1700315010
transform 1 0 2550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1126_
timestamp 1700315010
transform -1 0 450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1127_
timestamp 1700315010
transform 1 0 8250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1128_
timestamp 1700315010
transform -1 0 4650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1129_
timestamp 1700315010
transform -1 0 2850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1130_
timestamp 1700315010
transform 1 0 4950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1131_
timestamp 1700315010
transform -1 0 4950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1132_
timestamp 1700315010
transform -1 0 11850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1133_
timestamp 1700315010
transform -1 0 450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1134_
timestamp 1700315010
transform -1 0 2850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1135_
timestamp 1700315010
transform 1 0 2550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1136_
timestamp 1700315010
transform -1 0 4350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1137_
timestamp 1700315010
transform -1 0 450 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1138_
timestamp 1700315010
transform 1 0 7050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1139_
timestamp 1700315010
transform 1 0 8550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1140_
timestamp 1700315010
transform 1 0 26550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1141_
timestamp 1700315010
transform 1 0 33750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1142_
timestamp 1700315010
transform 1 0 37350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1143_
timestamp 1700315010
transform 1 0 49350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1144_
timestamp 1700315010
transform 1 0 54450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1145_
timestamp 1700315010
transform 1 0 44850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1146_
timestamp 1700315010
transform -1 0 49950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1147_
timestamp 1700315010
transform -1 0 43350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1148_
timestamp 1700315010
transform 1 0 47250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1149_
timestamp 1700315010
transform -1 0 47550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1150_
timestamp 1700315010
transform 1 0 41850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1151_
timestamp 1700315010
transform 1 0 49650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1152_
timestamp 1700315010
transform -1 0 47250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1153_
timestamp 1700315010
transform 1 0 34950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1154_
timestamp 1700315010
transform 1 0 37350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1155_
timestamp 1700315010
transform 1 0 39450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1156_
timestamp 1700315010
transform -1 0 39450 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1157_
timestamp 1700315010
transform -1 0 16350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1158_
timestamp 1700315010
transform 1 0 17250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1159_
timestamp 1700315010
transform -1 0 25650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1160_
timestamp 1700315010
transform 1 0 6450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1161_
timestamp 1700315010
transform 1 0 10950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1162_
timestamp 1700315010
transform 1 0 19650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1163_
timestamp 1700315010
transform 1 0 49350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1164_
timestamp 1700315010
transform 1 0 55950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1165_
timestamp 1700315010
transform -1 0 58350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1166_
timestamp 1700315010
transform 1 0 61950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1167_
timestamp 1700315010
transform 1 0 64050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1168_
timestamp 1700315010
transform -1 0 51750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1169_
timestamp 1700315010
transform 1 0 59850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1170_
timestamp 1700315010
transform 1 0 52050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1171_
timestamp 1700315010
transform 1 0 60450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1172_
timestamp 1700315010
transform 1 0 58350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1173_
timestamp 1700315010
transform 1 0 60450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1174_
timestamp 1700315010
transform 1 0 53550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1175_
timestamp 1700315010
transform -1 0 56250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1176_
timestamp 1700315010
transform 1 0 54450 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1177_
timestamp 1700315010
transform -1 0 44550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1178_
timestamp 1700315010
transform -1 0 44250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1179_
timestamp 1700315010
transform 1 0 49950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1180_
timestamp 1700315010
transform 1 0 31350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1181_
timestamp 1700315010
transform 1 0 49050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1182_
timestamp 1700315010
transform -1 0 59250 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1183_
timestamp 1700315010
transform 1 0 56550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1184_
timestamp 1700315010
transform -1 0 54450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1185_
timestamp 1700315010
transform -1 0 56250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1186_
timestamp 1700315010
transform 1 0 60150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1187_
timestamp 1700315010
transform -1 0 49650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1188_
timestamp 1700315010
transform -1 0 66450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1189_
timestamp 1700315010
transform 1 0 55950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1190_
timestamp 1700315010
transform 1 0 57750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1191_
timestamp 1700315010
transform -1 0 62850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1192_
timestamp 1700315010
transform 1 0 66750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1193_
timestamp 1700315010
transform 1 0 64950 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1194_
timestamp 1700315010
transform 1 0 62850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1195_
timestamp 1700315010
transform 1 0 66750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1196_
timestamp 1700315010
transform 1 0 58350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1197_
timestamp 1700315010
transform -1 0 61050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1198_
timestamp 1700315010
transform 1 0 46350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1199_
timestamp 1700315010
transform 1 0 41550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1200_
timestamp 1700315010
transform 1 0 52050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1201_
timestamp 1700315010
transform -1 0 56250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1202_
timestamp 1700315010
transform 1 0 60450 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1203_
timestamp 1700315010
transform 1 0 52650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1204_
timestamp 1700315010
transform -1 0 55350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1205_
timestamp 1700315010
transform 1 0 39750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1206_
timestamp 1700315010
transform -1 0 450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1207_
timestamp 1700315010
transform 1 0 11250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1208_
timestamp 1700315010
transform -1 0 450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1209_
timestamp 1700315010
transform 1 0 35250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1210_
timestamp 1700315010
transform -1 0 22950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1211_
timestamp 1700315010
transform -1 0 32250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1212_
timestamp 1700315010
transform 1 0 27150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1213_
timestamp 1700315010
transform 1 0 31050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1214_
timestamp 1700315010
transform 1 0 32850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1215_
timestamp 1700315010
transform -1 0 20550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1216_
timestamp 1700315010
transform -1 0 29250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1217_
timestamp 1700315010
transform 1 0 29550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1218_
timestamp 1700315010
transform -1 0 26850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1219_
timestamp 1700315010
transform 1 0 18150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1220_
timestamp 1700315010
transform -1 0 2850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1221_
timestamp 1700315010
transform -1 0 22650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1222_
timestamp 1700315010
transform -1 0 28350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1223_
timestamp 1700315010
transform 1 0 26550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1224_
timestamp 1700315010
transform -1 0 31350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1225_
timestamp 1700315010
transform 1 0 28650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1226_
timestamp 1700315010
transform -1 0 24750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1227_
timestamp 1700315010
transform 1 0 23250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1228_
timestamp 1700315010
transform 1 0 29250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1229_
timestamp 1700315010
transform 1 0 33150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1230_
timestamp 1700315010
transform 1 0 27450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1231_
timestamp 1700315010
transform -1 0 25350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1232_
timestamp 1700315010
transform 1 0 11250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1233_
timestamp 1700315010
transform 1 0 4350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1234_
timestamp 1700315010
transform 1 0 16350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1235_
timestamp 1700315010
transform 1 0 13650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1236_
timestamp 1700315010
transform -1 0 4050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1237_
timestamp 1700315010
transform 1 0 8250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1238_
timestamp 1700315010
transform 1 0 10950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1239_
timestamp 1700315010
transform -1 0 7350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1240_
timestamp 1700315010
transform -1 0 6150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1241_
timestamp 1700315010
transform -1 0 3150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1242_
timestamp 1700315010
transform 1 0 9150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1243_
timestamp 1700315010
transform 1 0 4950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1244_
timestamp 1700315010
transform 1 0 2550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1245_
timestamp 1700315010
transform -1 0 2850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1246_
timestamp 1700315010
transform -1 0 450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1247_
timestamp 1700315010
transform -1 0 450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1248_
timestamp 1700315010
transform 1 0 8250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1249_
timestamp 1700315010
transform 1 0 150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1250_
timestamp 1700315010
transform -1 0 2850 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1251_
timestamp 1700315010
transform -1 0 16350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1252_
timestamp 1700315010
transform 1 0 6750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1253_
timestamp 1700315010
transform 1 0 150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1254_
timestamp 1700315010
transform -1 0 9450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1255_
timestamp 1700315010
transform -1 0 450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1256_
timestamp 1700315010
transform 1 0 4650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1257_
timestamp 1700315010
transform -1 0 13950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1258_
timestamp 1700315010
transform 1 0 4950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1259_
timestamp 1700315010
transform -1 0 12150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1260_
timestamp 1700315010
transform -1 0 12150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1261_
timestamp 1700315010
transform 1 0 13950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1262_
timestamp 1700315010
transform 1 0 2550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1263_
timestamp 1700315010
transform -1 0 10050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1264_
timestamp 1700315010
transform 1 0 7050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1265_
timestamp 1700315010
transform -1 0 9750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1266_
timestamp 1700315010
transform -1 0 9450 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1267_
timestamp 1700315010
transform -1 0 5250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1268_
timestamp 1700315010
transform 1 0 15750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1269_
timestamp 1700315010
transform 1 0 18150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1270_
timestamp 1700315010
transform 1 0 34950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1271_
timestamp 1700315010
transform -1 0 46050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1272_
timestamp 1700315010
transform 1 0 74550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1273_
timestamp 1700315010
transform -1 0 70950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1274_
timestamp 1700315010
transform 1 0 61950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1275_
timestamp 1700315010
transform 1 0 58950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1276_
timestamp 1700315010
transform -1 0 66750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1277_
timestamp 1700315010
transform 1 0 61350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1278_
timestamp 1700315010
transform 1 0 70950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1279_
timestamp 1700315010
transform 1 0 70350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1280_
timestamp 1700315010
transform -1 0 52950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1281_
timestamp 1700315010
transform -1 0 57450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1282_
timestamp 1700315010
transform -1 0 60750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1283_
timestamp 1700315010
transform -1 0 55050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1284_
timestamp 1700315010
transform -1 0 24450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1285_
timestamp 1700315010
transform -1 0 48750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1286_
timestamp 1700315010
transform -1 0 22350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1287_
timestamp 1700315010
transform 1 0 28050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1288_
timestamp 1700315010
transform 1 0 44550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1289_
timestamp 1700315010
transform 1 0 42150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1290_
timestamp 1700315010
transform -1 0 46950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1291_
timestamp 1700315010
transform -1 0 35550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1292_
timestamp 1700315010
transform -1 0 33450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1293_
timestamp 1700315010
transform -1 0 39150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1294_
timestamp 1700315010
transform 1 0 18450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1295_
timestamp 1700315010
transform 1 0 16350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1296_
timestamp 1700315010
transform -1 0 24450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1297_
timestamp 1700315010
transform 1 0 23850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1298_
timestamp 1700315010
transform 1 0 4650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1299_
timestamp 1700315010
transform 1 0 11250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1300_
timestamp 1700315010
transform -1 0 23850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1301_
timestamp 1700315010
transform 1 0 30450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1302_
timestamp 1700315010
transform -1 0 28350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1303_
timestamp 1700315010
transform -1 0 30750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1304_
timestamp 1700315010
transform -1 0 25950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1305_
timestamp 1700315010
transform -1 0 20850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1306_
timestamp 1700315010
transform 1 0 11250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1307_
timestamp 1700315010
transform 1 0 4950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1308_
timestamp 1700315010
transform -1 0 450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1309_
timestamp 1700315010
transform 1 0 19350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1310_
timestamp 1700315010
transform 1 0 23850 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1311_
timestamp 1700315010
transform 1 0 16050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1312_
timestamp 1700315010
transform -1 0 25950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1313_
timestamp 1700315010
transform -1 0 19950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1314_
timestamp 1700315010
transform -1 0 18150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1315_
timestamp 1700315010
transform 1 0 19050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1316_
timestamp 1700315010
transform -1 0 11250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1317_
timestamp 1700315010
transform 1 0 13950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1318_
timestamp 1700315010
transform 1 0 41250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1319_
timestamp 1700315010
transform -1 0 30450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1320_
timestamp 1700315010
transform -1 0 26250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1321_
timestamp 1700315010
transform -1 0 23850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1322_
timestamp 1700315010
transform -1 0 16950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1323_
timestamp 1700315010
transform -1 0 21750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1324_
timestamp 1700315010
transform -1 0 11850 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1325_
timestamp 1700315010
transform -1 0 14850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1326_
timestamp 1700315010
transform -1 0 9750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1327_
timestamp 1700315010
transform -1 0 450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1328_
timestamp 1700315010
transform -1 0 450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1329_
timestamp 1700315010
transform 1 0 9150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1330_
timestamp 1700315010
transform -1 0 7050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1331_
timestamp 1700315010
transform 1 0 2250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1332_
timestamp 1700315010
transform 1 0 6750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1333_
timestamp 1700315010
transform 1 0 11550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1334_
timestamp 1700315010
transform 1 0 7050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1335_
timestamp 1700315010
transform -1 0 450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1336_
timestamp 1700315010
transform 1 0 6750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1337_
timestamp 1700315010
transform 1 0 16350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1338_
timestamp 1700315010
transform 1 0 150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1339_
timestamp 1700315010
transform 1 0 10350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1340_
timestamp 1700315010
transform 1 0 9150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1341_
timestamp 1700315010
transform 1 0 1950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1342_
timestamp 1700315010
transform -1 0 2550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1343_
timestamp 1700315010
transform 1 0 4350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1344_
timestamp 1700315010
transform -1 0 12750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1345_
timestamp 1700315010
transform -1 0 22050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1346_
timestamp 1700315010
transform 1 0 13050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1347_
timestamp 1700315010
transform 1 0 14850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1348_
timestamp 1700315010
transform -1 0 19950 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1349_
timestamp 1700315010
transform -1 0 20550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1350_
timestamp 1700315010
transform 1 0 7350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1351_
timestamp 1700315010
transform 1 0 14250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1352_
timestamp 1700315010
transform 1 0 25650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1353_
timestamp 1700315010
transform -1 0 17550 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1354_
timestamp 1700315010
transform 1 0 25050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1355_
timestamp 1700315010
transform -1 0 31950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1356_
timestamp 1700315010
transform 1 0 48750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1357_
timestamp 1700315010
transform 1 0 51150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1358_
timestamp 1700315010
transform 1 0 53250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1359_
timestamp 1700315010
transform 1 0 67950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_0__1360_
timestamp 1700315010
transform 1 0 67050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1361_
timestamp 1700315010
transform -1 0 62850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1362_
timestamp 1700315010
transform 1 0 64650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1363_
timestamp 1700315010
transform -1 0 60450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1364_
timestamp 1700315010
transform 1 0 58050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1365_
timestamp 1700315010
transform -1 0 71850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1366_
timestamp 1700315010
transform -1 0 22950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1367_
timestamp 1700315010
transform 1 0 20550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1368_
timestamp 1700315010
transform 1 0 31050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1369_
timestamp 1700315010
transform 1 0 43350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1370_
timestamp 1700315010
transform 1 0 33750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1371_
timestamp 1700315010
transform 1 0 37050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1372_
timestamp 1700315010
transform -1 0 18750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1373_
timestamp 1700315010
transform 1 0 14250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1374_
timestamp 1700315010
transform -1 0 7350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1375_
timestamp 1700315010
transform -1 0 4650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1376_
timestamp 1700315010
transform -1 0 19050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1377_
timestamp 1700315010
transform -1 0 12750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1378_
timestamp 1700315010
transform -1 0 17250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1379_
timestamp 1700315010
transform -1 0 15150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1380_
timestamp 1700315010
transform -1 0 16950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1381_
timestamp 1700315010
transform -1 0 14550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1382_
timestamp 1700315010
transform -1 0 10650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1383_
timestamp 1700315010
transform -1 0 14550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1384_
timestamp 1700315010
transform -1 0 16950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1385_
timestamp 1700315010
transform -1 0 12150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1386_
timestamp 1700315010
transform -1 0 3150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1387_
timestamp 1700315010
transform 1 0 8850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1388_
timestamp 1700315010
transform 1 0 23250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1389_
timestamp 1700315010
transform -1 0 26850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1390_
timestamp 1700315010
transform -1 0 24750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1391_
timestamp 1700315010
transform -1 0 22050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1392_
timestamp 1700315010
transform 1 0 30150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1393_
timestamp 1700315010
transform 1 0 27750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1394_
timestamp 1700315010
transform 1 0 20250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1395_
timestamp 1700315010
transform 1 0 5850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1396_
timestamp 1700315010
transform -1 0 8250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1397_
timestamp 1700315010
transform -1 0 450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1398_
timestamp 1700315010
transform -1 0 4650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1399_
timestamp 1700315010
transform -1 0 9750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1400_
timestamp 1700315010
transform -1 0 4050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1401_
timestamp 1700315010
transform -1 0 450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1402_
timestamp 1700315010
transform -1 0 1950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1403_
timestamp 1700315010
transform 1 0 4650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1404_
timestamp 1700315010
transform -1 0 7050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1405_
timestamp 1700315010
transform 1 0 4650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1406_
timestamp 1700315010
transform -1 0 450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1407_
timestamp 1700315010
transform -1 0 450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1408_
timestamp 1700315010
transform -1 0 5250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1409_
timestamp 1700315010
transform -1 0 2850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1410_
timestamp 1700315010
transform 1 0 2550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1411_
timestamp 1700315010
transform -1 0 5250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1412_
timestamp 1700315010
transform 1 0 8850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1413_
timestamp 1700315010
transform -1 0 450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1414_
timestamp 1700315010
transform -1 0 9150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1415_
timestamp 1700315010
transform -1 0 19050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1416_
timestamp 1700315010
transform 1 0 28050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1417_
timestamp 1700315010
transform 1 0 15450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1418_
timestamp 1700315010
transform -1 0 17850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1419_
timestamp 1700315010
transform 1 0 19950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1420_
timestamp 1700315010
transform -1 0 36750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1421_
timestamp 1700315010
transform -1 0 36450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1422_
timestamp 1700315010
transform 1 0 41250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1423_
timestamp 1700315010
transform -1 0 38850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1424_
timestamp 1700315010
transform 1 0 42450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1425_
timestamp 1700315010
transform -1 0 44550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1426_
timestamp 1700315010
transform 1 0 46350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1427_
timestamp 1700315010
transform 1 0 68550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1428_
timestamp 1700315010
transform -1 0 64050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1429_
timestamp 1700315010
transform 1 0 64650 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1430_
timestamp 1700315010
transform 1 0 67050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1431_
timestamp 1700315010
transform -1 0 70350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1432_
timestamp 1700315010
transform 1 0 70650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1433_
timestamp 1700315010
transform -1 0 64950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1434_
timestamp 1700315010
transform 1 0 69150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_0__1435_
timestamp 1700315010
transform 1 0 88650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1436_
timestamp 1700315010
transform -1 0 86250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1437_
timestamp 1700315010
transform -1 0 57750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1438_
timestamp 1700315010
transform 1 0 39450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1439_
timestamp 1700315010
transform 1 0 18750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1440_
timestamp 1700315010
transform -1 0 17550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1441_
timestamp 1700315010
transform 1 0 7050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1442_
timestamp 1700315010
transform 1 0 26850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1443_
timestamp 1700315010
transform -1 0 30750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1444_
timestamp 1700315010
transform -1 0 20850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1445_
timestamp 1700315010
transform -1 0 25650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1446_
timestamp 1700315010
transform 1 0 22650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1447_
timestamp 1700315010
transform 1 0 24750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1448_
timestamp 1700315010
transform 1 0 26550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1449_
timestamp 1700315010
transform -1 0 28350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1450_
timestamp 1700315010
transform -1 0 22950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1451_
timestamp 1700315010
transform 1 0 24450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1452_
timestamp 1700315010
transform 1 0 28050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1453_
timestamp 1700315010
transform 1 0 30750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1454_
timestamp 1700315010
transform 1 0 28350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1455_
timestamp 1700315010
transform 1 0 42750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1456_
timestamp 1700315010
transform -1 0 31950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1457_
timestamp 1700315010
transform -1 0 28950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1458_
timestamp 1700315010
transform -1 0 23850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1459_
timestamp 1700315010
transform -1 0 6750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1460_
timestamp 1700315010
transform 1 0 25650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1461_
timestamp 1700315010
transform 1 0 10650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1462_
timestamp 1700315010
transform -1 0 2250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1463_
timestamp 1700315010
transform -1 0 21150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1464_
timestamp 1700315010
transform -1 0 13050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1465_
timestamp 1700315010
transform -1 0 15150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1466_
timestamp 1700315010
transform -1 0 8550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1467_
timestamp 1700315010
transform -1 0 19350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1468_
timestamp 1700315010
transform 1 0 21150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1469_
timestamp 1700315010
transform -1 0 16350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1470_
timestamp 1700315010
transform -1 0 13050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1471_
timestamp 1700315010
transform 1 0 11250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1472_
timestamp 1700315010
transform 1 0 13650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1473_
timestamp 1700315010
transform 1 0 18150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1474_
timestamp 1700315010
transform 1 0 41250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1475_
timestamp 1700315010
transform 1 0 40650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1476_
timestamp 1700315010
transform 1 0 44250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1477_
timestamp 1700315010
transform 1 0 46650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1478_
timestamp 1700315010
transform 1 0 48150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1479_
timestamp 1700315010
transform 1 0 52350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1480_
timestamp 1700315010
transform -1 0 63150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1481_
timestamp 1700315010
transform -1 0 64950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1482_
timestamp 1700315010
transform 1 0 69150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1483_
timestamp 1700315010
transform 1 0 80250 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1484_
timestamp 1700315010
transform -1 0 82350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1485_
timestamp 1700315010
transform 1 0 82050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1486_
timestamp 1700315010
transform -1 0 84750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1487_
timestamp 1700315010
transform 1 0 86850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1488_
timestamp 1700315010
transform 1 0 32250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1489_
timestamp 1700315010
transform 1 0 34650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1490_
timestamp 1700315010
transform -1 0 34950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1491_
timestamp 1700315010
transform -1 0 42750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1492_
timestamp 1700315010
transform -1 0 31350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1493_
timestamp 1700315010
transform -1 0 33450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1494_
timestamp 1700315010
transform 1 0 37950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1495_
timestamp 1700315010
transform 1 0 44250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1496_
timestamp 1700315010
transform 1 0 35550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1497_
timestamp 1700315010
transform 1 0 38550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1498_
timestamp 1700315010
transform 1 0 40650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1499_
timestamp 1700315010
transform 1 0 32850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1500_
timestamp 1700315010
transform 1 0 36150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1501_
timestamp 1700315010
transform 1 0 40350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1502_
timestamp 1700315010
transform 1 0 40650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1503_
timestamp 1700315010
transform 1 0 41250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1504_
timestamp 1700315010
transform 1 0 42450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1505_
timestamp 1700315010
transform -1 0 36450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1506_
timestamp 1700315010
transform -1 0 39150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1507_
timestamp 1700315010
transform -1 0 36750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1508_
timestamp 1700315010
transform -1 0 32850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1509_
timestamp 1700315010
transform 1 0 30150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1510_
timestamp 1700315010
transform -1 0 28350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1511_
timestamp 1700315010
transform 1 0 34350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1512_
timestamp 1700315010
transform -1 0 40350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1513_
timestamp 1700315010
transform 1 0 49350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1514_
timestamp 1700315010
transform -1 0 45450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1515_
timestamp 1700315010
transform 1 0 46950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1516_
timestamp 1700315010
transform -1 0 37650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1517_
timestamp 1700315010
transform 1 0 42750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1518_
timestamp 1700315010
transform -1 0 47850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1519_
timestamp 1700315010
transform 1 0 43350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1520_
timestamp 1700315010
transform 1 0 45450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1521_
timestamp 1700315010
transform 1 0 37950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1522_
timestamp 1700315010
transform 1 0 40350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1523_
timestamp 1700315010
transform 1 0 42150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1524_
timestamp 1700315010
transform 1 0 49050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1525_
timestamp 1700315010
transform -1 0 81750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1526_
timestamp 1700315010
transform -1 0 74250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1527_
timestamp 1700315010
transform 1 0 66750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1528_
timestamp 1700315010
transform 1 0 64350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1529_
timestamp 1700315010
transform 1 0 68250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1530_
timestamp 1700315010
transform -1 0 72450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1531_
timestamp 1700315010
transform -1 0 75750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1532_
timestamp 1700315010
transform 1 0 77850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1533_
timestamp 1700315010
transform -1 0 79950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1534_
timestamp 1700315010
transform -1 0 76950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1535_
timestamp 1700315010
transform -1 0 55950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1536_
timestamp 1700315010
transform 1 0 47250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1537_
timestamp 1700315010
transform 1 0 41550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1538_
timestamp 1700315010
transform 1 0 38250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1539_
timestamp 1700315010
transform 1 0 34050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1540_
timestamp 1700315010
transform -1 0 39150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1541_
timestamp 1700315010
transform -1 0 41550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1542_
timestamp 1700315010
transform -1 0 36750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1543_
timestamp 1700315010
transform 1 0 39150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1544_
timestamp 1700315010
transform 1 0 36150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1545_
timestamp 1700315010
transform -1 0 36750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1546_
timestamp 1700315010
transform -1 0 37050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1547_
timestamp 1700315010
transform -1 0 39750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1548_
timestamp 1700315010
transform -1 0 45150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1549_
timestamp 1700315010
transform -1 0 41850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1550_
timestamp 1700315010
transform 1 0 51450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1551_
timestamp 1700315010
transform 1 0 58050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1552_
timestamp 1700315010
transform 1 0 62250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1553_
timestamp 1700315010
transform -1 0 75450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1554_
timestamp 1700315010
transform 1 0 77850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1555_
timestamp 1700315010
transform 1 0 77550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1556_
timestamp 1700315010
transform -1 0 74250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1557_
timestamp 1700315010
transform -1 0 72450 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1558_
timestamp 1700315010
transform 1 0 37350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1559_
timestamp 1700315010
transform 1 0 52350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1560_
timestamp 1700315010
transform 1 0 54150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1561_
timestamp 1700315010
transform -1 0 40050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1562_
timestamp 1700315010
transform 1 0 39750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1563_
timestamp 1700315010
transform 1 0 55050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1564_
timestamp 1700315010
transform -1 0 30450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1565_
timestamp 1700315010
transform -1 0 31950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1566_
timestamp 1700315010
transform -1 0 34050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1567_
timestamp 1700315010
transform 1 0 43050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1568_
timestamp 1700315010
transform 1 0 49350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1569_
timestamp 1700315010
transform 1 0 58650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1570_
timestamp 1700315010
transform 1 0 49950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1571_
timestamp 1700315010
transform -1 0 53850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1572_
timestamp 1700315010
transform 1 0 51150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1573_
timestamp 1700315010
transform 1 0 61050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1574_
timestamp 1700315010
transform -1 0 60450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1575_
timestamp 1700315010
transform 1 0 64350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1576_
timestamp 1700315010
transform 1 0 61950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1577_
timestamp 1700315010
transform 1 0 66450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1578_
timestamp 1700315010
transform 1 0 85050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1579_
timestamp 1700315010
transform -1 0 76350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1580_
timestamp 1700315010
transform -1 0 75750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1581_
timestamp 1700315010
transform 1 0 72750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1582_
timestamp 1700315010
transform -1 0 67050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1583_
timestamp 1700315010
transform -1 0 56850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1584_
timestamp 1700315010
transform 1 0 43650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1585_
timestamp 1700315010
transform 1 0 46050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1586_
timestamp 1700315010
transform 1 0 53850 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1587_
timestamp 1700315010
transform 1 0 37650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1588_
timestamp 1700315010
transform -1 0 57450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1589_
timestamp 1700315010
transform 1 0 73650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1590_
timestamp 1700315010
transform 1 0 71250 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0__1591_
timestamp 1700315010
transform -1 0 70650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_0__1592_
timestamp 1700315010
transform -1 0 64650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1593_
timestamp 1700315010
transform -1 0 64650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0__1594_
timestamp 1700315010
transform 1 0 64050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1595_
timestamp 1700315010
transform 1 0 59250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1596_
timestamp 1700315010
transform -1 0 61650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1597_
timestamp 1700315010
transform 1 0 59550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1598_
timestamp 1700315010
transform -1 0 61950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1599_
timestamp 1700315010
transform -1 0 58050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1600_
timestamp 1700315010
transform -1 0 59850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1601_
timestamp 1700315010
transform 1 0 49050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1602_
timestamp 1700315010
transform -1 0 49650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1603_
timestamp 1700315010
transform 1 0 43650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1604_
timestamp 1700315010
transform -1 0 46050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1605_
timestamp 1700315010
transform -1 0 66750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1606_
timestamp 1700315010
transform -1 0 76950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1607_
timestamp 1700315010
transform 1 0 65850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1608_
timestamp 1700315010
transform -1 0 68250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1636_
timestamp 1700315010
transform -1 0 88050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1637_
timestamp 1700315010
transform 1 0 88050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1638_
timestamp 1700315010
transform -1 0 79950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1639_
timestamp 1700315010
transform 1 0 77550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1640_
timestamp 1700315010
transform 1 0 77550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1641_
timestamp 1700315010
transform -1 0 55950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1642_
timestamp 1700315010
transform -1 0 46950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1643_
timestamp 1700315010
transform -1 0 44550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1644_
timestamp 1700315010
transform -1 0 57450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1645_
timestamp 1700315010
transform -1 0 65550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1646_
timestamp 1700315010
transform -1 0 61050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1647_
timestamp 1700315010
transform 1 0 46950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1648_
timestamp 1700315010
transform 1 0 86250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1649_
timestamp 1700315010
transform -1 0 63750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1650_
timestamp 1700315010
transform -1 0 66150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1651_
timestamp 1700315010
transform 1 0 64050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1652_
timestamp 1700315010
transform -1 0 53850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1653_
timestamp 1700315010
transform 1 0 61650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1654_
timestamp 1700315010
transform 1 0 86550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1655_
timestamp 1700315010
transform -1 0 84450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1656_
timestamp 1700315010
transform 1 0 88350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1657_
timestamp 1700315010
transform 1 0 86250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1658_
timestamp 1700315010
transform 1 0 83850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1659_
timestamp 1700315010
transform -1 0 79650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1660_
timestamp 1700315010
transform -1 0 82350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1661_
timestamp 1700315010
transform 1 0 79650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1662_
timestamp 1700315010
transform -1 0 51450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1663_
timestamp 1700315010
transform -1 0 49050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1664_
timestamp 1700315010
transform -1 0 51150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1665_
timestamp 1700315010
transform -1 0 54150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1666_
timestamp 1700315010
transform -1 0 56850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1667_
timestamp 1700315010
transform 1 0 57150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1668_
timestamp 1700315010
transform 1 0 55050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1669_
timestamp 1700315010
transform -1 0 60150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1670_
timestamp 1700315010
transform 1 0 62250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1671_
timestamp 1700315010
transform 1 0 77850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1672_
timestamp 1700315010
transform -1 0 84450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1673_
timestamp 1700315010
transform 1 0 81750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1674_
timestamp 1700315010
transform -1 0 79950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1675_
timestamp 1700315010
transform -1 0 82650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1676_
timestamp 1700315010
transform 1 0 81750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1677_
timestamp 1700315010
transform -1 0 72750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1678_
timestamp 1700315010
transform -1 0 73350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1679_
timestamp 1700315010
transform -1 0 67350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1680_
timestamp 1700315010
transform 1 0 68850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1681_
timestamp 1700315010
transform -1 0 59550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1682_
timestamp 1700315010
transform 1 0 68250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1683_
timestamp 1700315010
transform 1 0 70050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1684_
timestamp 1700315010
transform 1 0 74850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1685_
timestamp 1700315010
transform -1 0 62250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1686_
timestamp 1700315010
transform 1 0 64050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1687_
timestamp 1700315010
transform -1 0 76050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1688_
timestamp 1700315010
transform 1 0 77850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1689_
timestamp 1700315010
transform 1 0 72750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1690_
timestamp 1700315010
transform 1 0 75750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1691_
timestamp 1700315010
transform -1 0 73650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1692_
timestamp 1700315010
transform 1 0 53250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1693_
timestamp 1700315010
transform 1 0 46050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1694_
timestamp 1700315010
transform -1 0 48750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1695_
timestamp 1700315010
transform -1 0 43650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1696_
timestamp 1700315010
transform -1 0 45150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1697_
timestamp 1700315010
transform -1 0 49050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1698_
timestamp 1700315010
transform 1 0 51150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1699_
timestamp 1700315010
transform -1 0 57750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1700_
timestamp 1700315010
transform -1 0 58050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1701_
timestamp 1700315010
transform -1 0 53550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1702_
timestamp 1700315010
transform 1 0 55350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1703_
timestamp 1700315010
transform -1 0 68250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1704_
timestamp 1700315010
transform -1 0 71550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1705_
timestamp 1700315010
transform 1 0 60150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1706_
timestamp 1700315010
transform -1 0 64650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1707_
timestamp 1700315010
transform -1 0 66750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1708_
timestamp 1700315010
transform 1 0 66750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1709_
timestamp 1700315010
transform -1 0 54450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1710_
timestamp 1700315010
transform -1 0 57750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1711_
timestamp 1700315010
transform -1 0 52950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1712_
timestamp 1700315010
transform -1 0 55050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1713_
timestamp 1700315010
transform -1 0 50550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1714_
timestamp 1700315010
transform 1 0 56250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1715_
timestamp 1700315010
transform -1 0 58650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1716_
timestamp 1700315010
transform 1 0 60750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1717_
timestamp 1700315010
transform -1 0 66150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1718_
timestamp 1700315010
transform 1 0 67950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1719_
timestamp 1700315010
transform 1 0 70350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1720_
timestamp 1700315010
transform 1 0 63150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1721_
timestamp 1700315010
transform 1 0 69450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1722_
timestamp 1700315010
transform 1 0 70950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1723_
timestamp 1700315010
transform 1 0 71550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0__1724_
timestamp 1700315010
transform -1 0 71550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1725_
timestamp 1700315010
transform 1 0 65850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1726_
timestamp 1700315010
transform -1 0 63750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1727_
timestamp 1700315010
transform -1 0 65250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1728_
timestamp 1700315010
transform -1 0 44850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0__1729_
timestamp 1700315010
transform 1 0 45750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1730_
timestamp 1700315010
transform -1 0 48150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1731_
timestamp 1700315010
transform -1 0 50250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1732_
timestamp 1700315010
transform 1 0 52650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1733_
timestamp 1700315010
transform 1 0 54750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1734_
timestamp 1700315010
transform 1 0 73950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1735_
timestamp 1700315010
transform 1 0 73350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1736_
timestamp 1700315010
transform -1 0 78150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1737_
timestamp 1700315010
transform 1 0 75450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1738_
timestamp 1700315010
transform 1 0 76050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1739_
timestamp 1700315010
transform 1 0 73350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1740_
timestamp 1700315010
transform -1 0 76950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1741_
timestamp 1700315010
transform 1 0 77850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1742_
timestamp 1700315010
transform 1 0 52350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1743_
timestamp 1700315010
transform -1 0 41250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1744_
timestamp 1700315010
transform -1 0 43650 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1745_
timestamp 1700315010
transform -1 0 48150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1746_
timestamp 1700315010
transform 1 0 45450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1747_
timestamp 1700315010
transform 1 0 49950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1748_
timestamp 1700315010
transform -1 0 76050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1749_
timestamp 1700315010
transform 1 0 77850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1750_
timestamp 1700315010
transform 1 0 81150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1751_
timestamp 1700315010
transform 1 0 80250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1752_
timestamp 1700315010
transform -1 0 78750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1753_
timestamp 1700315010
transform 1 0 80250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1754_
timestamp 1700315010
transform 1 0 76950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_0__1755_
timestamp 1700315010
transform 1 0 80250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1756_
timestamp 1700315010
transform 1 0 72150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1757_
timestamp 1700315010
transform -1 0 65550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1758_
timestamp 1700315010
transform 1 0 63150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1759_
timestamp 1700315010
transform 1 0 59550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1760_
timestamp 1700315010
transform 1 0 67350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1761_
timestamp 1700315010
transform -1 0 70050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1762_
timestamp 1700315010
transform -1 0 76650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1763_
timestamp 1700315010
transform 1 0 78750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1764_
timestamp 1700315010
transform 1 0 83550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1765_
timestamp 1700315010
transform 1 0 85650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1766_
timestamp 1700315010
transform 1 0 87150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1767_
timestamp 1700315010
transform 1 0 73050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1768_
timestamp 1700315010
transform -1 0 70950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1769_
timestamp 1700315010
transform -1 0 68550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1770_
timestamp 1700315010
transform -1 0 74850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1771_
timestamp 1700315010
transform 1 0 82350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1772_
timestamp 1700315010
transform 1 0 82650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1773_
timestamp 1700315010
transform -1 0 86850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_0__1774_
timestamp 1700315010
transform -1 0 83550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1775_
timestamp 1700315010
transform -1 0 85350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1776_
timestamp 1700315010
transform 1 0 85350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1777_
timestamp 1700315010
transform 1 0 73650 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1778_
timestamp 1700315010
transform 1 0 66750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1779_
timestamp 1700315010
transform 1 0 64950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1780_
timestamp 1700315010
transform 1 0 62250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1781_
timestamp 1700315010
transform 1 0 69150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1782_
timestamp 1700315010
transform 1 0 71550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1783_
timestamp 1700315010
transform 1 0 83850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1784_
timestamp 1700315010
transform 1 0 81750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1785_
timestamp 1700315010
transform -1 0 86850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1786_
timestamp 1700315010
transform 1 0 88950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1787_
timestamp 1700315010
transform -1 0 88050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1788_
timestamp 1700315010
transform 1 0 85350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1789_
timestamp 1700315010
transform 1 0 89550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1790_
timestamp 1700315010
transform 1 0 89550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1791_
timestamp 1700315010
transform 1 0 89250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0__1792_
timestamp 1700315010
transform 1 0 69450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1793_
timestamp 1700315010
transform 1 0 67350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1794_
timestamp 1700315010
transform 1 0 72750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1795_
timestamp 1700315010
transform -1 0 83250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1796_
timestamp 1700315010
transform 1 0 80850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1797_
timestamp 1700315010
transform -1 0 75150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1798_
timestamp 1700315010
transform -1 0 87750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0__1799_
timestamp 1700315010
transform -1 0 87750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0__1800_
timestamp 1700315010
transform -1 0 87450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1801_
timestamp 1700315010
transform 1 0 80850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1802_
timestamp 1700315010
transform 1 0 70950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0__1803_
timestamp 1700315010
transform 1 0 87750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1804_
timestamp 1700315010
transform -1 0 88050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1805_
timestamp 1700315010
transform 1 0 89550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1806_
timestamp 1700315010
transform -1 0 85050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0__1807_
timestamp 1700315010
transform 1 0 84750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1808_
timestamp 1700315010
transform 1 0 82650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1809_
timestamp 1700315010
transform 1 0 84150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_0__1810_
timestamp 1700315010
transform 1 0 88050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_0__1811_
timestamp 1700315010
transform 1 0 85650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_0__1812_
timestamp 1700315010
transform 1 0 89250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0__1813_
timestamp 1700315010
transform -1 0 89550 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0__1814_
timestamp 1700315010
transform -1 0 89850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1815_
timestamp 1700315010
transform 1 0 87150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0__1816_
timestamp 1700315010
transform -1 0 89550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1817_
timestamp 1700315010
transform -1 0 87750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0__1818_
timestamp 1700315010
transform -1 0 48750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1819_
timestamp 1700315010
transform -1 0 38550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0__1820_
timestamp 1700315010
transform -1 0 68850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_0__1821_
timestamp 1700315010
transform -1 0 84150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1822_
timestamp 1700315010
transform 1 0 81750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1823_
timestamp 1700315010
transform 1 0 79950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1824_
timestamp 1700315010
transform 1 0 74250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1825_
timestamp 1700315010
transform 1 0 68550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0__1826_
timestamp 1700315010
transform 1 0 85950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert0
timestamp 1700315010
transform 1 0 58650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert1
timestamp 1700315010
transform -1 0 32850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert2
timestamp 1700315010
transform -1 0 34650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert3
timestamp 1700315010
transform -1 0 33750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert4
timestamp 1700315010
transform -1 0 65850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert5
timestamp 1700315010
transform -1 0 56250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert6
timestamp 1700315010
transform -1 0 40650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert7
timestamp 1700315010
transform -1 0 50850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert13
timestamp 1700315010
transform 1 0 77550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert14
timestamp 1700315010
transform -1 0 57150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert15
timestamp 1700315010
transform -1 0 64950 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert16
timestamp 1700315010
transform -1 0 60150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert17
timestamp 1700315010
transform 1 0 37650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert18
timestamp 1700315010
transform -1 0 34950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert19
timestamp 1700315010
transform 1 0 45150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert20
timestamp 1700315010
transform -1 0 36150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert21
timestamp 1700315010
transform 1 0 79650 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert22
timestamp 1700315010
transform -1 0 62850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert23
timestamp 1700315010
transform 1 0 63450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert24
timestamp 1700315010
transform 1 0 79050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert25
timestamp 1700315010
transform -1 0 34950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert26
timestamp 1700315010
transform -1 0 39450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert27
timestamp 1700315010
transform -1 0 35850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert28
timestamp 1700315010
transform 1 0 47250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert29
timestamp 1700315010
transform -1 0 32550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert30
timestamp 1700315010
transform 1 0 50550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert31
timestamp 1700315010
transform -1 0 32850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert32
timestamp 1700315010
transform 1 0 52350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert33
timestamp 1700315010
transform -1 0 76050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert34
timestamp 1700315010
transform -1 0 89850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert35
timestamp 1700315010
transform -1 0 73950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_0_BUFX2_insert36
timestamp 1700315010
transform -1 0 88950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1700315010
transform -1 0 67950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 73950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 86850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1700315010
transform -1 0 77550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 74250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__889_
timestamp 1700315010
transform 1 0 80250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__890_
timestamp 1700315010
transform -1 0 74550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__891_
timestamp 1700315010
transform -1 0 76650 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__892_
timestamp 1700315010
transform 1 0 80550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__893_
timestamp 1700315010
transform -1 0 78450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__894_
timestamp 1700315010
transform 1 0 82350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__895_
timestamp 1700315010
transform -1 0 78750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__896_
timestamp 1700315010
transform -1 0 76650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__897_
timestamp 1700315010
transform 1 0 76650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__898_
timestamp 1700315010
transform -1 0 82350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__899_
timestamp 1700315010
transform 1 0 78750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__900_
timestamp 1700315010
transform -1 0 87750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__901_
timestamp 1700315010
transform -1 0 85650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__902_
timestamp 1700315010
transform 1 0 86850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__903_
timestamp 1700315010
transform 1 0 73350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__904_
timestamp 1700315010
transform -1 0 80250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__905_
timestamp 1700315010
transform -1 0 85350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__906_
timestamp 1700315010
transform -1 0 63150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__907_
timestamp 1700315010
transform 1 0 74850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__908_
timestamp 1700315010
transform 1 0 89250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__909_
timestamp 1700315010
transform 1 0 83850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__910_
timestamp 1700315010
transform 1 0 82950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__911_
timestamp 1700315010
transform 1 0 81150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__912_
timestamp 1700315010
transform 1 0 86250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__913_
timestamp 1700315010
transform -1 0 83550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__914_
timestamp 1700315010
transform -1 0 78750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__915_
timestamp 1700315010
transform 1 0 78450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__916_
timestamp 1700315010
transform -1 0 84450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__917_
timestamp 1700315010
transform 1 0 87450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__918_
timestamp 1700315010
transform -1 0 80850 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__919_
timestamp 1700315010
transform 1 0 80850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__920_
timestamp 1700315010
transform -1 0 83550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__921_
timestamp 1700315010
transform 1 0 84750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__922_
timestamp 1700315010
transform 1 0 80550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__923_
timestamp 1700315010
transform 1 0 88650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__924_
timestamp 1700315010
transform 1 0 88350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__925_
timestamp 1700315010
transform -1 0 89550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__926_
timestamp 1700315010
transform -1 0 64950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__927_
timestamp 1700315010
transform 1 0 72750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__928_
timestamp 1700315010
transform 1 0 70350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__929_
timestamp 1700315010
transform 1 0 63150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__930_
timestamp 1700315010
transform 1 0 55050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__931_
timestamp 1700315010
transform -1 0 57450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__932_
timestamp 1700315010
transform 1 0 61950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__933_
timestamp 1700315010
transform -1 0 66150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__934_
timestamp 1700315010
transform 1 0 67950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__935_
timestamp 1700315010
transform -1 0 80850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__936_
timestamp 1700315010
transform 1 0 61050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__937_
timestamp 1700315010
transform -1 0 59850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__938_
timestamp 1700315010
transform -1 0 59850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__939_
timestamp 1700315010
transform 1 0 54750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__940_
timestamp 1700315010
transform 1 0 51750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__941_
timestamp 1700315010
transform -1 0 48750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__942_
timestamp 1700315010
transform 1 0 54450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__943_
timestamp 1700315010
transform 1 0 52050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__944_
timestamp 1700315010
transform -1 0 79650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__945_
timestamp 1700315010
transform 1 0 83550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__946_
timestamp 1700315010
transform 1 0 81150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__947_
timestamp 1700315010
transform 1 0 84750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__948_
timestamp 1700315010
transform 1 0 78750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__949_
timestamp 1700315010
transform 1 0 76350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__950_
timestamp 1700315010
transform -1 0 69750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__951_
timestamp 1700315010
transform 1 0 58650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__952_
timestamp 1700315010
transform 1 0 34950 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__953_
timestamp 1700315010
transform 1 0 39450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__954_
timestamp 1700315010
transform -1 0 37350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__955_
timestamp 1700315010
transform 1 0 41250 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__956_
timestamp 1700315010
transform 1 0 47550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__957_
timestamp 1700315010
transform 1 0 52350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__958_
timestamp 1700315010
transform 1 0 54150 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__959_
timestamp 1700315010
transform 1 0 54150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__960_
timestamp 1700315010
transform 1 0 47550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__961_
timestamp 1700315010
transform -1 0 52050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__962_
timestamp 1700315010
transform 1 0 56550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__963_
timestamp 1700315010
transform 1 0 43650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__964_
timestamp 1700315010
transform -1 0 39750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__965_
timestamp 1700315010
transform 1 0 37350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__966_
timestamp 1700315010
transform 1 0 49950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__967_
timestamp 1700315010
transform -1 0 43950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__968_
timestamp 1700315010
transform 1 0 38550 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__969_
timestamp 1700315010
transform -1 0 41550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__970_
timestamp 1700315010
transform 1 0 45450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__971_
timestamp 1700315010
transform 1 0 45450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__972_
timestamp 1700315010
transform -1 0 47850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__973_
timestamp 1700315010
transform 1 0 45450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__974_
timestamp 1700315010
transform -1 0 52350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__975_
timestamp 1700315010
transform 1 0 45750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__976_
timestamp 1700315010
transform 1 0 39150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__977_
timestamp 1700315010
transform 1 0 31650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__978_
timestamp 1700315010
transform 1 0 37350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__979_
timestamp 1700315010
transform 1 0 31350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__980_
timestamp 1700315010
transform 1 0 43350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__981_
timestamp 1700315010
transform 1 0 54450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__982_
timestamp 1700315010
transform -1 0 52050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__983_
timestamp 1700315010
transform -1 0 41250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__984_
timestamp 1700315010
transform -1 0 36450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__985_
timestamp 1700315010
transform -1 0 35250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__986_
timestamp 1700315010
transform -1 0 25950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__987_
timestamp 1700315010
transform -1 0 23850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__988_
timestamp 1700315010
transform -1 0 20550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__989_
timestamp 1700315010
transform -1 0 27150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__990_
timestamp 1700315010
transform 1 0 27750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__991_
timestamp 1700315010
transform 1 0 35850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__992_
timestamp 1700315010
transform -1 0 35850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__993_
timestamp 1700315010
transform 1 0 30150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__994_
timestamp 1700315010
transform 1 0 38850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__995_
timestamp 1700315010
transform -1 0 41850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__996_
timestamp 1700315010
transform 1 0 25350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__997_
timestamp 1700315010
transform -1 0 21450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__998_
timestamp 1700315010
transform 1 0 24150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__999_
timestamp 1700315010
transform 1 0 32850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1000_
timestamp 1700315010
transform 1 0 33450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1001_
timestamp 1700315010
transform 1 0 41550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1002_
timestamp 1700315010
transform 1 0 34950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1003_
timestamp 1700315010
transform -1 0 44250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1004_
timestamp 1700315010
transform 1 0 37050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1005_
timestamp 1700315010
transform -1 0 34950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1006_
timestamp 1700315010
transform 1 0 30450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1007_
timestamp 1700315010
transform -1 0 25050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1008_
timestamp 1700315010
transform 1 0 26550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1009_
timestamp 1700315010
transform -1 0 29250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1010_
timestamp 1700315010
transform 1 0 34650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1011_
timestamp 1700315010
transform -1 0 33150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1012_
timestamp 1700315010
transform -1 0 22050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1013_
timestamp 1700315010
transform -1 0 37050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1014_
timestamp 1700315010
transform -1 0 32850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1015_
timestamp 1700315010
transform -1 0 30750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1016_
timestamp 1700315010
transform -1 0 31050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1017_
timestamp 1700315010
transform 1 0 32850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1018_
timestamp 1700315010
transform -1 0 35550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1019_
timestamp 1700315010
transform -1 0 26550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1020_
timestamp 1700315010
transform -1 0 22650 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1021_
timestamp 1700315010
transform -1 0 21450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1022_
timestamp 1700315010
transform -1 0 20850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1023_
timestamp 1700315010
transform 1 0 16950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1024_
timestamp 1700315010
transform 1 0 22350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1025_
timestamp 1700315010
transform 1 0 21750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1026_
timestamp 1700315010
transform 1 0 18750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1027_
timestamp 1700315010
transform 1 0 22350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1028_
timestamp 1700315010
transform 1 0 15750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1029_
timestamp 1700315010
transform -1 0 13650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1030_
timestamp 1700315010
transform -1 0 23850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1031_
timestamp 1700315010
transform 1 0 19350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1032_
timestamp 1700315010
transform -1 0 18450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1033_
timestamp 1700315010
transform -1 0 16050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1034_
timestamp 1700315010
transform -1 0 24750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1035_
timestamp 1700315010
transform -1 0 16350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1036_
timestamp 1700315010
transform -1 0 17550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1037_
timestamp 1700315010
transform -1 0 15750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1038_
timestamp 1700315010
transform 1 0 24450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1039_
timestamp 1700315010
transform -1 0 19950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1040_
timestamp 1700315010
transform -1 0 30750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1041_
timestamp 1700315010
transform -1 0 39750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1042_
timestamp 1700315010
transform 1 0 28350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1043_
timestamp 1700315010
transform 1 0 34350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1044_
timestamp 1700315010
transform 1 0 33750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1045_
timestamp 1700315010
transform 1 0 31350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1046_
timestamp 1700315010
transform -1 0 24150 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1047_
timestamp 1700315010
transform 1 0 26250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1048_
timestamp 1700315010
transform -1 0 29250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1049_
timestamp 1700315010
transform -1 0 21750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1050_
timestamp 1700315010
transform 1 0 22350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1051_
timestamp 1700315010
transform -1 0 10350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1052_
timestamp 1700315010
transform 1 0 17850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1053_
timestamp 1700315010
transform 1 0 18150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1054_
timestamp 1700315010
transform -1 0 20550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1055_
timestamp 1700315010
transform -1 0 14250 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1056_
timestamp 1700315010
transform 1 0 14850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1057_
timestamp 1700315010
transform -1 0 28650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1058_
timestamp 1700315010
transform 1 0 18750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1059_
timestamp 1700315010
transform 1 0 16350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1060_
timestamp 1700315010
transform -1 0 17550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1061_
timestamp 1700315010
transform -1 0 43950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1062_
timestamp 1700315010
transform -1 0 28650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1063_
timestamp 1700315010
transform 1 0 32550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1064_
timestamp 1700315010
transform 1 0 20550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1065_
timestamp 1700315010
transform -1 0 13950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1066_
timestamp 1700315010
transform 1 0 15450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1067_
timestamp 1700315010
transform 1 0 19350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1068_
timestamp 1700315010
transform -1 0 12750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1069_
timestamp 1700315010
transform 1 0 18450 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1070_
timestamp 1700315010
transform 1 0 29250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1071_
timestamp 1700315010
transform 1 0 23550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1072_
timestamp 1700315010
transform -1 0 3150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1073_
timestamp 1700315010
transform -1 0 14250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1074_
timestamp 1700315010
transform -1 0 11850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1075_
timestamp 1700315010
transform -1 0 11850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1076_
timestamp 1700315010
transform -1 0 14550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1077_
timestamp 1700315010
transform 1 0 16650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1078_
timestamp 1700315010
transform -1 0 7350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1079_
timestamp 1700315010
transform -1 0 13350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1080_
timestamp 1700315010
transform -1 0 12750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1081_
timestamp 1700315010
transform -1 0 3150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1082_
timestamp 1700315010
transform -1 0 15450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1083_
timestamp 1700315010
transform -1 0 11250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1084_
timestamp 1700315010
transform -1 0 5550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1085_
timestamp 1700315010
transform -1 0 5250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1086_
timestamp 1700315010
transform 1 0 10050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1087_
timestamp 1700315010
transform 1 0 7650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1088_
timestamp 1700315010
transform -1 0 9450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1089_
timestamp 1700315010
transform 1 0 29250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1090_
timestamp 1700315010
transform 1 0 23250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1091_
timestamp 1700315010
transform -1 0 28350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1092_
timestamp 1700315010
transform -1 0 30450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1093_
timestamp 1700315010
transform 1 0 28050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1094_
timestamp 1700315010
transform 1 0 32550 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1095_
timestamp 1700315010
transform -1 0 27750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1096_
timestamp 1700315010
transform -1 0 25350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1097_
timestamp 1700315010
transform -1 0 23850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1098_
timestamp 1700315010
transform -1 0 25950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1099_
timestamp 1700315010
transform -1 0 21450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1100_
timestamp 1700315010
transform -1 0 750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1101_
timestamp 1700315010
transform -1 0 750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1102_
timestamp 1700315010
transform -1 0 13950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1103_
timestamp 1700315010
transform 1 0 9150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1104_
timestamp 1700315010
transform 1 0 7050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1105_
timestamp 1700315010
transform 1 0 2550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1106_
timestamp 1700315010
transform -1 0 750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1107_
timestamp 1700315010
transform 1 0 2850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1108_
timestamp 1700315010
transform 1 0 13050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1109_
timestamp 1700315010
transform -1 0 5250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1110_
timestamp 1700315010
transform -1 0 3150 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1111_
timestamp 1700315010
transform -1 0 750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1112_
timestamp 1700315010
transform -1 0 30450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1113_
timestamp 1700315010
transform 1 0 7050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1114_
timestamp 1700315010
transform -1 0 26550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1115_
timestamp 1700315010
transform -1 0 7650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1116_
timestamp 1700315010
transform -1 0 9450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1117_
timestamp 1700315010
transform 1 0 11250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1118_
timestamp 1700315010
transform -1 0 5250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1119_
timestamp 1700315010
transform 1 0 7350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1120_
timestamp 1700315010
transform 1 0 7050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1121_
timestamp 1700315010
transform 1 0 13350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1122_
timestamp 1700315010
transform -1 0 11250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1123_
timestamp 1700315010
transform -1 0 9750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1124_
timestamp 1700315010
transform 1 0 7650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1125_
timestamp 1700315010
transform 1 0 2850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1126_
timestamp 1700315010
transform -1 0 750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1127_
timestamp 1700315010
transform 1 0 8550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1128_
timestamp 1700315010
transform -1 0 4950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1129_
timestamp 1700315010
transform -1 0 3150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1130_
timestamp 1700315010
transform 1 0 5250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1131_
timestamp 1700315010
transform -1 0 5250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1132_
timestamp 1700315010
transform -1 0 12150 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1133_
timestamp 1700315010
transform -1 0 750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1134_
timestamp 1700315010
transform -1 0 3150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1135_
timestamp 1700315010
transform 1 0 2850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1136_
timestamp 1700315010
transform -1 0 4650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1137_
timestamp 1700315010
transform -1 0 750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1138_
timestamp 1700315010
transform 1 0 7350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1139_
timestamp 1700315010
transform 1 0 8850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1140_
timestamp 1700315010
transform 1 0 26850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1141_
timestamp 1700315010
transform 1 0 34050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1142_
timestamp 1700315010
transform 1 0 37650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1143_
timestamp 1700315010
transform 1 0 49650 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1144_
timestamp 1700315010
transform 1 0 54750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1145_
timestamp 1700315010
transform 1 0 45150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1146_
timestamp 1700315010
transform -1 0 50250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1147_
timestamp 1700315010
transform -1 0 43650 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1148_
timestamp 1700315010
transform 1 0 47550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1149_
timestamp 1700315010
transform -1 0 47850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1150_
timestamp 1700315010
transform 1 0 42150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1151_
timestamp 1700315010
transform 1 0 49950 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1152_
timestamp 1700315010
transform -1 0 47550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1153_
timestamp 1700315010
transform 1 0 35250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1154_
timestamp 1700315010
transform 1 0 37650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1155_
timestamp 1700315010
transform 1 0 39750 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1156_
timestamp 1700315010
transform -1 0 39750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1157_
timestamp 1700315010
transform -1 0 16650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1158_
timestamp 1700315010
transform 1 0 17550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1159_
timestamp 1700315010
transform -1 0 25950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1160_
timestamp 1700315010
transform 1 0 6750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1161_
timestamp 1700315010
transform 1 0 11250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1162_
timestamp 1700315010
transform 1 0 19950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1163_
timestamp 1700315010
transform 1 0 49650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1164_
timestamp 1700315010
transform 1 0 56250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1165_
timestamp 1700315010
transform -1 0 58650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1166_
timestamp 1700315010
transform 1 0 62250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1167_
timestamp 1700315010
transform 1 0 64350 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1168_
timestamp 1700315010
transform -1 0 52050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1169_
timestamp 1700315010
transform 1 0 60150 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1170_
timestamp 1700315010
transform 1 0 52350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1171_
timestamp 1700315010
transform 1 0 60750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1172_
timestamp 1700315010
transform 1 0 58650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1173_
timestamp 1700315010
transform 1 0 60750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1174_
timestamp 1700315010
transform 1 0 53850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1175_
timestamp 1700315010
transform -1 0 56550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1176_
timestamp 1700315010
transform 1 0 54750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1177_
timestamp 1700315010
transform -1 0 44850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1178_
timestamp 1700315010
transform -1 0 44550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1179_
timestamp 1700315010
transform 1 0 50250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1180_
timestamp 1700315010
transform 1 0 31650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1181_
timestamp 1700315010
transform 1 0 49350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1182_
timestamp 1700315010
transform -1 0 59550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1183_
timestamp 1700315010
transform 1 0 56850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1184_
timestamp 1700315010
transform -1 0 54750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1185_
timestamp 1700315010
transform -1 0 56550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1186_
timestamp 1700315010
transform 1 0 60450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1187_
timestamp 1700315010
transform -1 0 49950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1188_
timestamp 1700315010
transform -1 0 66750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1189_
timestamp 1700315010
transform 1 0 56250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1190_
timestamp 1700315010
transform 1 0 58050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1191_
timestamp 1700315010
transform -1 0 63150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1192_
timestamp 1700315010
transform 1 0 67050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1193_
timestamp 1700315010
transform 1 0 65250 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1194_
timestamp 1700315010
transform 1 0 63150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1195_
timestamp 1700315010
transform 1 0 67050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1196_
timestamp 1700315010
transform 1 0 58650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1197_
timestamp 1700315010
transform -1 0 61350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1198_
timestamp 1700315010
transform 1 0 46650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1199_
timestamp 1700315010
transform 1 0 41850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1200_
timestamp 1700315010
transform 1 0 52350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1201_
timestamp 1700315010
transform -1 0 56550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1202_
timestamp 1700315010
transform 1 0 60750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1203_
timestamp 1700315010
transform 1 0 52950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1204_
timestamp 1700315010
transform -1 0 55650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1205_
timestamp 1700315010
transform 1 0 40050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1206_
timestamp 1700315010
transform -1 0 750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1207_
timestamp 1700315010
transform 1 0 11550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1208_
timestamp 1700315010
transform -1 0 750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1209_
timestamp 1700315010
transform 1 0 35550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1210_
timestamp 1700315010
transform -1 0 23250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1211_
timestamp 1700315010
transform -1 0 32550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1212_
timestamp 1700315010
transform 1 0 27450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1213_
timestamp 1700315010
transform 1 0 31350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1214_
timestamp 1700315010
transform 1 0 33150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1215_
timestamp 1700315010
transform -1 0 20850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1216_
timestamp 1700315010
transform -1 0 29550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1217_
timestamp 1700315010
transform 1 0 29850 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1218_
timestamp 1700315010
transform -1 0 27150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1219_
timestamp 1700315010
transform 1 0 18450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1220_
timestamp 1700315010
transform -1 0 3150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1221_
timestamp 1700315010
transform -1 0 22950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1222_
timestamp 1700315010
transform -1 0 28650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1223_
timestamp 1700315010
transform 1 0 26850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1224_
timestamp 1700315010
transform -1 0 31650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1225_
timestamp 1700315010
transform 1 0 28950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1226_
timestamp 1700315010
transform -1 0 25050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1227_
timestamp 1700315010
transform 1 0 23550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1228_
timestamp 1700315010
transform 1 0 29550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1229_
timestamp 1700315010
transform 1 0 33450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1230_
timestamp 1700315010
transform 1 0 27750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1231_
timestamp 1700315010
transform -1 0 25650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1232_
timestamp 1700315010
transform 1 0 11550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1233_
timestamp 1700315010
transform 1 0 4650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1234_
timestamp 1700315010
transform 1 0 16650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1235_
timestamp 1700315010
transform 1 0 13950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1236_
timestamp 1700315010
transform -1 0 4350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1237_
timestamp 1700315010
transform 1 0 8550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1238_
timestamp 1700315010
transform 1 0 11250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1239_
timestamp 1700315010
transform -1 0 7650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1240_
timestamp 1700315010
transform -1 0 6450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1241_
timestamp 1700315010
transform -1 0 3450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1242_
timestamp 1700315010
transform 1 0 9450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1243_
timestamp 1700315010
transform 1 0 5250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1244_
timestamp 1700315010
transform 1 0 2850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1245_
timestamp 1700315010
transform -1 0 3150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1246_
timestamp 1700315010
transform -1 0 750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1247_
timestamp 1700315010
transform -1 0 750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1248_
timestamp 1700315010
transform 1 0 8550 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1249_
timestamp 1700315010
transform 1 0 450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1250_
timestamp 1700315010
transform -1 0 3150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1251_
timestamp 1700315010
transform -1 0 16650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1252_
timestamp 1700315010
transform 1 0 7050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1253_
timestamp 1700315010
transform 1 0 450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1254_
timestamp 1700315010
transform -1 0 9750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1255_
timestamp 1700315010
transform -1 0 750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1256_
timestamp 1700315010
transform 1 0 4950 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1257_
timestamp 1700315010
transform -1 0 14250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1258_
timestamp 1700315010
transform 1 0 5250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1259_
timestamp 1700315010
transform -1 0 12450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1260_
timestamp 1700315010
transform -1 0 12450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1261_
timestamp 1700315010
transform 1 0 14250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1262_
timestamp 1700315010
transform 1 0 2850 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1263_
timestamp 1700315010
transform -1 0 10350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1264_
timestamp 1700315010
transform 1 0 7350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1265_
timestamp 1700315010
transform -1 0 10050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1266_
timestamp 1700315010
transform -1 0 9750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1267_
timestamp 1700315010
transform -1 0 5550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1268_
timestamp 1700315010
transform 1 0 16050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1269_
timestamp 1700315010
transform 1 0 18450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1270_
timestamp 1700315010
transform 1 0 35250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1271_
timestamp 1700315010
transform -1 0 46350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1272_
timestamp 1700315010
transform 1 0 74850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1273_
timestamp 1700315010
transform -1 0 71250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1274_
timestamp 1700315010
transform 1 0 62250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1275_
timestamp 1700315010
transform 1 0 59250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1276_
timestamp 1700315010
transform -1 0 67050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1277_
timestamp 1700315010
transform 1 0 61650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1278_
timestamp 1700315010
transform 1 0 71250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1279_
timestamp 1700315010
transform 1 0 70650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1280_
timestamp 1700315010
transform -1 0 53250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1281_
timestamp 1700315010
transform -1 0 57750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1282_
timestamp 1700315010
transform -1 0 61050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1283_
timestamp 1700315010
transform -1 0 55350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1284_
timestamp 1700315010
transform -1 0 24750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1285_
timestamp 1700315010
transform -1 0 49050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1286_
timestamp 1700315010
transform -1 0 22650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1287_
timestamp 1700315010
transform 1 0 28350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1288_
timestamp 1700315010
transform 1 0 44850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1289_
timestamp 1700315010
transform 1 0 42450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1290_
timestamp 1700315010
transform -1 0 47250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1291_
timestamp 1700315010
transform -1 0 35850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1292_
timestamp 1700315010
transform -1 0 33750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1293_
timestamp 1700315010
transform -1 0 39450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1294_
timestamp 1700315010
transform 1 0 18750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1295_
timestamp 1700315010
transform 1 0 16650 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1296_
timestamp 1700315010
transform -1 0 24750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1297_
timestamp 1700315010
transform 1 0 24150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1298_
timestamp 1700315010
transform 1 0 4950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1299_
timestamp 1700315010
transform 1 0 11550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1300_
timestamp 1700315010
transform -1 0 24150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1301_
timestamp 1700315010
transform 1 0 30750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1302_
timestamp 1700315010
transform -1 0 28650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1303_
timestamp 1700315010
transform -1 0 31050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1304_
timestamp 1700315010
transform -1 0 26250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1305_
timestamp 1700315010
transform -1 0 21150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1306_
timestamp 1700315010
transform 1 0 11550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1307_
timestamp 1700315010
transform 1 0 5250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1308_
timestamp 1700315010
transform -1 0 750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1309_
timestamp 1700315010
transform 1 0 19650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1310_
timestamp 1700315010
transform 1 0 24150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1311_
timestamp 1700315010
transform 1 0 16350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1312_
timestamp 1700315010
transform -1 0 26250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1313_
timestamp 1700315010
transform -1 0 20250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1314_
timestamp 1700315010
transform -1 0 18450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1315_
timestamp 1700315010
transform 1 0 19350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1316_
timestamp 1700315010
transform -1 0 11550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1317_
timestamp 1700315010
transform 1 0 14250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1318_
timestamp 1700315010
transform 1 0 41550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1319_
timestamp 1700315010
transform -1 0 30750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1320_
timestamp 1700315010
transform -1 0 26550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1321_
timestamp 1700315010
transform -1 0 24150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1322_
timestamp 1700315010
transform -1 0 17250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1323_
timestamp 1700315010
transform -1 0 22050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1324_
timestamp 1700315010
transform -1 0 12150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1325_
timestamp 1700315010
transform -1 0 15150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1326_
timestamp 1700315010
transform -1 0 10050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1327_
timestamp 1700315010
transform -1 0 750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1328_
timestamp 1700315010
transform -1 0 750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1329_
timestamp 1700315010
transform 1 0 9450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1330_
timestamp 1700315010
transform -1 0 7350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1331_
timestamp 1700315010
transform 1 0 2550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1332_
timestamp 1700315010
transform 1 0 7050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1333_
timestamp 1700315010
transform 1 0 11850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1334_
timestamp 1700315010
transform 1 0 7350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1335_
timestamp 1700315010
transform -1 0 750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1336_
timestamp 1700315010
transform 1 0 7050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1337_
timestamp 1700315010
transform 1 0 16650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1338_
timestamp 1700315010
transform 1 0 450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1339_
timestamp 1700315010
transform 1 0 10650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1340_
timestamp 1700315010
transform 1 0 9450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1341_
timestamp 1700315010
transform 1 0 2250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1342_
timestamp 1700315010
transform -1 0 2850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1343_
timestamp 1700315010
transform 1 0 4650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1344_
timestamp 1700315010
transform -1 0 13050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1345_
timestamp 1700315010
transform -1 0 22350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1346_
timestamp 1700315010
transform 1 0 13350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1347_
timestamp 1700315010
transform 1 0 15150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1348_
timestamp 1700315010
transform -1 0 20250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1349_
timestamp 1700315010
transform -1 0 20850 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1350_
timestamp 1700315010
transform 1 0 7650 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1351_
timestamp 1700315010
transform 1 0 14550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1352_
timestamp 1700315010
transform 1 0 25950 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1353_
timestamp 1700315010
transform -1 0 17850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1354_
timestamp 1700315010
transform 1 0 25350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1355_
timestamp 1700315010
transform -1 0 32250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1356_
timestamp 1700315010
transform 1 0 49050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1357_
timestamp 1700315010
transform 1 0 51450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1358_
timestamp 1700315010
transform 1 0 53550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1359_
timestamp 1700315010
transform 1 0 68250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_1__1360_
timestamp 1700315010
transform 1 0 67350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1361_
timestamp 1700315010
transform -1 0 63150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1362_
timestamp 1700315010
transform 1 0 64950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1363_
timestamp 1700315010
transform -1 0 60750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1364_
timestamp 1700315010
transform 1 0 58350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1365_
timestamp 1700315010
transform -1 0 72150 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1366_
timestamp 1700315010
transform -1 0 23250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1367_
timestamp 1700315010
transform 1 0 20850 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1368_
timestamp 1700315010
transform 1 0 31350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1369_
timestamp 1700315010
transform 1 0 43650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1370_
timestamp 1700315010
transform 1 0 34050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1371_
timestamp 1700315010
transform 1 0 37350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1372_
timestamp 1700315010
transform -1 0 19050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1373_
timestamp 1700315010
transform 1 0 14550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1374_
timestamp 1700315010
transform -1 0 7650 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1375_
timestamp 1700315010
transform -1 0 4950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1376_
timestamp 1700315010
transform -1 0 19350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1377_
timestamp 1700315010
transform -1 0 13050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1378_
timestamp 1700315010
transform -1 0 17550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1379_
timestamp 1700315010
transform -1 0 15450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1380_
timestamp 1700315010
transform -1 0 17250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1381_
timestamp 1700315010
transform -1 0 14850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1382_
timestamp 1700315010
transform -1 0 10950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1383_
timestamp 1700315010
transform -1 0 14850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1384_
timestamp 1700315010
transform -1 0 17250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1385_
timestamp 1700315010
transform -1 0 12450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1386_
timestamp 1700315010
transform -1 0 3450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1387_
timestamp 1700315010
transform 1 0 9150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1388_
timestamp 1700315010
transform 1 0 23550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1389_
timestamp 1700315010
transform -1 0 27150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1390_
timestamp 1700315010
transform -1 0 25050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1391_
timestamp 1700315010
transform -1 0 22350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1392_
timestamp 1700315010
transform 1 0 30450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1393_
timestamp 1700315010
transform 1 0 28050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1394_
timestamp 1700315010
transform 1 0 20550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1395_
timestamp 1700315010
transform 1 0 6150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1396_
timestamp 1700315010
transform -1 0 8550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1397_
timestamp 1700315010
transform -1 0 750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1398_
timestamp 1700315010
transform -1 0 4950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1399_
timestamp 1700315010
transform -1 0 10050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1400_
timestamp 1700315010
transform -1 0 4350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1401_
timestamp 1700315010
transform -1 0 750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1402_
timestamp 1700315010
transform -1 0 2250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1403_
timestamp 1700315010
transform 1 0 4950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1404_
timestamp 1700315010
transform -1 0 7350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1405_
timestamp 1700315010
transform 1 0 4950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1406_
timestamp 1700315010
transform -1 0 750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1407_
timestamp 1700315010
transform -1 0 750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1408_
timestamp 1700315010
transform -1 0 5550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1409_
timestamp 1700315010
transform -1 0 3150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1410_
timestamp 1700315010
transform 1 0 2850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1411_
timestamp 1700315010
transform -1 0 5550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1412_
timestamp 1700315010
transform 1 0 9150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1413_
timestamp 1700315010
transform -1 0 750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1414_
timestamp 1700315010
transform -1 0 9450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1415_
timestamp 1700315010
transform -1 0 19350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1416_
timestamp 1700315010
transform 1 0 28350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1417_
timestamp 1700315010
transform 1 0 15750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1418_
timestamp 1700315010
transform -1 0 18150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1419_
timestamp 1700315010
transform 1 0 20250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1420_
timestamp 1700315010
transform -1 0 37050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1421_
timestamp 1700315010
transform -1 0 36750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1422_
timestamp 1700315010
transform 1 0 41550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1423_
timestamp 1700315010
transform -1 0 39150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1424_
timestamp 1700315010
transform 1 0 42750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1425_
timestamp 1700315010
transform -1 0 44850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1426_
timestamp 1700315010
transform 1 0 46650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1427_
timestamp 1700315010
transform 1 0 68850 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1428_
timestamp 1700315010
transform -1 0 64350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1429_
timestamp 1700315010
transform 1 0 64950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1430_
timestamp 1700315010
transform 1 0 67350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1431_
timestamp 1700315010
transform -1 0 70650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1432_
timestamp 1700315010
transform 1 0 70950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1433_
timestamp 1700315010
transform -1 0 65250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1434_
timestamp 1700315010
transform 1 0 69450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_1__1435_
timestamp 1700315010
transform 1 0 88950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1436_
timestamp 1700315010
transform -1 0 86550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1437_
timestamp 1700315010
transform -1 0 58050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1438_
timestamp 1700315010
transform 1 0 39750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1439_
timestamp 1700315010
transform 1 0 19050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1440_
timestamp 1700315010
transform -1 0 17850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1441_
timestamp 1700315010
transform 1 0 7350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1442_
timestamp 1700315010
transform 1 0 27150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1443_
timestamp 1700315010
transform -1 0 31050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1444_
timestamp 1700315010
transform -1 0 21150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1445_
timestamp 1700315010
transform -1 0 25950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1446_
timestamp 1700315010
transform 1 0 22950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1447_
timestamp 1700315010
transform 1 0 25050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1448_
timestamp 1700315010
transform 1 0 26850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1449_
timestamp 1700315010
transform -1 0 28650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1450_
timestamp 1700315010
transform -1 0 23250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1451_
timestamp 1700315010
transform 1 0 24750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1452_
timestamp 1700315010
transform 1 0 28350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1453_
timestamp 1700315010
transform 1 0 31050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1454_
timestamp 1700315010
transform 1 0 28650 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1455_
timestamp 1700315010
transform 1 0 43050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1456_
timestamp 1700315010
transform -1 0 32250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1457_
timestamp 1700315010
transform -1 0 29250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1458_
timestamp 1700315010
transform -1 0 24150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1459_
timestamp 1700315010
transform -1 0 7050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1460_
timestamp 1700315010
transform 1 0 25950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1461_
timestamp 1700315010
transform 1 0 10950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1462_
timestamp 1700315010
transform -1 0 2550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1463_
timestamp 1700315010
transform -1 0 21450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1464_
timestamp 1700315010
transform -1 0 13350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1465_
timestamp 1700315010
transform -1 0 15450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1466_
timestamp 1700315010
transform -1 0 8850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1467_
timestamp 1700315010
transform -1 0 19650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1468_
timestamp 1700315010
transform 1 0 21450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1469_
timestamp 1700315010
transform -1 0 16650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1470_
timestamp 1700315010
transform -1 0 13350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1471_
timestamp 1700315010
transform 1 0 11550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1472_
timestamp 1700315010
transform 1 0 13950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1473_
timestamp 1700315010
transform 1 0 18450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1474_
timestamp 1700315010
transform 1 0 41550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1475_
timestamp 1700315010
transform 1 0 40950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1476_
timestamp 1700315010
transform 1 0 44550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1477_
timestamp 1700315010
transform 1 0 46950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1478_
timestamp 1700315010
transform 1 0 48450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1479_
timestamp 1700315010
transform 1 0 52650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1480_
timestamp 1700315010
transform -1 0 63450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1481_
timestamp 1700315010
transform -1 0 65250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1482_
timestamp 1700315010
transform 1 0 69450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1483_
timestamp 1700315010
transform 1 0 80550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1484_
timestamp 1700315010
transform -1 0 82650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1485_
timestamp 1700315010
transform 1 0 82350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1486_
timestamp 1700315010
transform -1 0 85050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1487_
timestamp 1700315010
transform 1 0 87150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1488_
timestamp 1700315010
transform 1 0 32550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1489_
timestamp 1700315010
transform 1 0 34950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1490_
timestamp 1700315010
transform -1 0 35250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1491_
timestamp 1700315010
transform -1 0 43050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1492_
timestamp 1700315010
transform -1 0 31650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1493_
timestamp 1700315010
transform -1 0 33750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1494_
timestamp 1700315010
transform 1 0 38250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1495_
timestamp 1700315010
transform 1 0 44550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1496_
timestamp 1700315010
transform 1 0 35850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1497_
timestamp 1700315010
transform 1 0 38850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1498_
timestamp 1700315010
transform 1 0 40950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1499_
timestamp 1700315010
transform 1 0 33150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1500_
timestamp 1700315010
transform 1 0 36450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1501_
timestamp 1700315010
transform 1 0 40650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1502_
timestamp 1700315010
transform 1 0 40950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1503_
timestamp 1700315010
transform 1 0 41550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1504_
timestamp 1700315010
transform 1 0 42750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1505_
timestamp 1700315010
transform -1 0 36750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1506_
timestamp 1700315010
transform -1 0 39450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1507_
timestamp 1700315010
transform -1 0 37050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1508_
timestamp 1700315010
transform -1 0 33150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1509_
timestamp 1700315010
transform 1 0 30450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1510_
timestamp 1700315010
transform -1 0 28650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1511_
timestamp 1700315010
transform 1 0 34650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1512_
timestamp 1700315010
transform -1 0 40650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1513_
timestamp 1700315010
transform 1 0 49650 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1514_
timestamp 1700315010
transform -1 0 45750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1515_
timestamp 1700315010
transform 1 0 47250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1516_
timestamp 1700315010
transform -1 0 37950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1517_
timestamp 1700315010
transform 1 0 43050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1518_
timestamp 1700315010
transform -1 0 48150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1519_
timestamp 1700315010
transform 1 0 43650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1520_
timestamp 1700315010
transform 1 0 45750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1521_
timestamp 1700315010
transform 1 0 38250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1522_
timestamp 1700315010
transform 1 0 40650 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1523_
timestamp 1700315010
transform 1 0 42450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1524_
timestamp 1700315010
transform 1 0 49350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1525_
timestamp 1700315010
transform -1 0 82050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1526_
timestamp 1700315010
transform -1 0 74550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1527_
timestamp 1700315010
transform 1 0 67050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1528_
timestamp 1700315010
transform 1 0 64650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1529_
timestamp 1700315010
transform 1 0 68550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1530_
timestamp 1700315010
transform -1 0 72750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1531_
timestamp 1700315010
transform -1 0 76050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1532_
timestamp 1700315010
transform 1 0 78150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1533_
timestamp 1700315010
transform -1 0 80250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1534_
timestamp 1700315010
transform -1 0 77250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1535_
timestamp 1700315010
transform -1 0 56250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1536_
timestamp 1700315010
transform 1 0 47550 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1537_
timestamp 1700315010
transform 1 0 41850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1538_
timestamp 1700315010
transform 1 0 38550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1539_
timestamp 1700315010
transform 1 0 34350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1540_
timestamp 1700315010
transform -1 0 39450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1541_
timestamp 1700315010
transform -1 0 41850 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1542_
timestamp 1700315010
transform -1 0 37050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1543_
timestamp 1700315010
transform 1 0 39450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1544_
timestamp 1700315010
transform 1 0 36450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1545_
timestamp 1700315010
transform -1 0 37050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1546_
timestamp 1700315010
transform -1 0 37350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1547_
timestamp 1700315010
transform -1 0 40050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1548_
timestamp 1700315010
transform -1 0 45450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1549_
timestamp 1700315010
transform -1 0 42150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1550_
timestamp 1700315010
transform 1 0 51750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1551_
timestamp 1700315010
transform 1 0 58350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1552_
timestamp 1700315010
transform 1 0 62550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1553_
timestamp 1700315010
transform -1 0 75750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1554_
timestamp 1700315010
transform 1 0 78150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1555_
timestamp 1700315010
transform 1 0 77850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1556_
timestamp 1700315010
transform -1 0 74550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1557_
timestamp 1700315010
transform -1 0 72750 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1558_
timestamp 1700315010
transform 1 0 37650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1559_
timestamp 1700315010
transform 1 0 52650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1560_
timestamp 1700315010
transform 1 0 54450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1561_
timestamp 1700315010
transform -1 0 40350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1562_
timestamp 1700315010
transform 1 0 40050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1563_
timestamp 1700315010
transform 1 0 55350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1564_
timestamp 1700315010
transform -1 0 30750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1565_
timestamp 1700315010
transform -1 0 32250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1566_
timestamp 1700315010
transform -1 0 34350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1567_
timestamp 1700315010
transform 1 0 43350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1568_
timestamp 1700315010
transform 1 0 49650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1569_
timestamp 1700315010
transform 1 0 58950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1570_
timestamp 1700315010
transform 1 0 50250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1571_
timestamp 1700315010
transform -1 0 54150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1572_
timestamp 1700315010
transform 1 0 51450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1573_
timestamp 1700315010
transform 1 0 61350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1574_
timestamp 1700315010
transform -1 0 60750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1575_
timestamp 1700315010
transform 1 0 64650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1576_
timestamp 1700315010
transform 1 0 62250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1577_
timestamp 1700315010
transform 1 0 66750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1578_
timestamp 1700315010
transform 1 0 85350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1579_
timestamp 1700315010
transform -1 0 76650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1580_
timestamp 1700315010
transform -1 0 76050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1581_
timestamp 1700315010
transform 1 0 73050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1582_
timestamp 1700315010
transform -1 0 67350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1583_
timestamp 1700315010
transform -1 0 57150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1584_
timestamp 1700315010
transform 1 0 43950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1585_
timestamp 1700315010
transform 1 0 46350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1586_
timestamp 1700315010
transform 1 0 54150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1587_
timestamp 1700315010
transform 1 0 37950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1588_
timestamp 1700315010
transform -1 0 57750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1589_
timestamp 1700315010
transform 1 0 73950 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1590_
timestamp 1700315010
transform 1 0 71550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1__1591_
timestamp 1700315010
transform -1 0 70950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_1__1592_
timestamp 1700315010
transform -1 0 64950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1593_
timestamp 1700315010
transform -1 0 64950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1__1594_
timestamp 1700315010
transform 1 0 64350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1595_
timestamp 1700315010
transform 1 0 59550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1596_
timestamp 1700315010
transform -1 0 61950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1597_
timestamp 1700315010
transform 1 0 59850 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1598_
timestamp 1700315010
transform -1 0 62250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1599_
timestamp 1700315010
transform -1 0 58350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1600_
timestamp 1700315010
transform -1 0 60150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1601_
timestamp 1700315010
transform 1 0 49350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1602_
timestamp 1700315010
transform -1 0 49950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1603_
timestamp 1700315010
transform 1 0 43950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1604_
timestamp 1700315010
transform -1 0 46350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1605_
timestamp 1700315010
transform -1 0 67050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1606_
timestamp 1700315010
transform -1 0 77250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1607_
timestamp 1700315010
transform 1 0 66150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1608_
timestamp 1700315010
transform -1 0 68550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1636_
timestamp 1700315010
transform -1 0 88350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1637_
timestamp 1700315010
transform 1 0 88350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1638_
timestamp 1700315010
transform -1 0 80250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1639_
timestamp 1700315010
transform 1 0 77850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1640_
timestamp 1700315010
transform 1 0 77850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1641_
timestamp 1700315010
transform -1 0 56250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1642_
timestamp 1700315010
transform -1 0 47250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1643_
timestamp 1700315010
transform -1 0 44850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1644_
timestamp 1700315010
transform -1 0 57750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1645_
timestamp 1700315010
transform -1 0 65850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1646_
timestamp 1700315010
transform -1 0 61350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1647_
timestamp 1700315010
transform 1 0 47250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1648_
timestamp 1700315010
transform 1 0 86550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1649_
timestamp 1700315010
transform -1 0 64050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1650_
timestamp 1700315010
transform -1 0 66450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1651_
timestamp 1700315010
transform 1 0 64350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1652_
timestamp 1700315010
transform -1 0 54150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1653_
timestamp 1700315010
transform 1 0 61950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1654_
timestamp 1700315010
transform 1 0 86850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1655_
timestamp 1700315010
transform -1 0 84750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1656_
timestamp 1700315010
transform 1 0 88650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1657_
timestamp 1700315010
transform 1 0 86550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1658_
timestamp 1700315010
transform 1 0 84150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1659_
timestamp 1700315010
transform -1 0 79950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1660_
timestamp 1700315010
transform -1 0 82650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1661_
timestamp 1700315010
transform 1 0 79950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1662_
timestamp 1700315010
transform -1 0 51750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1663_
timestamp 1700315010
transform -1 0 49350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1664_
timestamp 1700315010
transform -1 0 51450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1665_
timestamp 1700315010
transform -1 0 54450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1666_
timestamp 1700315010
transform -1 0 57150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1667_
timestamp 1700315010
transform 1 0 57450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1668_
timestamp 1700315010
transform 1 0 55350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1669_
timestamp 1700315010
transform -1 0 60450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1670_
timestamp 1700315010
transform 1 0 62550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1671_
timestamp 1700315010
transform 1 0 78150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1672_
timestamp 1700315010
transform -1 0 84750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1673_
timestamp 1700315010
transform 1 0 82050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1674_
timestamp 1700315010
transform -1 0 80250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1675_
timestamp 1700315010
transform -1 0 82950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1676_
timestamp 1700315010
transform 1 0 82050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1677_
timestamp 1700315010
transform -1 0 73050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1678_
timestamp 1700315010
transform -1 0 73650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1679_
timestamp 1700315010
transform -1 0 67650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1680_
timestamp 1700315010
transform 1 0 69150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1681_
timestamp 1700315010
transform -1 0 59850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1682_
timestamp 1700315010
transform 1 0 68550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1683_
timestamp 1700315010
transform 1 0 70350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1684_
timestamp 1700315010
transform 1 0 75150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1685_
timestamp 1700315010
transform -1 0 62550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1686_
timestamp 1700315010
transform 1 0 64350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1687_
timestamp 1700315010
transform -1 0 76350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1688_
timestamp 1700315010
transform 1 0 78150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1689_
timestamp 1700315010
transform 1 0 73050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1690_
timestamp 1700315010
transform 1 0 76050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1691_
timestamp 1700315010
transform -1 0 73950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1692_
timestamp 1700315010
transform 1 0 53550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1693_
timestamp 1700315010
transform 1 0 46350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1694_
timestamp 1700315010
transform -1 0 49050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1695_
timestamp 1700315010
transform -1 0 43950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1696_
timestamp 1700315010
transform -1 0 45450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1697_
timestamp 1700315010
transform -1 0 49350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1698_
timestamp 1700315010
transform 1 0 51450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1699_
timestamp 1700315010
transform -1 0 58050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1700_
timestamp 1700315010
transform -1 0 58350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1701_
timestamp 1700315010
transform -1 0 53850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1702_
timestamp 1700315010
transform 1 0 55650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1703_
timestamp 1700315010
transform -1 0 68550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1704_
timestamp 1700315010
transform -1 0 71850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1705_
timestamp 1700315010
transform 1 0 60450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1706_
timestamp 1700315010
transform -1 0 64950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1707_
timestamp 1700315010
transform -1 0 67050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1708_
timestamp 1700315010
transform 1 0 67050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1709_
timestamp 1700315010
transform -1 0 54750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1710_
timestamp 1700315010
transform -1 0 58050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1711_
timestamp 1700315010
transform -1 0 53250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1712_
timestamp 1700315010
transform -1 0 55350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1713_
timestamp 1700315010
transform -1 0 50850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1714_
timestamp 1700315010
transform 1 0 56550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1715_
timestamp 1700315010
transform -1 0 58950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1716_
timestamp 1700315010
transform 1 0 61050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1717_
timestamp 1700315010
transform -1 0 66450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1718_
timestamp 1700315010
transform 1 0 68250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1719_
timestamp 1700315010
transform 1 0 70650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1720_
timestamp 1700315010
transform 1 0 63450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1721_
timestamp 1700315010
transform 1 0 69750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1722_
timestamp 1700315010
transform 1 0 71250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1723_
timestamp 1700315010
transform 1 0 71850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1__1724_
timestamp 1700315010
transform -1 0 71850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1725_
timestamp 1700315010
transform 1 0 66150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1726_
timestamp 1700315010
transform -1 0 64050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1727_
timestamp 1700315010
transform -1 0 65550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1728_
timestamp 1700315010
transform -1 0 45150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1__1729_
timestamp 1700315010
transform 1 0 46050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1730_
timestamp 1700315010
transform -1 0 48450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1731_
timestamp 1700315010
transform -1 0 50550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1732_
timestamp 1700315010
transform 1 0 52950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1733_
timestamp 1700315010
transform 1 0 55050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1734_
timestamp 1700315010
transform 1 0 74250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1735_
timestamp 1700315010
transform 1 0 73650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1736_
timestamp 1700315010
transform -1 0 78450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1737_
timestamp 1700315010
transform 1 0 75750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1738_
timestamp 1700315010
transform 1 0 76350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1739_
timestamp 1700315010
transform 1 0 73650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1740_
timestamp 1700315010
transform -1 0 77250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1741_
timestamp 1700315010
transform 1 0 78150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1742_
timestamp 1700315010
transform 1 0 52650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1743_
timestamp 1700315010
transform -1 0 41550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1744_
timestamp 1700315010
transform -1 0 43950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1745_
timestamp 1700315010
transform -1 0 48450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1746_
timestamp 1700315010
transform 1 0 45750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1747_
timestamp 1700315010
transform 1 0 50250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1748_
timestamp 1700315010
transform -1 0 76350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1749_
timestamp 1700315010
transform 1 0 78150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1750_
timestamp 1700315010
transform 1 0 81450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1751_
timestamp 1700315010
transform 1 0 80550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1752_
timestamp 1700315010
transform -1 0 79050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1753_
timestamp 1700315010
transform 1 0 80550 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1754_
timestamp 1700315010
transform 1 0 77250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_1__1755_
timestamp 1700315010
transform 1 0 80550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1756_
timestamp 1700315010
transform 1 0 72450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1757_
timestamp 1700315010
transform -1 0 65850 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1758_
timestamp 1700315010
transform 1 0 63450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1759_
timestamp 1700315010
transform 1 0 59850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1760_
timestamp 1700315010
transform 1 0 67650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1761_
timestamp 1700315010
transform -1 0 70350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1762_
timestamp 1700315010
transform -1 0 76950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1763_
timestamp 1700315010
transform 1 0 79050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1764_
timestamp 1700315010
transform 1 0 83850 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1765_
timestamp 1700315010
transform 1 0 85950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1766_
timestamp 1700315010
transform 1 0 87450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1767_
timestamp 1700315010
transform 1 0 73350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1768_
timestamp 1700315010
transform -1 0 71250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1769_
timestamp 1700315010
transform -1 0 68850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1770_
timestamp 1700315010
transform -1 0 75150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1771_
timestamp 1700315010
transform 1 0 82650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1772_
timestamp 1700315010
transform 1 0 82950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1773_
timestamp 1700315010
transform -1 0 87150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_1__1774_
timestamp 1700315010
transform -1 0 83850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1775_
timestamp 1700315010
transform -1 0 85650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1776_
timestamp 1700315010
transform 1 0 85650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1777_
timestamp 1700315010
transform 1 0 73950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1778_
timestamp 1700315010
transform 1 0 67050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1779_
timestamp 1700315010
transform 1 0 65250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1780_
timestamp 1700315010
transform 1 0 62550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1781_
timestamp 1700315010
transform 1 0 69450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1782_
timestamp 1700315010
transform 1 0 71850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1783_
timestamp 1700315010
transform 1 0 84150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1784_
timestamp 1700315010
transform 1 0 82050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1785_
timestamp 1700315010
transform -1 0 87150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1786_
timestamp 1700315010
transform 1 0 89250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1787_
timestamp 1700315010
transform -1 0 88350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1788_
timestamp 1700315010
transform 1 0 85650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1789_
timestamp 1700315010
transform 1 0 89850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1790_
timestamp 1700315010
transform 1 0 89850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1791_
timestamp 1700315010
transform 1 0 89550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1__1792_
timestamp 1700315010
transform 1 0 69750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1793_
timestamp 1700315010
transform 1 0 67650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1794_
timestamp 1700315010
transform 1 0 73050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1795_
timestamp 1700315010
transform -1 0 83550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1796_
timestamp 1700315010
transform 1 0 81150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1797_
timestamp 1700315010
transform -1 0 75450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1798_
timestamp 1700315010
transform -1 0 88050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1__1799_
timestamp 1700315010
transform -1 0 88050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1__1800_
timestamp 1700315010
transform -1 0 87750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1801_
timestamp 1700315010
transform 1 0 81150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1802_
timestamp 1700315010
transform 1 0 71250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1__1803_
timestamp 1700315010
transform 1 0 88050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1804_
timestamp 1700315010
transform -1 0 88350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1805_
timestamp 1700315010
transform 1 0 89850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1806_
timestamp 1700315010
transform -1 0 85350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1__1807_
timestamp 1700315010
transform 1 0 85050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1808_
timestamp 1700315010
transform 1 0 82950 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1809_
timestamp 1700315010
transform 1 0 84450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_1__1810_
timestamp 1700315010
transform 1 0 88350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_1__1811_
timestamp 1700315010
transform 1 0 85950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_1__1812_
timestamp 1700315010
transform 1 0 89550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1__1813_
timestamp 1700315010
transform -1 0 89850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1__1814_
timestamp 1700315010
transform -1 0 90150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1815_
timestamp 1700315010
transform 1 0 87450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1__1816_
timestamp 1700315010
transform -1 0 89850 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1817_
timestamp 1700315010
transform -1 0 88050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1__1818_
timestamp 1700315010
transform -1 0 49050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1819_
timestamp 1700315010
transform -1 0 38850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1__1820_
timestamp 1700315010
transform -1 0 69150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_1__1821_
timestamp 1700315010
transform -1 0 84450 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1822_
timestamp 1700315010
transform 1 0 82050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1823_
timestamp 1700315010
transform 1 0 80250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1824_
timestamp 1700315010
transform 1 0 74550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1825_
timestamp 1700315010
transform 1 0 68850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1__1826_
timestamp 1700315010
transform 1 0 86250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert0
timestamp 1700315010
transform 1 0 58950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert1
timestamp 1700315010
transform -1 0 33150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert2
timestamp 1700315010
transform -1 0 34950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert3
timestamp 1700315010
transform -1 0 34050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert4
timestamp 1700315010
transform -1 0 66150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert5
timestamp 1700315010
transform -1 0 56550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert6
timestamp 1700315010
transform -1 0 40950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert7
timestamp 1700315010
transform -1 0 51150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert13
timestamp 1700315010
transform 1 0 77850 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert14
timestamp 1700315010
transform -1 0 57450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert15
timestamp 1700315010
transform -1 0 65250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert16
timestamp 1700315010
transform -1 0 60450 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert17
timestamp 1700315010
transform 1 0 37950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert18
timestamp 1700315010
transform -1 0 35250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert19
timestamp 1700315010
transform 1 0 45450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert20
timestamp 1700315010
transform -1 0 36450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert21
timestamp 1700315010
transform 1 0 79950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert22
timestamp 1700315010
transform -1 0 63150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert23
timestamp 1700315010
transform 1 0 63750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert24
timestamp 1700315010
transform 1 0 79350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert25
timestamp 1700315010
transform -1 0 35250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert26
timestamp 1700315010
transform -1 0 39750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert27
timestamp 1700315010
transform -1 0 36150 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert28
timestamp 1700315010
transform 1 0 47550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert29
timestamp 1700315010
transform -1 0 32850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert30
timestamp 1700315010
transform 1 0 50850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert31
timestamp 1700315010
transform -1 0 33150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert32
timestamp 1700315010
transform 1 0 52650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert33
timestamp 1700315010
transform -1 0 76350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert34
timestamp 1700315010
transform -1 0 90150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert35
timestamp 1700315010
transform -1 0 74250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_1_BUFX2_insert36
timestamp 1700315010
transform -1 0 89250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1700315010
transform -1 0 68250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 74250 0 1 43050
box -180 -120 480 4080
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 87150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1700315010
transform -1 0 77850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 74550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__889_
timestamp 1700315010
transform 1 0 80550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__890_
timestamp 1700315010
transform -1 0 74850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__892_
timestamp 1700315010
transform 1 0 80850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__893_
timestamp 1700315010
transform -1 0 78750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__894_
timestamp 1700315010
transform 1 0 82650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__896_
timestamp 1700315010
transform -1 0 76950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__897_
timestamp 1700315010
transform 1 0 76950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__899_
timestamp 1700315010
transform 1 0 79050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__900_
timestamp 1700315010
transform -1 0 88050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__902_
timestamp 1700315010
transform 1 0 87150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__903_
timestamp 1700315010
transform 1 0 73650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__905_
timestamp 1700315010
transform -1 0 85650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__906_
timestamp 1700315010
transform -1 0 63450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__908_
timestamp 1700315010
transform 1 0 89550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__909_
timestamp 1700315010
transform 1 0 84150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__911_
timestamp 1700315010
transform 1 0 81450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__912_
timestamp 1700315010
transform 1 0 86550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__914_
timestamp 1700315010
transform -1 0 79050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__915_
timestamp 1700315010
transform 1 0 78750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__916_
timestamp 1700315010
transform -1 0 84750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__918_
timestamp 1700315010
transform -1 0 81150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__919_
timestamp 1700315010
transform 1 0 81150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__921_
timestamp 1700315010
transform 1 0 85050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__922_
timestamp 1700315010
transform 1 0 80850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__924_
timestamp 1700315010
transform 1 0 88650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__925_
timestamp 1700315010
transform -1 0 89850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__927_
timestamp 1700315010
transform 1 0 73050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__928_
timestamp 1700315010
transform 1 0 70650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__930_
timestamp 1700315010
transform 1 0 55350 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__931_
timestamp 1700315010
transform -1 0 57750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__933_
timestamp 1700315010
transform -1 0 66450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__934_
timestamp 1700315010
transform 1 0 68250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__936_
timestamp 1700315010
transform 1 0 61350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__937_
timestamp 1700315010
transform -1 0 60150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__939_
timestamp 1700315010
transform 1 0 55050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__940_
timestamp 1700315010
transform 1 0 52050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__941_
timestamp 1700315010
transform -1 0 49050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__943_
timestamp 1700315010
transform 1 0 52350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__944_
timestamp 1700315010
transform -1 0 79950 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__946_
timestamp 1700315010
transform 1 0 81450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__947_
timestamp 1700315010
transform 1 0 85050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__949_
timestamp 1700315010
transform 1 0 76650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__950_
timestamp 1700315010
transform -1 0 70050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__952_
timestamp 1700315010
transform 1 0 35250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__953_
timestamp 1700315010
transform 1 0 39750 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__955_
timestamp 1700315010
transform 1 0 41550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__956_
timestamp 1700315010
transform 1 0 47850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__958_
timestamp 1700315010
transform 1 0 54450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__959_
timestamp 1700315010
transform 1 0 54450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__961_
timestamp 1700315010
transform -1 0 52350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__962_
timestamp 1700315010
transform 1 0 56850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__963_
timestamp 1700315010
transform 1 0 43950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__965_
timestamp 1700315010
transform 1 0 37650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__966_
timestamp 1700315010
transform 1 0 50250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__968_
timestamp 1700315010
transform 1 0 38850 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__969_
timestamp 1700315010
transform -1 0 41850 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__971_
timestamp 1700315010
transform 1 0 45750 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__972_
timestamp 1700315010
transform -1 0 48150 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__974_
timestamp 1700315010
transform -1 0 52650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__975_
timestamp 1700315010
transform 1 0 46050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__977_
timestamp 1700315010
transform 1 0 31950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__978_
timestamp 1700315010
transform 1 0 37650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__980_
timestamp 1700315010
transform 1 0 43650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__981_
timestamp 1700315010
transform 1 0 54750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__983_
timestamp 1700315010
transform -1 0 41550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__984_
timestamp 1700315010
transform -1 0 36750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__985_
timestamp 1700315010
transform -1 0 35550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__987_
timestamp 1700315010
transform -1 0 24150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__988_
timestamp 1700315010
transform -1 0 20850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__990_
timestamp 1700315010
transform 1 0 28050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__991_
timestamp 1700315010
transform 1 0 36150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__993_
timestamp 1700315010
transform 1 0 30450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__994_
timestamp 1700315010
transform 1 0 39150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__996_
timestamp 1700315010
transform 1 0 25650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__997_
timestamp 1700315010
transform -1 0 21750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__999_
timestamp 1700315010
transform 1 0 33150 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1001_
timestamp 1700315010
transform 1 0 41850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1002_
timestamp 1700315010
transform 1 0 35250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1004_
timestamp 1700315010
transform 1 0 37350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1005_
timestamp 1700315010
transform -1 0 35250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1007_
timestamp 1700315010
transform -1 0 25350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1008_
timestamp 1700315010
transform 1 0 26850 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1009_
timestamp 1700315010
transform -1 0 29550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1011_
timestamp 1700315010
transform -1 0 33450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1012_
timestamp 1700315010
transform -1 0 22350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1014_
timestamp 1700315010
transform -1 0 33150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1015_
timestamp 1700315010
transform -1 0 31050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1017_
timestamp 1700315010
transform 1 0 33150 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1018_
timestamp 1700315010
transform -1 0 35850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1020_
timestamp 1700315010
transform -1 0 22950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1021_
timestamp 1700315010
transform -1 0 21750 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1023_
timestamp 1700315010
transform 1 0 17250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1024_
timestamp 1700315010
transform 1 0 22650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1026_
timestamp 1700315010
transform 1 0 19050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1027_
timestamp 1700315010
transform 1 0 22650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1029_
timestamp 1700315010
transform -1 0 13950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1030_
timestamp 1700315010
transform -1 0 24150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1032_
timestamp 1700315010
transform -1 0 18750 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1033_
timestamp 1700315010
transform -1 0 16350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1034_
timestamp 1700315010
transform -1 0 25050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1036_
timestamp 1700315010
transform -1 0 17850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1037_
timestamp 1700315010
transform -1 0 16050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1039_
timestamp 1700315010
transform -1 0 20250 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1040_
timestamp 1700315010
transform -1 0 31050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1042_
timestamp 1700315010
transform 1 0 28650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1043_
timestamp 1700315010
transform 1 0 34650 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1045_
timestamp 1700315010
transform 1 0 31650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1046_
timestamp 1700315010
transform -1 0 24450 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1048_
timestamp 1700315010
transform -1 0 29550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1049_
timestamp 1700315010
transform -1 0 22050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1051_
timestamp 1700315010
transform -1 0 10650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1052_
timestamp 1700315010
transform 1 0 18150 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1054_
timestamp 1700315010
transform -1 0 20850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1055_
timestamp 1700315010
transform -1 0 14550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1056_
timestamp 1700315010
transform 1 0 15150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1058_
timestamp 1700315010
transform 1 0 19050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1059_
timestamp 1700315010
transform 1 0 16650 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1061_
timestamp 1700315010
transform -1 0 44250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1062_
timestamp 1700315010
transform -1 0 28950 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1064_
timestamp 1700315010
transform 1 0 20850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1065_
timestamp 1700315010
transform -1 0 14250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1067_
timestamp 1700315010
transform 1 0 19650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1068_
timestamp 1700315010
transform -1 0 13050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1070_
timestamp 1700315010
transform 1 0 29550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1071_
timestamp 1700315010
transform 1 0 23850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1073_
timestamp 1700315010
transform -1 0 14550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1074_
timestamp 1700315010
transform -1 0 12150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1076_
timestamp 1700315010
transform -1 0 14850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1077_
timestamp 1700315010
transform 1 0 16950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1079_
timestamp 1700315010
transform -1 0 13650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1080_
timestamp 1700315010
transform -1 0 13050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1081_
timestamp 1700315010
transform -1 0 3450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1083_
timestamp 1700315010
transform -1 0 11550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1084_
timestamp 1700315010
transform -1 0 5850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1086_
timestamp 1700315010
transform 1 0 10350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1087_
timestamp 1700315010
transform 1 0 7950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1089_
timestamp 1700315010
transform 1 0 29550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1090_
timestamp 1700315010
transform 1 0 23550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1092_
timestamp 1700315010
transform -1 0 30750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1093_
timestamp 1700315010
transform 1 0 28350 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1095_
timestamp 1700315010
transform -1 0 28050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1096_
timestamp 1700315010
transform -1 0 25650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1098_
timestamp 1700315010
transform -1 0 26250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1099_
timestamp 1700315010
transform -1 0 21750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1101_
timestamp 1700315010
transform -1 0 1050 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1102_
timestamp 1700315010
transform -1 0 14250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1103_
timestamp 1700315010
transform 1 0 9450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1105_
timestamp 1700315010
transform 1 0 2850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1106_
timestamp 1700315010
transform -1 0 1050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1108_
timestamp 1700315010
transform 1 0 13350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1109_
timestamp 1700315010
transform -1 0 5550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1111_
timestamp 1700315010
transform -1 0 1050 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1112_
timestamp 1700315010
transform -1 0 30750 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1114_
timestamp 1700315010
transform -1 0 26850 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1115_
timestamp 1700315010
transform -1 0 7950 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1117_
timestamp 1700315010
transform 1 0 11550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1118_
timestamp 1700315010
transform -1 0 5550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1120_
timestamp 1700315010
transform 1 0 7350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1121_
timestamp 1700315010
transform 1 0 13650 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1123_
timestamp 1700315010
transform -1 0 10050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1124_
timestamp 1700315010
transform 1 0 7950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1126_
timestamp 1700315010
transform -1 0 1050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1127_
timestamp 1700315010
transform 1 0 8850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1128_
timestamp 1700315010
transform -1 0 5250 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1130_
timestamp 1700315010
transform 1 0 5550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1131_
timestamp 1700315010
transform -1 0 5550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1133_
timestamp 1700315010
transform -1 0 1050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1134_
timestamp 1700315010
transform -1 0 3450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1136_
timestamp 1700315010
transform -1 0 4950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1137_
timestamp 1700315010
transform -1 0 1050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1139_
timestamp 1700315010
transform 1 0 9150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1140_
timestamp 1700315010
transform 1 0 27150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1142_
timestamp 1700315010
transform 1 0 37950 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1143_
timestamp 1700315010
transform 1 0 49950 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1145_
timestamp 1700315010
transform 1 0 45450 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1146_
timestamp 1700315010
transform -1 0 50550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1148_
timestamp 1700315010
transform 1 0 47850 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1149_
timestamp 1700315010
transform -1 0 48150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1150_
timestamp 1700315010
transform 1 0 42450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1152_
timestamp 1700315010
transform -1 0 47850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1153_
timestamp 1700315010
transform 1 0 35550 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1155_
timestamp 1700315010
transform 1 0 40050 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1156_
timestamp 1700315010
transform -1 0 40050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1158_
timestamp 1700315010
transform 1 0 17850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1159_
timestamp 1700315010
transform -1 0 26250 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1161_
timestamp 1700315010
transform 1 0 11550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1162_
timestamp 1700315010
transform 1 0 20250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1164_
timestamp 1700315010
transform 1 0 56550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1165_
timestamp 1700315010
transform -1 0 58950 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1167_
timestamp 1700315010
transform 1 0 64650 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1168_
timestamp 1700315010
transform -1 0 52350 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1170_
timestamp 1700315010
transform 1 0 52650 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1171_
timestamp 1700315010
transform 1 0 61050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1173_
timestamp 1700315010
transform 1 0 61050 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1174_
timestamp 1700315010
transform 1 0 54150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1175_
timestamp 1700315010
transform -1 0 56850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1177_
timestamp 1700315010
transform -1 0 45150 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1178_
timestamp 1700315010
transform -1 0 44850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1180_
timestamp 1700315010
transform 1 0 31950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1181_
timestamp 1700315010
transform 1 0 49650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1183_
timestamp 1700315010
transform 1 0 57150 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1184_
timestamp 1700315010
transform -1 0 55050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1186_
timestamp 1700315010
transform 1 0 60750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1187_
timestamp 1700315010
transform -1 0 50250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1189_
timestamp 1700315010
transform 1 0 56550 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1190_
timestamp 1700315010
transform 1 0 58350 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1192_
timestamp 1700315010
transform 1 0 67350 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1193_
timestamp 1700315010
transform 1 0 65550 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1195_
timestamp 1700315010
transform 1 0 67350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1196_
timestamp 1700315010
transform 1 0 58950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1197_
timestamp 1700315010
transform -1 0 61650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1199_
timestamp 1700315010
transform 1 0 42150 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1200_
timestamp 1700315010
transform 1 0 52650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1202_
timestamp 1700315010
transform 1 0 61050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1203_
timestamp 1700315010
transform 1 0 53250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1205_
timestamp 1700315010
transform 1 0 40350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1206_
timestamp 1700315010
transform -1 0 1050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1208_
timestamp 1700315010
transform -1 0 1050 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1209_
timestamp 1700315010
transform 1 0 35850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1211_
timestamp 1700315010
transform -1 0 32850 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1212_
timestamp 1700315010
transform 1 0 27750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1214_
timestamp 1700315010
transform 1 0 33450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1215_
timestamp 1700315010
transform -1 0 21150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1217_
timestamp 1700315010
transform 1 0 30150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1218_
timestamp 1700315010
transform -1 0 27450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1219_
timestamp 1700315010
transform 1 0 18750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1221_
timestamp 1700315010
transform -1 0 23250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1222_
timestamp 1700315010
transform -1 0 28950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1224_
timestamp 1700315010
transform -1 0 31950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1225_
timestamp 1700315010
transform 1 0 29250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1227_
timestamp 1700315010
transform 1 0 23850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1228_
timestamp 1700315010
transform 1 0 29850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1230_
timestamp 1700315010
transform 1 0 28050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1231_
timestamp 1700315010
transform -1 0 25950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1233_
timestamp 1700315010
transform 1 0 4950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1234_
timestamp 1700315010
transform 1 0 16950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1236_
timestamp 1700315010
transform -1 0 4650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1237_
timestamp 1700315010
transform 1 0 8850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1239_
timestamp 1700315010
transform -1 0 7950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1240_
timestamp 1700315010
transform -1 0 6750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1242_
timestamp 1700315010
transform 1 0 9750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1243_
timestamp 1700315010
transform 1 0 5550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1244_
timestamp 1700315010
transform 1 0 3150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1246_
timestamp 1700315010
transform -1 0 1050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1247_
timestamp 1700315010
transform -1 0 1050 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1249_
timestamp 1700315010
transform 1 0 750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1250_
timestamp 1700315010
transform -1 0 3450 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1252_
timestamp 1700315010
transform 1 0 7350 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1253_
timestamp 1700315010
transform 1 0 750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1255_
timestamp 1700315010
transform -1 0 1050 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1256_
timestamp 1700315010
transform 1 0 5250 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1258_
timestamp 1700315010
transform 1 0 5550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1259_
timestamp 1700315010
transform -1 0 12750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1261_
timestamp 1700315010
transform 1 0 14550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1262_
timestamp 1700315010
transform 1 0 3150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1264_
timestamp 1700315010
transform 1 0 7650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1265_
timestamp 1700315010
transform -1 0 10350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1266_
timestamp 1700315010
transform -1 0 10050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1268_
timestamp 1700315010
transform 1 0 16350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1269_
timestamp 1700315010
transform 1 0 18750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1271_
timestamp 1700315010
transform -1 0 46650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1272_
timestamp 1700315010
transform 1 0 75150 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1274_
timestamp 1700315010
transform 1 0 62550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1275_
timestamp 1700315010
transform 1 0 59550 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1277_
timestamp 1700315010
transform 1 0 61950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1278_
timestamp 1700315010
transform 1 0 71550 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1280_
timestamp 1700315010
transform -1 0 53550 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1281_
timestamp 1700315010
transform -1 0 58050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1283_
timestamp 1700315010
transform -1 0 55650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1284_
timestamp 1700315010
transform -1 0 25050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1286_
timestamp 1700315010
transform -1 0 22950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1287_
timestamp 1700315010
transform 1 0 28650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1289_
timestamp 1700315010
transform 1 0 42750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1290_
timestamp 1700315010
transform -1 0 47550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1291_
timestamp 1700315010
transform -1 0 36150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1293_
timestamp 1700315010
transform -1 0 39750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1294_
timestamp 1700315010
transform 1 0 19050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1296_
timestamp 1700315010
transform -1 0 25050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1297_
timestamp 1700315010
transform 1 0 24450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1299_
timestamp 1700315010
transform 1 0 11850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1300_
timestamp 1700315010
transform -1 0 24450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1302_
timestamp 1700315010
transform -1 0 28950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1303_
timestamp 1700315010
transform -1 0 31350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1305_
timestamp 1700315010
transform -1 0 21450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1306_
timestamp 1700315010
transform 1 0 11850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1308_
timestamp 1700315010
transform -1 0 1050 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1309_
timestamp 1700315010
transform 1 0 19950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1311_
timestamp 1700315010
transform 1 0 16650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1312_
timestamp 1700315010
transform -1 0 26550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1313_
timestamp 1700315010
transform -1 0 20550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1315_
timestamp 1700315010
transform 1 0 19650 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1316_
timestamp 1700315010
transform -1 0 11850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1318_
timestamp 1700315010
transform 1 0 41850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1319_
timestamp 1700315010
transform -1 0 31050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1321_
timestamp 1700315010
transform -1 0 24450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1322_
timestamp 1700315010
transform -1 0 17550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1324_
timestamp 1700315010
transform -1 0 12450 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1325_
timestamp 1700315010
transform -1 0 15450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1327_
timestamp 1700315010
transform -1 0 1050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1328_
timestamp 1700315010
transform -1 0 1050 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1330_
timestamp 1700315010
transform -1 0 7650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1331_
timestamp 1700315010
transform 1 0 2850 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1333_
timestamp 1700315010
transform 1 0 12150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1334_
timestamp 1700315010
transform 1 0 7650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1336_
timestamp 1700315010
transform 1 0 7350 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1337_
timestamp 1700315010
transform 1 0 16950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1338_
timestamp 1700315010
transform 1 0 750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1340_
timestamp 1700315010
transform 1 0 9750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1341_
timestamp 1700315010
transform 1 0 2550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1343_
timestamp 1700315010
transform 1 0 4950 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1344_
timestamp 1700315010
transform -1 0 13350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1346_
timestamp 1700315010
transform 1 0 13650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1347_
timestamp 1700315010
transform 1 0 15450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1349_
timestamp 1700315010
transform -1 0 21150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1350_
timestamp 1700315010
transform 1 0 7950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1352_
timestamp 1700315010
transform 1 0 26250 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1353_
timestamp 1700315010
transform -1 0 18150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1355_
timestamp 1700315010
transform -1 0 32550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1356_
timestamp 1700315010
transform 1 0 49350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1358_
timestamp 1700315010
transform 1 0 53850 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1359_
timestamp 1700315010
transform 1 0 68550 0 -1 27450
box -180 -120 480 4080
use FILL  FILL_2__1360_
timestamp 1700315010
transform 1 0 67650 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1362_
timestamp 1700315010
transform 1 0 65250 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1363_
timestamp 1700315010
transform -1 0 61050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1365_
timestamp 1700315010
transform -1 0 72450 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1366_
timestamp 1700315010
transform -1 0 23550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1368_
timestamp 1700315010
transform 1 0 31650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1369_
timestamp 1700315010
transform 1 0 43950 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1371_
timestamp 1700315010
transform 1 0 37650 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1372_
timestamp 1700315010
transform -1 0 19350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1374_
timestamp 1700315010
transform -1 0 7950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1375_
timestamp 1700315010
transform -1 0 5250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1377_
timestamp 1700315010
transform -1 0 13350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1378_
timestamp 1700315010
transform -1 0 17850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1380_
timestamp 1700315010
transform -1 0 17550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1381_
timestamp 1700315010
transform -1 0 15150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1383_
timestamp 1700315010
transform -1 0 15150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1384_
timestamp 1700315010
transform -1 0 17550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1385_
timestamp 1700315010
transform -1 0 12750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1387_
timestamp 1700315010
transform 1 0 9450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1388_
timestamp 1700315010
transform 1 0 23850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1390_
timestamp 1700315010
transform -1 0 25350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1391_
timestamp 1700315010
transform -1 0 22650 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1393_
timestamp 1700315010
transform 1 0 28350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1394_
timestamp 1700315010
transform 1 0 20850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1396_
timestamp 1700315010
transform -1 0 8850 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1397_
timestamp 1700315010
transform -1 0 1050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1399_
timestamp 1700315010
transform -1 0 10350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1400_
timestamp 1700315010
transform -1 0 4650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1402_
timestamp 1700315010
transform -1 0 2550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1403_
timestamp 1700315010
transform 1 0 5250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1405_
timestamp 1700315010
transform 1 0 5250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1406_
timestamp 1700315010
transform -1 0 1050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1407_
timestamp 1700315010
transform -1 0 1050 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1409_
timestamp 1700315010
transform -1 0 3450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1410_
timestamp 1700315010
transform 1 0 3150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1412_
timestamp 1700315010
transform 1 0 9450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1413_
timestamp 1700315010
transform -1 0 1050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1415_
timestamp 1700315010
transform -1 0 19650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1416_
timestamp 1700315010
transform 1 0 28650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1418_
timestamp 1700315010
transform -1 0 18450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1419_
timestamp 1700315010
transform 1 0 20550 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1421_
timestamp 1700315010
transform -1 0 37050 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1422_
timestamp 1700315010
transform 1 0 41850 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1424_
timestamp 1700315010
transform 1 0 43050 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1425_
timestamp 1700315010
transform -1 0 45150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1427_
timestamp 1700315010
transform 1 0 69150 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1428_
timestamp 1700315010
transform -1 0 64650 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1429_
timestamp 1700315010
transform 1 0 65250 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1431_
timestamp 1700315010
transform -1 0 70950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1432_
timestamp 1700315010
transform 1 0 71250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1434_
timestamp 1700315010
transform 1 0 69750 0 1 19650
box -180 -120 480 4080
use FILL  FILL_2__1435_
timestamp 1700315010
transform 1 0 89250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1437_
timestamp 1700315010
transform -1 0 58350 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1438_
timestamp 1700315010
transform 1 0 40050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1440_
timestamp 1700315010
transform -1 0 18150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1441_
timestamp 1700315010
transform 1 0 7650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1443_
timestamp 1700315010
transform -1 0 31350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1444_
timestamp 1700315010
transform -1 0 21450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1446_
timestamp 1700315010
transform 1 0 23250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1447_
timestamp 1700315010
transform 1 0 25350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1449_
timestamp 1700315010
transform -1 0 28950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1450_
timestamp 1700315010
transform -1 0 23550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1452_
timestamp 1700315010
transform 1 0 28650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1453_
timestamp 1700315010
transform 1 0 31350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1454_
timestamp 1700315010
transform 1 0 28950 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1456_
timestamp 1700315010
transform -1 0 32550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1457_
timestamp 1700315010
transform -1 0 29550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1459_
timestamp 1700315010
transform -1 0 7350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1460_
timestamp 1700315010
transform 1 0 26250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1462_
timestamp 1700315010
transform -1 0 2850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1463_
timestamp 1700315010
transform -1 0 21750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1465_
timestamp 1700315010
transform -1 0 15750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1466_
timestamp 1700315010
transform -1 0 9150 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1468_
timestamp 1700315010
transform 1 0 21750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1469_
timestamp 1700315010
transform -1 0 16950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1471_
timestamp 1700315010
transform 1 0 11850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1472_
timestamp 1700315010
transform 1 0 14250 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1474_
timestamp 1700315010
transform 1 0 41850 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1475_
timestamp 1700315010
transform 1 0 41250 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1476_
timestamp 1700315010
transform 1 0 44850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1478_
timestamp 1700315010
transform 1 0 48750 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1479_
timestamp 1700315010
transform 1 0 52950 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1481_
timestamp 1700315010
transform -1 0 65550 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1482_
timestamp 1700315010
transform 1 0 69750 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1484_
timestamp 1700315010
transform -1 0 82950 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1485_
timestamp 1700315010
transform 1 0 82650 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1487_
timestamp 1700315010
transform 1 0 87450 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1488_
timestamp 1700315010
transform 1 0 32850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1490_
timestamp 1700315010
transform -1 0 35550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1491_
timestamp 1700315010
transform -1 0 43350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1493_
timestamp 1700315010
transform -1 0 34050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1494_
timestamp 1700315010
transform 1 0 38550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1496_
timestamp 1700315010
transform 1 0 36150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1497_
timestamp 1700315010
transform 1 0 39150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1499_
timestamp 1700315010
transform 1 0 33450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1500_
timestamp 1700315010
transform 1 0 36750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1501_
timestamp 1700315010
transform 1 0 40950 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1503_
timestamp 1700315010
transform 1 0 41850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1504_
timestamp 1700315010
transform 1 0 43050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1506_
timestamp 1700315010
transform -1 0 39750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1507_
timestamp 1700315010
transform -1 0 37350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1509_
timestamp 1700315010
transform 1 0 30750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1510_
timestamp 1700315010
transform -1 0 28950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1512_
timestamp 1700315010
transform -1 0 40950 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1513_
timestamp 1700315010
transform 1 0 49950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1515_
timestamp 1700315010
transform 1 0 47550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1516_
timestamp 1700315010
transform -1 0 38250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1518_
timestamp 1700315010
transform -1 0 48450 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1519_
timestamp 1700315010
transform 1 0 43950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1521_
timestamp 1700315010
transform 1 0 38550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1522_
timestamp 1700315010
transform 1 0 40950 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1523_
timestamp 1700315010
transform 1 0 42750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1525_
timestamp 1700315010
transform -1 0 82350 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1526_
timestamp 1700315010
transform -1 0 74850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1528_
timestamp 1700315010
transform 1 0 64950 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1529_
timestamp 1700315010
transform 1 0 68850 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1531_
timestamp 1700315010
transform -1 0 76350 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1532_
timestamp 1700315010
transform 1 0 78450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1534_
timestamp 1700315010
transform -1 0 77550 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1535_
timestamp 1700315010
transform -1 0 56550 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1537_
timestamp 1700315010
transform 1 0 42150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1538_
timestamp 1700315010
transform 1 0 38850 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1540_
timestamp 1700315010
transform -1 0 39750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1541_
timestamp 1700315010
transform -1 0 42150 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1543_
timestamp 1700315010
transform 1 0 39750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1544_
timestamp 1700315010
transform 1 0 36750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1546_
timestamp 1700315010
transform -1 0 37650 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1547_
timestamp 1700315010
transform -1 0 40350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1548_
timestamp 1700315010
transform -1 0 45750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1550_
timestamp 1700315010
transform 1 0 52050 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1551_
timestamp 1700315010
transform 1 0 58650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1553_
timestamp 1700315010
transform -1 0 76050 0 1 27450
box -180 -120 480 4080
use FILL  FILL_2__1554_
timestamp 1700315010
transform 1 0 78450 0 -1 19650
box -180 -120 480 4080
use FILL  FILL_2__1556_
timestamp 1700315010
transform -1 0 74850 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1557_
timestamp 1700315010
transform -1 0 73050 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1559_
timestamp 1700315010
transform 1 0 52950 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1560_
timestamp 1700315010
transform 1 0 54750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1562_
timestamp 1700315010
transform 1 0 40350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1563_
timestamp 1700315010
transform 1 0 55650 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1565_
timestamp 1700315010
transform -1 0 32550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1566_
timestamp 1700315010
transform -1 0 34650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1568_
timestamp 1700315010
transform 1 0 49950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1569_
timestamp 1700315010
transform 1 0 59250 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1570_
timestamp 1700315010
transform 1 0 50550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1572_
timestamp 1700315010
transform 1 0 51750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1573_
timestamp 1700315010
transform 1 0 61650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1575_
timestamp 1700315010
transform 1 0 64950 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1576_
timestamp 1700315010
transform 1 0 62550 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1578_
timestamp 1700315010
transform 1 0 85650 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1579_
timestamp 1700315010
transform -1 0 76950 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1581_
timestamp 1700315010
transform 1 0 73350 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1582_
timestamp 1700315010
transform -1 0 67650 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1584_
timestamp 1700315010
transform 1 0 44250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1585_
timestamp 1700315010
transform 1 0 46650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1587_
timestamp 1700315010
transform 1 0 38250 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1588_
timestamp 1700315010
transform -1 0 58050 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1590_
timestamp 1700315010
transform 1 0 71850 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2__1591_
timestamp 1700315010
transform -1 0 71250 0 -1 11850
box -180 -120 480 4080
use FILL  FILL_2__1593_
timestamp 1700315010
transform -1 0 65250 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2__1594_
timestamp 1700315010
transform 1 0 64650 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1595_
timestamp 1700315010
transform 1 0 59850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1597_
timestamp 1700315010
transform 1 0 60150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1598_
timestamp 1700315010
transform -1 0 62550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1600_
timestamp 1700315010
transform -1 0 60450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1601_
timestamp 1700315010
transform 1 0 49650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1603_
timestamp 1700315010
transform 1 0 44250 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1604_
timestamp 1700315010
transform -1 0 46650 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1606_
timestamp 1700315010
transform -1 0 77550 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1607_
timestamp 1700315010
transform 1 0 66450 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1636_
timestamp 1700315010
transform -1 0 88650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1637_
timestamp 1700315010
transform 1 0 88650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1639_
timestamp 1700315010
transform 1 0 78150 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1640_
timestamp 1700315010
transform 1 0 78150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1642_
timestamp 1700315010
transform -1 0 47550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1643_
timestamp 1700315010
transform -1 0 45150 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1644_
timestamp 1700315010
transform -1 0 58050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1646_
timestamp 1700315010
transform -1 0 61650 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1647_
timestamp 1700315010
transform 1 0 47550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1649_
timestamp 1700315010
transform -1 0 64350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1650_
timestamp 1700315010
transform -1 0 66750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1652_
timestamp 1700315010
transform -1 0 54450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1653_
timestamp 1700315010
transform 1 0 62250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1655_
timestamp 1700315010
transform -1 0 85050 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1656_
timestamp 1700315010
transform 1 0 88950 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1658_
timestamp 1700315010
transform 1 0 84450 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1659_
timestamp 1700315010
transform -1 0 80250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1661_
timestamp 1700315010
transform 1 0 80250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1662_
timestamp 1700315010
transform -1 0 52050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1664_
timestamp 1700315010
transform -1 0 51750 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1665_
timestamp 1700315010
transform -1 0 54750 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1666_
timestamp 1700315010
transform -1 0 57450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1668_
timestamp 1700315010
transform 1 0 55650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1669_
timestamp 1700315010
transform -1 0 60750 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1671_
timestamp 1700315010
transform 1 0 78450 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1672_
timestamp 1700315010
transform -1 0 85050 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1674_
timestamp 1700315010
transform -1 0 80550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1675_
timestamp 1700315010
transform -1 0 83250 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1677_
timestamp 1700315010
transform -1 0 73350 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1678_
timestamp 1700315010
transform -1 0 73950 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1680_
timestamp 1700315010
transform 1 0 69450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1681_
timestamp 1700315010
transform -1 0 60150 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1683_
timestamp 1700315010
transform 1 0 70650 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1684_
timestamp 1700315010
transform 1 0 75450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1686_
timestamp 1700315010
transform 1 0 64650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1687_
timestamp 1700315010
transform -1 0 76650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1689_
timestamp 1700315010
transform 1 0 73350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1690_
timestamp 1700315010
transform 1 0 76350 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1691_
timestamp 1700315010
transform -1 0 74250 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1693_
timestamp 1700315010
transform 1 0 46650 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1694_
timestamp 1700315010
transform -1 0 49350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1696_
timestamp 1700315010
transform -1 0 45750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1697_
timestamp 1700315010
transform -1 0 49650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1699_
timestamp 1700315010
transform -1 0 58350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1700_
timestamp 1700315010
transform -1 0 58650 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1702_
timestamp 1700315010
transform 1 0 55950 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1703_
timestamp 1700315010
transform -1 0 68850 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1705_
timestamp 1700315010
transform 1 0 60750 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1706_
timestamp 1700315010
transform -1 0 65250 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1708_
timestamp 1700315010
transform 1 0 67350 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1709_
timestamp 1700315010
transform -1 0 55050 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1711_
timestamp 1700315010
transform -1 0 53550 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1712_
timestamp 1700315010
transform -1 0 55650 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1713_
timestamp 1700315010
transform -1 0 51150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1715_
timestamp 1700315010
transform -1 0 59250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1716_
timestamp 1700315010
transform 1 0 61350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1718_
timestamp 1700315010
transform 1 0 68550 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1719_
timestamp 1700315010
transform 1 0 70950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1721_
timestamp 1700315010
transform 1 0 70050 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2__1722_
timestamp 1700315010
transform 1 0 71550 0 1 89850
box -180 -120 480 4080
use FILL  FILL_2__1724_
timestamp 1700315010
transform -1 0 72150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1725_
timestamp 1700315010
transform 1 0 66450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1727_
timestamp 1700315010
transform -1 0 65850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1728_
timestamp 1700315010
transform -1 0 45450 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2__1730_
timestamp 1700315010
transform -1 0 48750 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1731_
timestamp 1700315010
transform -1 0 50850 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1733_
timestamp 1700315010
transform 1 0 55350 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1734_
timestamp 1700315010
transform 1 0 74550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1736_
timestamp 1700315010
transform -1 0 78750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1737_
timestamp 1700315010
transform 1 0 76050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1738_
timestamp 1700315010
transform 1 0 76650 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1740_
timestamp 1700315010
transform -1 0 77550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1741_
timestamp 1700315010
transform 1 0 78450 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1743_
timestamp 1700315010
transform -1 0 41850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1744_
timestamp 1700315010
transform -1 0 44250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1746_
timestamp 1700315010
transform 1 0 46050 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1747_
timestamp 1700315010
transform 1 0 50550 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1749_
timestamp 1700315010
transform 1 0 78450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1750_
timestamp 1700315010
transform 1 0 81750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1752_
timestamp 1700315010
transform -1 0 79350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1753_
timestamp 1700315010
transform 1 0 80850 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1755_
timestamp 1700315010
transform 1 0 80850 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1756_
timestamp 1700315010
transform 1 0 72750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1758_
timestamp 1700315010
transform 1 0 63750 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1759_
timestamp 1700315010
transform 1 0 60150 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1760_
timestamp 1700315010
transform 1 0 67950 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1762_
timestamp 1700315010
transform -1 0 77250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1763_
timestamp 1700315010
transform 1 0 79350 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1765_
timestamp 1700315010
transform 1 0 86250 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1766_
timestamp 1700315010
transform 1 0 87750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1768_
timestamp 1700315010
transform -1 0 71550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1769_
timestamp 1700315010
transform -1 0 69150 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1771_
timestamp 1700315010
transform 1 0 82950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1772_
timestamp 1700315010
transform 1 0 83250 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1774_
timestamp 1700315010
transform -1 0 84150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1775_
timestamp 1700315010
transform -1 0 85950 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1777_
timestamp 1700315010
transform 1 0 74250 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1778_
timestamp 1700315010
transform 1 0 67350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1780_
timestamp 1700315010
transform 1 0 62850 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1781_
timestamp 1700315010
transform 1 0 69750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1783_
timestamp 1700315010
transform 1 0 84450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1784_
timestamp 1700315010
transform 1 0 82350 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1785_
timestamp 1700315010
transform -1 0 87450 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1787_
timestamp 1700315010
transform -1 0 88650 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1788_
timestamp 1700315010
transform 1 0 85950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1790_
timestamp 1700315010
transform 1 0 90150 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1791_
timestamp 1700315010
transform 1 0 89850 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2__1793_
timestamp 1700315010
transform 1 0 67950 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2__1794_
timestamp 1700315010
transform 1 0 73350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1796_
timestamp 1700315010
transform 1 0 81450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1797_
timestamp 1700315010
transform -1 0 75750 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1799_
timestamp 1700315010
transform -1 0 88350 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2__1800_
timestamp 1700315010
transform -1 0 88050 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1802_
timestamp 1700315010
transform 1 0 71550 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2__1803_
timestamp 1700315010
transform 1 0 88350 0 1 4050
box -180 -120 480 4080
use FILL  FILL_2__1805_
timestamp 1700315010
transform 1 0 90150 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1806_
timestamp 1700315010
transform -1 0 85650 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2__1807_
timestamp 1700315010
transform 1 0 85350 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1809_
timestamp 1700315010
transform 1 0 84750 0 1 74250
box -180 -120 480 4080
use FILL  FILL_2__1810_
timestamp 1700315010
transform 1 0 88650 0 -1 74250
box -180 -120 480 4080
use FILL  FILL_2__1812_
timestamp 1700315010
transform 1 0 89850 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2__1813_
timestamp 1700315010
transform -1 0 90150 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2__1815_
timestamp 1700315010
transform 1 0 87750 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2__1816_
timestamp 1700315010
transform -1 0 90150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2__1818_
timestamp 1700315010
transform -1 0 49350 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1819_
timestamp 1700315010
transform -1 0 39150 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2__1821_
timestamp 1700315010
transform -1 0 84750 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1822_
timestamp 1700315010
transform 1 0 82350 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1824_
timestamp 1700315010
transform 1 0 74850 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2__1825_
timestamp 1700315010
transform 1 0 69150 0 -1 4050
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert0
timestamp 1700315010
transform 1 0 59250 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert1
timestamp 1700315010
transform -1 0 33450 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert3
timestamp 1700315010
transform -1 0 34350 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert4
timestamp 1700315010
transform -1 0 66450 0 -1 58650
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert6
timestamp 1700315010
transform -1 0 41250 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert7
timestamp 1700315010
transform -1 0 51450 0 -1 35250
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert13
timestamp 1700315010
transform 1 0 78150 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert14
timestamp 1700315010
transform -1 0 57750 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert16
timestamp 1700315010
transform -1 0 60750 0 -1 43050
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert17
timestamp 1700315010
transform 1 0 38250 0 1 58650
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert19
timestamp 1700315010
transform 1 0 45750 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert20
timestamp 1700315010
transform -1 0 36750 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert22
timestamp 1700315010
transform -1 0 63450 0 1 50850
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert23
timestamp 1700315010
transform 1 0 64050 0 -1 50850
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert25
timestamp 1700315010
transform -1 0 35550 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert26
timestamp 1700315010
transform -1 0 40050 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert28
timestamp 1700315010
transform 1 0 47850 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert29
timestamp 1700315010
transform -1 0 33150 0 1 35250
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert31
timestamp 1700315010
transform -1 0 33450 0 -1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert32
timestamp 1700315010
transform 1 0 52950 0 1 66450
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert34
timestamp 1700315010
transform -1 0 90450 0 -1 82050
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert35
timestamp 1700315010
transform -1 0 74550 0 -1 89850
box -180 -120 480 4080
use FILL  FILL_2_BUFX2_insert36
timestamp 1700315010
transform -1 0 89550 0 1 82050
box -180 -120 480 4080
use FILL  FILL_2_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 74550 0 1 43050
box -180 -120 480 4080
use FILL  FILL_2_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 87450 0 1 11850
box -180 -120 480 4080
use FILL  FILL_2_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 74850 0 -1 19650
box -180 -120 480 4080
<< labels >>
flabel metal1 s 92145 30 93045 30 3 FreeSans 240 270 0 0 gnd
port 0 nsew
flabel metal1 s -945 30 -45 30 7 FreeSans 240 270 0 0 vdd
port 1 nsew
flabel metal2 s 50040 94440 50160 94560 3 FreeSans 240 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal2 s 72840 94440 72960 94560 3 FreeSans 240 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal2 s 74340 94440 74460 94560 3 FreeSans 240 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal2 s 76740 94440 76860 94560 3 FreeSans 240 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal2 s 87240 94440 87360 94560 3 FreeSans 240 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal3 s 92640 81540 92760 81660 3 FreeSans 240 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal2 s 75540 -360 75660 -240 7 FreeSans 240 270 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 80940 -360 81060 -240 7 FreeSans 240 270 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 83040 -360 83160 -240 7 FreeSans 240 270 0 0 ACC_o[4]
port 13 nsew
flabel metal2 s 85140 -360 85260 -240 7 FreeSans 240 270 0 0 ACC_o[3]
port 14 nsew
flabel metal3 s -360 17640 -240 17760 7 FreeSans 240 0 0 0 ACC_o[2]
port 15 nsew
flabel metal3 s -360 33840 -240 33960 7 FreeSans 240 0 0 0 ACC_o[0]
port 17 nsew
flabel metal2 s 86940 -360 87060 -240 7 FreeSans 240 270 0 0 Done_o
port 18 nsew
flabel metal2 s 87840 94440 87960 94560 3 FreeSans 240 90 0 0 LoadCmd_i
port 21 nsew
flabel metal3 s 92640 13740 92760 13860 3 FreeSans 240 0 0 0 clk
port 22 nsew
flabel metal3 s 93045 79140 93165 79260 3 FreeSans 240 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal3 s 93045 77640 93165 77760 3 FreeSans 240 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal3 s 93045 20940 93165 21060 3 FreeSans 240 0 0 0 reset
port 23 nsew
flabel metal3 s -360 32940 -240 33060 7 FreeSans 240 0 0 0 ACC_o[1]
port 16 nsew
flabel metal2 s 69840 -360 69960 -240 7 FreeSans 240 270 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 90040 94440 90160 94560 3 FreeSans 240 90 0 0 LoadA_i
port 19 nsew
flabel metal2 s 88735 94440 88855 94560 3 FreeSans 240 90 0 0 LoadB_i
port 20 nsew
<< properties >>
string FIXED_BBOX -600 -600 92700 94500
<< end >>
