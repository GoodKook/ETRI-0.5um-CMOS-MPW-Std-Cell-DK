magic
tech scmos
magscale 1 2
timestamp 1728304916
<< nwell >>
rect -12 134 133 252
<< ntransistor >>
rect 21 14 25 54
rect 41 14 45 54
rect 61 14 65 54
rect 81 14 85 54
<< ptransistor >>
rect 21 146 25 226
rect 41 146 45 226
rect 61 146 65 226
rect 81 146 85 226
<< ndiffusion >>
rect 19 14 21 54
rect 25 14 27 54
rect 39 14 41 54
rect 45 14 47 54
rect 59 14 61 54
rect 65 14 67 54
rect 79 14 81 54
rect 85 14 87 54
<< pdiffusion >>
rect 19 146 21 226
rect 25 146 27 226
rect 39 146 41 226
rect 45 146 47 226
rect 59 146 61 226
rect 65 146 67 226
rect 79 146 81 226
rect 85 146 87 226
<< ndcontact >>
rect 7 14 19 54
rect 27 14 39 54
rect 47 14 59 54
rect 67 14 79 54
rect 87 14 99 54
<< pdcontact >>
rect 7 146 19 226
rect 27 146 39 226
rect 47 146 59 226
rect 67 146 79 226
rect 87 146 99 226
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 234 126 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 61 226 65 230
rect 81 226 85 230
rect 21 142 25 146
rect 41 142 45 146
rect 61 142 65 146
rect 81 142 85 146
rect 21 138 85 142
rect 21 123 27 138
rect 21 111 24 123
rect 21 62 27 111
rect 21 58 85 62
rect 21 54 25 58
rect 41 54 45 58
rect 61 54 65 58
rect 81 54 85 58
rect 21 10 25 14
rect 41 10 45 14
rect 61 10 65 14
rect 81 10 85 14
<< polycontact >>
rect 24 111 36 123
<< metal1 >>
rect -6 246 126 248
rect -6 232 126 234
rect 7 226 19 232
rect 47 226 59 232
rect 87 226 99 232
rect 27 140 39 146
rect 67 140 75 146
rect 27 134 75 140
rect 67 111 75 134
rect 67 68 75 97
rect 27 60 75 68
rect 27 54 35 60
rect 67 54 75 60
rect 7 8 19 14
rect 47 8 59 14
rect 87 8 99 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 23 97 37 111
rect 63 97 77 111
<< metal2 >>
rect 23 83 37 97
rect 63 83 77 97
<< m1p >>
rect -6 232 126 248
rect -6 -8 126 8
<< m2p >>
rect 23 83 37 97
rect 63 83 77 97
<< labels >>
rlabel metal1 -6 -8 126 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 -6 232 126 248 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal2 23 83 37 97 0 A
port 0 nsew signal input
rlabel metal2 63 83 77 97 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
