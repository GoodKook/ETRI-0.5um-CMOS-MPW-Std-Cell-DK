VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU_wrapper
  CLASS BLOCK ;
  FOREIGN ALU_wrapper ;
  ORIGIN 6.000 6.000 ;
  SIZE 933.000 BY 951.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 16.800 899.700 18.600 903.600 ;
        RECT 37.800 899.700 39.600 904.800 ;
        RECT 58.800 899.700 60.600 904.800 ;
        RECT 79.800 899.700 81.600 903.600 ;
        RECT 103.800 899.700 105.600 909.600 ;
        RECT 113.400 899.700 115.200 909.600 ;
        RECT 142.800 899.700 144.600 904.800 ;
        RECT 169.800 899.700 171.600 909.600 ;
        RECT 187.800 899.700 189.600 903.600 ;
        RECT 205.800 899.700 207.600 904.800 ;
        RECT 221.400 899.700 223.200 909.600 ;
        RECT 245.700 899.700 247.500 903.600 ;
        RECT 253.200 899.700 255.000 906.600 ;
        RECT 266.400 899.700 268.200 909.600 ;
        RECT 298.500 899.700 300.300 906.600 ;
        RECT 311.400 899.700 313.200 909.600 ;
        RECT 340.500 899.700 342.300 906.600 ;
        RECT 350.400 899.700 352.200 909.600 ;
        RECT 385.800 899.700 387.600 909.600 ;
        RECT 403.800 899.700 405.600 903.600 ;
        RECT 409.800 900.600 411.600 903.600 ;
        RECT 410.400 899.700 411.600 900.600 ;
        RECT 422.700 899.700 424.500 906.600 ;
        RECT 445.800 899.700 447.600 903.600 ;
        RECT 460.800 899.700 462.600 903.600 ;
        RECT 466.800 899.700 468.600 903.600 ;
        RECT 479.400 899.700 481.200 906.600 ;
        RECT 505.800 899.700 507.600 904.800 ;
        RECT 529.500 899.700 531.300 906.600 ;
        RECT 547.800 899.700 549.600 904.800 ;
        RECT 566.400 899.700 568.200 904.800 ;
        RECT 590.700 899.700 592.500 903.600 ;
        RECT 598.200 899.700 600.000 906.600 ;
        RECT 611.400 899.700 613.200 903.600 ;
        RECT 634.800 899.700 636.600 904.800 ;
        RECT 653.400 899.700 655.200 904.800 ;
        RECT 676.800 899.700 678.600 903.600 ;
        RECT 694.800 899.700 696.600 905.700 ;
        RECT 703.800 899.700 705.600 905.700 ;
        RECT 719.400 899.700 721.200 909.600 ;
        RECT 751.800 899.700 753.600 904.800 ;
        RECT 767.400 899.700 769.200 903.600 ;
        RECT 773.400 899.700 775.200 903.600 ;
        RECT 788.400 899.700 790.200 903.600 ;
        RECT 814.500 899.700 816.300 906.600 ;
        RECT 827.400 899.700 829.200 904.800 ;
        RECT 836.400 899.700 838.200 907.800 ;
        RECT 859.800 899.700 861.600 904.800 ;
        RECT 877.800 899.700 879.600 903.600 ;
        RECT 890.400 899.700 892.200 906.600 ;
        RECT 896.400 899.700 898.200 906.600 ;
        RECT 921.450 899.700 930.450 938.700 ;
        RECT 0.600 897.300 930.450 899.700 ;
        RECT 16.500 890.400 18.300 897.300 ;
        RECT 25.500 890.400 27.300 897.300 ;
        RECT 43.500 890.400 45.300 897.300 ;
        RECT 56.400 887.400 58.200 897.300 ;
        RECT 81.000 890.400 82.800 897.300 ;
        RECT 88.500 893.400 90.300 897.300 ;
        RECT 111.300 890.400 113.100 897.300 ;
        RECT 136.800 892.200 138.600 897.300 ;
        RECT 159.300 890.400 161.100 897.300 ;
        RECT 178.800 893.400 180.600 897.300 ;
        RECT 184.800 893.400 186.600 897.300 ;
        RECT 197.400 892.200 199.200 897.300 ;
        RECT 223.800 893.400 225.600 897.300 ;
        RECT 241.800 893.400 243.600 897.300 ;
        RECT 254.400 892.200 256.200 897.300 ;
        RECT 272.400 893.400 274.200 897.300 ;
        RECT 301.800 887.400 303.600 897.300 ;
        RECT 319.800 893.400 321.600 897.300 ;
        RECT 335.400 892.200 337.200 897.300 ;
        RECT 353.400 893.400 355.200 897.300 ;
        RECT 376.800 892.200 378.600 897.300 ;
        RECT 393.000 890.400 394.800 897.300 ;
        RECT 400.500 893.400 402.300 897.300 ;
        RECT 413.400 893.400 415.200 897.300 ;
        RECT 419.400 893.400 421.200 897.300 ;
        RECT 434.400 893.400 436.200 897.300 ;
        RECT 457.800 890.400 459.600 897.300 ;
        RECT 470.400 887.400 472.200 897.300 ;
        RECT 499.500 890.400 501.300 897.300 ;
        RECT 508.500 890.400 510.300 897.300 ;
        RECT 521.400 892.200 523.200 897.300 ;
        RECT 539.700 890.400 541.500 897.300 ;
        RECT 563.400 892.200 565.200 897.300 ;
        RECT 592.800 892.200 594.600 897.300 ;
        RECT 616.800 892.200 618.600 897.300 ;
        RECT 630.000 890.400 631.800 897.300 ;
        RECT 637.500 893.400 639.300 897.300 ;
        RECT 661.800 892.200 663.600 897.300 ;
        RECT 677.700 890.400 679.500 897.300 ;
        RECT 686.700 890.400 688.500 897.300 ;
        RECT 704.700 890.400 706.500 897.300 ;
        RECT 722.400 887.400 724.200 897.300 ;
        RECT 751.800 893.400 753.600 897.300 ;
        RECT 775.500 890.400 777.300 897.300 ;
        RECT 785.700 890.400 787.500 897.300 ;
        RECT 809.400 892.200 811.200 897.300 ;
        RECT 829.800 893.400 831.600 897.300 ;
        RECT 835.800 893.400 837.600 897.300 ;
        RECT 851.400 892.200 853.200 897.300 ;
        RECT 872.400 892.200 874.200 897.300 ;
        RECT 893.400 893.400 895.200 897.300 ;
        RECT 899.400 893.400 901.200 897.300 ;
        RECT 13.800 821.700 15.600 825.600 ;
        RECT 34.500 821.700 36.300 828.600 ;
        RECT 55.500 821.700 57.300 828.600 ;
        RECT 66.000 821.700 67.800 828.600 ;
        RECT 73.500 821.700 75.300 825.600 ;
        RECT 100.800 821.700 102.600 831.600 ;
        RECT 121.800 821.700 123.600 831.600 ;
        RECT 139.800 821.700 141.600 825.600 ;
        RECT 157.800 821.700 159.600 825.600 ;
        RECT 163.800 822.600 165.600 825.600 ;
        RECT 164.400 821.700 165.600 822.600 ;
        RECT 184.500 821.700 186.300 828.600 ;
        RECT 202.500 821.700 204.300 828.600 ;
        RECT 217.800 821.700 219.600 825.600 ;
        RECT 223.800 821.700 225.600 825.600 ;
        RECT 236.700 821.700 238.500 828.600 ;
        RECT 257.400 821.700 259.200 825.600 ;
        RECT 263.400 821.700 265.200 825.600 ;
        RECT 275.700 821.700 277.500 828.600 ;
        RECT 303.300 821.700 305.100 828.600 ;
        RECT 325.800 821.700 327.600 826.800 ;
        RECT 349.800 821.700 351.600 826.800 ;
        RECT 368.400 821.700 370.200 826.800 ;
        RECT 389.400 822.600 391.200 825.600 ;
        RECT 389.400 821.700 390.600 822.600 ;
        RECT 395.400 821.700 397.200 825.600 ;
        RECT 413.700 821.700 415.500 828.600 ;
        RECT 442.500 821.700 444.300 828.600 ;
        RECT 463.500 821.700 465.300 828.600 ;
        RECT 484.500 821.700 486.300 828.600 ;
        RECT 505.800 821.700 507.600 831.600 ;
        RECT 523.500 821.700 525.300 828.600 ;
        RECT 532.500 821.700 534.300 828.600 ;
        RECT 553.500 821.700 555.300 828.600 ;
        RECT 568.800 821.700 570.600 828.600 ;
        RECT 589.500 821.700 591.300 828.600 ;
        RECT 605.700 821.700 607.500 825.600 ;
        RECT 613.200 821.700 615.000 828.600 ;
        RECT 629.400 821.700 631.200 826.800 ;
        RECT 647.700 821.700 649.500 828.600 ;
        RECT 676.800 821.700 678.600 826.800 ;
        RECT 689.700 821.700 691.500 828.600 ;
        RECT 710.400 821.700 712.200 831.600 ;
        RECT 742.800 821.700 744.600 826.800 ;
        RECT 758.700 821.700 760.500 828.600 ;
        RECT 767.700 821.700 769.500 828.600 ;
        RECT 785.400 821.700 787.200 825.600 ;
        RECT 808.800 821.700 810.600 827.700 ;
        RECT 817.800 821.700 819.600 827.700 ;
        RECT 838.800 821.700 840.600 825.600 ;
        RECT 854.700 821.700 856.500 825.600 ;
        RECT 862.200 821.700 864.000 828.600 ;
        RECT 875.400 821.700 877.200 826.800 ;
        RECT 901.800 821.700 903.600 825.600 ;
        RECT 921.450 821.700 930.450 897.300 ;
        RECT 0.600 819.300 930.450 821.700 ;
        RECT 16.800 815.400 18.600 819.300 ;
        RECT 23.400 818.400 24.600 819.300 ;
        RECT 22.800 815.400 24.600 818.400 ;
        RECT 38.700 815.400 40.500 819.300 ;
        RECT 46.200 812.400 48.000 819.300 ;
        RECT 64.500 812.400 66.300 819.300 ;
        RECT 85.800 809.400 87.600 819.300 ;
        RECT 98.400 809.400 100.200 819.300 ;
        RECT 123.000 812.400 124.800 819.300 ;
        RECT 130.500 815.400 132.300 819.300 ;
        RECT 149.400 814.200 151.200 819.300 ;
        RECT 178.500 812.400 180.300 819.300 ;
        RECT 188.400 809.400 190.200 819.300 ;
        RECT 215.400 813.300 217.200 819.300 ;
        RECT 224.100 813.300 225.900 819.300 ;
        RECT 242.700 812.400 244.500 819.300 ;
        RECT 271.800 813.900 273.600 819.300 ;
        RECT 290.400 814.200 292.200 819.300 ;
        RECT 308.400 815.400 310.200 819.300 ;
        RECT 334.800 814.200 336.600 819.300 ;
        RECT 350.400 814.200 352.200 819.300 ;
        RECT 371.400 809.400 373.200 819.300 ;
        RECT 395.700 812.400 397.500 819.300 ;
        RECT 416.400 814.200 418.200 819.300 ;
        RECT 434.400 815.400 436.200 819.300 ;
        RECT 449.400 815.400 451.200 819.300 ;
        RECT 468.900 812.400 470.700 819.300 ;
        RECT 496.500 812.400 498.300 819.300 ;
        RECT 514.500 812.400 516.300 819.300 ;
        RECT 523.500 812.400 525.300 819.300 ;
        RECT 536.400 814.200 538.200 819.300 ;
        RECT 560.400 814.200 562.200 819.300 ;
        RECT 581.400 814.200 583.200 819.300 ;
        RECT 604.800 815.400 606.600 819.300 ;
        RECT 622.500 812.400 624.300 819.300 ;
        RECT 631.500 812.400 633.300 819.300 ;
        RECT 649.800 815.400 651.600 819.300 ;
        RECT 667.500 812.400 669.300 819.300 ;
        RECT 685.500 812.400 687.300 819.300 ;
        RECT 698.700 812.400 700.500 819.300 ;
        RECT 719.400 815.400 721.200 819.300 ;
        RECT 725.400 815.400 727.200 819.300 ;
        RECT 742.800 811.200 744.600 819.300 ;
        RECT 751.800 814.200 753.600 819.300 ;
        RECT 769.800 815.400 771.600 819.300 ;
        RECT 785.400 815.400 787.200 819.300 ;
        RECT 791.400 815.400 793.200 819.300 ;
        RECT 811.800 814.200 813.600 819.300 ;
        RECT 827.400 814.200 829.200 819.300 ;
        RECT 851.400 814.200 853.200 819.300 ;
        RECT 869.400 815.400 871.200 819.300 ;
        RECT 892.800 815.400 894.600 819.300 ;
        RECT 910.800 815.400 912.600 819.300 ;
        RECT 19.800 743.700 21.600 748.800 ;
        RECT 38.400 743.700 40.200 748.800 ;
        RECT 67.800 743.700 69.600 753.600 ;
        RECT 85.800 743.700 87.600 747.600 ;
        RECT 106.800 743.700 108.600 753.600 ;
        RECT 124.800 743.700 126.600 747.600 ;
        RECT 145.800 743.700 147.600 753.600 ;
        RECT 163.800 743.700 165.600 748.800 ;
        RECT 181.800 743.700 183.600 747.600 ;
        RECT 187.800 743.700 189.600 747.600 ;
        RECT 200.700 743.700 202.500 750.600 ;
        RECT 209.700 743.700 211.500 750.600 ;
        RECT 232.500 743.700 234.300 750.600 ;
        RECT 241.500 743.700 243.300 750.600 ;
        RECT 262.500 743.700 264.300 750.600 ;
        RECT 280.500 743.700 282.300 750.600 ;
        RECT 293.400 744.600 295.200 747.600 ;
        RECT 293.400 743.700 294.600 744.600 ;
        RECT 299.400 743.700 301.200 747.600 ;
        RECT 317.700 743.700 319.500 750.600 ;
        RECT 338.400 743.700 340.200 747.600 ;
        RECT 361.800 743.700 363.600 747.600 ;
        RECT 382.800 743.700 384.600 749.100 ;
        RECT 400.800 743.700 402.600 747.600 ;
        RECT 406.800 743.700 408.600 747.600 ;
        RECT 426.300 743.700 428.100 750.600 ;
        RECT 451.500 743.700 453.300 750.600 ;
        RECT 467.400 743.700 469.200 748.800 ;
        RECT 490.500 743.700 492.300 750.600 ;
        RECT 499.500 743.700 501.300 750.600 ;
        RECT 520.800 743.700 522.600 748.800 ;
        RECT 544.500 743.700 546.300 750.600 ;
        RECT 562.500 743.700 564.300 750.600 ;
        RECT 571.500 743.700 573.300 750.600 ;
        RECT 588.300 743.700 590.100 750.600 ;
        RECT 605.700 743.700 607.500 750.600 ;
        RECT 614.700 743.700 616.500 750.600 ;
        RECT 632.700 743.700 634.500 750.600 ;
        RECT 641.700 743.700 643.500 750.600 ;
        RECT 656.700 743.700 658.500 750.600 ;
        RECT 681.900 743.700 683.700 750.600 ;
        RECT 704.400 743.700 706.200 748.800 ;
        RECT 725.400 743.700 727.200 748.800 ;
        RECT 746.700 743.700 748.500 750.600 ;
        RECT 772.800 743.700 774.600 748.800 ;
        RECT 789.000 743.700 790.800 750.600 ;
        RECT 796.500 743.700 798.300 747.600 ;
        RECT 814.800 743.700 816.600 747.600 ;
        RECT 828.000 743.700 829.800 750.600 ;
        RECT 835.500 743.700 837.300 747.600 ;
        RECT 852.000 743.700 853.800 750.600 ;
        RECT 859.500 743.700 861.300 747.600 ;
        RECT 883.800 743.700 885.600 748.800 ;
        RECT 899.400 743.700 901.200 748.800 ;
        RECT 921.450 743.700 930.450 819.300 ;
        RECT 0.600 741.300 930.450 743.700 ;
        RECT 19.500 734.400 21.300 741.300 ;
        RECT 33.000 734.400 34.800 741.300 ;
        RECT 40.500 737.400 42.300 741.300 ;
        RECT 59.400 736.200 61.200 741.300 ;
        RECT 80.400 731.400 82.200 741.300 ;
        RECT 112.800 731.400 114.600 741.300 ;
        RECT 136.800 731.400 138.600 741.300 ;
        RECT 147.000 734.400 148.800 741.300 ;
        RECT 154.500 737.400 156.300 741.300 ;
        RECT 170.400 737.400 172.200 741.300 ;
        RECT 193.500 734.400 195.300 741.300 ;
        RECT 213.300 734.400 215.100 741.300 ;
        RECT 230.400 734.400 232.200 741.300 ;
        RECT 245.700 734.400 247.500 741.300 ;
        RECT 273.300 734.400 275.100 741.300 ;
        RECT 290.700 734.400 292.500 741.300 ;
        RECT 313.800 737.400 315.600 741.300 ;
        RECT 334.500 734.400 336.300 741.300 ;
        RECT 355.800 736.200 357.600 741.300 ;
        RECT 374.400 735.300 376.200 741.300 ;
        RECT 383.100 735.300 384.900 741.300 ;
        RECT 401.700 734.400 403.500 741.300 ;
        RECT 433.800 731.400 435.600 741.300 ;
        RECT 446.400 731.400 448.200 741.300 ;
        RECT 470.700 734.400 472.500 741.300 ;
        RECT 496.800 737.400 498.600 741.300 ;
        RECT 512.400 736.200 514.200 741.300 ;
        RECT 530.700 734.400 532.500 741.300 ;
        RECT 559.500 734.400 561.300 741.300 ;
        RECT 572.400 736.200 574.200 741.300 ;
        RECT 601.800 736.200 603.600 741.300 ;
        RECT 618.000 734.400 619.800 741.300 ;
        RECT 625.500 737.400 627.300 741.300 ;
        RECT 641.700 734.400 643.500 741.300 ;
        RECT 666.300 734.400 668.100 741.300 ;
        RECT 686.400 736.200 688.200 741.300 ;
        RECT 715.800 735.900 717.600 741.300 ;
        RECT 731.400 737.400 733.200 741.300 ;
        RECT 752.400 736.200 754.200 741.300 ;
        RECT 781.800 736.200 783.600 741.300 ;
        RECT 798.000 734.400 799.800 741.300 ;
        RECT 805.500 737.400 807.300 741.300 ;
        RECT 824.400 736.200 826.200 741.300 ;
        RECT 845.400 736.200 847.200 741.300 ;
        RECT 869.400 736.200 871.200 741.300 ;
        RECT 893.400 735.300 895.200 741.300 ;
        RECT 902.400 735.300 904.200 741.300 ;
        RECT 16.500 665.700 18.300 672.600 ;
        RECT 29.400 665.700 31.200 675.600 ;
        RECT 56.700 665.700 58.500 669.600 ;
        RECT 64.200 665.700 66.000 672.600 ;
        RECT 77.400 665.700 79.200 675.600 ;
        RECT 102.000 665.700 103.800 672.600 ;
        RECT 109.500 665.700 111.300 669.600 ;
        RECT 128.400 665.700 130.200 671.700 ;
        RECT 137.400 665.700 139.200 671.700 ;
        RECT 157.800 665.700 159.600 669.600 ;
        RECT 163.800 665.700 165.600 669.600 ;
        RECT 187.800 665.700 189.600 671.100 ;
        RECT 203.700 665.700 205.500 672.600 ;
        RECT 232.800 665.700 234.600 675.600 ;
        RECT 248.700 665.700 250.500 669.600 ;
        RECT 256.200 665.700 258.000 672.600 ;
        RECT 274.800 665.700 276.600 670.800 ;
        RECT 298.500 665.700 300.300 672.600 ;
        RECT 319.800 665.700 321.600 670.800 ;
        RECT 340.800 665.700 342.600 669.600 ;
        RECT 358.800 665.700 360.600 669.600 ;
        RECT 376.800 665.700 378.600 671.700 ;
        RECT 385.800 665.700 387.600 671.700 ;
        RECT 406.800 665.700 408.600 669.600 ;
        RECT 422.400 665.700 424.200 672.600 ;
        RECT 440.400 665.700 442.200 670.800 ;
        RECT 464.400 665.700 466.200 669.600 ;
        RECT 485.400 665.700 487.200 669.600 ;
        RECT 506.400 665.700 508.200 671.700 ;
        RECT 515.400 665.700 517.200 671.700 ;
        RECT 536.400 665.700 538.200 669.600 ;
        RECT 554.700 665.700 556.500 672.600 ;
        RECT 577.800 665.700 579.600 669.600 ;
        RECT 583.800 665.700 585.600 669.600 ;
        RECT 599.400 665.700 601.200 669.600 ;
        RECT 617.700 665.700 619.500 672.600 ;
        RECT 635.400 665.700 637.200 669.600 ;
        RECT 655.800 665.700 657.600 669.600 ;
        RECT 673.800 665.700 675.600 670.800 ;
        RECT 692.400 665.700 694.200 670.800 ;
        RECT 716.400 665.700 718.200 671.700 ;
        RECT 725.400 665.700 727.200 671.700 ;
        RECT 741.000 665.700 742.800 672.600 ;
        RECT 748.500 665.700 750.300 669.600 ;
        RECT 767.400 665.700 769.200 670.800 ;
        RECT 796.800 665.700 798.600 670.800 ;
        RECT 812.400 665.700 814.200 670.800 ;
        RECT 833.400 666.600 835.200 669.600 ;
        RECT 833.400 665.700 834.600 666.600 ;
        RECT 839.400 665.700 841.200 669.600 ;
        RECT 862.800 665.700 864.600 671.700 ;
        RECT 871.800 665.700 873.600 671.700 ;
        RECT 886.800 665.700 888.600 669.600 ;
        RECT 892.800 665.700 894.600 669.600 ;
        RECT 906.000 665.700 907.800 672.600 ;
        RECT 913.500 665.700 915.300 669.600 ;
        RECT 921.450 665.700 930.450 741.300 ;
        RECT 0.600 663.300 930.450 665.700 ;
        RECT 13.800 659.400 15.600 663.300 ;
        RECT 19.800 659.400 21.600 663.300 ;
        RECT 37.800 658.200 39.600 663.300 ;
        RECT 54.000 656.400 55.800 663.300 ;
        RECT 61.500 659.400 63.300 663.300 ;
        RECT 77.400 658.200 79.200 663.300 ;
        RECT 98.400 662.400 99.600 663.300 ;
        RECT 98.400 659.400 100.200 662.400 ;
        RECT 104.400 659.400 106.200 663.300 ;
        RECT 125.400 657.300 127.200 663.300 ;
        RECT 134.100 657.300 135.900 663.300 ;
        RECT 152.400 658.200 154.200 663.300 ;
        RECT 173.700 656.400 175.500 663.300 ;
        RECT 202.500 656.400 204.300 663.300 ;
        RECT 221.100 657.300 222.900 663.300 ;
        RECT 229.800 657.300 231.600 663.300 ;
        RECT 253.500 656.400 255.300 663.300 ;
        RECT 274.800 657.900 276.600 663.300 ;
        RECT 297.300 656.400 299.100 663.300 ;
        RECT 322.500 656.400 324.300 663.300 ;
        RECT 340.800 659.400 342.600 663.300 ;
        RECT 361.800 659.400 363.600 663.300 ;
        RECT 382.800 657.300 384.600 663.300 ;
        RECT 391.800 657.300 393.600 663.300 ;
        RECT 410.400 658.200 412.200 663.300 ;
        RECT 425.850 659.400 427.650 663.300 ;
        RECT 434.850 659.400 436.650 663.300 ;
        RECT 441.750 659.400 443.550 663.300 ;
        RECT 451.050 659.400 452.850 663.300 ;
        RECT 461.850 659.400 463.650 663.300 ;
        RECT 470.850 659.400 472.650 663.300 ;
        RECT 477.750 659.400 479.550 663.300 ;
        RECT 487.050 659.400 488.850 663.300 ;
        RECT 508.800 658.200 510.600 663.300 ;
        RECT 527.400 658.200 529.200 663.300 ;
        RECT 553.800 659.400 555.600 663.300 ;
        RECT 560.850 659.400 562.650 663.300 ;
        RECT 569.850 659.400 571.650 663.300 ;
        RECT 576.750 659.400 578.550 663.300 ;
        RECT 586.050 659.400 587.850 663.300 ;
        RECT 610.800 658.200 612.600 663.300 ;
        RECT 623.400 659.400 625.200 663.300 ;
        RECT 641.400 657.300 643.200 663.300 ;
        RECT 650.100 657.300 651.900 663.300 ;
        RECT 671.400 658.200 673.200 663.300 ;
        RECT 695.700 659.400 697.500 663.300 ;
        RECT 703.200 656.400 705.000 663.300 ;
        RECT 719.700 659.400 721.500 663.300 ;
        RECT 727.200 656.400 729.000 663.300 ;
        RECT 737.400 659.400 739.200 663.300 ;
        RECT 760.800 658.200 762.600 663.300 ;
        RECT 781.800 659.400 783.600 663.300 ;
        RECT 799.800 659.400 801.600 663.300 ;
        RECT 815.400 658.200 817.200 663.300 ;
        RECT 836.700 656.400 838.500 663.300 ;
        RECT 845.700 656.400 847.500 663.300 ;
        RECT 863.400 658.200 865.200 663.300 ;
        RECT 892.500 656.400 894.300 663.300 ;
        RECT 902.400 659.400 904.200 663.300 ;
        RECT 14.700 587.700 16.500 591.600 ;
        RECT 22.200 587.700 24.000 594.600 ;
        RECT 35.400 587.700 37.200 597.600 ;
        RECT 56.400 587.700 58.200 591.600 ;
        RECT 62.400 587.700 64.200 591.600 ;
        RECT 85.800 587.700 87.600 592.800 ;
        RECT 98.400 587.700 100.200 591.600 ;
        RECT 104.400 587.700 106.200 591.600 ;
        RECT 119.400 587.700 121.200 593.700 ;
        RECT 128.100 587.700 129.900 593.700 ;
        RECT 146.400 587.700 148.200 593.700 ;
        RECT 155.400 587.700 157.200 593.700 ;
        RECT 173.400 587.700 175.200 597.600 ;
        RECT 205.500 587.700 207.300 594.600 ;
        RECT 225.300 587.700 227.100 594.600 ;
        RECT 242.400 587.700 244.200 591.600 ;
        RECT 271.800 587.700 273.600 597.600 ;
        RECT 284.400 587.700 286.200 591.600 ;
        RECT 302.700 587.700 304.500 594.600 ;
        RECT 323.400 587.700 325.200 594.600 ;
        RECT 338.700 587.700 340.500 594.600 ;
        RECT 347.700 587.700 349.500 594.600 ;
        RECT 365.700 587.700 367.500 594.600 ;
        RECT 389.400 587.700 391.200 591.600 ;
        RECT 412.500 587.700 414.300 594.600 ;
        RECT 425.400 587.700 427.200 591.600 ;
        RECT 445.800 587.700 447.600 594.600 ;
        RECT 451.800 587.700 453.600 594.600 ;
        RECT 458.850 587.700 460.650 591.600 ;
        RECT 467.850 587.700 469.650 591.600 ;
        RECT 474.750 587.700 476.550 591.600 ;
        RECT 484.050 587.700 485.850 591.600 ;
        RECT 500.700 587.700 502.500 594.600 ;
        RECT 515.850 587.700 517.650 591.600 ;
        RECT 524.850 587.700 526.650 591.600 ;
        RECT 531.750 587.700 533.550 591.600 ;
        RECT 541.050 587.700 542.850 591.600 ;
        RECT 557.700 587.700 559.500 594.600 ;
        RECT 586.800 587.700 588.600 592.800 ;
        RECT 602.700 587.700 604.500 594.600 ;
        RECT 628.800 587.700 630.600 592.800 ;
        RECT 646.800 587.700 648.600 591.600 ;
        RECT 667.800 587.700 669.600 592.800 ;
        RECT 683.700 587.700 685.500 594.600 ;
        RECT 701.400 587.700 703.200 591.600 ;
        RECT 707.400 587.700 709.200 591.600 ;
        RECT 730.500 587.700 732.300 594.600 ;
        RECT 743.400 587.700 745.200 593.700 ;
        RECT 752.400 587.700 754.200 593.700 ;
        RECT 770.400 587.700 772.200 591.600 ;
        RECT 789.000 587.700 790.800 594.600 ;
        RECT 796.500 587.700 798.300 591.600 ;
        RECT 815.400 587.700 817.200 593.700 ;
        RECT 824.400 587.700 826.200 593.700 ;
        RECT 850.500 587.700 852.300 594.600 ;
        RECT 863.700 587.700 865.500 594.600 ;
        RECT 892.800 587.700 894.600 597.600 ;
        RECT 905.400 587.700 907.200 597.600 ;
        RECT 921.450 587.700 930.450 663.300 ;
        RECT 0.600 585.300 930.450 587.700 ;
        RECT 16.500 578.400 18.300 585.300 ;
        RECT 25.500 578.400 27.300 585.300 ;
        RECT 42.300 578.400 44.100 585.300 ;
        RECT 59.700 578.400 61.500 585.300 ;
        RECT 88.500 578.400 90.300 585.300 ;
        RECT 101.700 578.400 103.500 585.300 ;
        RECT 119.700 578.400 121.500 585.300 ;
        RECT 140.400 575.400 142.200 585.300 ;
        RECT 162.000 578.400 163.800 585.300 ;
        RECT 169.500 581.400 171.300 585.300 ;
        RECT 193.800 580.200 195.600 585.300 ;
        RECT 209.400 575.400 211.200 585.300 ;
        RECT 241.500 578.400 243.300 585.300 ;
        RECT 262.800 575.400 264.600 585.300 ;
        RECT 275.400 580.200 277.200 585.300 ;
        RECT 299.400 580.200 301.200 585.300 ;
        RECT 327.300 578.400 329.100 585.300 ;
        RECT 349.800 581.400 351.600 585.300 ;
        RECT 367.800 581.400 369.600 585.300 ;
        RECT 380.400 575.400 382.200 585.300 ;
        RECT 406.800 581.400 408.600 585.300 ;
        RECT 412.800 581.400 414.600 585.300 ;
        RECT 430.800 580.200 432.600 585.300 ;
        RECT 446.700 578.400 448.500 585.300 ;
        RECT 475.800 580.200 477.600 585.300 ;
        RECT 485.850 581.400 487.650 585.300 ;
        RECT 494.850 581.400 496.650 585.300 ;
        RECT 501.750 581.400 503.550 585.300 ;
        RECT 511.050 581.400 512.850 585.300 ;
        RECT 530.400 580.200 532.200 585.300 ;
        RECT 548.700 578.400 550.500 585.300 ;
        RECT 571.800 581.400 573.600 585.300 ;
        RECT 592.500 578.400 594.300 585.300 ;
        RECT 613.800 580.200 615.600 585.300 ;
        RECT 623.850 581.400 625.650 585.300 ;
        RECT 632.850 581.400 634.650 585.300 ;
        RECT 639.750 581.400 641.550 585.300 ;
        RECT 649.050 581.400 650.850 585.300 ;
        RECT 670.800 581.400 672.600 585.300 ;
        RECT 685.800 578.400 687.600 585.300 ;
        RECT 691.800 578.400 693.600 585.300 ;
        RECT 697.800 578.400 699.600 585.300 ;
        RECT 703.800 578.400 705.600 585.300 ;
        RECT 709.800 578.400 711.600 585.300 ;
        RECT 724.800 581.400 726.600 585.300 ;
        RECT 737.400 581.400 739.200 585.300 ;
        RECT 743.400 581.400 745.200 585.300 ;
        RECT 765.300 578.400 767.100 585.300 ;
        RECT 781.800 578.400 783.600 585.300 ;
        RECT 787.800 578.400 789.600 585.300 ;
        RECT 793.800 578.400 795.600 585.300 ;
        RECT 799.800 578.400 801.600 585.300 ;
        RECT 805.800 578.400 807.600 585.300 ;
        RECT 818.400 581.400 820.200 585.300 ;
        RECT 824.400 581.400 826.200 585.300 ;
        RECT 847.800 575.400 849.600 585.300 ;
        RECT 868.500 578.400 870.300 585.300 ;
        RECT 881.700 578.400 883.500 585.300 ;
        RECT 902.400 581.400 904.200 585.300 ;
        RECT 14.100 509.700 16.200 513.600 ;
        RECT 20.400 509.700 22.200 513.600 ;
        RECT 55.500 509.700 57.300 516.600 ;
        RECT 79.800 509.700 81.600 519.600 ;
        RECT 90.000 509.700 91.800 516.600 ;
        RECT 97.500 509.700 99.300 513.600 ;
        RECT 111.000 509.700 112.800 516.600 ;
        RECT 118.500 509.700 120.300 513.600 ;
        RECT 142.800 509.700 144.600 514.800 ;
        RECT 161.400 509.700 163.200 514.800 ;
        RECT 193.800 509.700 195.600 519.600 ;
        RECT 214.800 509.700 216.600 519.600 ;
        RECT 235.800 509.700 237.600 519.600 ;
        RECT 248.400 509.700 250.200 513.600 ;
        RECT 266.400 509.700 268.200 519.600 ;
        RECT 290.400 509.700 292.200 519.600 ;
        RECT 311.400 509.700 313.200 513.600 ;
        RECT 317.400 509.700 319.200 513.600 ;
        RECT 329.700 509.700 331.500 516.600 ;
        RECT 338.700 509.700 340.500 516.600 ;
        RECT 356.400 509.700 358.200 516.600 ;
        RECT 379.500 509.700 381.300 516.600 ;
        RECT 392.400 509.700 394.200 513.600 ;
        RECT 418.500 509.700 420.300 516.600 ;
        RECT 431.700 509.700 433.500 516.600 ;
        RECT 440.700 509.700 442.500 516.600 ;
        RECT 466.800 509.700 468.600 514.800 ;
        RECT 479.700 509.700 481.500 516.600 ;
        RECT 500.400 509.700 502.200 514.800 ;
        RECT 524.400 509.700 526.200 514.800 ;
        RECT 547.800 509.700 549.600 513.600 ;
        RECT 560.400 509.700 562.200 513.600 ;
        RECT 583.800 509.700 585.600 513.600 ;
        RECT 593.850 509.700 595.650 513.600 ;
        RECT 602.850 509.700 604.650 513.600 ;
        RECT 609.750 509.700 611.550 513.600 ;
        RECT 619.050 509.700 620.850 513.600 ;
        RECT 640.800 509.700 642.600 513.600 ;
        RECT 658.800 509.700 660.600 513.600 ;
        RECT 679.500 509.700 681.300 516.600 ;
        RECT 686.850 509.700 688.650 513.600 ;
        RECT 695.850 509.700 697.650 513.600 ;
        RECT 702.750 509.700 704.550 513.600 ;
        RECT 712.050 509.700 713.850 513.600 ;
        RECT 722.850 509.700 724.650 513.600 ;
        RECT 731.850 509.700 733.650 513.600 ;
        RECT 738.750 509.700 740.550 513.600 ;
        RECT 748.050 509.700 749.850 513.600 ;
        RECT 758.850 509.700 760.650 513.600 ;
        RECT 767.850 509.700 769.650 513.600 ;
        RECT 774.750 509.700 776.550 513.600 ;
        RECT 784.050 509.700 785.850 513.600 ;
        RECT 805.800 509.700 807.600 513.600 ;
        RECT 815.700 509.700 817.500 516.600 ;
        RECT 833.400 509.700 835.200 519.600 ;
        RECT 860.400 509.700 862.200 514.800 ;
        RECT 889.500 509.700 891.300 516.600 ;
        RECT 913.800 509.700 915.600 519.600 ;
        RECT 921.450 509.700 930.450 585.300 ;
        RECT 0.600 507.300 930.450 509.700 ;
        RECT 14.400 502.200 16.200 507.300 ;
        RECT 43.800 497.400 45.600 507.300 ;
        RECT 54.000 500.400 55.800 507.300 ;
        RECT 61.500 503.400 63.300 507.300 ;
        RECT 77.400 497.400 79.200 507.300 ;
        RECT 109.800 497.400 111.600 507.300 ;
        RECT 125.400 502.200 127.200 507.300 ;
        RECT 148.500 500.400 150.300 507.300 ;
        RECT 157.500 500.400 159.300 507.300 ;
        RECT 174.300 500.400 176.100 507.300 ;
        RECT 191.700 500.400 193.500 507.300 ;
        RECT 223.800 497.400 225.600 507.300 ;
        RECT 238.800 503.400 240.600 507.300 ;
        RECT 259.800 502.200 261.600 507.300 ;
        RECT 283.800 502.200 285.600 507.300 ;
        RECT 303.300 500.400 305.100 507.300 ;
        RECT 317.700 500.400 319.500 507.300 ;
        RECT 338.400 506.400 339.600 507.300 ;
        RECT 338.400 503.400 340.200 506.400 ;
        RECT 344.400 503.400 346.200 507.300 ;
        RECT 362.700 500.400 364.500 507.300 ;
        RECT 391.500 500.400 393.300 507.300 ;
        RECT 404.400 503.400 406.200 507.300 ;
        RECT 422.700 500.400 424.500 507.300 ;
        RECT 443.700 500.400 445.500 507.300 ;
        RECT 464.400 502.200 466.200 507.300 ;
        RECT 488.700 503.400 490.500 507.300 ;
        RECT 496.200 500.400 498.000 507.300 ;
        RECT 510.000 500.400 511.800 507.300 ;
        RECT 517.500 503.400 519.300 507.300 ;
        RECT 533.400 503.400 535.200 507.300 ;
        RECT 551.400 497.400 553.200 507.300 ;
        RECT 575.700 503.400 577.500 507.300 ;
        RECT 583.200 500.400 585.000 507.300 ;
        RECT 596.400 497.400 598.200 507.300 ;
        RECT 620.400 497.400 622.200 507.300 ;
        RECT 647.400 503.400 649.200 507.300 ;
        RECT 673.500 500.400 675.300 507.300 ;
        RECT 689.400 502.200 691.200 507.300 ;
        RECT 713.400 502.200 715.200 507.300 ;
        RECT 734.700 500.400 736.500 507.300 ;
        RECT 755.400 503.400 757.200 507.300 ;
        RECT 761.400 503.400 763.200 507.300 ;
        RECT 784.800 502.200 786.600 507.300 ;
        RECT 800.400 503.400 802.200 507.300 ;
        RECT 821.400 502.200 823.200 507.300 ;
        RECT 839.700 500.400 841.500 507.300 ;
        RECT 860.400 503.400 862.200 507.300 ;
        RECT 866.400 503.400 868.200 507.300 ;
        RECT 881.400 497.400 883.200 507.300 ;
        RECT 910.500 500.400 912.300 507.300 ;
        RECT 14.400 431.700 16.200 436.800 ;
        RECT 46.800 431.700 48.600 441.600 ;
        RECT 60.000 431.700 61.800 438.600 ;
        RECT 67.500 431.700 69.300 435.600 ;
        RECT 84.000 431.700 85.800 438.600 ;
        RECT 91.500 431.700 93.300 435.600 ;
        RECT 112.800 431.700 114.600 436.800 ;
        RECT 136.800 431.700 138.600 436.800 ;
        RECT 152.400 431.700 154.200 436.800 ;
        RECT 171.000 431.700 172.800 438.600 ;
        RECT 178.500 431.700 180.300 435.600 ;
        RECT 194.400 431.700 196.200 435.600 ;
        RECT 223.800 431.700 225.600 441.600 ;
        RECT 239.700 431.700 241.500 435.600 ;
        RECT 247.200 431.700 249.000 438.600 ;
        RECT 257.400 431.700 259.200 441.600 ;
        RECT 284.400 431.700 286.200 436.800 ;
        RECT 305.400 431.700 307.200 435.600 ;
        RECT 311.400 431.700 313.200 435.600 ;
        RECT 334.500 431.700 336.300 438.600 ;
        RECT 345.000 431.700 346.800 438.600 ;
        RECT 352.500 431.700 354.300 435.600 ;
        RECT 373.800 431.700 375.600 435.600 ;
        RECT 390.000 431.700 391.800 438.600 ;
        RECT 397.500 431.700 399.300 435.600 ;
        RECT 416.400 431.700 418.200 436.800 ;
        RECT 434.700 431.700 436.500 438.600 ;
        RECT 443.700 431.700 445.500 438.600 ;
        RECT 460.800 431.700 462.600 435.600 ;
        RECT 466.800 431.700 468.600 435.600 ;
        RECT 479.400 431.700 481.200 441.600 ;
        RECT 503.400 431.700 505.200 435.600 ;
        RECT 509.400 431.700 511.200 435.600 ;
        RECT 524.400 431.700 526.200 441.600 ;
        RECT 548.400 431.700 550.200 436.800 ;
        RECT 563.850 431.700 565.650 435.600 ;
        RECT 572.850 431.700 574.650 435.600 ;
        RECT 579.750 431.700 581.550 435.600 ;
        RECT 589.050 431.700 590.850 435.600 ;
        RECT 605.700 431.700 607.500 438.600 ;
        RECT 634.800 431.700 636.600 436.800 ;
        RECT 653.400 431.700 655.200 436.800 ;
        RECT 668.850 431.700 670.650 435.600 ;
        RECT 677.850 431.700 679.650 435.600 ;
        RECT 684.750 431.700 686.550 435.600 ;
        RECT 694.050 431.700 695.850 435.600 ;
        RECT 704.850 431.700 706.650 435.600 ;
        RECT 713.850 431.700 715.650 435.600 ;
        RECT 720.750 431.700 722.550 435.600 ;
        RECT 730.050 431.700 731.850 435.600 ;
        RECT 748.800 431.700 750.600 438.600 ;
        RECT 754.800 431.700 756.600 438.600 ;
        RECT 760.800 431.700 762.600 438.600 ;
        RECT 766.800 431.700 768.600 438.600 ;
        RECT 772.800 431.700 774.600 438.600 ;
        RECT 788.400 431.700 790.200 435.600 ;
        RECT 806.400 431.700 808.200 435.600 ;
        RECT 829.800 431.700 831.600 435.600 ;
        RECT 835.800 432.600 837.600 435.600 ;
        RECT 836.400 431.700 837.600 432.600 ;
        RECT 850.800 431.700 852.600 435.600 ;
        RECT 856.800 431.700 858.600 435.600 ;
        RECT 871.800 431.700 873.600 435.600 ;
        RECT 889.500 431.700 891.300 438.600 ;
        RECT 913.800 431.700 915.600 441.600 ;
        RECT 921.450 431.700 930.450 507.300 ;
        RECT 0.600 429.300 930.450 431.700 ;
        RECT 22.800 419.400 24.600 429.300 ;
        RECT 35.400 419.400 37.200 429.300 ;
        RECT 67.800 419.400 69.600 429.300 ;
        RECT 81.000 422.400 82.800 429.300 ;
        RECT 88.500 425.400 90.300 429.300 ;
        RECT 112.800 424.200 114.600 429.300 ;
        RECT 128.700 425.400 130.500 429.300 ;
        RECT 136.200 422.400 138.000 429.300 ;
        RECT 149.400 425.400 151.200 429.300 ;
        RECT 167.400 419.400 169.200 429.300 ;
        RECT 191.400 419.400 193.200 429.300 ;
        RECT 212.700 422.400 214.500 429.300 ;
        RECT 221.700 422.400 223.500 429.300 ;
        RECT 239.400 425.400 241.200 429.300 ;
        RECT 268.800 419.400 270.600 429.300 ;
        RECT 286.800 425.400 288.600 429.300 ;
        RECT 299.700 422.400 301.500 429.300 ;
        RECT 320.400 425.400 322.200 429.300 ;
        RECT 326.400 425.400 328.200 429.300 ;
        RECT 346.500 422.400 348.300 429.300 ;
        RECT 360.900 422.400 362.700 429.300 ;
        RECT 380.400 425.400 382.200 429.300 ;
        RECT 406.800 424.200 408.600 429.300 ;
        RECT 422.700 422.400 424.500 429.300 ;
        RECT 443.400 419.400 445.200 429.300 ;
        RECT 472.800 423.300 474.600 429.300 ;
        RECT 481.800 423.300 483.600 429.300 ;
        RECT 501.900 422.400 503.700 429.300 ;
        RECT 521.400 424.200 523.200 429.300 ;
        RECT 545.400 424.200 547.200 429.300 ;
        RECT 571.800 425.400 573.600 429.300 ;
        RECT 592.800 424.200 594.600 429.300 ;
        RECT 613.800 425.400 615.600 429.300 ;
        RECT 632.400 424.200 634.200 429.300 ;
        RECT 661.500 422.400 663.300 429.300 ;
        RECT 679.800 424.200 681.600 429.300 ;
        RECT 695.400 425.400 697.200 429.300 ;
        RECT 701.400 425.400 703.200 429.300 ;
        RECT 715.800 425.400 717.600 429.300 ;
        RECT 721.800 425.400 723.600 429.300 ;
        RECT 729.150 425.400 730.950 429.300 ;
        RECT 738.450 425.400 740.250 429.300 ;
        RECT 745.350 425.400 747.150 429.300 ;
        RECT 754.350 425.400 756.150 429.300 ;
        RECT 773.400 424.200 775.200 429.300 ;
        RECT 791.700 422.400 793.500 429.300 ;
        RECT 823.800 423.900 825.600 429.300 ;
        RECT 841.800 425.400 843.600 429.300 ;
        RECT 854.700 422.400 856.500 429.300 ;
        RECT 863.700 422.400 865.500 429.300 ;
        RECT 878.400 425.400 880.200 429.300 ;
        RECT 884.400 425.400 886.200 429.300 ;
        RECT 899.400 425.400 901.200 429.300 ;
        RECT 15.300 353.700 17.100 360.600 ;
        RECT 32.700 353.700 34.500 360.600 ;
        RECT 54.000 353.700 55.800 360.600 ;
        RECT 61.500 353.700 63.300 357.600 ;
        RECT 79.800 353.700 81.600 357.600 ;
        RECT 95.400 353.700 97.200 358.800 ;
        RECT 118.800 353.700 120.600 357.600 ;
        RECT 124.800 353.700 126.600 357.600 ;
        RECT 145.500 353.700 147.300 360.600 ;
        RECT 163.500 353.700 165.300 360.600 ;
        RECT 176.400 353.700 178.200 357.600 ;
        RECT 197.400 353.700 199.200 358.800 ;
        RECT 229.800 353.700 231.600 363.600 ;
        RECT 247.800 353.700 249.600 358.800 ;
        RECT 271.800 353.700 273.600 358.800 ;
        RECT 287.700 353.700 289.500 360.600 ;
        RECT 315.300 353.700 317.100 360.600 ;
        RECT 337.800 353.700 339.600 357.600 ;
        RECT 355.800 353.700 357.600 357.600 ;
        RECT 374.700 353.700 376.500 357.600 ;
        RECT 382.200 353.700 384.000 360.600 ;
        RECT 400.800 353.700 402.600 358.800 ;
        RECT 419.100 353.700 421.200 357.600 ;
        RECT 425.400 353.700 427.200 357.600 ;
        RECT 453.000 353.700 454.800 360.600 ;
        RECT 460.500 353.700 462.300 357.600 ;
        RECT 473.400 353.700 475.200 357.600 ;
        RECT 494.400 353.700 496.200 358.800 ;
        RECT 515.400 353.700 517.200 357.600 ;
        RECT 536.400 353.700 538.200 358.800 ;
        RECT 565.800 353.700 567.600 358.800 ;
        RECT 586.800 353.700 588.600 357.600 ;
        RECT 600.000 353.700 601.800 360.600 ;
        RECT 607.500 353.700 609.300 357.600 ;
        RECT 626.400 353.700 628.200 358.800 ;
        RECT 649.800 353.700 651.600 357.600 ;
        RECT 655.800 353.700 657.600 357.600 ;
        RECT 668.700 353.700 670.500 360.600 ;
        RECT 694.800 353.700 696.600 358.800 ;
        RECT 712.800 353.700 714.600 357.600 ;
        RECT 718.800 353.700 720.600 357.600 ;
        RECT 736.500 353.700 738.300 360.600 ;
        RECT 760.800 353.700 762.600 363.600 ;
        RECT 773.400 353.700 775.200 357.600 ;
        RECT 799.800 353.700 801.600 358.800 ;
        RECT 815.400 354.600 817.200 357.600 ;
        RECT 815.400 353.700 816.600 354.600 ;
        RECT 821.400 353.700 823.200 357.600 ;
        RECT 844.800 353.700 846.600 358.800 ;
        RECT 865.800 353.700 867.600 358.800 ;
        RECT 883.800 353.700 885.600 357.600 ;
        RECT 889.800 353.700 891.600 357.600 ;
        RECT 902.700 353.700 904.500 360.600 ;
        RECT 921.450 353.700 930.450 429.300 ;
        RECT 0.600 351.300 930.450 353.700 ;
        RECT 19.800 346.200 21.600 351.300 ;
        RECT 46.800 341.400 48.600 351.300 ;
        RECT 67.800 346.200 69.600 351.300 ;
        RECT 83.400 341.400 85.200 351.300 ;
        RECT 110.400 346.200 112.200 351.300 ;
        RECT 136.800 347.400 138.600 351.300 ;
        RECT 160.800 341.400 162.600 351.300 ;
        RECT 173.700 344.400 175.500 351.300 ;
        RECT 182.700 344.400 184.500 351.300 ;
        RECT 197.700 344.400 199.500 351.300 ;
        RECT 206.700 344.400 208.500 351.300 ;
        RECT 221.700 344.400 223.500 351.300 ;
        RECT 244.800 347.400 246.600 351.300 ;
        RECT 250.800 347.400 252.600 351.300 ;
        RECT 265.500 344.400 267.300 351.300 ;
        RECT 274.500 344.400 276.300 351.300 ;
        RECT 291.300 344.400 293.100 351.300 ;
        RECT 316.500 344.400 318.300 351.300 ;
        RECT 331.800 347.400 333.600 351.300 ;
        RECT 337.800 347.400 339.600 351.300 ;
        RECT 350.400 344.400 352.200 351.300 ;
        RECT 375.300 344.400 377.100 351.300 ;
        RECT 397.800 347.400 399.600 351.300 ;
        RECT 418.800 347.400 420.600 351.300 ;
        RECT 434.400 347.400 436.200 351.300 ;
        RECT 454.800 347.400 456.600 351.300 ;
        RECT 460.800 347.400 462.600 351.300 ;
        RECT 473.400 346.200 475.200 351.300 ;
        RECT 499.800 347.400 501.600 351.300 ;
        RECT 520.800 347.400 522.600 351.300 ;
        RECT 541.800 347.400 543.600 351.300 ;
        RECT 548.850 347.400 550.650 351.300 ;
        RECT 557.850 347.400 559.650 351.300 ;
        RECT 564.750 347.400 566.550 351.300 ;
        RECT 574.050 347.400 575.850 351.300 ;
        RECT 587.700 344.400 589.500 351.300 ;
        RECT 596.700 344.400 598.500 351.300 ;
        RECT 619.800 346.200 621.600 351.300 ;
        RECT 637.800 347.400 639.600 351.300 ;
        RECT 643.800 347.400 645.600 351.300 ;
        RECT 658.500 344.400 660.300 351.300 ;
        RECT 667.500 344.400 669.300 351.300 ;
        RECT 674.850 347.400 676.650 351.300 ;
        RECT 683.850 347.400 685.650 351.300 ;
        RECT 690.750 347.400 692.550 351.300 ;
        RECT 700.050 347.400 701.850 351.300 ;
        RECT 716.400 347.400 718.200 351.300 ;
        RECT 722.400 347.400 724.200 351.300 ;
        RECT 737.400 347.400 739.200 351.300 ;
        RECT 752.400 347.400 754.200 351.300 ;
        RECT 772.800 347.400 774.600 351.300 ;
        RECT 778.800 347.400 780.600 351.300 ;
        RECT 791.700 344.400 793.500 351.300 ;
        RECT 812.400 341.400 814.200 351.300 ;
        RECT 836.400 346.200 838.200 351.300 ;
        RECT 862.800 347.400 864.600 351.300 ;
        RECT 875.400 347.400 877.200 351.300 ;
        RECT 894.900 344.400 896.700 351.300 ;
        RECT 22.800 275.700 24.600 285.600 ;
        RECT 35.700 275.700 37.500 279.600 ;
        RECT 43.200 275.700 45.000 282.600 ;
        RECT 56.700 275.700 58.500 279.600 ;
        RECT 64.200 275.700 66.000 282.600 ;
        RECT 74.400 275.700 76.200 285.600 ;
        RECT 98.400 275.700 100.200 285.600 ;
        RECT 127.800 275.700 129.600 280.800 ;
        RECT 146.700 275.700 148.500 279.600 ;
        RECT 154.200 275.700 156.000 282.600 ;
        RECT 172.800 275.700 174.600 280.800 ;
        RECT 196.800 275.700 198.600 280.800 ;
        RECT 217.500 275.700 219.300 282.600 ;
        RECT 230.700 275.700 232.500 282.600 ;
        RECT 248.700 275.700 250.500 282.600 ;
        RECT 269.400 275.700 271.200 280.800 ;
        RECT 290.700 275.700 292.500 282.600 ;
        RECT 318.300 275.700 320.100 282.600 ;
        RECT 335.700 275.700 337.500 282.600 ;
        RECT 367.800 275.700 369.600 285.600 ;
        RECT 380.700 275.700 382.500 282.600 ;
        RECT 406.500 275.700 408.300 282.600 ;
        RECT 427.800 275.700 429.600 280.800 ;
        RECT 445.800 275.700 447.600 279.600 ;
        RECT 461.400 275.700 463.200 280.800 ;
        RECT 482.700 275.700 484.500 282.600 ;
        RECT 511.500 275.700 513.300 282.600 ;
        RECT 529.500 275.700 531.300 282.600 ;
        RECT 538.500 275.700 540.300 282.600 ;
        RECT 556.800 275.700 558.600 279.600 ;
        RECT 574.800 275.700 576.600 280.800 ;
        RECT 598.500 275.700 600.300 282.600 ;
        RECT 614.700 275.700 616.500 279.600 ;
        RECT 622.200 275.700 624.000 282.600 ;
        RECT 640.800 275.700 642.600 280.800 ;
        RECT 659.400 275.700 661.200 280.800 ;
        RECT 680.700 275.700 682.500 282.600 ;
        RECT 706.800 275.700 708.600 279.600 ;
        RECT 719.700 275.700 721.500 282.600 ;
        RECT 740.400 275.700 742.200 282.600 ;
        RECT 746.400 275.700 748.200 282.600 ;
        RECT 766.800 275.700 768.600 279.600 ;
        RECT 776.400 275.700 778.200 279.600 ;
        RECT 795.000 275.700 796.800 282.600 ;
        RECT 802.500 275.700 804.300 279.600 ;
        RECT 818.700 275.700 820.500 282.600 ;
        RECT 827.700 275.700 829.500 282.600 ;
        RECT 848.400 275.700 850.200 280.800 ;
        RECT 869.700 275.700 871.500 282.600 ;
        RECT 893.400 275.700 895.200 280.800 ;
        RECT 921.450 275.700 930.450 351.300 ;
        RECT 0.600 273.300 930.450 275.700 ;
        RECT 19.800 268.200 21.600 273.300 ;
        RECT 40.800 268.200 42.600 273.300 ;
        RECT 67.800 263.400 69.600 273.300 ;
        RECT 85.800 269.400 87.600 273.300 ;
        RECT 100.500 266.400 102.300 273.300 ;
        RECT 109.500 266.400 111.300 273.300 ;
        RECT 119.700 266.400 121.500 273.300 ;
        RECT 151.800 263.400 153.600 273.300 ;
        RECT 161.400 269.400 163.200 273.300 ;
        RECT 190.800 263.400 192.600 273.300 ;
        RECT 208.800 269.400 210.600 273.300 ;
        RECT 232.800 263.400 234.600 273.300 ;
        RECT 256.800 263.400 258.600 273.300 ;
        RECT 274.500 266.400 276.300 273.300 ;
        RECT 283.500 266.400 285.300 273.300 ;
        RECT 304.800 268.200 306.600 273.300 ;
        RECT 323.400 268.200 325.200 273.300 ;
        RECT 341.700 266.400 343.500 273.300 ;
        RECT 361.800 269.400 363.600 273.300 ;
        RECT 367.800 269.400 369.600 273.300 ;
        RECT 380.700 266.400 382.500 273.300 ;
        RECT 405.300 266.400 407.100 273.300 ;
        RECT 426.900 266.400 428.700 273.300 ;
        RECT 448.800 269.400 450.600 273.300 ;
        RECT 461.400 269.400 463.200 273.300 ;
        RECT 467.400 269.400 469.200 273.300 ;
        RECT 489.300 266.400 491.100 273.300 ;
        RECT 506.400 272.400 507.600 273.300 ;
        RECT 506.400 269.400 508.200 272.400 ;
        RECT 512.400 269.400 514.200 273.300 ;
        RECT 527.700 266.400 529.500 273.300 ;
        RECT 548.400 272.400 549.600 273.300 ;
        RECT 548.400 269.400 550.200 272.400 ;
        RECT 554.400 269.400 556.200 273.300 ;
        RECT 572.700 266.400 574.500 273.300 ;
        RECT 590.400 269.400 592.200 273.300 ;
        RECT 608.400 268.200 610.200 273.300 ;
        RECT 626.400 272.400 627.600 273.300 ;
        RECT 626.400 269.400 628.200 272.400 ;
        RECT 632.400 269.400 634.200 273.300 ;
        RECT 650.700 266.400 652.500 273.300 ;
        RECT 670.800 269.400 672.600 273.300 ;
        RECT 676.800 269.400 678.600 273.300 ;
        RECT 693.900 266.400 695.700 273.300 ;
        RECT 713.400 268.200 715.200 273.300 ;
        RECT 728.850 269.400 730.650 273.300 ;
        RECT 737.850 269.400 739.650 273.300 ;
        RECT 744.750 269.400 746.550 273.300 ;
        RECT 754.050 269.400 755.850 273.300 ;
        RECT 778.500 266.400 780.300 273.300 ;
        RECT 790.800 269.400 792.600 273.300 ;
        RECT 796.800 269.400 798.600 273.300 ;
        RECT 809.400 269.400 811.200 273.300 ;
        RECT 826.800 269.400 828.600 273.300 ;
        RECT 832.800 269.400 834.600 273.300 ;
        RECT 838.200 269.400 840.000 273.300 ;
        RECT 850.500 266.400 852.300 273.300 ;
        RECT 873.000 269.400 874.800 273.300 ;
        RECT 880.500 269.400 882.300 273.300 ;
        RECT 899.100 266.400 900.900 273.300 ;
        RECT 22.800 197.700 24.600 207.600 ;
        RECT 33.000 197.700 34.800 204.600 ;
        RECT 40.500 197.700 42.300 201.600 ;
        RECT 64.500 197.700 66.300 204.600 ;
        RECT 77.700 197.700 79.500 204.600 ;
        RECT 103.800 197.700 105.600 202.800 ;
        RECT 119.400 197.700 121.200 201.600 ;
        RECT 125.400 197.700 127.200 201.600 ;
        RECT 143.400 197.700 145.200 202.800 ;
        RECT 167.700 197.700 169.500 201.600 ;
        RECT 175.200 197.700 177.000 204.600 ;
        RECT 185.400 197.700 187.200 207.600 ;
        RECT 217.500 197.700 219.300 204.600 ;
        RECT 238.800 197.700 240.600 202.800 ;
        RECT 259.800 197.700 261.600 201.600 ;
        RECT 275.400 197.700 277.200 202.800 ;
        RECT 307.800 197.700 309.600 207.600 ;
        RECT 320.400 197.700 322.200 202.800 ;
        RECT 338.400 197.700 340.200 201.600 ;
        RECT 356.700 197.700 358.500 204.600 ;
        RECT 381.300 197.700 383.100 204.600 ;
        RECT 395.700 197.700 397.500 204.600 ;
        RECT 424.800 197.700 426.600 202.800 ;
        RECT 445.800 197.700 447.600 202.800 ;
        RECT 461.400 197.700 463.200 202.800 ;
        RECT 483.900 197.700 485.700 204.600 ;
        RECT 503.400 197.700 505.200 201.600 ;
        RECT 509.400 197.700 511.200 201.600 ;
        RECT 532.800 197.700 534.600 202.800 ;
        RECT 548.700 197.700 550.500 204.600 ;
        RECT 569.400 197.700 571.200 201.600 ;
        RECT 590.400 197.700 592.200 202.800 ;
        RECT 611.400 198.600 613.200 201.600 ;
        RECT 611.400 197.700 612.600 198.600 ;
        RECT 617.400 197.700 619.200 201.600 ;
        RECT 643.800 197.700 645.600 207.600 ;
        RECT 657.000 197.700 658.800 204.600 ;
        RECT 664.500 197.700 666.300 201.600 ;
        RECT 680.400 197.700 682.200 202.800 ;
        RECT 704.400 197.700 706.200 202.800 ;
        RECT 733.800 197.700 735.600 202.800 ;
        RECT 751.800 197.700 753.600 201.600 ;
        RECT 757.800 197.700 759.600 201.600 ;
        RECT 775.500 197.700 777.300 204.600 ;
        RECT 793.800 197.700 795.600 201.600 ;
        RECT 811.800 197.700 813.600 202.800 ;
        RECT 820.200 197.700 822.000 201.600 ;
        RECT 832.500 197.700 834.300 204.600 ;
        RECT 855.000 197.700 856.800 201.600 ;
        RECT 862.500 197.700 864.300 201.600 ;
        RECT 881.100 197.700 882.900 204.600 ;
        RECT 904.800 197.700 906.600 201.600 ;
        RECT 921.450 197.700 930.450 273.300 ;
        RECT 0.600 195.300 930.450 197.700 ;
        RECT 19.800 190.200 21.600 195.300 ;
        RECT 40.500 188.400 42.300 195.300 ;
        RECT 64.800 185.400 66.600 195.300 ;
        RECT 74.400 191.400 76.200 195.300 ;
        RECT 92.400 185.400 94.200 195.300 ;
        RECT 124.800 185.400 126.600 195.300 ;
        RECT 140.400 190.200 142.200 195.300 ;
        RECT 164.700 191.400 166.500 195.300 ;
        RECT 172.200 188.400 174.000 195.300 ;
        RECT 185.400 185.400 187.200 195.300 ;
        RECT 217.500 188.400 219.300 195.300 ;
        RECT 231.900 188.400 233.700 195.300 ;
        RECT 254.700 191.400 256.500 195.300 ;
        RECT 262.200 188.400 264.000 195.300 ;
        RECT 277.800 191.400 279.600 195.300 ;
        RECT 292.800 191.400 294.600 195.300 ;
        RECT 298.800 191.400 300.600 195.300 ;
        RECT 311.400 190.200 313.200 195.300 ;
        RECT 332.400 190.200 334.200 195.300 ;
        RECT 364.800 185.400 366.600 195.300 ;
        RECT 380.400 190.200 382.200 195.300 ;
        RECT 401.400 191.400 403.200 195.300 ;
        RECT 407.400 191.400 409.200 195.300 ;
        RECT 422.700 191.400 424.500 195.300 ;
        RECT 430.200 188.400 432.000 195.300 ;
        RECT 443.400 191.400 445.200 195.300 ;
        RECT 458.400 185.400 460.200 195.300 ;
        RECT 482.400 185.400 484.200 195.300 ;
        RECT 509.700 191.400 511.500 195.300 ;
        RECT 517.200 188.400 519.000 195.300 ;
        RECT 533.400 190.200 535.200 195.300 ;
        RECT 551.400 191.400 553.200 195.300 ;
        RECT 569.400 185.400 571.200 195.300 ;
        RECT 591.000 188.400 592.800 195.300 ;
        RECT 598.500 191.400 600.300 195.300 ;
        RECT 614.400 185.400 616.200 195.300 ;
        RECT 643.500 188.400 645.300 195.300 ;
        RECT 664.500 188.400 666.300 195.300 ;
        RECT 677.400 191.400 679.200 195.300 ;
        RECT 697.800 191.400 699.600 195.300 ;
        RECT 707.850 191.400 709.650 195.300 ;
        RECT 716.850 191.400 718.650 195.300 ;
        RECT 723.750 191.400 725.550 195.300 ;
        RECT 733.050 191.400 734.850 195.300 ;
        RECT 751.800 188.400 753.600 195.300 ;
        RECT 757.800 188.400 759.600 195.300 ;
        RECT 763.800 188.400 765.600 195.300 ;
        RECT 769.800 188.400 771.600 195.300 ;
        RECT 775.800 188.400 777.600 195.300 ;
        RECT 789.000 188.400 790.800 195.300 ;
        RECT 796.500 191.400 798.300 195.300 ;
        RECT 812.400 191.400 814.200 195.300 ;
        RECT 830.400 188.400 832.200 195.300 ;
        RECT 841.200 191.400 843.000 195.300 ;
        RECT 853.500 188.400 855.300 195.300 ;
        RECT 876.000 191.400 877.800 195.300 ;
        RECT 883.500 191.400 885.300 195.300 ;
        RECT 902.100 188.400 903.900 195.300 ;
        RECT 14.700 119.700 16.500 123.600 ;
        RECT 22.200 119.700 24.000 126.600 ;
        RECT 32.400 119.700 34.200 129.600 ;
        RECT 57.000 119.700 58.800 126.600 ;
        RECT 64.500 119.700 66.300 123.600 ;
        RECT 77.400 119.700 79.200 129.600 ;
        RECT 109.500 119.700 111.300 126.600 ;
        RECT 125.700 119.700 127.500 123.600 ;
        RECT 133.200 119.700 135.000 126.600 ;
        RECT 157.800 119.700 159.600 129.600 ;
        RECT 173.400 119.700 175.200 124.800 ;
        RECT 194.400 119.700 196.200 129.600 ;
        RECT 229.800 119.700 231.600 129.600 ;
        RECT 247.800 119.700 249.600 123.600 ;
        RECT 263.400 119.700 265.200 124.800 ;
        RECT 284.400 119.700 286.200 129.600 ;
        RECT 311.400 119.700 313.200 124.800 ;
        RECT 340.500 119.700 342.300 126.600 ;
        RECT 354.900 119.700 356.700 126.600 ;
        RECT 374.700 119.700 376.500 123.600 ;
        RECT 382.200 119.700 384.000 126.600 ;
        RECT 395.400 119.700 397.200 129.600 ;
        RECT 419.700 119.700 421.500 126.600 ;
        RECT 443.400 119.700 445.200 124.800 ;
        RECT 464.400 119.700 466.200 123.600 ;
        RECT 485.700 119.700 487.500 123.600 ;
        RECT 493.200 119.700 495.000 126.600 ;
        RECT 503.400 119.700 505.200 129.600 ;
        RECT 538.800 119.700 540.600 129.600 ;
        RECT 552.000 119.700 553.800 126.600 ;
        RECT 559.500 119.700 561.300 123.600 ;
        RECT 575.400 119.700 577.200 129.600 ;
        RECT 601.800 119.700 603.600 123.600 ;
        RECT 617.400 119.700 619.200 124.800 ;
        RECT 638.400 119.700 640.200 124.800 ;
        RECT 659.400 119.700 661.200 123.600 ;
        RECT 677.400 119.700 679.200 129.600 ;
        RECT 701.700 119.700 703.500 126.600 ;
        RECT 725.400 119.700 727.200 124.800 ;
        RECT 743.700 119.700 745.500 126.600 ;
        RECT 772.800 119.700 774.600 124.800 ;
        RECT 789.000 119.700 790.800 126.600 ;
        RECT 796.500 119.700 798.300 123.600 ;
        RECT 809.700 119.700 811.500 126.600 ;
        RECT 838.800 119.700 840.600 124.800 ;
        RECT 854.400 119.700 856.200 126.600 ;
        RECT 860.400 119.700 862.200 126.600 ;
        RECT 877.800 119.700 879.600 126.600 ;
        RECT 883.800 119.700 885.600 126.600 ;
        RECT 889.800 119.700 891.600 126.600 ;
        RECT 895.800 119.700 897.600 126.600 ;
        RECT 901.800 119.700 903.600 126.600 ;
        RECT 921.450 119.700 930.450 195.300 ;
        RECT 0.600 117.300 930.450 119.700 ;
        RECT 19.800 112.200 21.600 117.300 ;
        RECT 46.800 107.400 48.600 117.300 ;
        RECT 62.400 112.200 64.200 117.300 ;
        RECT 83.400 107.400 85.200 117.300 ;
        RECT 115.800 112.200 117.600 117.300 ;
        RECT 134.700 113.400 136.500 117.300 ;
        RECT 142.200 110.400 144.000 117.300 ;
        RECT 155.400 107.400 157.200 117.300 ;
        RECT 187.800 107.400 189.600 117.300 ;
        RECT 201.000 110.400 202.800 117.300 ;
        RECT 208.500 113.400 210.300 117.300 ;
        RECT 227.700 113.400 229.500 117.300 ;
        RECT 235.200 110.400 237.000 117.300 ;
        RECT 245.400 107.400 247.200 117.300 ;
        RECT 269.700 113.400 271.500 117.300 ;
        RECT 277.200 110.400 279.000 117.300 ;
        RECT 295.800 112.200 297.600 117.300 ;
        RECT 319.800 112.200 321.600 117.300 ;
        RECT 346.800 107.400 348.600 117.300 ;
        RECT 362.400 112.200 364.200 117.300 ;
        RECT 380.400 107.400 382.200 117.300 ;
        RECT 404.400 107.400 406.200 117.300 ;
        RECT 432.900 110.400 434.700 117.300 ;
        RECT 457.500 110.400 459.300 117.300 ;
        RECT 466.500 110.400 468.300 117.300 ;
        RECT 482.700 113.400 484.500 117.300 ;
        RECT 490.200 110.400 492.000 117.300 ;
        RECT 500.400 107.400 502.200 117.300 ;
        RECT 529.800 112.200 531.600 117.300 ;
        RECT 548.400 112.200 550.200 117.300 ;
        RECT 580.800 107.400 582.600 117.300 ;
        RECT 594.000 110.400 595.800 117.300 ;
        RECT 601.500 113.400 603.300 117.300 ;
        RECT 631.800 113.400 633.600 117.300 ;
        RECT 637.800 113.400 639.900 117.300 ;
        RECT 656.400 112.200 658.200 117.300 ;
        RECT 674.400 113.400 676.200 117.300 ;
        RECT 692.700 110.400 694.500 117.300 ;
        RECT 716.700 113.400 718.500 117.300 ;
        RECT 724.200 110.400 726.000 117.300 ;
        RECT 737.700 110.400 739.500 117.300 ;
        RECT 746.700 110.400 748.500 117.300 ;
        RECT 764.700 113.400 766.500 117.300 ;
        RECT 772.200 110.400 774.000 117.300 ;
        RECT 783.000 110.400 784.800 117.300 ;
        RECT 790.500 113.400 792.300 117.300 ;
        RECT 808.500 110.400 810.300 117.300 ;
        RECT 817.500 110.400 819.300 117.300 ;
        RECT 831.000 110.400 832.800 117.300 ;
        RECT 838.500 113.400 840.300 117.300 ;
        RECT 856.500 110.400 858.300 117.300 ;
        RECT 865.500 110.400 867.300 117.300 ;
        RECT 878.400 113.400 880.200 117.300 ;
        RECT 896.400 113.400 898.200 117.300 ;
        RECT 22.800 41.700 24.600 51.600 ;
        RECT 33.000 41.700 34.800 48.600 ;
        RECT 40.500 41.700 42.300 45.600 ;
        RECT 59.700 41.700 61.500 45.600 ;
        RECT 67.200 41.700 69.000 48.600 ;
        RECT 77.400 41.700 79.200 51.600 ;
        RECT 109.800 41.700 111.600 46.800 ;
        RECT 125.700 41.700 127.500 45.600 ;
        RECT 133.200 41.700 135.000 48.600 ;
        RECT 154.800 41.700 156.600 46.800 ;
        RECT 175.800 41.700 177.600 46.800 ;
        RECT 191.400 41.700 193.200 46.800 ;
        RECT 215.400 41.700 217.200 47.700 ;
        RECT 224.100 41.700 225.900 47.700 ;
        RECT 242.700 41.700 244.500 48.600 ;
        RECT 268.500 41.700 270.300 48.600 ;
        RECT 277.500 41.700 279.300 48.600 ;
        RECT 290.400 41.700 292.200 51.600 ;
        RECT 322.800 41.700 324.600 51.600 ;
        RECT 336.000 41.700 337.800 48.600 ;
        RECT 343.500 41.700 345.300 45.600 ;
        RECT 367.800 41.700 369.600 46.800 ;
        RECT 383.400 41.700 385.200 45.600 ;
        RECT 412.800 41.700 414.600 51.600 ;
        RECT 425.400 41.700 427.200 51.600 ;
        RECT 457.800 41.700 459.600 46.800 ;
        RECT 473.400 41.700 475.200 46.800 ;
        RECT 496.800 41.700 498.600 45.600 ;
        RECT 506.400 41.700 508.200 51.600 ;
        RECT 530.400 41.700 532.200 51.600 ;
        RECT 551.400 41.700 553.200 45.600 ;
        RECT 577.800 41.700 579.600 51.600 ;
        RECT 591.000 41.700 592.800 48.600 ;
        RECT 598.500 41.700 600.300 45.600 ;
        RECT 614.400 41.700 616.200 45.600 ;
        RECT 632.400 41.700 634.200 46.800 ;
        RECT 655.500 41.700 657.300 48.600 ;
        RECT 664.500 41.700 666.300 48.600 ;
        RECT 682.800 41.700 684.600 45.600 ;
        RECT 689.850 41.700 691.650 45.600 ;
        RECT 698.850 41.700 700.650 45.600 ;
        RECT 705.750 41.700 707.550 45.600 ;
        RECT 715.050 41.700 716.850 45.600 ;
        RECT 736.800 41.700 738.600 45.600 ;
        RECT 754.500 41.700 756.300 48.600 ;
        RECT 763.500 41.700 765.300 48.600 ;
        RECT 781.800 41.700 783.600 45.600 ;
        RECT 788.850 41.700 790.650 45.600 ;
        RECT 797.850 41.700 799.650 45.600 ;
        RECT 804.750 41.700 806.550 45.600 ;
        RECT 814.050 41.700 815.850 45.600 ;
        RECT 825.150 41.700 826.950 45.600 ;
        RECT 834.450 41.700 836.250 45.600 ;
        RECT 841.350 41.700 843.150 45.600 ;
        RECT 850.350 41.700 852.150 45.600 ;
        RECT 863.400 41.700 865.200 51.600 ;
        RECT 890.400 41.700 892.200 46.800 ;
        RECT 921.450 41.700 930.450 117.300 ;
        RECT 0.600 39.300 930.450 41.700 ;
        RECT 14.700 35.400 16.500 39.300 ;
        RECT 22.200 32.400 24.000 39.300 ;
        RECT 37.800 35.400 39.600 39.300 ;
        RECT 58.800 34.200 60.600 39.300 ;
        RECT 71.400 29.400 73.200 39.300 ;
        RECT 95.400 29.400 97.200 39.300 ;
        RECT 122.400 34.200 124.200 39.300 ;
        RECT 148.800 35.400 150.600 39.300 ;
        RECT 158.400 29.400 160.200 39.300 ;
        RECT 182.400 29.400 184.200 39.300 ;
        RECT 207.000 32.400 208.800 39.300 ;
        RECT 214.500 35.400 216.300 39.300 ;
        RECT 238.500 32.400 240.300 39.300 ;
        RECT 262.800 29.400 264.600 39.300 ;
        RECT 276.000 32.400 277.800 39.300 ;
        RECT 283.500 35.400 285.300 39.300 ;
        RECT 299.400 29.400 301.200 39.300 ;
        RECT 324.000 32.400 325.800 39.300 ;
        RECT 331.500 35.400 333.300 39.300 ;
        RECT 344.400 35.400 346.200 39.300 ;
        RECT 365.700 35.400 367.500 39.300 ;
        RECT 373.200 32.400 375.000 39.300 ;
        RECT 386.700 32.400 388.500 39.300 ;
        RECT 410.400 34.200 412.200 39.300 ;
        RECT 432.000 32.400 433.800 39.300 ;
        RECT 439.500 35.400 441.300 39.300 ;
        RECT 452.400 29.400 454.200 39.300 ;
        RECT 484.800 34.200 486.600 39.300 ;
        RECT 503.100 35.400 505.200 39.300 ;
        RECT 509.400 35.400 511.200 39.300 ;
        RECT 539.400 34.200 541.200 39.300 ;
        RECT 560.700 35.400 562.500 39.300 ;
        RECT 568.200 32.400 570.000 39.300 ;
        RECT 587.100 33.300 588.900 39.300 ;
        RECT 595.800 33.300 597.600 39.300 ;
        RECT 616.500 32.400 618.300 39.300 ;
        RECT 630.000 32.400 631.800 39.300 ;
        RECT 637.500 35.400 639.300 39.300 ;
        RECT 653.400 35.400 655.200 39.300 ;
        RECT 659.400 35.400 661.200 39.300 ;
        RECT 674.400 34.200 676.200 39.300 ;
        RECT 698.400 35.400 700.200 39.300 ;
        RECT 711.150 35.400 712.950 39.300 ;
        RECT 720.450 35.400 722.250 39.300 ;
        RECT 727.350 35.400 729.150 39.300 ;
        RECT 736.350 35.400 738.150 39.300 ;
        RECT 755.400 35.400 757.200 39.300 ;
        RECT 768.150 35.400 769.950 39.300 ;
        RECT 777.450 35.400 779.250 39.300 ;
        RECT 784.350 35.400 786.150 39.300 ;
        RECT 793.350 35.400 795.150 39.300 ;
        RECT 809.400 35.400 811.200 39.300 ;
        RECT 830.400 35.400 832.200 39.300 ;
        RECT 853.800 35.400 855.600 39.300 ;
        RECT 869.400 35.400 871.200 39.300 ;
        RECT 895.500 32.400 897.300 39.300 ;
        RECT 921.450 0.300 930.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 936.300 920.400 938.700 ;
        RECT -9.450 860.700 -0.450 936.300 ;
        RECT 16.800 929.400 18.600 936.300 ;
        RECT 32.400 929.400 34.200 936.300 ;
        RECT 40.500 923.400 42.300 936.300 ;
        RECT 53.400 929.400 55.200 936.300 ;
        RECT 61.500 923.400 63.300 936.300 ;
        RECT 79.800 929.400 81.600 936.300 ;
        RECT 97.800 930.000 99.600 936.300 ;
        RECT 103.800 929.400 105.600 936.300 ;
        RECT 113.400 929.400 115.200 936.300 ;
        RECT 119.400 930.000 121.200 936.300 ;
        RECT 137.400 929.400 139.200 936.300 ;
        RECT 145.500 923.400 147.300 936.300 ;
        RECT 163.800 930.000 165.600 936.300 ;
        RECT 169.800 929.400 171.600 936.300 ;
        RECT 187.800 929.400 189.600 936.300 ;
        RECT 200.400 929.400 202.200 936.300 ;
        RECT 208.500 923.400 210.300 936.300 ;
        RECT 221.400 929.400 223.200 936.300 ;
        RECT 227.400 930.000 229.200 936.300 ;
        RECT 250.800 925.200 252.600 936.300 ;
        RECT 266.400 929.400 268.200 936.300 ;
        RECT 272.400 930.000 274.200 936.300 ;
        RECT 292.800 929.400 294.600 936.300 ;
        RECT 298.800 929.400 300.600 936.300 ;
        RECT 311.400 929.400 313.200 936.300 ;
        RECT 317.400 930.000 319.200 936.300 ;
        RECT 334.800 929.400 336.600 936.300 ;
        RECT 340.800 929.400 342.600 936.300 ;
        RECT 350.400 929.400 352.200 936.300 ;
        RECT 356.400 930.000 358.200 936.300 ;
        RECT 379.800 930.000 381.600 936.300 ;
        RECT 385.800 929.400 387.600 936.300 ;
        RECT 405.300 923.400 407.100 936.300 ;
        RECT 422.400 929.400 424.200 936.300 ;
        RECT 428.400 929.400 430.200 936.300 ;
        RECT 445.800 929.400 447.600 936.300 ;
        RECT 466.800 923.400 468.600 936.300 ;
        RECT 479.400 923.400 481.200 936.300 ;
        RECT 500.400 929.400 502.200 936.300 ;
        RECT 508.500 923.400 510.300 936.300 ;
        RECT 523.800 929.400 525.600 936.300 ;
        RECT 529.800 929.400 531.600 936.300 ;
        RECT 542.400 929.400 544.200 936.300 ;
        RECT 550.500 923.400 552.300 936.300 ;
        RECT 563.700 923.400 565.500 936.300 ;
        RECT 571.800 929.400 573.600 936.300 ;
        RECT 595.800 925.200 597.600 936.300 ;
        RECT 611.400 929.400 613.200 936.300 ;
        RECT 629.400 929.400 631.200 936.300 ;
        RECT 637.500 923.400 639.300 936.300 ;
        RECT 650.700 923.400 652.500 936.300 ;
        RECT 658.800 929.400 660.600 936.300 ;
        RECT 676.800 929.400 678.600 936.300 ;
        RECT 694.800 925.500 696.600 936.300 ;
        RECT 703.800 925.500 705.600 936.300 ;
        RECT 719.400 929.400 721.200 936.300 ;
        RECT 725.400 930.000 727.200 936.300 ;
        RECT 746.400 929.400 748.200 936.300 ;
        RECT 754.500 923.400 756.300 936.300 ;
        RECT 767.400 923.400 769.200 936.300 ;
        RECT 788.400 929.400 790.200 936.300 ;
        RECT 808.800 929.400 810.600 936.300 ;
        RECT 814.800 929.400 816.600 936.300 ;
        RECT 827.400 928.200 829.200 936.300 ;
        RECT 836.400 923.400 838.200 936.300 ;
        RECT 854.400 929.400 856.200 936.300 ;
        RECT 862.500 923.400 864.300 936.300 ;
        RECT 877.800 929.400 879.600 936.300 ;
        RECT 890.400 923.400 892.200 936.300 ;
        RECT 896.400 923.400 898.200 936.300 ;
        RECT 22.800 860.700 24.600 871.500 ;
        RECT 37.800 860.700 39.600 867.600 ;
        RECT 43.800 860.700 45.600 867.600 ;
        RECT 56.400 860.700 58.200 867.600 ;
        RECT 62.400 860.700 64.200 867.000 ;
        RECT 83.400 860.700 85.200 871.800 ;
        RECT 109.800 860.700 111.600 867.600 ;
        RECT 115.800 860.700 117.600 867.600 ;
        RECT 131.400 860.700 133.200 867.600 ;
        RECT 139.500 860.700 141.300 873.600 ;
        RECT 157.800 860.700 159.600 867.600 ;
        RECT 163.800 860.700 165.600 867.600 ;
        RECT 184.800 860.700 186.600 873.600 ;
        RECT 194.700 860.700 196.500 873.600 ;
        RECT 202.800 860.700 204.600 867.600 ;
        RECT 223.800 860.700 225.600 867.600 ;
        RECT 241.800 860.700 243.600 867.600 ;
        RECT 251.700 860.700 253.500 873.600 ;
        RECT 259.800 860.700 261.600 867.600 ;
        RECT 272.400 860.700 274.200 867.600 ;
        RECT 295.800 860.700 297.600 867.000 ;
        RECT 301.800 860.700 303.600 867.600 ;
        RECT 319.800 860.700 321.600 867.600 ;
        RECT 332.700 860.700 334.500 873.600 ;
        RECT 340.800 860.700 342.600 867.600 ;
        RECT 353.400 860.700 355.200 867.600 ;
        RECT 371.400 860.700 373.200 867.600 ;
        RECT 379.500 860.700 381.300 873.600 ;
        RECT 395.400 860.700 397.200 871.800 ;
        RECT 413.400 860.700 415.200 873.600 ;
        RECT 434.400 860.700 436.200 867.600 ;
        RECT 457.800 860.700 459.600 873.600 ;
        RECT 470.400 860.700 472.200 867.600 ;
        RECT 476.400 860.700 478.200 867.000 ;
        RECT 505.800 860.700 507.600 871.500 ;
        RECT 518.700 860.700 520.500 873.600 ;
        RECT 526.800 860.700 528.600 867.600 ;
        RECT 539.400 860.700 541.200 867.600 ;
        RECT 545.400 860.700 547.200 867.600 ;
        RECT 560.700 860.700 562.500 873.600 ;
        RECT 568.800 860.700 570.600 867.600 ;
        RECT 587.400 860.700 589.200 867.600 ;
        RECT 595.500 860.700 597.300 873.600 ;
        RECT 611.400 860.700 613.200 867.600 ;
        RECT 619.500 860.700 621.300 873.600 ;
        RECT 632.400 860.700 634.200 871.800 ;
        RECT 656.400 860.700 658.200 867.600 ;
        RECT 664.500 860.700 666.300 873.600 ;
        RECT 680.400 860.700 682.200 871.500 ;
        RECT 704.400 860.700 706.200 867.600 ;
        RECT 710.400 860.700 712.200 867.600 ;
        RECT 722.400 860.700 724.200 867.600 ;
        RECT 728.400 860.700 730.200 867.000 ;
        RECT 751.800 860.700 753.600 867.600 ;
        RECT 769.800 860.700 771.600 867.600 ;
        RECT 775.800 860.700 777.600 867.600 ;
        RECT 785.400 860.700 787.200 867.600 ;
        RECT 791.400 860.700 793.200 867.600 ;
        RECT 806.700 860.700 808.500 873.600 ;
        RECT 814.800 860.700 816.600 867.600 ;
        RECT 835.800 860.700 837.600 873.600 ;
        RECT 848.700 860.700 850.500 873.600 ;
        RECT 856.800 860.700 858.600 867.600 ;
        RECT 869.700 860.700 871.500 873.600 ;
        RECT 877.800 860.700 879.600 867.600 ;
        RECT 893.400 860.700 895.200 873.600 ;
        RECT -9.450 858.300 920.400 860.700 ;
        RECT -9.450 782.700 -0.450 858.300 ;
        RECT 13.800 851.400 15.600 858.300 ;
        RECT 28.800 851.400 30.600 858.300 ;
        RECT 34.800 851.400 36.600 858.300 ;
        RECT 49.800 851.400 51.600 858.300 ;
        RECT 55.800 851.400 57.600 858.300 ;
        RECT 68.400 847.200 70.200 858.300 ;
        RECT 94.800 852.000 96.600 858.300 ;
        RECT 100.800 851.400 102.600 858.300 ;
        RECT 115.800 852.000 117.600 858.300 ;
        RECT 121.800 851.400 123.600 858.300 ;
        RECT 139.800 851.400 141.600 858.300 ;
        RECT 159.300 845.400 161.100 858.300 ;
        RECT 178.800 851.400 180.600 858.300 ;
        RECT 184.800 851.400 186.600 858.300 ;
        RECT 196.800 851.400 198.600 858.300 ;
        RECT 202.800 851.400 204.600 858.300 ;
        RECT 223.800 845.400 225.600 858.300 ;
        RECT 236.400 851.400 238.200 858.300 ;
        RECT 242.400 851.400 244.200 858.300 ;
        RECT 257.400 845.400 259.200 858.300 ;
        RECT 275.400 851.400 277.200 858.300 ;
        RECT 281.400 851.400 283.200 858.300 ;
        RECT 301.800 851.400 303.600 858.300 ;
        RECT 307.800 851.400 309.600 858.300 ;
        RECT 320.400 851.400 322.200 858.300 ;
        RECT 328.500 845.400 330.300 858.300 ;
        RECT 344.400 851.400 346.200 858.300 ;
        RECT 352.500 845.400 354.300 858.300 ;
        RECT 365.700 845.400 367.500 858.300 ;
        RECT 373.800 851.400 375.600 858.300 ;
        RECT 393.900 845.400 395.700 858.300 ;
        RECT 413.400 851.400 415.200 858.300 ;
        RECT 419.400 851.400 421.200 858.300 ;
        RECT 436.800 851.400 438.600 858.300 ;
        RECT 442.800 851.400 444.600 858.300 ;
        RECT 457.800 851.400 459.600 858.300 ;
        RECT 463.800 851.400 465.600 858.300 ;
        RECT 478.800 851.400 480.600 858.300 ;
        RECT 484.800 851.400 486.600 858.300 ;
        RECT 499.800 852.000 501.600 858.300 ;
        RECT 505.800 851.400 507.600 858.300 ;
        RECT 529.800 847.500 531.600 858.300 ;
        RECT 547.800 851.400 549.600 858.300 ;
        RECT 553.800 851.400 555.600 858.300 ;
        RECT 568.800 845.400 570.600 858.300 ;
        RECT 583.800 851.400 585.600 858.300 ;
        RECT 589.800 851.400 591.600 858.300 ;
        RECT 610.800 847.200 612.600 858.300 ;
        RECT 626.700 845.400 628.500 858.300 ;
        RECT 634.800 851.400 636.600 858.300 ;
        RECT 647.400 851.400 649.200 858.300 ;
        RECT 653.400 851.400 655.200 858.300 ;
        RECT 671.400 851.400 673.200 858.300 ;
        RECT 679.500 845.400 681.300 858.300 ;
        RECT 689.400 851.400 691.200 858.300 ;
        RECT 695.400 851.400 697.200 858.300 ;
        RECT 710.400 851.400 712.200 858.300 ;
        RECT 716.400 852.000 718.200 858.300 ;
        RECT 737.400 851.400 739.200 858.300 ;
        RECT 745.500 845.400 747.300 858.300 ;
        RECT 761.400 847.500 763.200 858.300 ;
        RECT 785.400 851.400 787.200 858.300 ;
        RECT 808.800 847.500 810.600 858.300 ;
        RECT 817.800 847.500 819.600 858.300 ;
        RECT 838.800 851.400 840.600 858.300 ;
        RECT 859.800 847.200 861.600 858.300 ;
        RECT 872.700 845.400 874.500 858.300 ;
        RECT 880.800 851.400 882.600 858.300 ;
        RECT 901.800 851.400 903.600 858.300 ;
        RECT 18.300 782.700 20.100 795.600 ;
        RECT 43.800 782.700 45.600 793.800 ;
        RECT 58.800 782.700 60.600 789.600 ;
        RECT 64.800 782.700 66.600 789.600 ;
        RECT 79.800 782.700 81.600 789.000 ;
        RECT 85.800 782.700 87.600 789.600 ;
        RECT 98.400 782.700 100.200 789.600 ;
        RECT 104.400 782.700 106.200 789.000 ;
        RECT 125.400 782.700 127.200 793.800 ;
        RECT 146.700 782.700 148.500 795.600 ;
        RECT 154.800 782.700 156.600 789.600 ;
        RECT 172.800 782.700 174.600 789.600 ;
        RECT 178.800 782.700 180.600 789.600 ;
        RECT 188.400 782.700 190.200 789.600 ;
        RECT 194.400 782.700 196.200 789.000 ;
        RECT 215.400 782.700 217.200 793.500 ;
        RECT 224.100 782.700 226.200 793.500 ;
        RECT 242.400 782.700 244.200 789.600 ;
        RECT 248.400 782.700 250.200 789.600 ;
        RECT 264.300 782.700 266.100 795.600 ;
        RECT 274.800 782.700 276.600 795.600 ;
        RECT 287.700 782.700 289.500 795.600 ;
        RECT 295.800 782.700 297.600 789.600 ;
        RECT 308.400 782.700 310.200 789.600 ;
        RECT 329.400 782.700 331.200 789.600 ;
        RECT 337.500 782.700 339.300 795.600 ;
        RECT 347.700 782.700 349.500 795.600 ;
        RECT 355.800 782.700 357.600 789.600 ;
        RECT 371.400 782.700 373.200 789.600 ;
        RECT 377.400 782.700 379.200 789.000 ;
        RECT 395.400 782.700 397.200 789.600 ;
        RECT 401.400 782.700 403.200 789.600 ;
        RECT 413.700 782.700 415.500 795.600 ;
        RECT 421.800 782.700 423.600 789.600 ;
        RECT 434.400 782.700 436.200 789.600 ;
        RECT 449.400 782.700 451.200 789.600 ;
        RECT 464.400 782.700 466.200 789.600 ;
        RECT 470.400 782.700 472.200 789.600 ;
        RECT 490.800 782.700 492.600 789.600 ;
        RECT 496.800 782.700 498.600 789.600 ;
        RECT 520.800 782.700 522.600 793.500 ;
        RECT 533.700 782.700 535.500 795.600 ;
        RECT 541.800 782.700 543.600 789.600 ;
        RECT 557.700 782.700 559.500 795.600 ;
        RECT 565.800 782.700 567.600 789.600 ;
        RECT 578.700 782.700 580.500 795.600 ;
        RECT 586.800 782.700 588.600 789.600 ;
        RECT 604.800 782.700 606.600 789.600 ;
        RECT 628.800 782.700 630.600 793.500 ;
        RECT 649.800 782.700 651.600 789.600 ;
        RECT 661.800 782.700 663.600 789.600 ;
        RECT 667.800 782.700 669.600 789.600 ;
        RECT 679.800 782.700 681.600 789.600 ;
        RECT 685.800 782.700 687.600 789.600 ;
        RECT 698.400 782.700 700.200 789.600 ;
        RECT 704.400 782.700 706.200 789.600 ;
        RECT 719.400 782.700 721.200 795.600 ;
        RECT 742.800 782.700 744.600 795.600 ;
        RECT 751.800 782.700 753.600 790.800 ;
        RECT 769.800 782.700 771.600 789.600 ;
        RECT 785.400 782.700 787.200 795.600 ;
        RECT 806.400 782.700 808.200 789.600 ;
        RECT 814.500 782.700 816.300 795.600 ;
        RECT 824.700 782.700 826.500 795.600 ;
        RECT 832.800 782.700 834.600 789.600 ;
        RECT 848.700 782.700 850.500 795.600 ;
        RECT 856.800 782.700 858.600 789.600 ;
        RECT 869.400 782.700 871.200 789.600 ;
        RECT 892.800 782.700 894.600 789.600 ;
        RECT 910.800 782.700 912.600 789.600 ;
        RECT -9.450 780.300 920.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT 14.400 773.400 16.200 780.300 ;
        RECT 22.500 767.400 24.300 780.300 ;
        RECT 35.700 767.400 37.500 780.300 ;
        RECT 43.800 773.400 45.600 780.300 ;
        RECT 61.800 774.000 63.600 780.300 ;
        RECT 67.800 773.400 69.600 780.300 ;
        RECT 85.800 773.400 87.600 780.300 ;
        RECT 100.800 774.000 102.600 780.300 ;
        RECT 106.800 773.400 108.600 780.300 ;
        RECT 124.800 773.400 126.600 780.300 ;
        RECT 139.800 774.000 141.600 780.300 ;
        RECT 145.800 773.400 147.600 780.300 ;
        RECT 158.400 773.400 160.200 780.300 ;
        RECT 166.500 767.400 168.300 780.300 ;
        RECT 187.800 767.400 189.600 780.300 ;
        RECT 203.400 769.500 205.200 780.300 ;
        RECT 238.800 769.500 240.600 780.300 ;
        RECT 256.800 773.400 258.600 780.300 ;
        RECT 262.800 773.400 264.600 780.300 ;
        RECT 274.800 773.400 276.600 780.300 ;
        RECT 280.800 773.400 282.600 780.300 ;
        RECT 297.900 767.400 299.700 780.300 ;
        RECT 317.400 773.400 319.200 780.300 ;
        RECT 323.400 773.400 325.200 780.300 ;
        RECT 338.400 773.400 340.200 780.300 ;
        RECT 361.800 773.400 363.600 780.300 ;
        RECT 375.300 767.400 377.100 780.300 ;
        RECT 385.800 767.400 387.600 780.300 ;
        RECT 406.800 767.400 408.600 780.300 ;
        RECT 424.800 773.400 426.600 780.300 ;
        RECT 430.800 773.400 432.600 780.300 ;
        RECT 445.800 773.400 447.600 780.300 ;
        RECT 451.800 773.400 453.600 780.300 ;
        RECT 464.700 767.400 466.500 780.300 ;
        RECT 472.800 773.400 474.600 780.300 ;
        RECT 496.800 769.500 498.600 780.300 ;
        RECT 515.400 773.400 517.200 780.300 ;
        RECT 523.500 767.400 525.300 780.300 ;
        RECT 538.800 773.400 540.600 780.300 ;
        RECT 544.800 773.400 546.600 780.300 ;
        RECT 568.800 769.500 570.600 780.300 ;
        RECT 586.800 773.400 588.600 780.300 ;
        RECT 592.800 773.400 594.600 780.300 ;
        RECT 608.400 769.500 610.200 780.300 ;
        RECT 635.400 769.500 637.200 780.300 ;
        RECT 656.400 773.400 658.200 780.300 ;
        RECT 662.400 773.400 664.200 780.300 ;
        RECT 677.400 773.400 679.200 780.300 ;
        RECT 683.400 773.400 685.200 780.300 ;
        RECT 701.700 767.400 703.500 780.300 ;
        RECT 709.800 773.400 711.600 780.300 ;
        RECT 722.700 767.400 724.500 780.300 ;
        RECT 730.800 773.400 732.600 780.300 ;
        RECT 746.400 773.400 748.200 780.300 ;
        RECT 752.400 773.400 754.200 780.300 ;
        RECT 767.400 773.400 769.200 780.300 ;
        RECT 775.500 767.400 777.300 780.300 ;
        RECT 791.400 769.200 793.200 780.300 ;
        RECT 814.800 773.400 816.600 780.300 ;
        RECT 830.400 769.200 832.200 780.300 ;
        RECT 854.400 769.200 856.200 780.300 ;
        RECT 878.400 773.400 880.200 780.300 ;
        RECT 886.500 767.400 888.300 780.300 ;
        RECT 896.700 767.400 898.500 780.300 ;
        RECT 904.800 773.400 906.600 780.300 ;
        RECT 13.800 704.700 15.600 711.600 ;
        RECT 19.800 704.700 21.600 711.600 ;
        RECT 35.400 704.700 37.200 715.800 ;
        RECT 56.700 704.700 58.500 717.600 ;
        RECT 64.800 704.700 66.600 711.600 ;
        RECT 80.400 704.700 82.200 711.600 ;
        RECT 86.400 704.700 88.200 711.000 ;
        RECT 106.800 704.700 108.600 711.000 ;
        RECT 112.800 704.700 114.600 711.600 ;
        RECT 130.800 704.700 132.600 711.000 ;
        RECT 136.800 704.700 138.600 711.600 ;
        RECT 149.400 704.700 151.200 715.800 ;
        RECT 170.400 704.700 172.200 711.600 ;
        RECT 187.800 704.700 189.600 711.600 ;
        RECT 193.800 704.700 195.600 711.600 ;
        RECT 211.800 704.700 213.600 711.600 ;
        RECT 217.800 704.700 219.600 711.600 ;
        RECT 230.400 704.700 232.200 717.600 ;
        RECT 245.400 704.700 247.200 711.600 ;
        RECT 251.400 704.700 253.200 711.600 ;
        RECT 271.800 704.700 273.600 711.600 ;
        RECT 277.800 704.700 279.600 711.600 ;
        RECT 290.400 704.700 292.200 711.600 ;
        RECT 296.400 704.700 298.200 711.600 ;
        RECT 313.800 704.700 315.600 711.600 ;
        RECT 328.800 704.700 330.600 711.600 ;
        RECT 334.800 704.700 336.600 711.600 ;
        RECT 350.400 704.700 352.200 711.600 ;
        RECT 358.500 704.700 360.300 717.600 ;
        RECT 374.400 704.700 376.200 715.500 ;
        RECT 383.100 704.700 385.200 715.500 ;
        RECT 401.400 704.700 403.200 711.600 ;
        RECT 407.400 704.700 409.200 711.600 ;
        RECT 427.800 704.700 429.600 711.000 ;
        RECT 433.800 704.700 435.600 711.600 ;
        RECT 446.400 704.700 448.200 711.600 ;
        RECT 452.400 704.700 454.200 711.000 ;
        RECT 470.400 704.700 472.200 711.600 ;
        RECT 476.400 704.700 478.200 711.600 ;
        RECT 496.800 704.700 498.600 711.600 ;
        RECT 509.700 704.700 511.500 717.600 ;
        RECT 517.800 704.700 519.600 711.600 ;
        RECT 530.400 704.700 532.200 711.600 ;
        RECT 536.400 704.700 538.200 711.600 ;
        RECT 553.800 704.700 555.600 711.600 ;
        RECT 559.800 704.700 561.600 711.600 ;
        RECT 569.700 704.700 571.500 717.600 ;
        RECT 577.800 704.700 579.600 711.600 ;
        RECT 596.400 704.700 598.200 711.600 ;
        RECT 604.500 704.700 606.300 717.600 ;
        RECT 620.400 704.700 622.200 715.800 ;
        RECT 641.400 704.700 643.200 711.600 ;
        RECT 647.400 704.700 649.200 711.600 ;
        RECT 664.800 704.700 666.600 711.600 ;
        RECT 670.800 704.700 672.600 711.600 ;
        RECT 683.700 704.700 685.500 717.600 ;
        RECT 691.800 704.700 693.600 711.600 ;
        RECT 708.300 704.700 710.100 717.600 ;
        RECT 718.800 704.700 720.600 717.600 ;
        RECT 731.400 704.700 733.200 711.600 ;
        RECT 749.700 704.700 751.500 717.600 ;
        RECT 757.800 704.700 759.600 711.600 ;
        RECT 776.400 704.700 778.200 711.600 ;
        RECT 784.500 704.700 786.300 717.600 ;
        RECT 800.400 704.700 802.200 715.800 ;
        RECT 821.700 704.700 823.500 717.600 ;
        RECT 829.800 704.700 831.600 711.600 ;
        RECT 842.700 704.700 844.500 717.600 ;
        RECT 850.800 704.700 852.600 711.600 ;
        RECT 866.700 704.700 868.500 717.600 ;
        RECT 874.800 704.700 876.600 711.600 ;
        RECT 893.400 704.700 895.200 715.500 ;
        RECT 902.400 704.700 904.200 715.500 ;
        RECT -9.450 702.300 920.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT 10.800 695.400 12.600 702.300 ;
        RECT 16.800 695.400 18.600 702.300 ;
        RECT 29.400 695.400 31.200 702.300 ;
        RECT 35.400 696.000 37.200 702.300 ;
        RECT 61.800 691.200 63.600 702.300 ;
        RECT 77.400 695.400 79.200 702.300 ;
        RECT 83.400 696.000 85.200 702.300 ;
        RECT 104.400 691.200 106.200 702.300 ;
        RECT 128.400 691.500 130.200 702.300 ;
        RECT 137.400 691.500 139.200 702.300 ;
        RECT 163.800 689.400 165.600 702.300 ;
        RECT 180.300 689.400 182.100 702.300 ;
        RECT 190.800 689.400 192.600 702.300 ;
        RECT 203.400 695.400 205.200 702.300 ;
        RECT 209.400 695.400 211.200 702.300 ;
        RECT 226.800 696.000 228.600 702.300 ;
        RECT 232.800 695.400 234.600 702.300 ;
        RECT 253.800 691.200 255.600 702.300 ;
        RECT 269.400 695.400 271.200 702.300 ;
        RECT 277.500 689.400 279.300 702.300 ;
        RECT 292.800 695.400 294.600 702.300 ;
        RECT 298.800 695.400 300.600 702.300 ;
        RECT 314.400 695.400 316.200 702.300 ;
        RECT 322.500 689.400 324.300 702.300 ;
        RECT 340.800 695.400 342.600 702.300 ;
        RECT 358.800 695.400 360.600 702.300 ;
        RECT 376.800 691.500 378.600 702.300 ;
        RECT 385.800 691.500 387.600 702.300 ;
        RECT 406.800 695.400 408.600 702.300 ;
        RECT 422.400 689.400 424.200 702.300 ;
        RECT 437.700 689.400 439.500 702.300 ;
        RECT 445.800 695.400 447.600 702.300 ;
        RECT 464.400 695.400 466.200 702.300 ;
        RECT 485.400 695.400 487.200 702.300 ;
        RECT 506.400 691.500 508.200 702.300 ;
        RECT 515.400 691.500 517.200 702.300 ;
        RECT 536.400 695.400 538.200 702.300 ;
        RECT 554.400 695.400 556.200 702.300 ;
        RECT 560.400 695.400 562.200 702.300 ;
        RECT 583.800 689.400 585.600 702.300 ;
        RECT 599.400 695.400 601.200 702.300 ;
        RECT 617.400 695.400 619.200 702.300 ;
        RECT 623.400 695.400 625.200 702.300 ;
        RECT 635.400 695.400 637.200 702.300 ;
        RECT 655.800 695.400 657.600 702.300 ;
        RECT 668.400 695.400 670.200 702.300 ;
        RECT 676.500 689.400 678.300 702.300 ;
        RECT 689.700 689.400 691.500 702.300 ;
        RECT 697.800 695.400 699.600 702.300 ;
        RECT 716.400 691.500 718.200 702.300 ;
        RECT 725.400 691.500 727.200 702.300 ;
        RECT 743.400 691.200 745.200 702.300 ;
        RECT 764.700 689.400 766.500 702.300 ;
        RECT 772.800 695.400 774.600 702.300 ;
        RECT 791.400 695.400 793.200 702.300 ;
        RECT 799.500 689.400 801.300 702.300 ;
        RECT 809.700 689.400 811.500 702.300 ;
        RECT 817.800 695.400 819.600 702.300 ;
        RECT 837.900 689.400 839.700 702.300 ;
        RECT 862.800 691.500 864.600 702.300 ;
        RECT 871.800 691.500 873.600 702.300 ;
        RECT 892.800 689.400 894.600 702.300 ;
        RECT 908.400 691.200 910.200 702.300 ;
        RECT 19.800 626.700 21.600 639.600 ;
        RECT 32.400 626.700 34.200 633.600 ;
        RECT 40.500 626.700 42.300 639.600 ;
        RECT 56.400 626.700 58.200 637.800 ;
        RECT 74.700 626.700 76.500 639.600 ;
        RECT 82.800 626.700 84.600 633.600 ;
        RECT 102.900 626.700 104.700 639.600 ;
        RECT 125.400 626.700 127.200 637.500 ;
        RECT 134.100 626.700 136.200 637.500 ;
        RECT 149.700 626.700 151.500 639.600 ;
        RECT 157.800 626.700 159.600 633.600 ;
        RECT 173.400 626.700 175.200 633.600 ;
        RECT 179.400 626.700 181.200 633.600 ;
        RECT 196.800 626.700 198.600 633.600 ;
        RECT 202.800 626.700 204.600 633.600 ;
        RECT 220.800 626.700 222.900 637.500 ;
        RECT 229.800 626.700 231.600 637.500 ;
        RECT 247.800 626.700 249.600 633.600 ;
        RECT 253.800 626.700 255.600 633.600 ;
        RECT 267.300 626.700 269.100 639.600 ;
        RECT 277.800 626.700 279.600 639.600 ;
        RECT 295.800 626.700 297.600 633.600 ;
        RECT 301.800 626.700 303.600 633.600 ;
        RECT 316.800 626.700 318.600 633.600 ;
        RECT 322.800 626.700 324.600 633.600 ;
        RECT 340.800 626.700 342.600 633.600 ;
        RECT 361.800 626.700 363.600 633.600 ;
        RECT 382.800 626.700 384.600 637.500 ;
        RECT 391.800 626.700 393.600 637.500 ;
        RECT 407.700 626.700 409.500 639.600 ;
        RECT 415.800 626.700 417.600 633.600 ;
        RECT 425.550 626.700 427.350 630.600 ;
        RECT 434.250 626.700 436.050 633.600 ;
        RECT 440.850 626.700 442.650 633.600 ;
        RECT 451.050 626.700 452.850 633.600 ;
        RECT 461.550 626.700 463.350 630.600 ;
        RECT 470.250 626.700 472.050 633.600 ;
        RECT 476.850 626.700 478.650 633.600 ;
        RECT 487.050 626.700 488.850 633.600 ;
        RECT 503.400 626.700 505.200 633.600 ;
        RECT 511.500 626.700 513.300 639.600 ;
        RECT 524.700 626.700 526.500 639.600 ;
        RECT 532.800 626.700 534.600 633.600 ;
        RECT 553.800 626.700 555.600 633.600 ;
        RECT 560.550 626.700 562.350 630.600 ;
        RECT 569.250 626.700 571.050 633.600 ;
        RECT 575.850 626.700 577.650 633.600 ;
        RECT 586.050 626.700 587.850 633.600 ;
        RECT 605.400 626.700 607.200 633.600 ;
        RECT 613.500 626.700 615.300 639.600 ;
        RECT 623.400 626.700 625.200 633.600 ;
        RECT 641.400 626.700 643.200 637.500 ;
        RECT 650.100 626.700 652.200 637.500 ;
        RECT 668.700 626.700 670.500 639.600 ;
        RECT 676.800 626.700 678.600 633.600 ;
        RECT 700.800 626.700 702.600 637.800 ;
        RECT 724.800 626.700 726.600 637.800 ;
        RECT 737.400 626.700 739.200 633.600 ;
        RECT 755.400 626.700 757.200 633.600 ;
        RECT 763.500 626.700 765.300 639.600 ;
        RECT 781.800 626.700 783.600 633.600 ;
        RECT 799.800 626.700 801.600 633.600 ;
        RECT 812.700 626.700 814.500 639.600 ;
        RECT 820.800 626.700 822.600 633.600 ;
        RECT 839.400 626.700 841.200 637.500 ;
        RECT 860.700 626.700 862.500 639.600 ;
        RECT 868.800 626.700 870.600 633.600 ;
        RECT 886.800 626.700 888.600 633.600 ;
        RECT 892.800 626.700 894.600 633.600 ;
        RECT 902.400 626.700 904.200 633.600 ;
        RECT -9.450 624.300 920.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT 19.800 613.200 21.600 624.300 ;
        RECT 35.400 617.400 37.200 624.300 ;
        RECT 41.400 618.000 43.200 624.300 ;
        RECT 56.400 611.400 58.200 624.300 ;
        RECT 80.400 617.400 82.200 624.300 ;
        RECT 88.500 611.400 90.300 624.300 ;
        RECT 98.400 611.400 100.200 624.300 ;
        RECT 119.400 613.500 121.200 624.300 ;
        RECT 128.100 613.500 130.200 624.300 ;
        RECT 146.400 613.500 148.200 624.300 ;
        RECT 155.400 613.500 157.200 624.300 ;
        RECT 173.400 617.400 175.200 624.300 ;
        RECT 179.400 618.000 181.200 624.300 ;
        RECT 199.800 617.400 201.600 624.300 ;
        RECT 205.800 617.400 207.600 624.300 ;
        RECT 223.800 617.400 225.600 624.300 ;
        RECT 229.800 617.400 231.600 624.300 ;
        RECT 242.400 617.400 244.200 624.300 ;
        RECT 265.800 618.000 267.600 624.300 ;
        RECT 271.800 617.400 273.600 624.300 ;
        RECT 284.400 617.400 286.200 624.300 ;
        RECT 302.400 617.400 304.200 624.300 ;
        RECT 308.400 617.400 310.200 624.300 ;
        RECT 323.400 611.400 325.200 624.300 ;
        RECT 341.400 613.500 343.200 624.300 ;
        RECT 365.400 617.400 367.200 624.300 ;
        RECT 371.400 617.400 373.200 624.300 ;
        RECT 389.400 617.400 391.200 624.300 ;
        RECT 406.800 617.400 408.600 624.300 ;
        RECT 412.800 617.400 414.600 624.300 ;
        RECT 425.400 617.400 427.200 624.300 ;
        RECT 445.800 611.400 447.600 624.300 ;
        RECT 451.800 611.400 453.600 624.300 ;
        RECT 458.550 620.400 460.350 624.300 ;
        RECT 467.250 617.400 469.050 624.300 ;
        RECT 473.850 617.400 475.650 624.300 ;
        RECT 484.050 617.400 485.850 624.300 ;
        RECT 500.400 617.400 502.200 624.300 ;
        RECT 506.400 617.400 508.200 624.300 ;
        RECT 515.550 620.400 517.350 624.300 ;
        RECT 524.250 617.400 526.050 624.300 ;
        RECT 530.850 617.400 532.650 624.300 ;
        RECT 541.050 617.400 542.850 624.300 ;
        RECT 557.400 617.400 559.200 624.300 ;
        RECT 563.400 617.400 565.200 624.300 ;
        RECT 581.400 617.400 583.200 624.300 ;
        RECT 589.500 611.400 591.300 624.300 ;
        RECT 602.400 617.400 604.200 624.300 ;
        RECT 608.400 617.400 610.200 624.300 ;
        RECT 623.400 617.400 625.200 624.300 ;
        RECT 631.500 611.400 633.300 624.300 ;
        RECT 646.800 617.400 648.600 624.300 ;
        RECT 662.400 617.400 664.200 624.300 ;
        RECT 670.500 611.400 672.300 624.300 ;
        RECT 683.400 617.400 685.200 624.300 ;
        RECT 689.400 617.400 691.200 624.300 ;
        RECT 701.400 611.400 703.200 624.300 ;
        RECT 724.800 617.400 726.600 624.300 ;
        RECT 730.800 617.400 732.600 624.300 ;
        RECT 743.400 613.500 745.200 624.300 ;
        RECT 752.400 613.500 754.200 624.300 ;
        RECT 770.400 617.400 772.200 624.300 ;
        RECT 791.400 613.200 793.200 624.300 ;
        RECT 815.400 613.500 817.200 624.300 ;
        RECT 824.400 613.500 826.200 624.300 ;
        RECT 844.800 617.400 846.600 624.300 ;
        RECT 850.800 617.400 852.600 624.300 ;
        RECT 863.400 617.400 865.200 624.300 ;
        RECT 869.400 617.400 871.200 624.300 ;
        RECT 886.800 618.000 888.600 624.300 ;
        RECT 892.800 617.400 894.600 624.300 ;
        RECT 905.400 617.400 907.200 624.300 ;
        RECT 911.400 618.000 913.200 624.300 ;
        RECT 22.800 548.700 24.600 559.500 ;
        RECT 40.800 548.700 42.600 555.600 ;
        RECT 46.800 548.700 48.600 555.600 ;
        RECT 59.400 548.700 61.200 555.600 ;
        RECT 65.400 548.700 67.200 555.600 ;
        RECT 82.800 548.700 84.600 555.600 ;
        RECT 88.800 548.700 90.600 555.600 ;
        RECT 101.400 548.700 103.200 555.600 ;
        RECT 107.400 548.700 109.200 555.600 ;
        RECT 119.400 548.700 121.200 555.600 ;
        RECT 125.400 548.700 127.200 555.600 ;
        RECT 140.400 548.700 142.200 555.600 ;
        RECT 146.400 548.700 148.200 555.000 ;
        RECT 164.400 548.700 166.200 559.800 ;
        RECT 188.400 548.700 190.200 555.600 ;
        RECT 196.500 548.700 198.300 561.600 ;
        RECT 209.400 548.700 211.200 555.600 ;
        RECT 215.400 548.700 217.200 555.000 ;
        RECT 235.800 548.700 237.600 555.600 ;
        RECT 241.800 548.700 243.600 555.600 ;
        RECT 256.800 548.700 258.600 555.000 ;
        RECT 262.800 548.700 264.600 555.600 ;
        RECT 272.700 548.700 274.500 561.600 ;
        RECT 280.800 548.700 282.600 555.600 ;
        RECT 296.700 548.700 298.500 561.600 ;
        RECT 304.800 548.700 306.600 555.600 ;
        RECT 325.800 548.700 327.600 555.600 ;
        RECT 331.800 548.700 333.600 555.600 ;
        RECT 349.800 548.700 351.600 555.600 ;
        RECT 367.800 548.700 369.600 555.600 ;
        RECT 380.400 548.700 382.200 555.600 ;
        RECT 386.400 548.700 388.200 555.000 ;
        RECT 412.800 548.700 414.600 561.600 ;
        RECT 425.400 548.700 427.200 555.600 ;
        RECT 433.500 548.700 435.300 561.600 ;
        RECT 446.400 548.700 448.200 555.600 ;
        RECT 452.400 548.700 454.200 555.600 ;
        RECT 470.400 548.700 472.200 555.600 ;
        RECT 478.500 548.700 480.300 561.600 ;
        RECT 485.550 548.700 487.350 552.600 ;
        RECT 494.250 548.700 496.050 555.600 ;
        RECT 500.850 548.700 502.650 555.600 ;
        RECT 511.050 548.700 512.850 555.600 ;
        RECT 527.700 548.700 529.500 561.600 ;
        RECT 535.800 548.700 537.600 555.600 ;
        RECT 548.400 548.700 550.200 555.600 ;
        RECT 554.400 548.700 556.200 555.600 ;
        RECT 571.800 548.700 573.600 555.600 ;
        RECT 586.800 548.700 588.600 555.600 ;
        RECT 592.800 548.700 594.600 555.600 ;
        RECT 608.400 548.700 610.200 555.600 ;
        RECT 616.500 548.700 618.300 561.600 ;
        RECT 623.550 548.700 625.350 552.600 ;
        RECT 632.250 548.700 634.050 555.600 ;
        RECT 638.850 548.700 640.650 555.600 ;
        RECT 649.050 548.700 650.850 555.600 ;
        RECT 670.800 548.700 672.600 555.600 ;
        RECT 685.800 548.700 687.600 561.600 ;
        RECT 691.800 548.700 693.600 561.600 ;
        RECT 697.800 548.700 699.600 561.600 ;
        RECT 703.800 548.700 705.600 561.600 ;
        RECT 709.800 548.700 711.600 561.600 ;
        RECT 724.800 548.700 726.600 555.600 ;
        RECT 737.400 548.700 739.200 561.600 ;
        RECT 763.800 548.700 765.600 555.600 ;
        RECT 769.800 548.700 771.600 555.600 ;
        RECT 781.800 548.700 783.600 561.600 ;
        RECT 787.800 548.700 789.600 561.600 ;
        RECT 793.800 548.700 795.600 561.600 ;
        RECT 799.800 548.700 801.600 561.600 ;
        RECT 805.800 548.700 807.600 561.600 ;
        RECT 818.400 548.700 820.200 561.600 ;
        RECT 841.800 548.700 843.600 555.000 ;
        RECT 847.800 548.700 849.600 555.600 ;
        RECT 862.800 548.700 864.600 555.600 ;
        RECT 868.800 548.700 870.600 555.600 ;
        RECT 881.400 548.700 883.200 555.600 ;
        RECT 887.400 548.700 889.200 555.600 ;
        RECT 902.400 548.700 904.200 555.600 ;
        RECT -9.450 546.300 920.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT 14.400 536.400 16.200 546.300 ;
        RECT 49.800 539.400 51.600 546.300 ;
        RECT 55.800 539.400 57.600 546.300 ;
        RECT 73.800 540.000 75.600 546.300 ;
        RECT 79.800 539.400 81.600 546.300 ;
        RECT 92.400 535.200 94.200 546.300 ;
        RECT 113.400 535.200 115.200 546.300 ;
        RECT 137.400 539.400 139.200 546.300 ;
        RECT 145.500 533.400 147.300 546.300 ;
        RECT 158.700 533.400 160.500 546.300 ;
        RECT 166.800 539.400 168.600 546.300 ;
        RECT 187.800 540.000 189.600 546.300 ;
        RECT 193.800 539.400 195.600 546.300 ;
        RECT 208.800 540.000 210.600 546.300 ;
        RECT 214.800 539.400 216.600 546.300 ;
        RECT 229.800 540.000 231.600 546.300 ;
        RECT 235.800 539.400 237.600 546.300 ;
        RECT 248.400 539.400 250.200 546.300 ;
        RECT 266.400 539.400 268.200 546.300 ;
        RECT 272.400 540.000 274.200 546.300 ;
        RECT 290.400 539.400 292.200 546.300 ;
        RECT 296.400 540.000 298.200 546.300 ;
        RECT 311.400 533.400 313.200 546.300 ;
        RECT 332.400 535.500 334.200 546.300 ;
        RECT 356.400 533.400 358.200 546.300 ;
        RECT 373.800 539.400 375.600 546.300 ;
        RECT 379.800 539.400 381.600 546.300 ;
        RECT 392.400 539.400 394.200 546.300 ;
        RECT 412.800 539.400 414.600 546.300 ;
        RECT 418.800 539.400 420.600 546.300 ;
        RECT 434.400 535.500 436.200 546.300 ;
        RECT 461.400 539.400 463.200 546.300 ;
        RECT 469.500 533.400 471.300 546.300 ;
        RECT 479.400 539.400 481.200 546.300 ;
        RECT 485.400 539.400 487.200 546.300 ;
        RECT 497.700 533.400 499.500 546.300 ;
        RECT 505.800 539.400 507.600 546.300 ;
        RECT 521.700 533.400 523.500 546.300 ;
        RECT 529.800 539.400 531.600 546.300 ;
        RECT 547.800 539.400 549.600 546.300 ;
        RECT 560.400 539.400 562.200 546.300 ;
        RECT 583.800 539.400 585.600 546.300 ;
        RECT 593.550 542.400 595.350 546.300 ;
        RECT 602.250 539.400 604.050 546.300 ;
        RECT 608.850 539.400 610.650 546.300 ;
        RECT 619.050 539.400 620.850 546.300 ;
        RECT 640.800 539.400 642.600 546.300 ;
        RECT 658.800 539.400 660.600 546.300 ;
        RECT 673.800 539.400 675.600 546.300 ;
        RECT 679.800 539.400 681.600 546.300 ;
        RECT 686.550 542.400 688.350 546.300 ;
        RECT 695.250 539.400 697.050 546.300 ;
        RECT 701.850 539.400 703.650 546.300 ;
        RECT 712.050 539.400 713.850 546.300 ;
        RECT 722.550 542.400 724.350 546.300 ;
        RECT 731.250 539.400 733.050 546.300 ;
        RECT 737.850 539.400 739.650 546.300 ;
        RECT 748.050 539.400 749.850 546.300 ;
        RECT 758.550 542.400 760.350 546.300 ;
        RECT 767.250 539.400 769.050 546.300 ;
        RECT 773.850 539.400 775.650 546.300 ;
        RECT 784.050 539.400 785.850 546.300 ;
        RECT 805.800 539.400 807.600 546.300 ;
        RECT 815.400 539.400 817.200 546.300 ;
        RECT 821.400 539.400 823.200 546.300 ;
        RECT 833.400 539.400 835.200 546.300 ;
        RECT 839.400 540.000 841.200 546.300 ;
        RECT 857.700 533.400 859.500 546.300 ;
        RECT 865.800 539.400 867.600 546.300 ;
        RECT 883.800 539.400 885.600 546.300 ;
        RECT 889.800 539.400 891.600 546.300 ;
        RECT 907.800 540.000 909.600 546.300 ;
        RECT 913.800 539.400 915.600 546.300 ;
        RECT 11.700 470.700 13.500 483.600 ;
        RECT 19.800 470.700 21.600 477.600 ;
        RECT 37.800 470.700 39.600 477.000 ;
        RECT 43.800 470.700 45.600 477.600 ;
        RECT 56.400 470.700 58.200 481.800 ;
        RECT 77.400 470.700 79.200 477.600 ;
        RECT 83.400 470.700 85.200 477.000 ;
        RECT 103.800 470.700 105.600 477.000 ;
        RECT 109.800 470.700 111.600 477.600 ;
        RECT 122.700 470.700 124.500 483.600 ;
        RECT 130.800 470.700 132.600 477.600 ;
        RECT 154.800 470.700 156.600 481.500 ;
        RECT 172.800 470.700 174.600 477.600 ;
        RECT 178.800 470.700 180.600 477.600 ;
        RECT 191.400 470.700 193.200 477.600 ;
        RECT 197.400 470.700 199.200 477.600 ;
        RECT 217.800 470.700 219.600 477.000 ;
        RECT 223.800 470.700 225.600 477.600 ;
        RECT 238.800 470.700 240.600 477.600 ;
        RECT 254.400 470.700 256.200 477.600 ;
        RECT 262.500 470.700 264.300 483.600 ;
        RECT 278.400 470.700 280.200 477.600 ;
        RECT 286.500 470.700 288.300 483.600 ;
        RECT 301.800 470.700 303.600 477.600 ;
        RECT 307.800 470.700 309.600 477.600 ;
        RECT 317.400 470.700 319.200 477.600 ;
        RECT 323.400 470.700 325.200 477.600 ;
        RECT 342.900 470.700 344.700 483.600 ;
        RECT 362.400 470.700 364.200 477.600 ;
        RECT 368.400 470.700 370.200 477.600 ;
        RECT 385.800 470.700 387.600 477.600 ;
        RECT 391.800 470.700 393.600 477.600 ;
        RECT 404.400 470.700 406.200 477.600 ;
        RECT 422.400 470.700 424.200 477.600 ;
        RECT 428.400 470.700 430.200 477.600 ;
        RECT 443.400 470.700 445.200 477.600 ;
        RECT 449.400 470.700 451.200 477.600 ;
        RECT 461.700 470.700 463.500 483.600 ;
        RECT 469.800 470.700 471.600 477.600 ;
        RECT 493.800 470.700 495.600 481.800 ;
        RECT 512.400 470.700 514.200 481.800 ;
        RECT 533.400 470.700 535.200 477.600 ;
        RECT 551.400 470.700 553.200 477.600 ;
        RECT 557.400 470.700 559.200 477.000 ;
        RECT 580.800 470.700 582.600 481.800 ;
        RECT 596.400 470.700 598.200 477.600 ;
        RECT 602.400 470.700 604.200 477.000 ;
        RECT 620.400 470.700 622.200 477.600 ;
        RECT 626.400 470.700 628.200 477.000 ;
        RECT 647.400 470.700 649.200 477.600 ;
        RECT 667.800 470.700 669.600 477.600 ;
        RECT 673.800 470.700 675.600 477.600 ;
        RECT 686.700 470.700 688.500 483.600 ;
        RECT 694.800 470.700 696.600 477.600 ;
        RECT 710.700 470.700 712.500 483.600 ;
        RECT 718.800 470.700 720.600 477.600 ;
        RECT 734.400 470.700 736.200 477.600 ;
        RECT 740.400 470.700 742.200 477.600 ;
        RECT 755.400 470.700 757.200 483.600 ;
        RECT 779.400 470.700 781.200 477.600 ;
        RECT 787.500 470.700 789.300 483.600 ;
        RECT 800.400 470.700 802.200 477.600 ;
        RECT 818.700 470.700 820.500 483.600 ;
        RECT 826.800 470.700 828.600 477.600 ;
        RECT 839.400 470.700 841.200 477.600 ;
        RECT 845.400 470.700 847.200 477.600 ;
        RECT 860.400 470.700 862.200 483.600 ;
        RECT 881.400 470.700 883.200 477.600 ;
        RECT 887.400 470.700 889.200 477.000 ;
        RECT 904.800 470.700 906.600 477.600 ;
        RECT 910.800 470.700 912.600 477.600 ;
        RECT -9.450 468.300 920.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT 11.700 455.400 13.500 468.300 ;
        RECT 19.800 461.400 21.600 468.300 ;
        RECT 40.800 462.000 42.600 468.300 ;
        RECT 46.800 461.400 48.600 468.300 ;
        RECT 62.400 457.200 64.200 468.300 ;
        RECT 86.400 457.200 88.200 468.300 ;
        RECT 107.400 461.400 109.200 468.300 ;
        RECT 115.500 455.400 117.300 468.300 ;
        RECT 131.400 461.400 133.200 468.300 ;
        RECT 139.500 455.400 141.300 468.300 ;
        RECT 149.700 455.400 151.500 468.300 ;
        RECT 157.800 461.400 159.600 468.300 ;
        RECT 173.400 457.200 175.200 468.300 ;
        RECT 194.400 461.400 196.200 468.300 ;
        RECT 217.800 462.000 219.600 468.300 ;
        RECT 223.800 461.400 225.600 468.300 ;
        RECT 244.800 457.200 246.600 468.300 ;
        RECT 257.400 461.400 259.200 468.300 ;
        RECT 263.400 462.000 265.200 468.300 ;
        RECT 281.700 455.400 283.500 468.300 ;
        RECT 289.800 461.400 291.600 468.300 ;
        RECT 305.400 455.400 307.200 468.300 ;
        RECT 328.800 461.400 330.600 468.300 ;
        RECT 334.800 461.400 336.600 468.300 ;
        RECT 347.400 457.200 349.200 468.300 ;
        RECT 373.800 461.400 375.600 468.300 ;
        RECT 392.400 457.200 394.200 468.300 ;
        RECT 413.700 455.400 415.500 468.300 ;
        RECT 421.800 461.400 423.600 468.300 ;
        RECT 437.400 457.500 439.200 468.300 ;
        RECT 466.800 455.400 468.600 468.300 ;
        RECT 479.400 461.400 481.200 468.300 ;
        RECT 485.400 462.000 487.200 468.300 ;
        RECT 503.400 455.400 505.200 468.300 ;
        RECT 524.400 461.400 526.200 468.300 ;
        RECT 530.400 462.000 532.200 468.300 ;
        RECT 545.700 455.400 547.500 468.300 ;
        RECT 553.800 461.400 555.600 468.300 ;
        RECT 563.550 464.400 565.350 468.300 ;
        RECT 572.250 461.400 574.050 468.300 ;
        RECT 578.850 461.400 580.650 468.300 ;
        RECT 589.050 461.400 590.850 468.300 ;
        RECT 605.400 461.400 607.200 468.300 ;
        RECT 611.400 461.400 613.200 468.300 ;
        RECT 629.400 461.400 631.200 468.300 ;
        RECT 637.500 455.400 639.300 468.300 ;
        RECT 650.700 455.400 652.500 468.300 ;
        RECT 658.800 461.400 660.600 468.300 ;
        RECT 668.550 464.400 670.350 468.300 ;
        RECT 677.250 461.400 679.050 468.300 ;
        RECT 683.850 461.400 685.650 468.300 ;
        RECT 694.050 461.400 695.850 468.300 ;
        RECT 704.550 464.400 706.350 468.300 ;
        RECT 713.250 461.400 715.050 468.300 ;
        RECT 719.850 461.400 721.650 468.300 ;
        RECT 730.050 461.400 731.850 468.300 ;
        RECT 748.800 455.400 750.600 468.300 ;
        RECT 754.800 455.400 756.600 468.300 ;
        RECT 760.800 455.400 762.600 468.300 ;
        RECT 766.800 455.400 768.600 468.300 ;
        RECT 772.800 455.400 774.600 468.300 ;
        RECT 788.400 461.400 790.200 468.300 ;
        RECT 806.400 461.400 808.200 468.300 ;
        RECT 831.300 455.400 833.100 468.300 ;
        RECT 856.800 455.400 858.600 468.300 ;
        RECT 871.800 461.400 873.600 468.300 ;
        RECT 883.800 461.400 885.600 468.300 ;
        RECT 889.800 461.400 891.600 468.300 ;
        RECT 907.800 462.000 909.600 468.300 ;
        RECT 913.800 461.400 915.600 468.300 ;
        RECT 16.800 392.700 18.600 399.000 ;
        RECT 22.800 392.700 24.600 399.600 ;
        RECT 35.400 392.700 37.200 399.600 ;
        RECT 41.400 392.700 43.200 399.000 ;
        RECT 61.800 392.700 63.600 399.000 ;
        RECT 67.800 392.700 69.600 399.600 ;
        RECT 83.400 392.700 85.200 403.800 ;
        RECT 107.400 392.700 109.200 399.600 ;
        RECT 115.500 392.700 117.300 405.600 ;
        RECT 133.800 392.700 135.600 403.800 ;
        RECT 149.400 392.700 151.200 399.600 ;
        RECT 167.400 392.700 169.200 399.600 ;
        RECT 173.400 392.700 175.200 399.000 ;
        RECT 191.400 392.700 193.200 399.600 ;
        RECT 197.400 392.700 199.200 399.000 ;
        RECT 215.400 392.700 217.200 403.500 ;
        RECT 239.400 392.700 241.200 399.600 ;
        RECT 262.800 392.700 264.600 399.000 ;
        RECT 268.800 392.700 270.600 399.600 ;
        RECT 286.800 392.700 288.600 399.600 ;
        RECT 299.400 392.700 301.200 399.600 ;
        RECT 305.400 392.700 307.200 399.600 ;
        RECT 320.400 392.700 322.200 405.600 ;
        RECT 340.800 392.700 342.600 399.600 ;
        RECT 346.800 392.700 348.600 399.600 ;
        RECT 356.400 392.700 358.200 399.600 ;
        RECT 362.400 392.700 364.200 399.600 ;
        RECT 380.400 392.700 382.200 399.600 ;
        RECT 401.400 392.700 403.200 399.600 ;
        RECT 409.500 392.700 411.300 405.600 ;
        RECT 422.400 392.700 424.200 399.600 ;
        RECT 428.400 392.700 430.200 399.600 ;
        RECT 443.400 392.700 445.200 399.600 ;
        RECT 449.400 392.700 451.200 399.000 ;
        RECT 472.800 392.700 474.600 403.500 ;
        RECT 481.800 392.700 483.600 403.500 ;
        RECT 497.400 392.700 499.200 399.600 ;
        RECT 503.400 392.700 505.200 399.600 ;
        RECT 518.700 392.700 520.500 405.600 ;
        RECT 526.800 392.700 528.600 399.600 ;
        RECT 542.700 392.700 544.500 405.600 ;
        RECT 550.800 392.700 552.600 399.600 ;
        RECT 571.800 392.700 573.600 399.600 ;
        RECT 587.400 392.700 589.200 399.600 ;
        RECT 595.500 392.700 597.300 405.600 ;
        RECT 613.800 392.700 615.600 399.600 ;
        RECT 629.700 392.700 631.500 405.600 ;
        RECT 637.800 392.700 639.600 399.600 ;
        RECT 655.800 392.700 657.600 399.600 ;
        RECT 661.800 392.700 663.600 399.600 ;
        RECT 674.400 392.700 676.200 399.600 ;
        RECT 682.500 392.700 684.300 405.600 ;
        RECT 695.400 392.700 697.200 405.600 ;
        RECT 721.800 392.700 723.600 405.600 ;
        RECT 729.150 392.700 730.950 399.600 ;
        RECT 739.350 392.700 741.150 399.600 ;
        RECT 745.950 392.700 747.750 399.600 ;
        RECT 754.650 392.700 756.450 396.600 ;
        RECT 770.700 392.700 772.500 405.600 ;
        RECT 778.800 392.700 780.600 399.600 ;
        RECT 791.400 392.700 793.200 399.600 ;
        RECT 797.400 392.700 799.200 399.600 ;
        RECT 816.300 392.700 818.100 405.600 ;
        RECT 826.800 392.700 828.600 405.600 ;
        RECT 841.800 392.700 843.600 399.600 ;
        RECT 857.400 392.700 859.200 403.500 ;
        RECT 878.400 392.700 880.200 405.600 ;
        RECT 899.400 392.700 901.200 399.600 ;
        RECT -9.450 390.300 920.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT 13.800 383.400 15.600 390.300 ;
        RECT 19.800 383.400 21.600 390.300 ;
        RECT 32.400 383.400 34.200 390.300 ;
        RECT 38.400 383.400 40.200 390.300 ;
        RECT 56.400 379.200 58.200 390.300 ;
        RECT 79.800 383.400 81.600 390.300 ;
        RECT 92.700 377.400 94.500 390.300 ;
        RECT 100.800 383.400 102.600 390.300 ;
        RECT 124.800 377.400 126.600 390.300 ;
        RECT 139.800 383.400 141.600 390.300 ;
        RECT 145.800 383.400 147.600 390.300 ;
        RECT 157.800 383.400 159.600 390.300 ;
        RECT 163.800 383.400 165.600 390.300 ;
        RECT 176.400 383.400 178.200 390.300 ;
        RECT 194.700 377.400 196.500 390.300 ;
        RECT 202.800 383.400 204.600 390.300 ;
        RECT 223.800 384.000 225.600 390.300 ;
        RECT 229.800 383.400 231.600 390.300 ;
        RECT 242.400 383.400 244.200 390.300 ;
        RECT 250.500 377.400 252.300 390.300 ;
        RECT 266.400 383.400 268.200 390.300 ;
        RECT 274.500 377.400 276.300 390.300 ;
        RECT 287.400 383.400 289.200 390.300 ;
        RECT 293.400 383.400 295.200 390.300 ;
        RECT 313.800 383.400 315.600 390.300 ;
        RECT 319.800 383.400 321.600 390.300 ;
        RECT 337.800 383.400 339.600 390.300 ;
        RECT 355.800 383.400 357.600 390.300 ;
        RECT 379.800 379.200 381.600 390.300 ;
        RECT 395.400 383.400 397.200 390.300 ;
        RECT 403.500 377.400 405.300 390.300 ;
        RECT 419.400 380.400 421.200 390.300 ;
        RECT 455.400 379.200 457.200 390.300 ;
        RECT 473.400 383.400 475.200 390.300 ;
        RECT 491.700 377.400 493.500 390.300 ;
        RECT 499.800 383.400 501.600 390.300 ;
        RECT 515.400 383.400 517.200 390.300 ;
        RECT 533.700 377.400 535.500 390.300 ;
        RECT 541.800 383.400 543.600 390.300 ;
        RECT 560.400 383.400 562.200 390.300 ;
        RECT 568.500 377.400 570.300 390.300 ;
        RECT 586.800 383.400 588.600 390.300 ;
        RECT 602.400 379.200 604.200 390.300 ;
        RECT 623.700 377.400 625.500 390.300 ;
        RECT 631.800 383.400 633.600 390.300 ;
        RECT 655.800 377.400 657.600 390.300 ;
        RECT 668.400 383.400 670.200 390.300 ;
        RECT 674.400 383.400 676.200 390.300 ;
        RECT 689.400 383.400 691.200 390.300 ;
        RECT 697.500 377.400 699.300 390.300 ;
        RECT 718.800 377.400 720.600 390.300 ;
        RECT 730.800 383.400 732.600 390.300 ;
        RECT 736.800 383.400 738.600 390.300 ;
        RECT 754.800 384.000 756.600 390.300 ;
        RECT 760.800 383.400 762.600 390.300 ;
        RECT 773.400 383.400 775.200 390.300 ;
        RECT 794.400 383.400 796.200 390.300 ;
        RECT 802.500 377.400 804.300 390.300 ;
        RECT 819.900 377.400 821.700 390.300 ;
        RECT 839.400 383.400 841.200 390.300 ;
        RECT 847.500 377.400 849.300 390.300 ;
        RECT 860.400 383.400 862.200 390.300 ;
        RECT 868.500 377.400 870.300 390.300 ;
        RECT 889.800 377.400 891.600 390.300 ;
        RECT 902.400 383.400 904.200 390.300 ;
        RECT 908.400 383.400 910.200 390.300 ;
        RECT 14.400 314.700 16.200 321.600 ;
        RECT 22.500 314.700 24.300 327.600 ;
        RECT 40.800 314.700 42.600 321.000 ;
        RECT 46.800 314.700 48.600 321.600 ;
        RECT 62.400 314.700 64.200 321.600 ;
        RECT 70.500 314.700 72.300 327.600 ;
        RECT 83.400 314.700 85.200 321.600 ;
        RECT 89.400 314.700 91.200 321.000 ;
        RECT 107.700 314.700 109.500 327.600 ;
        RECT 115.800 314.700 117.600 321.600 ;
        RECT 136.800 314.700 138.600 321.600 ;
        RECT 154.800 314.700 156.600 321.000 ;
        RECT 160.800 314.700 162.600 321.600 ;
        RECT 176.400 314.700 178.200 325.500 ;
        RECT 200.400 314.700 202.200 325.500 ;
        RECT 221.400 314.700 223.200 321.600 ;
        RECT 227.400 314.700 229.200 321.600 ;
        RECT 250.800 314.700 252.600 327.600 ;
        RECT 271.800 314.700 273.600 325.500 ;
        RECT 289.800 314.700 291.600 321.600 ;
        RECT 295.800 314.700 297.600 321.600 ;
        RECT 310.800 314.700 312.600 321.600 ;
        RECT 316.800 314.700 318.600 321.600 ;
        RECT 337.800 314.700 339.600 327.600 ;
        RECT 350.400 314.700 352.200 327.600 ;
        RECT 373.800 314.700 375.600 321.600 ;
        RECT 379.800 314.700 381.600 321.600 ;
        RECT 397.800 314.700 399.600 321.600 ;
        RECT 418.800 314.700 420.600 321.600 ;
        RECT 434.400 314.700 436.200 321.600 ;
        RECT 460.800 314.700 462.600 327.600 ;
        RECT 470.700 314.700 472.500 327.600 ;
        RECT 478.800 314.700 480.600 321.600 ;
        RECT 499.800 314.700 501.600 321.600 ;
        RECT 520.800 314.700 522.600 321.600 ;
        RECT 541.800 314.700 543.600 321.600 ;
        RECT 548.550 314.700 550.350 318.600 ;
        RECT 557.250 314.700 559.050 321.600 ;
        RECT 563.850 314.700 565.650 321.600 ;
        RECT 574.050 314.700 575.850 321.600 ;
        RECT 590.400 314.700 592.200 325.500 ;
        RECT 614.400 314.700 616.200 321.600 ;
        RECT 622.500 314.700 624.300 327.600 ;
        RECT 643.800 314.700 645.600 327.600 ;
        RECT 664.800 314.700 666.600 325.500 ;
        RECT 674.550 314.700 676.350 318.600 ;
        RECT 683.250 314.700 685.050 321.600 ;
        RECT 689.850 314.700 691.650 321.600 ;
        RECT 700.050 314.700 701.850 321.600 ;
        RECT 716.400 314.700 718.200 327.600 ;
        RECT 737.400 314.700 739.200 321.600 ;
        RECT 752.400 314.700 754.200 321.600 ;
        RECT 778.800 314.700 780.600 327.600 ;
        RECT 791.400 314.700 793.200 321.600 ;
        RECT 797.400 314.700 799.200 321.600 ;
        RECT 812.400 314.700 814.200 321.600 ;
        RECT 818.400 314.700 820.200 321.000 ;
        RECT 833.700 314.700 835.500 327.600 ;
        RECT 841.800 314.700 843.600 321.600 ;
        RECT 862.800 314.700 864.600 321.600 ;
        RECT 875.400 314.700 877.200 321.600 ;
        RECT 890.400 314.700 892.200 321.600 ;
        RECT 896.400 314.700 898.200 321.600 ;
        RECT -9.450 312.300 920.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT 16.800 306.000 18.600 312.300 ;
        RECT 22.800 305.400 24.600 312.300 ;
        RECT 40.800 301.200 42.600 312.300 ;
        RECT 61.800 301.200 63.600 312.300 ;
        RECT 74.400 305.400 76.200 312.300 ;
        RECT 80.400 306.000 82.200 312.300 ;
        RECT 98.400 305.400 100.200 312.300 ;
        RECT 104.400 306.000 106.200 312.300 ;
        RECT 122.400 305.400 124.200 312.300 ;
        RECT 130.500 299.400 132.300 312.300 ;
        RECT 151.800 301.200 153.600 312.300 ;
        RECT 167.400 305.400 169.200 312.300 ;
        RECT 175.500 299.400 177.300 312.300 ;
        RECT 191.400 305.400 193.200 312.300 ;
        RECT 199.500 299.400 201.300 312.300 ;
        RECT 211.800 305.400 213.600 312.300 ;
        RECT 217.800 305.400 219.600 312.300 ;
        RECT 230.400 305.400 232.200 312.300 ;
        RECT 236.400 305.400 238.200 312.300 ;
        RECT 248.400 305.400 250.200 312.300 ;
        RECT 254.400 305.400 256.200 312.300 ;
        RECT 266.700 299.400 268.500 312.300 ;
        RECT 274.800 305.400 276.600 312.300 ;
        RECT 290.400 305.400 292.200 312.300 ;
        RECT 296.400 305.400 298.200 312.300 ;
        RECT 316.800 305.400 318.600 312.300 ;
        RECT 322.800 305.400 324.600 312.300 ;
        RECT 335.400 305.400 337.200 312.300 ;
        RECT 341.400 305.400 343.200 312.300 ;
        RECT 361.800 306.000 363.600 312.300 ;
        RECT 367.800 305.400 369.600 312.300 ;
        RECT 380.400 305.400 382.200 312.300 ;
        RECT 386.400 305.400 388.200 312.300 ;
        RECT 400.800 305.400 402.600 312.300 ;
        RECT 406.800 305.400 408.600 312.300 ;
        RECT 422.400 305.400 424.200 312.300 ;
        RECT 430.500 299.400 432.300 312.300 ;
        RECT 445.800 305.400 447.600 312.300 ;
        RECT 458.700 299.400 460.500 312.300 ;
        RECT 466.800 305.400 468.600 312.300 ;
        RECT 482.400 305.400 484.200 312.300 ;
        RECT 488.400 305.400 490.200 312.300 ;
        RECT 505.800 305.400 507.600 312.300 ;
        RECT 511.800 305.400 513.600 312.300 ;
        RECT 535.800 301.500 537.600 312.300 ;
        RECT 556.800 305.400 558.600 312.300 ;
        RECT 569.400 305.400 571.200 312.300 ;
        RECT 577.500 299.400 579.300 312.300 ;
        RECT 592.800 305.400 594.600 312.300 ;
        RECT 598.800 305.400 600.600 312.300 ;
        RECT 619.800 301.200 621.600 312.300 ;
        RECT 635.400 305.400 637.200 312.300 ;
        RECT 643.500 299.400 645.300 312.300 ;
        RECT 656.700 299.400 658.500 312.300 ;
        RECT 664.800 305.400 666.600 312.300 ;
        RECT 680.400 305.400 682.200 312.300 ;
        RECT 686.400 305.400 688.200 312.300 ;
        RECT 706.800 305.400 708.600 312.300 ;
        RECT 719.400 305.400 721.200 312.300 ;
        RECT 725.400 305.400 727.200 312.300 ;
        RECT 740.400 299.400 742.200 312.300 ;
        RECT 746.400 299.400 748.200 312.300 ;
        RECT 766.800 305.400 768.600 312.300 ;
        RECT 776.400 305.400 778.200 312.300 ;
        RECT 797.400 301.200 799.200 312.300 ;
        RECT 821.400 301.500 823.200 312.300 ;
        RECT 845.700 299.400 847.500 312.300 ;
        RECT 853.800 305.400 855.600 312.300 ;
        RECT 869.400 305.400 871.200 312.300 ;
        RECT 875.400 305.400 877.200 312.300 ;
        RECT 890.700 299.400 892.500 312.300 ;
        RECT 898.800 305.400 900.600 312.300 ;
        RECT 14.400 236.700 16.200 243.600 ;
        RECT 22.500 236.700 24.300 249.600 ;
        RECT 35.400 236.700 37.200 243.600 ;
        RECT 43.500 236.700 45.300 249.600 ;
        RECT 61.800 236.700 63.600 243.000 ;
        RECT 67.800 236.700 69.600 243.600 ;
        RECT 85.800 236.700 87.600 243.600 ;
        RECT 106.800 236.700 108.600 247.500 ;
        RECT 119.400 236.700 121.200 243.600 ;
        RECT 125.400 236.700 127.200 243.600 ;
        RECT 145.800 236.700 147.600 243.000 ;
        RECT 151.800 236.700 153.600 243.600 ;
        RECT 161.400 236.700 163.200 243.600 ;
        RECT 184.800 236.700 186.600 243.000 ;
        RECT 190.800 236.700 192.600 243.600 ;
        RECT 208.800 236.700 210.600 243.600 ;
        RECT 226.800 236.700 228.600 243.000 ;
        RECT 232.800 236.700 234.600 243.600 ;
        RECT 250.800 236.700 252.600 243.000 ;
        RECT 256.800 236.700 258.600 243.600 ;
        RECT 280.800 236.700 282.600 247.500 ;
        RECT 299.400 236.700 301.200 243.600 ;
        RECT 307.500 236.700 309.300 249.600 ;
        RECT 320.700 236.700 322.500 249.600 ;
        RECT 328.800 236.700 330.600 243.600 ;
        RECT 341.400 236.700 343.200 243.600 ;
        RECT 347.400 236.700 349.200 243.600 ;
        RECT 367.800 236.700 369.600 249.600 ;
        RECT 380.400 236.700 382.200 243.600 ;
        RECT 386.400 236.700 388.200 243.600 ;
        RECT 403.800 236.700 405.600 243.600 ;
        RECT 409.800 236.700 411.600 243.600 ;
        RECT 422.400 236.700 424.200 243.600 ;
        RECT 428.400 236.700 430.200 243.600 ;
        RECT 448.800 236.700 450.600 243.600 ;
        RECT 461.400 236.700 463.200 249.600 ;
        RECT 487.800 236.700 489.600 243.600 ;
        RECT 493.800 236.700 495.600 243.600 ;
        RECT 510.900 236.700 512.700 249.600 ;
        RECT 527.400 236.700 529.200 243.600 ;
        RECT 533.400 236.700 535.200 243.600 ;
        RECT 552.900 236.700 554.700 249.600 ;
        RECT 572.400 236.700 574.200 243.600 ;
        RECT 578.400 236.700 580.200 243.600 ;
        RECT 590.400 236.700 592.200 243.600 ;
        RECT 605.700 236.700 607.500 249.600 ;
        RECT 613.800 236.700 615.600 243.600 ;
        RECT 630.900 236.700 632.700 249.600 ;
        RECT 650.400 236.700 652.200 243.600 ;
        RECT 656.400 236.700 658.200 243.600 ;
        RECT 676.800 236.700 678.600 249.600 ;
        RECT 689.400 236.700 691.200 243.600 ;
        RECT 695.400 236.700 697.200 243.600 ;
        RECT 710.700 236.700 712.500 249.600 ;
        RECT 718.800 236.700 720.600 243.600 ;
        RECT 728.550 236.700 730.350 240.600 ;
        RECT 737.250 236.700 739.050 243.600 ;
        RECT 743.850 236.700 745.650 243.600 ;
        RECT 754.050 236.700 755.850 243.600 ;
        RECT 772.800 236.700 774.600 243.600 ;
        RECT 778.800 236.700 780.600 243.600 ;
        RECT 796.800 236.700 798.600 249.600 ;
        RECT 809.400 236.700 811.200 243.600 ;
        RECT 832.800 236.700 834.600 249.600 ;
        RECT 838.200 236.700 840.000 243.600 ;
        RECT 844.800 236.700 846.600 243.600 ;
        RECT 850.800 241.050 852.600 243.600 ;
        RECT 850.650 238.950 852.750 241.050 ;
        RECT 850.800 236.700 852.600 238.950 ;
        RECT 856.800 236.700 858.600 243.600 ;
        RECT 873.000 236.700 874.800 243.600 ;
        RECT 879.900 236.700 881.700 243.600 ;
        RECT 892.500 236.700 894.300 242.400 ;
        RECT 898.500 236.700 900.300 243.600 ;
        RECT 904.500 236.700 906.300 243.600 ;
        RECT -9.450 234.300 920.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT 16.800 228.000 18.600 234.300 ;
        RECT 22.800 227.400 24.600 234.300 ;
        RECT 35.400 223.200 37.200 234.300 ;
        RECT 58.800 227.400 60.600 234.300 ;
        RECT 64.800 227.400 66.600 234.300 ;
        RECT 77.400 227.400 79.200 234.300 ;
        RECT 83.400 227.400 85.200 234.300 ;
        RECT 98.400 227.400 100.200 234.300 ;
        RECT 106.500 221.400 108.300 234.300 ;
        RECT 119.400 221.400 121.200 234.300 ;
        RECT 140.700 221.400 142.500 234.300 ;
        RECT 148.800 227.400 150.600 234.300 ;
        RECT 172.800 223.200 174.600 234.300 ;
        RECT 185.400 227.400 187.200 234.300 ;
        RECT 191.400 228.000 193.200 234.300 ;
        RECT 211.800 227.400 213.600 234.300 ;
        RECT 217.800 227.400 219.600 234.300 ;
        RECT 233.400 227.400 235.200 234.300 ;
        RECT 241.500 221.400 243.300 234.300 ;
        RECT 259.800 227.400 261.600 234.300 ;
        RECT 272.700 221.400 274.500 234.300 ;
        RECT 280.800 227.400 282.600 234.300 ;
        RECT 301.800 228.000 303.600 234.300 ;
        RECT 307.800 227.400 309.600 234.300 ;
        RECT 317.700 221.400 319.500 234.300 ;
        RECT 325.800 227.400 327.600 234.300 ;
        RECT 338.400 227.400 340.200 234.300 ;
        RECT 356.400 227.400 358.200 234.300 ;
        RECT 362.400 227.400 364.200 234.300 ;
        RECT 379.800 227.400 381.600 234.300 ;
        RECT 385.800 227.400 387.600 234.300 ;
        RECT 395.400 227.400 397.200 234.300 ;
        RECT 401.400 227.400 403.200 234.300 ;
        RECT 419.400 227.400 421.200 234.300 ;
        RECT 427.500 221.400 429.300 234.300 ;
        RECT 440.400 227.400 442.200 234.300 ;
        RECT 448.500 221.400 450.300 234.300 ;
        RECT 458.700 221.400 460.500 234.300 ;
        RECT 466.800 227.400 468.600 234.300 ;
        RECT 479.400 227.400 481.200 234.300 ;
        RECT 485.400 227.400 487.200 234.300 ;
        RECT 503.400 221.400 505.200 234.300 ;
        RECT 527.400 227.400 529.200 234.300 ;
        RECT 535.500 221.400 537.300 234.300 ;
        RECT 548.400 227.400 550.200 234.300 ;
        RECT 554.400 227.400 556.200 234.300 ;
        RECT 569.400 227.400 571.200 234.300 ;
        RECT 587.700 221.400 589.500 234.300 ;
        RECT 595.800 227.400 597.600 234.300 ;
        RECT 615.900 221.400 617.700 234.300 ;
        RECT 637.800 228.000 639.600 234.300 ;
        RECT 643.800 227.400 645.600 234.300 ;
        RECT 659.400 223.200 661.200 234.300 ;
        RECT 677.700 221.400 679.500 234.300 ;
        RECT 685.800 227.400 687.600 234.300 ;
        RECT 701.700 221.400 703.500 234.300 ;
        RECT 709.800 227.400 711.600 234.300 ;
        RECT 728.400 227.400 730.200 234.300 ;
        RECT 736.500 221.400 738.300 234.300 ;
        RECT 757.800 221.400 759.600 234.300 ;
        RECT 769.800 227.400 771.600 234.300 ;
        RECT 775.800 227.400 777.600 234.300 ;
        RECT 793.800 227.400 795.600 234.300 ;
        RECT 806.400 227.400 808.200 234.300 ;
        RECT 814.500 221.400 816.300 234.300 ;
        RECT 820.200 227.400 822.000 234.300 ;
        RECT 826.800 227.400 828.600 234.300 ;
        RECT 832.800 227.400 834.600 234.300 ;
        RECT 838.800 227.400 840.600 234.300 ;
        RECT 855.000 227.400 856.800 234.300 ;
        RECT 861.900 227.400 863.700 234.300 ;
        RECT 874.500 228.600 876.300 234.300 ;
        RECT 880.500 227.400 882.300 234.300 ;
        RECT 886.500 229.650 888.300 234.300 ;
        RECT 886.500 227.550 889.050 229.650 ;
        RECT 886.500 227.400 888.300 227.550 ;
        RECT 904.800 227.400 906.600 234.300 ;
        RECT 14.400 158.700 16.200 165.600 ;
        RECT 22.500 158.700 24.300 171.600 ;
        RECT 34.800 158.700 36.600 165.600 ;
        RECT 40.800 158.700 42.600 165.600 ;
        RECT 58.800 158.700 60.600 165.000 ;
        RECT 64.800 158.700 66.600 165.600 ;
        RECT 74.400 158.700 76.200 165.600 ;
        RECT 92.400 158.700 94.200 165.600 ;
        RECT 98.400 158.700 100.200 165.000 ;
        RECT 118.800 158.700 120.600 165.000 ;
        RECT 124.800 158.700 126.600 165.600 ;
        RECT 137.700 158.700 139.500 171.600 ;
        RECT 145.800 158.700 147.600 165.600 ;
        RECT 169.800 158.700 171.600 169.800 ;
        RECT 185.400 158.700 187.200 165.600 ;
        RECT 191.400 158.700 193.200 165.000 ;
        RECT 211.800 158.700 213.600 165.600 ;
        RECT 217.800 158.700 219.600 165.600 ;
        RECT 227.400 158.700 229.200 165.600 ;
        RECT 233.400 158.700 235.200 165.600 ;
        RECT 259.800 158.700 261.600 169.800 ;
        RECT 277.800 158.700 279.600 165.600 ;
        RECT 298.800 158.700 300.600 171.600 ;
        RECT 308.700 158.700 310.500 171.600 ;
        RECT 316.800 158.700 318.600 165.600 ;
        RECT 329.700 158.700 331.500 171.600 ;
        RECT 337.800 158.700 339.600 165.600 ;
        RECT 358.800 158.700 360.600 165.000 ;
        RECT 364.800 158.700 366.600 165.600 ;
        RECT 377.700 158.700 379.500 171.600 ;
        RECT 385.800 158.700 387.600 165.600 ;
        RECT 401.400 158.700 403.200 171.600 ;
        RECT 427.800 158.700 429.600 169.800 ;
        RECT 443.400 158.700 445.200 165.600 ;
        RECT 458.400 158.700 460.200 165.600 ;
        RECT 464.400 158.700 466.200 165.000 ;
        RECT 482.400 158.700 484.200 165.600 ;
        RECT 488.400 158.700 490.200 165.000 ;
        RECT 514.800 158.700 516.600 169.800 ;
        RECT 530.700 158.700 532.500 171.600 ;
        RECT 538.800 158.700 540.600 165.600 ;
        RECT 551.400 158.700 553.200 165.600 ;
        RECT 569.400 158.700 571.200 165.600 ;
        RECT 575.400 158.700 577.200 165.000 ;
        RECT 593.400 158.700 595.200 169.800 ;
        RECT 614.400 158.700 616.200 165.600 ;
        RECT 620.400 158.700 622.200 165.000 ;
        RECT 637.800 158.700 639.600 165.600 ;
        RECT 643.800 158.700 645.600 165.600 ;
        RECT 658.800 158.700 660.600 165.600 ;
        RECT 664.800 158.700 666.600 165.600 ;
        RECT 677.400 158.700 679.200 165.600 ;
        RECT 697.800 158.700 699.600 165.600 ;
        RECT 707.550 158.700 709.350 162.600 ;
        RECT 716.250 158.700 718.050 165.600 ;
        RECT 722.850 158.700 724.650 165.600 ;
        RECT 733.050 158.700 734.850 165.600 ;
        RECT 751.800 158.700 753.600 171.600 ;
        RECT 757.800 158.700 759.600 171.600 ;
        RECT 763.800 158.700 765.600 171.600 ;
        RECT 769.800 158.700 771.600 171.600 ;
        RECT 775.800 158.700 777.600 171.600 ;
        RECT 791.400 158.700 793.200 169.800 ;
        RECT 812.400 158.700 814.200 165.600 ;
        RECT 830.400 158.700 832.200 171.600 ;
        RECT 841.200 158.700 843.000 165.600 ;
        RECT 847.800 158.700 849.600 165.600 ;
        RECT 853.800 158.700 855.600 165.600 ;
        RECT 859.800 158.700 861.600 165.600 ;
        RECT 876.000 158.700 877.800 165.600 ;
        RECT 882.900 158.700 884.700 165.600 ;
        RECT 895.500 158.700 897.300 164.400 ;
        RECT 901.350 163.950 903.450 166.050 ;
        RECT 901.500 158.700 903.300 163.950 ;
        RECT 907.500 158.700 909.300 165.600 ;
        RECT -9.450 156.300 920.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT 19.800 145.200 21.600 156.300 ;
        RECT 32.400 149.400 34.200 156.300 ;
        RECT 38.400 150.000 40.200 156.300 ;
        RECT 59.400 145.200 61.200 156.300 ;
        RECT 77.400 149.400 79.200 156.300 ;
        RECT 83.400 150.000 85.200 156.300 ;
        RECT 103.800 149.400 105.600 156.300 ;
        RECT 109.800 149.400 111.600 156.300 ;
        RECT 130.800 145.200 132.600 156.300 ;
        RECT 151.800 150.000 153.600 156.300 ;
        RECT 157.800 149.400 159.600 156.300 ;
        RECT 170.700 143.400 172.500 156.300 ;
        RECT 178.800 149.400 180.600 156.300 ;
        RECT 194.400 149.400 196.200 156.300 ;
        RECT 200.400 150.000 202.200 156.300 ;
        RECT 223.800 150.000 225.600 156.300 ;
        RECT 229.800 149.400 231.600 156.300 ;
        RECT 247.800 149.400 249.600 156.300 ;
        RECT 260.700 143.400 262.500 156.300 ;
        RECT 268.800 149.400 270.600 156.300 ;
        RECT 284.400 149.400 286.200 156.300 ;
        RECT 290.400 150.000 292.200 156.300 ;
        RECT 308.700 143.400 310.500 156.300 ;
        RECT 316.800 149.400 318.600 156.300 ;
        RECT 334.800 149.400 336.600 156.300 ;
        RECT 340.800 149.400 342.600 156.300 ;
        RECT 350.400 149.400 352.200 156.300 ;
        RECT 356.400 149.400 358.200 156.300 ;
        RECT 379.800 145.200 381.600 156.300 ;
        RECT 395.400 149.400 397.200 156.300 ;
        RECT 401.400 150.000 403.200 156.300 ;
        RECT 419.400 149.400 421.200 156.300 ;
        RECT 425.400 149.400 427.200 156.300 ;
        RECT 440.700 143.400 442.500 156.300 ;
        RECT 448.800 149.400 450.600 156.300 ;
        RECT 464.400 149.400 466.200 156.300 ;
        RECT 490.800 145.200 492.600 156.300 ;
        RECT 503.400 149.400 505.200 156.300 ;
        RECT 509.400 150.000 511.200 156.300 ;
        RECT 532.800 150.000 534.600 156.300 ;
        RECT 538.800 149.400 540.600 156.300 ;
        RECT 554.400 145.200 556.200 156.300 ;
        RECT 575.400 149.400 577.200 156.300 ;
        RECT 581.400 150.000 583.200 156.300 ;
        RECT 601.800 149.400 603.600 156.300 ;
        RECT 614.700 143.400 616.500 156.300 ;
        RECT 622.800 149.400 624.600 156.300 ;
        RECT 635.700 143.400 637.500 156.300 ;
        RECT 643.800 149.400 645.600 156.300 ;
        RECT 659.400 149.400 661.200 156.300 ;
        RECT 677.400 149.400 679.200 156.300 ;
        RECT 683.400 150.000 685.200 156.300 ;
        RECT 701.400 149.400 703.200 156.300 ;
        RECT 707.400 149.400 709.200 156.300 ;
        RECT 722.700 143.400 724.500 156.300 ;
        RECT 730.800 149.400 732.600 156.300 ;
        RECT 743.400 149.400 745.200 156.300 ;
        RECT 749.400 149.400 751.200 156.300 ;
        RECT 767.400 149.400 769.200 156.300 ;
        RECT 775.500 143.400 777.300 156.300 ;
        RECT 791.400 145.200 793.200 156.300 ;
        RECT 809.400 149.400 811.200 156.300 ;
        RECT 815.400 149.400 817.200 156.300 ;
        RECT 833.400 149.400 835.200 156.300 ;
        RECT 841.500 143.400 843.300 156.300 ;
        RECT 854.400 143.400 856.200 156.300 ;
        RECT 860.400 143.400 862.200 156.300 ;
        RECT 877.800 143.400 879.600 156.300 ;
        RECT 883.800 143.400 885.600 156.300 ;
        RECT 889.800 143.400 891.600 156.300 ;
        RECT 895.800 143.400 897.600 156.300 ;
        RECT 901.800 143.400 903.600 156.300 ;
        RECT 14.400 80.700 16.200 87.600 ;
        RECT 22.500 80.700 24.300 93.600 ;
        RECT 40.800 80.700 42.600 87.000 ;
        RECT 46.800 80.700 48.600 87.600 ;
        RECT 59.700 80.700 61.500 93.600 ;
        RECT 67.800 80.700 69.600 87.600 ;
        RECT 83.400 80.700 85.200 87.600 ;
        RECT 89.400 80.700 91.200 87.000 ;
        RECT 110.400 80.700 112.200 87.600 ;
        RECT 118.500 80.700 120.300 93.600 ;
        RECT 139.800 80.700 141.600 91.800 ;
        RECT 155.400 80.700 157.200 87.600 ;
        RECT 161.400 80.700 163.200 87.000 ;
        RECT 181.800 80.700 183.600 87.000 ;
        RECT 187.800 80.700 189.600 87.600 ;
        RECT 203.400 80.700 205.200 91.800 ;
        RECT 232.800 80.700 234.600 91.800 ;
        RECT 245.400 80.700 247.200 87.600 ;
        RECT 251.400 80.700 253.200 87.000 ;
        RECT 274.800 80.700 276.600 91.800 ;
        RECT 290.400 80.700 292.200 87.600 ;
        RECT 298.500 80.700 300.300 93.600 ;
        RECT 314.400 80.700 316.200 87.600 ;
        RECT 322.500 80.700 324.300 93.600 ;
        RECT 340.800 80.700 342.600 87.000 ;
        RECT 346.800 80.700 348.600 87.600 ;
        RECT 359.700 80.700 361.500 93.600 ;
        RECT 367.800 80.700 369.600 87.600 ;
        RECT 380.400 80.700 382.200 87.600 ;
        RECT 386.400 80.700 388.200 87.000 ;
        RECT 404.400 80.700 406.200 87.600 ;
        RECT 410.400 80.700 412.200 87.000 ;
        RECT 428.400 80.700 430.200 87.600 ;
        RECT 434.400 80.700 436.200 87.600 ;
        RECT 463.800 80.700 465.600 91.500 ;
        RECT 487.800 80.700 489.600 91.800 ;
        RECT 500.400 80.700 502.200 87.600 ;
        RECT 506.400 80.700 508.200 87.000 ;
        RECT 524.400 80.700 526.200 87.600 ;
        RECT 532.500 80.700 534.300 93.600 ;
        RECT 545.700 80.700 547.500 93.600 ;
        RECT 553.800 80.700 555.600 87.600 ;
        RECT 574.800 80.700 576.600 87.000 ;
        RECT 580.800 80.700 582.600 87.600 ;
        RECT 596.400 80.700 598.200 91.800 ;
        RECT 637.800 80.700 639.600 90.600 ;
        RECT 653.700 80.700 655.500 93.600 ;
        RECT 661.800 80.700 663.600 87.600 ;
        RECT 674.400 80.700 676.200 87.600 ;
        RECT 692.400 80.700 694.200 87.600 ;
        RECT 698.400 80.700 700.200 87.600 ;
        RECT 721.800 80.700 723.600 91.800 ;
        RECT 740.400 80.700 742.200 91.500 ;
        RECT 769.800 80.700 771.600 91.800 ;
        RECT 785.400 80.700 787.200 91.800 ;
        RECT 814.800 80.700 816.600 91.500 ;
        RECT 833.400 80.700 835.200 91.800 ;
        RECT 862.800 80.700 864.600 91.500 ;
        RECT 878.400 80.700 880.200 87.600 ;
        RECT 896.400 80.700 898.200 87.600 ;
        RECT -9.450 78.300 920.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT 16.800 72.000 18.600 78.300 ;
        RECT 22.800 71.400 24.600 78.300 ;
        RECT 35.400 67.200 37.200 78.300 ;
        RECT 64.800 67.200 66.600 78.300 ;
        RECT 77.400 71.400 79.200 78.300 ;
        RECT 83.400 72.000 85.200 78.300 ;
        RECT 104.400 71.400 106.200 78.300 ;
        RECT 112.500 65.400 114.300 78.300 ;
        RECT 130.800 67.200 132.600 78.300 ;
        RECT 149.400 71.400 151.200 78.300 ;
        RECT 157.500 65.400 159.300 78.300 ;
        RECT 170.400 71.400 172.200 78.300 ;
        RECT 178.500 65.400 180.300 78.300 ;
        RECT 188.700 65.400 190.500 78.300 ;
        RECT 196.800 71.400 198.600 78.300 ;
        RECT 215.400 67.500 217.200 78.300 ;
        RECT 224.100 67.500 226.200 78.300 ;
        RECT 242.400 71.400 244.200 78.300 ;
        RECT 248.400 71.400 250.200 78.300 ;
        RECT 274.800 67.500 276.600 78.300 ;
        RECT 290.400 71.400 292.200 78.300 ;
        RECT 296.400 72.000 298.200 78.300 ;
        RECT 316.800 72.000 318.600 78.300 ;
        RECT 322.800 71.400 324.600 78.300 ;
        RECT 338.400 67.200 340.200 78.300 ;
        RECT 362.400 71.400 364.200 78.300 ;
        RECT 370.500 65.400 372.300 78.300 ;
        RECT 383.400 71.400 385.200 78.300 ;
        RECT 406.800 72.000 408.600 78.300 ;
        RECT 412.800 71.400 414.600 78.300 ;
        RECT 425.400 71.400 427.200 78.300 ;
        RECT 431.400 72.000 433.200 78.300 ;
        RECT 452.400 71.400 454.200 78.300 ;
        RECT 460.500 65.400 462.300 78.300 ;
        RECT 470.700 65.400 472.500 78.300 ;
        RECT 478.800 71.400 480.600 78.300 ;
        RECT 496.800 71.400 498.600 78.300 ;
        RECT 506.400 71.400 508.200 78.300 ;
        RECT 512.400 72.000 514.200 78.300 ;
        RECT 530.400 71.400 532.200 78.300 ;
        RECT 536.400 72.000 538.200 78.300 ;
        RECT 551.400 71.400 553.200 78.300 ;
        RECT 571.800 72.000 573.600 78.300 ;
        RECT 577.800 71.400 579.600 78.300 ;
        RECT 593.400 67.200 595.200 78.300 ;
        RECT 614.400 71.400 616.200 78.300 ;
        RECT 629.700 65.400 631.500 78.300 ;
        RECT 637.800 71.400 639.600 78.300 ;
        RECT 661.800 67.500 663.600 78.300 ;
        RECT 682.800 71.400 684.600 78.300 ;
        RECT 689.550 74.400 691.350 78.300 ;
        RECT 698.250 71.400 700.050 78.300 ;
        RECT 704.850 71.400 706.650 78.300 ;
        RECT 715.050 71.400 716.850 78.300 ;
        RECT 736.800 71.400 738.600 78.300 ;
        RECT 760.800 67.500 762.600 78.300 ;
        RECT 781.800 71.400 783.600 78.300 ;
        RECT 788.550 74.400 790.350 78.300 ;
        RECT 797.250 71.400 799.050 78.300 ;
        RECT 803.850 71.400 805.650 78.300 ;
        RECT 814.050 71.400 815.850 78.300 ;
        RECT 825.150 71.400 826.950 78.300 ;
        RECT 835.350 71.400 837.150 78.300 ;
        RECT 841.950 71.400 843.750 78.300 ;
        RECT 850.650 74.400 852.450 78.300 ;
        RECT 863.400 71.400 865.200 78.300 ;
        RECT 869.400 72.000 871.200 78.300 ;
        RECT 887.700 65.400 889.500 78.300 ;
        RECT 895.800 71.400 897.600 78.300 ;
        RECT 19.800 2.700 21.600 13.800 ;
        RECT 37.800 2.700 39.600 9.600 ;
        RECT 53.400 2.700 55.200 9.600 ;
        RECT 61.500 2.700 63.300 15.600 ;
        RECT 71.400 2.700 73.200 9.600 ;
        RECT 77.400 2.700 79.200 9.000 ;
        RECT 95.400 2.700 97.200 9.600 ;
        RECT 101.400 2.700 103.200 9.000 ;
        RECT 119.700 2.700 121.500 15.600 ;
        RECT 127.800 2.700 129.600 9.600 ;
        RECT 148.800 2.700 150.600 9.600 ;
        RECT 158.400 2.700 160.200 9.600 ;
        RECT 164.400 2.700 166.200 9.000 ;
        RECT 182.400 2.700 184.200 9.600 ;
        RECT 188.400 2.700 190.200 9.000 ;
        RECT 209.400 2.700 211.200 13.800 ;
        RECT 232.800 2.700 234.600 9.600 ;
        RECT 238.800 2.700 240.600 9.600 ;
        RECT 256.800 2.700 258.600 9.000 ;
        RECT 262.800 2.700 264.600 9.600 ;
        RECT 278.400 2.700 280.200 13.800 ;
        RECT 299.400 2.700 301.200 9.600 ;
        RECT 305.400 2.700 307.200 9.000 ;
        RECT 326.400 2.700 328.200 13.800 ;
        RECT 344.400 2.700 346.200 9.600 ;
        RECT 370.800 2.700 372.600 13.800 ;
        RECT 386.400 2.700 388.200 9.600 ;
        RECT 392.400 2.700 394.200 9.600 ;
        RECT 407.700 2.700 409.500 15.600 ;
        RECT 415.800 2.700 417.600 9.600 ;
        RECT 434.400 2.700 436.200 13.800 ;
        RECT 452.400 2.700 454.200 9.600 ;
        RECT 458.400 2.700 460.200 9.000 ;
        RECT 479.400 2.700 481.200 9.600 ;
        RECT 487.500 2.700 489.300 15.600 ;
        RECT 503.400 2.700 505.200 12.600 ;
        RECT 536.700 2.700 538.500 15.600 ;
        RECT 544.800 2.700 546.600 9.600 ;
        RECT 565.800 2.700 567.600 13.800 ;
        RECT 586.800 2.700 588.900 13.500 ;
        RECT 595.800 2.700 597.600 13.500 ;
        RECT 610.800 2.700 612.600 9.600 ;
        RECT 616.800 2.700 618.600 9.600 ;
        RECT 632.400 2.700 634.200 13.800 ;
        RECT 653.400 2.700 655.200 15.600 ;
        RECT 671.700 2.700 673.500 15.600 ;
        RECT 679.800 2.700 681.600 9.600 ;
        RECT 698.400 2.700 700.200 9.600 ;
        RECT 711.150 2.700 712.950 9.600 ;
        RECT 721.350 2.700 723.150 9.600 ;
        RECT 727.950 2.700 729.750 9.600 ;
        RECT 736.650 2.700 738.450 6.600 ;
        RECT 755.400 2.700 757.200 9.600 ;
        RECT 768.150 2.700 769.950 9.600 ;
        RECT 778.350 2.700 780.150 9.600 ;
        RECT 784.950 2.700 786.750 9.600 ;
        RECT 793.650 2.700 795.450 6.600 ;
        RECT 809.400 2.700 811.200 9.600 ;
        RECT 830.400 2.700 832.200 9.600 ;
        RECT 853.800 2.700 855.600 9.600 ;
        RECT 869.400 2.700 871.200 9.600 ;
        RECT 889.800 2.700 891.600 9.600 ;
        RECT 895.800 2.700 897.600 9.600 ;
        RECT -9.450 0.300 920.400 2.700 ;
      LAYER metal2 ;
        RECT 892.950 258.600 897.000 259.050 ;
        RECT 892.950 256.950 897.600 258.600 ;
        RECT 896.400 256.050 897.600 256.950 ;
        RECT 895.950 253.950 898.050 256.050 ;
        RECT 850.650 250.950 852.750 253.050 ;
        RECT 851.100 241.050 852.300 250.950 ;
        RECT 850.650 238.950 852.750 241.050 ;
        RECT 886.950 228.600 889.050 229.650 ;
        RECT 884.400 227.550 889.050 228.600 ;
        RECT 884.400 227.400 888.600 227.550 ;
        RECT 884.400 217.050 885.600 227.400 ;
        RECT 883.950 214.950 886.050 217.050 ;
        RECT 895.950 180.600 900.000 181.050 ;
        RECT 895.950 178.950 900.600 180.600 ;
        RECT 899.400 178.050 900.600 178.950 ;
        RECT 898.950 175.950 901.050 178.050 ;
        RECT 901.350 169.950 903.450 172.050 ;
        RECT 901.800 166.050 903.000 169.950 ;
        RECT 901.350 163.950 903.450 166.050 ;
      LAYER metal3 ;
        RECT 892.950 258.600 895.050 259.050 ;
        RECT 881.400 257.400 895.050 258.600 ;
        RECT 881.400 255.600 882.600 257.400 ;
        RECT 892.950 256.950 895.050 257.400 ;
        RECT 851.400 255.000 882.600 255.600 ;
        RECT 850.950 254.400 882.600 255.000 ;
        RECT 850.950 253.050 853.050 254.400 ;
        RECT 850.650 252.000 853.050 253.050 ;
        RECT 850.650 250.950 852.750 252.000 ;
        RECT 895.950 178.950 898.050 181.050 ;
        RECT 896.400 171.600 897.600 178.950 ;
        RECT 901.350 171.600 903.450 172.050 ;
        RECT 896.400 170.400 903.600 171.600 ;
        RECT 901.350 169.950 903.450 170.400 ;
    END
  END vdd
  PIN ABCmd_i[7]
    PORT
      LAYER metal1 ;
        RECT 504.000 495.450 508.050 496.050 ;
        RECT 503.550 493.950 508.050 495.450 ;
        RECT 503.550 490.050 504.450 493.950 ;
        RECT 503.550 488.550 508.050 490.050 ;
        RECT 504.000 487.950 508.050 488.550 ;
        RECT 481.950 339.450 486.000 340.050 ;
        RECT 481.950 337.950 486.450 339.450 ;
        RECT 485.550 334.050 486.450 337.950 ;
        RECT 481.950 332.550 486.450 334.050 ;
        RECT 481.950 331.950 486.000 332.550 ;
        RECT 625.950 297.450 628.050 298.050 ;
        RECT 634.950 297.450 637.050 298.050 ;
        RECT 625.950 296.550 637.050 297.450 ;
        RECT 625.950 295.950 628.050 296.550 ;
        RECT 634.950 295.950 637.050 296.550 ;
      LAYER metal2 ;
        RECT 500.400 940.050 501.600 945.600 ;
        RECT 499.950 937.950 502.050 940.050 ;
        RECT 580.950 937.950 583.050 940.050 ;
        RECT 581.400 841.050 582.600 937.950 ;
        RECT 580.950 838.950 583.050 841.050 ;
        RECT 580.950 832.950 583.050 835.050 ;
        RECT 581.400 826.050 582.600 832.950 ;
        RECT 550.950 823.950 553.050 826.050 ;
        RECT 580.950 823.950 583.050 826.050 ;
        RECT 551.400 754.050 552.600 823.950 ;
        RECT 544.950 751.950 547.050 754.050 ;
        RECT 550.950 751.950 553.050 754.050 ;
        RECT 545.400 655.050 546.600 751.950 ;
        RECT 544.950 652.950 547.050 655.050 ;
        RECT 547.950 643.950 550.050 646.050 ;
        RECT 548.400 631.050 549.600 643.950 ;
        RECT 547.950 628.950 550.050 631.050 ;
        RECT 565.950 628.950 568.050 631.050 ;
        RECT 566.400 621.600 567.600 628.950 ;
        RECT 566.400 620.400 570.600 621.600 ;
        RECT 569.400 600.600 570.600 620.400 ;
        RECT 566.400 599.400 570.600 600.600 ;
        RECT 566.400 574.050 567.600 599.400 ;
        RECT 565.950 571.950 568.050 574.050 ;
        RECT 523.950 565.950 526.050 568.050 ;
        RECT 524.400 544.050 525.600 565.950 ;
        RECT 505.950 541.950 508.050 544.050 ;
        RECT 523.950 541.950 526.050 544.050 ;
        RECT 506.400 529.200 507.600 541.950 ;
        RECT 505.950 527.100 508.050 529.200 ;
        RECT 506.400 526.050 507.600 527.100 ;
        RECT 505.950 523.950 508.050 526.050 ;
        RECT 505.950 517.950 508.050 520.050 ;
        RECT 506.400 496.050 507.600 517.950 ;
        RECT 811.950 514.950 814.050 517.050 ;
        RECT 847.950 514.950 850.050 517.050 ;
        RECT 505.950 493.950 508.050 496.050 ;
        RECT 754.950 494.100 757.050 496.200 ;
        RECT 755.400 493.050 756.600 494.100 ;
        RECT 772.950 493.800 775.050 495.900 ;
        RECT 754.950 490.950 757.050 493.050 ;
        RECT 505.950 487.950 508.050 490.050 ;
        RECT 506.400 481.050 507.600 487.950 ;
        RECT 505.950 478.950 508.050 481.050 ;
        RECT 514.950 478.950 517.050 481.050 ;
        RECT 515.400 418.050 516.600 478.950 ;
        RECT 773.400 463.050 774.600 493.800 ;
        RECT 812.400 463.050 813.600 514.950 ;
        RECT 848.400 496.200 849.600 514.950 ;
        RECT 847.950 494.100 850.050 496.200 ;
        RECT 859.950 494.100 862.050 496.200 ;
        RECT 860.400 493.050 861.600 494.100 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 772.950 462.600 775.050 463.050 ;
        RECT 772.950 461.400 777.600 462.600 ;
        RECT 772.950 460.950 775.050 461.400 ;
        RECT 776.400 427.050 777.600 461.400 ;
        RECT 811.950 460.950 814.050 463.050 ;
        RECT 835.950 460.950 838.050 463.050 ;
        RECT 836.400 448.050 837.600 460.950 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 775.950 424.950 778.050 427.050 ;
        RECT 514.950 415.950 517.050 418.050 ;
        RECT 694.950 416.100 697.050 418.200 ;
        RECT 695.400 415.050 696.600 416.100 ;
        RECT 526.950 412.950 529.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 508.950 409.950 511.050 412.050 ;
        RECT 527.400 411.900 528.600 412.950 ;
        RECT 481.950 385.950 484.050 388.050 ;
        RECT 496.950 385.950 499.050 388.050 ;
        RECT 482.400 340.050 483.600 385.950 ;
        RECT 497.400 381.600 498.600 385.950 ;
        RECT 497.400 380.400 501.600 381.600 ;
        RECT 500.400 373.200 501.600 380.400 ;
        RECT 509.400 373.200 510.600 409.950 ;
        RECT 526.950 409.800 529.050 411.900 ;
        RECT 553.950 409.800 556.050 411.900 ;
        RECT 664.950 409.950 667.050 412.050 ;
        RECT 680.400 411.900 681.600 412.950 ;
        RECT 554.400 397.050 555.600 409.800 ;
        RECT 665.400 397.050 666.600 409.950 ;
        RECT 679.950 409.800 682.050 411.900 ;
        RECT 553.950 394.950 556.050 397.050 ;
        RECT 664.950 394.950 667.050 397.050 ;
        RECT 680.400 388.050 681.600 409.800 ;
        RECT 679.950 385.950 682.050 388.050 ;
        RECT 703.950 385.950 706.050 388.050 ;
        RECT 499.950 371.100 502.050 373.200 ;
        RECT 508.950 371.100 511.050 373.200 ;
        RECT 500.400 370.050 501.600 371.100 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 704.400 366.900 705.600 385.950 ;
        RECT 718.950 367.950 721.050 370.050 ;
        RECT 719.400 366.900 720.600 367.950 ;
        RECT 703.950 364.800 706.050 366.900 ;
        RECT 718.950 364.800 721.050 366.900 ;
        RECT 481.950 337.950 484.050 340.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 479.400 334.050 480.600 334.950 ;
        RECT 479.400 332.400 484.050 334.050 ;
        RECT 614.400 333.000 615.600 334.950 ;
        RECT 480.000 331.950 484.050 332.400 ;
        RECT 482.400 316.050 483.600 331.950 ;
        RECT 535.950 328.950 538.050 331.050 ;
        RECT 613.950 328.950 616.050 333.000 ;
        RECT 536.400 316.050 537.600 328.950 ;
        RECT 481.950 313.950 484.050 316.050 ;
        RECT 535.950 313.950 538.050 316.050 ;
        RECT 614.400 298.050 615.600 328.950 ;
        RECT 613.950 295.950 616.050 298.050 ;
        RECT 625.950 295.950 628.050 301.050 ;
        RECT 634.950 294.000 637.050 298.050 ;
        RECT 649.950 295.950 652.050 298.050 ;
        RECT 635.400 292.050 636.600 294.000 ;
        RECT 650.400 292.050 651.600 295.950 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 649.950 289.950 652.050 292.050 ;
        RECT 652.950 286.950 655.050 289.050 ;
        RECT 653.400 268.050 654.600 286.950 ;
        RECT 652.950 265.950 655.050 268.050 ;
        RECT 661.950 265.950 664.050 268.050 ;
        RECT 662.400 255.600 663.600 265.950 ;
        RECT 659.400 254.400 663.600 255.600 ;
        RECT 659.400 220.050 660.600 254.400 ;
        RECT 649.950 217.950 652.050 220.050 ;
        RECT 658.950 217.950 661.050 220.050 ;
        RECT 650.400 195.600 651.600 217.950 ;
        RECT 685.950 216.000 688.050 220.050 ;
        RECT 686.400 214.050 687.600 216.000 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 650.400 194.400 654.600 195.600 ;
        RECT 653.400 163.050 654.600 194.400 ;
        RECT 703.950 166.950 706.050 169.050 ;
        RECT 793.950 166.950 796.050 169.050 ;
        RECT 704.400 163.050 705.600 166.950 ;
        RECT 652.950 160.950 655.050 163.050 ;
        RECT 703.950 160.950 706.050 163.050 ;
        RECT 653.400 109.050 654.600 160.950 ;
        RECT 794.400 145.050 795.600 166.950 ;
        RECT 793.950 142.950 796.050 145.050 ;
        RECT 799.950 142.950 802.050 145.050 ;
        RECT 800.400 139.050 801.600 142.950 ;
        RECT 799.950 136.950 802.050 139.050 ;
        RECT 853.950 136.950 856.050 139.050 ;
        RECT 854.400 136.050 855.600 136.950 ;
        RECT 853.950 133.950 856.050 136.050 ;
        RECT 643.950 106.950 646.050 109.050 ;
        RECT 652.950 106.950 655.050 109.050 ;
        RECT 644.400 61.200 645.600 106.950 ;
        RECT 637.950 59.100 640.050 61.200 ;
        RECT 643.950 59.100 646.050 61.200 ;
        RECT 638.400 58.050 639.600 59.100 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 644.400 10.050 645.600 59.100 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 680.400 10.050 681.600 22.950 ;
        RECT 643.950 7.950 646.050 10.050 ;
        RECT 679.950 7.950 682.050 10.050 ;
      LAYER metal3 ;
        RECT 499.950 939.600 502.050 940.050 ;
        RECT 580.950 939.600 583.050 940.050 ;
        RECT 499.950 938.400 583.050 939.600 ;
        RECT 499.950 937.950 502.050 938.400 ;
        RECT 580.950 937.950 583.050 938.400 ;
        RECT 580.950 838.950 583.050 841.050 ;
        RECT 581.400 835.050 582.600 838.950 ;
        RECT 580.950 832.950 583.050 835.050 ;
        RECT 550.950 825.600 553.050 826.050 ;
        RECT 580.950 825.600 583.050 826.050 ;
        RECT 550.950 824.400 583.050 825.600 ;
        RECT 550.950 823.950 553.050 824.400 ;
        RECT 580.950 823.950 583.050 824.400 ;
        RECT 544.950 753.600 547.050 754.050 ;
        RECT 550.950 753.600 553.050 754.050 ;
        RECT 544.950 752.400 553.050 753.600 ;
        RECT 544.950 751.950 547.050 752.400 ;
        RECT 550.950 751.950 553.050 752.400 ;
        RECT 544.950 652.950 547.050 655.050 ;
        RECT 545.400 646.050 546.600 652.950 ;
        RECT 545.400 644.400 550.050 646.050 ;
        RECT 546.000 643.950 550.050 644.400 ;
        RECT 547.950 630.600 550.050 631.050 ;
        RECT 565.950 630.600 568.050 631.050 ;
        RECT 547.950 629.400 568.050 630.600 ;
        RECT 547.950 628.950 550.050 629.400 ;
        RECT 565.950 628.950 568.050 629.400 ;
        RECT 565.950 571.950 568.050 574.050 ;
        RECT 523.950 567.600 526.050 568.050 ;
        RECT 566.400 567.600 567.600 571.950 ;
        RECT 523.950 566.400 567.600 567.600 ;
        RECT 523.950 565.950 526.050 566.400 ;
        RECT 505.950 543.600 508.050 544.050 ;
        RECT 523.950 543.600 526.050 544.050 ;
        RECT 505.950 542.400 526.050 543.600 ;
        RECT 505.950 541.950 508.050 542.400 ;
        RECT 523.950 541.950 526.050 542.400 ;
        RECT 505.950 527.100 508.050 529.200 ;
        RECT 506.400 520.050 507.600 527.100 ;
        RECT 505.950 517.950 508.050 520.050 ;
        RECT 811.950 516.600 814.050 517.050 ;
        RECT 847.950 516.600 850.050 517.050 ;
        RECT 811.950 515.400 850.050 516.600 ;
        RECT 811.950 514.950 814.050 515.400 ;
        RECT 847.950 514.950 850.050 515.400 ;
        RECT 754.950 495.600 757.050 496.200 ;
        RECT 772.950 495.600 775.050 495.900 ;
        RECT 754.950 494.400 775.050 495.600 ;
        RECT 754.950 494.100 757.050 494.400 ;
        RECT 772.950 493.800 775.050 494.400 ;
        RECT 847.950 495.750 850.050 496.200 ;
        RECT 859.950 495.750 862.050 496.200 ;
        RECT 847.950 494.550 862.050 495.750 ;
        RECT 847.950 494.100 850.050 494.550 ;
        RECT 859.950 494.100 862.050 494.550 ;
        RECT 505.950 480.600 508.050 481.050 ;
        RECT 514.950 480.600 517.050 481.050 ;
        RECT 505.950 479.400 517.050 480.600 ;
        RECT 505.950 478.950 508.050 479.400 ;
        RECT 514.950 478.950 517.050 479.400 ;
        RECT 772.950 462.600 775.050 463.050 ;
        RECT 811.950 462.600 814.050 463.050 ;
        RECT 835.950 462.600 838.050 463.050 ;
        RECT 772.950 461.400 838.050 462.600 ;
        RECT 772.950 460.950 775.050 461.400 ;
        RECT 811.950 460.950 814.050 461.400 ;
        RECT 835.950 460.950 838.050 461.400 ;
        RECT 775.950 426.600 778.050 427.050 ;
        RECT 719.400 425.400 778.050 426.600 ;
        RECT 719.400 423.600 720.600 425.400 ;
        RECT 775.950 424.950 778.050 425.400 ;
        RECT 710.400 422.400 720.600 423.600 ;
        RECT 710.400 420.600 711.600 422.400 ;
        RECT 698.400 419.400 711.600 420.600 ;
        RECT 514.950 415.950 517.050 418.050 ;
        RECT 694.950 417.600 697.050 418.200 ;
        RECT 698.400 417.600 699.600 419.400 ;
        RECT 680.400 416.400 699.600 417.600 ;
        RECT 508.950 411.600 511.050 412.050 ;
        RECT 515.400 411.600 516.600 415.950 ;
        RECT 526.950 411.600 529.050 411.900 ;
        RECT 508.950 411.450 529.050 411.600 ;
        RECT 553.950 411.450 556.050 411.900 ;
        RECT 508.950 410.400 556.050 411.450 ;
        RECT 508.950 409.950 511.050 410.400 ;
        RECT 526.950 410.250 556.050 410.400 ;
        RECT 526.950 409.800 529.050 410.250 ;
        RECT 553.950 409.800 556.050 410.250 ;
        RECT 664.950 411.600 667.050 412.050 ;
        RECT 680.400 411.900 681.600 416.400 ;
        RECT 694.950 416.100 697.050 416.400 ;
        RECT 679.950 411.600 682.050 411.900 ;
        RECT 664.950 410.400 682.050 411.600 ;
        RECT 664.950 409.950 667.050 410.400 ;
        RECT 679.950 409.800 682.050 410.400 ;
        RECT 553.950 396.600 556.050 397.050 ;
        RECT 664.950 396.600 667.050 397.050 ;
        RECT 553.950 395.400 667.050 396.600 ;
        RECT 553.950 394.950 556.050 395.400 ;
        RECT 664.950 394.950 667.050 395.400 ;
        RECT 481.950 387.600 484.050 388.050 ;
        RECT 496.950 387.600 499.050 388.050 ;
        RECT 481.950 386.400 499.050 387.600 ;
        RECT 481.950 385.950 484.050 386.400 ;
        RECT 496.950 385.950 499.050 386.400 ;
        RECT 679.950 387.600 682.050 388.050 ;
        RECT 703.950 387.600 706.050 388.050 ;
        RECT 679.950 386.400 706.050 387.600 ;
        RECT 679.950 385.950 682.050 386.400 ;
        RECT 703.950 385.950 706.050 386.400 ;
        RECT 499.950 372.750 502.050 373.200 ;
        RECT 508.950 372.750 511.050 373.200 ;
        RECT 499.950 371.550 511.050 372.750 ;
        RECT 499.950 371.100 502.050 371.550 ;
        RECT 508.950 371.100 511.050 371.550 ;
        RECT 703.950 366.450 706.050 366.900 ;
        RECT 718.950 366.450 721.050 366.900 ;
        RECT 703.950 365.250 721.050 366.450 ;
        RECT 703.950 364.800 706.050 365.250 ;
        RECT 718.950 364.800 721.050 365.250 ;
        RECT 535.950 330.600 538.050 331.050 ;
        RECT 613.950 330.600 616.050 331.050 ;
        RECT 535.950 329.400 616.050 330.600 ;
        RECT 535.950 328.950 538.050 329.400 ;
        RECT 613.950 328.950 616.050 329.400 ;
        RECT 481.950 315.600 484.050 316.050 ;
        RECT 535.950 315.600 538.050 316.050 ;
        RECT 481.950 314.400 538.050 315.600 ;
        RECT 481.950 313.950 484.050 314.400 ;
        RECT 535.950 313.950 538.050 314.400 ;
        RECT 613.950 297.600 616.050 298.050 ;
        RECT 625.950 297.600 628.050 301.050 ;
        RECT 613.950 297.000 628.050 297.600 ;
        RECT 634.950 297.600 637.050 298.050 ;
        RECT 649.950 297.600 652.050 298.050 ;
        RECT 613.950 296.400 627.600 297.000 ;
        RECT 634.950 296.400 652.050 297.600 ;
        RECT 613.950 295.950 616.050 296.400 ;
        RECT 634.950 295.950 637.050 296.400 ;
        RECT 649.950 295.950 652.050 296.400 ;
        RECT 649.950 291.600 654.000 292.050 ;
        RECT 649.950 291.000 654.600 291.600 ;
        RECT 649.950 289.950 655.050 291.000 ;
        RECT 652.950 286.950 655.050 289.950 ;
        RECT 652.950 267.600 655.050 268.050 ;
        RECT 661.950 267.600 664.050 268.050 ;
        RECT 652.950 266.400 664.050 267.600 ;
        RECT 652.950 265.950 655.050 266.400 ;
        RECT 661.950 265.950 664.050 266.400 ;
        RECT 649.950 219.600 652.050 220.050 ;
        RECT 658.950 219.600 661.050 220.050 ;
        RECT 685.950 219.600 688.050 220.050 ;
        RECT 649.950 218.400 688.050 219.600 ;
        RECT 649.950 217.950 652.050 218.400 ;
        RECT 658.950 217.950 661.050 218.400 ;
        RECT 685.950 217.950 688.050 218.400 ;
        RECT 703.950 168.600 706.050 169.050 ;
        RECT 793.950 168.600 796.050 169.050 ;
        RECT 703.950 167.400 796.050 168.600 ;
        RECT 703.950 166.950 706.050 167.400 ;
        RECT 793.950 166.950 796.050 167.400 ;
        RECT 652.950 162.600 655.050 163.050 ;
        RECT 703.950 162.600 706.050 163.050 ;
        RECT 652.950 161.400 706.050 162.600 ;
        RECT 652.950 160.950 655.050 161.400 ;
        RECT 703.950 160.950 706.050 161.400 ;
        RECT 793.950 144.600 796.050 145.050 ;
        RECT 799.950 144.600 802.050 145.050 ;
        RECT 793.950 143.400 802.050 144.600 ;
        RECT 793.950 142.950 796.050 143.400 ;
        RECT 799.950 142.950 802.050 143.400 ;
        RECT 799.950 138.600 802.050 139.050 ;
        RECT 853.950 138.600 856.050 139.050 ;
        RECT 799.950 137.400 856.050 138.600 ;
        RECT 799.950 136.950 802.050 137.400 ;
        RECT 853.950 136.950 856.050 137.400 ;
        RECT 643.950 108.600 646.050 109.050 ;
        RECT 652.950 108.600 655.050 109.050 ;
        RECT 643.950 107.400 655.050 108.600 ;
        RECT 643.950 106.950 646.050 107.400 ;
        RECT 652.950 106.950 655.050 107.400 ;
        RECT 637.950 60.750 640.050 61.200 ;
        RECT 643.950 60.750 646.050 61.200 ;
        RECT 637.950 59.550 646.050 60.750 ;
        RECT 637.950 59.100 640.050 59.550 ;
        RECT 643.950 59.100 646.050 59.550 ;
        RECT 643.950 9.600 646.050 10.050 ;
        RECT 679.950 9.600 682.050 10.050 ;
        RECT 643.950 8.400 682.050 9.600 ;
        RECT 643.950 7.950 646.050 8.400 ;
        RECT 679.950 7.950 682.050 8.400 ;
    END
  END ABCmd_i[7]
  PIN ABCmd_i[6]
    PORT
      LAYER metal2 ;
        RECT 728.400 940.050 729.600 945.600 ;
        RECT 727.950 937.950 730.050 940.050 ;
        RECT 778.950 937.950 781.050 940.050 ;
        RECT 779.400 910.050 780.600 937.950 ;
        RECT 763.950 907.950 766.050 910.050 ;
        RECT 778.950 907.950 781.050 910.050 ;
        RECT 764.400 877.050 765.600 907.950 ;
        RECT 763.950 874.950 766.050 877.050 ;
        RECT 775.950 874.950 778.050 877.050 ;
        RECT 776.400 808.050 777.600 874.950 ;
        RECT 775.950 805.950 778.050 808.050 ;
        RECT 763.950 799.950 766.050 802.050 ;
        RECT 764.400 763.050 765.600 799.950 ;
        RECT 763.950 760.950 766.050 763.050 ;
        RECT 763.950 754.950 766.050 757.050 ;
        RECT 764.400 694.050 765.600 754.950 ;
        RECT 763.950 691.950 766.050 694.050 ;
        RECT 778.950 691.950 781.050 694.050 ;
        RECT 779.400 661.050 780.600 691.950 ;
        RECT 736.950 658.950 739.050 661.050 ;
        RECT 769.950 658.950 772.050 661.050 ;
        RECT 778.950 658.950 781.050 661.050 ;
        RECT 737.400 649.050 738.600 658.950 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 770.400 616.050 771.600 658.950 ;
        RECT 730.950 613.950 733.050 616.050 ;
        RECT 769.950 613.950 772.050 616.050 ;
        RECT 775.950 613.950 778.050 616.050 ;
        RECT 731.400 604.050 732.600 613.950 ;
        RECT 776.400 606.600 777.600 613.950 ;
        RECT 776.400 605.400 780.600 606.600 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 779.400 573.600 780.600 605.400 ;
        RECT 776.400 572.400 780.600 573.600 ;
        RECT 776.400 532.050 777.600 572.400 ;
        RECT 775.950 529.950 778.050 532.050 ;
        RECT 793.950 529.800 796.050 531.900 ;
        RECT 794.400 522.900 795.600 529.800 ;
        RECT 814.950 528.000 817.050 532.050 ;
        RECT 832.950 528.000 835.050 532.050 ;
        RECT 815.400 526.050 816.600 528.000 ;
        RECT 833.400 526.050 834.600 528.000 ;
        RECT 805.950 523.950 808.050 526.050 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 832.950 523.950 835.050 526.050 ;
        RECT 806.400 522.900 807.600 523.950 ;
        RECT 793.950 520.800 796.050 522.900 ;
        RECT 805.950 520.800 808.050 522.900 ;
      LAYER metal3 ;
        RECT 727.950 939.600 730.050 940.050 ;
        RECT 778.950 939.600 781.050 940.050 ;
        RECT 727.950 938.400 781.050 939.600 ;
        RECT 727.950 937.950 730.050 938.400 ;
        RECT 778.950 937.950 781.050 938.400 ;
        RECT 763.950 909.600 766.050 910.050 ;
        RECT 778.950 909.600 781.050 910.050 ;
        RECT 763.950 908.400 781.050 909.600 ;
        RECT 763.950 907.950 766.050 908.400 ;
        RECT 778.950 907.950 781.050 908.400 ;
        RECT 763.950 876.600 766.050 877.050 ;
        RECT 775.950 876.600 778.050 877.050 ;
        RECT 763.950 875.400 778.050 876.600 ;
        RECT 763.950 874.950 766.050 875.400 ;
        RECT 775.950 874.950 778.050 875.400 ;
        RECT 775.950 805.950 778.050 808.050 ;
        RECT 763.950 801.600 766.050 802.050 ;
        RECT 776.400 801.600 777.600 805.950 ;
        RECT 763.950 800.400 777.600 801.600 ;
        RECT 763.950 799.950 766.050 800.400 ;
        RECT 763.950 760.950 766.050 763.050 ;
        RECT 764.400 757.050 765.600 760.950 ;
        RECT 763.950 754.950 766.050 757.050 ;
        RECT 763.950 693.600 766.050 694.050 ;
        RECT 778.950 693.600 781.050 694.050 ;
        RECT 763.950 692.400 781.050 693.600 ;
        RECT 763.950 691.950 766.050 692.400 ;
        RECT 778.950 691.950 781.050 692.400 ;
        RECT 736.950 660.600 739.050 661.050 ;
        RECT 769.950 660.600 772.050 661.050 ;
        RECT 778.950 660.600 781.050 661.050 ;
        RECT 736.950 659.400 781.050 660.600 ;
        RECT 736.950 658.950 739.050 659.400 ;
        RECT 769.950 658.950 772.050 659.400 ;
        RECT 778.950 658.950 781.050 659.400 ;
        RECT 730.950 615.600 733.050 616.050 ;
        RECT 769.950 615.600 772.050 616.050 ;
        RECT 775.950 615.600 778.050 616.050 ;
        RECT 730.950 614.400 778.050 615.600 ;
        RECT 730.950 613.950 733.050 614.400 ;
        RECT 769.950 613.950 772.050 614.400 ;
        RECT 775.950 613.950 778.050 614.400 ;
        RECT 775.950 531.600 778.050 532.050 ;
        RECT 793.950 531.600 796.050 531.900 ;
        RECT 814.950 531.600 817.050 532.050 ;
        RECT 832.950 531.600 835.050 532.050 ;
        RECT 775.950 530.400 835.050 531.600 ;
        RECT 775.950 529.950 778.050 530.400 ;
        RECT 793.950 529.800 796.050 530.400 ;
        RECT 814.950 529.950 817.050 530.400 ;
        RECT 832.950 529.950 835.050 530.400 ;
        RECT 793.950 522.450 796.050 522.900 ;
        RECT 805.950 522.450 808.050 522.900 ;
        RECT 793.950 521.250 808.050 522.450 ;
        RECT 793.950 520.800 796.050 521.250 ;
        RECT 805.950 520.800 808.050 521.250 ;
    END
  END ABCmd_i[6]
  PIN ABCmd_i[5]
    PORT
      LAYER metal1 ;
        RECT 478.950 762.450 481.050 763.050 ;
        RECT 484.950 762.450 487.050 763.050 ;
        RECT 478.950 761.550 487.050 762.450 ;
        RECT 478.950 760.950 481.050 761.550 ;
        RECT 484.950 760.950 487.050 761.550 ;
      LAYER metal2 ;
        RECT 529.950 934.950 532.050 937.050 ;
        RECT 577.950 934.950 580.050 937.050 ;
        RECT 655.950 934.950 658.050 937.050 ;
        RECT 530.400 931.050 531.600 934.950 ;
        RECT 478.950 928.950 481.050 931.050 ;
        RECT 487.950 928.950 490.050 931.050 ;
        RECT 529.950 928.950 532.050 931.050 ;
        RECT 479.400 916.050 480.600 928.950 ;
        RECT 478.950 913.950 481.050 916.050 ;
        RECT 488.400 847.050 489.600 928.950 ;
        RECT 530.400 916.050 531.600 928.950 ;
        RECT 529.950 913.950 532.050 916.050 ;
        RECT 538.950 880.950 541.050 883.050 ;
        RECT 539.400 868.050 540.600 880.950 ;
        RECT 578.400 868.050 579.600 934.950 ;
        RECT 656.400 931.050 657.600 934.950 ;
        RECT 743.400 931.050 744.600 945.600 ;
        RECT 655.950 928.950 658.050 931.050 ;
        RECT 742.950 928.950 745.050 931.050 ;
        RECT 799.950 928.950 802.050 931.050 ;
        RECT 538.950 865.950 541.050 868.050 ;
        RECT 547.950 865.950 550.050 868.050 ;
        RECT 577.950 865.950 580.050 868.050 ;
        RECT 607.950 865.950 610.050 868.050 ;
        RECT 463.950 844.950 466.050 847.050 ;
        RECT 469.950 844.950 472.050 847.050 ;
        RECT 487.950 844.950 490.050 847.050 ;
        RECT 464.400 838.050 465.600 844.950 ;
        RECT 463.950 835.950 466.050 838.050 ;
        RECT 470.400 823.050 471.600 844.950 ;
        RECT 548.400 838.050 549.600 865.950 ;
        RECT 608.400 838.050 609.600 865.950 ;
        RECT 547.950 835.950 550.050 838.050 ;
        RECT 607.950 835.950 610.050 838.050 ;
        RECT 469.950 820.950 472.050 823.050 ;
        RECT 484.950 820.950 487.050 823.050 ;
        RECT 485.400 763.050 486.600 820.950 ;
        RECT 800.400 820.050 801.600 928.950 ;
        RECT 784.950 817.950 787.050 820.050 ;
        RECT 799.950 817.950 802.050 820.050 ;
        RECT 785.400 811.050 786.600 817.950 ;
        RECT 778.950 808.950 781.050 811.050 ;
        RECT 779.400 769.050 780.600 808.950 ;
        RECT 784.950 807.000 787.050 811.050 ;
        RECT 785.400 805.050 786.600 807.000 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 748.950 765.600 751.050 769.050 ;
        RECT 775.950 767.400 780.600 769.050 ;
        RECT 775.950 766.950 780.000 767.400 ;
        RECT 746.400 765.000 751.050 765.600 ;
        RECT 746.400 764.400 750.600 765.000 ;
        RECT 478.950 760.950 481.050 763.050 ;
        RECT 484.950 760.950 487.050 763.050 ;
        RECT 479.400 736.050 480.600 760.950 ;
        RECT 746.400 760.050 747.600 764.400 ;
        RECT 745.950 757.950 748.050 760.050 ;
        RECT 478.950 733.950 481.050 736.050 ;
        RECT 496.950 733.950 499.050 736.050 ;
        RECT 497.400 730.200 498.600 733.950 ;
        RECT 496.950 728.100 499.050 730.200 ;
        RECT 497.400 727.050 498.600 728.100 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 530.400 723.900 531.600 724.950 ;
        RECT 560.400 723.900 561.600 724.950 ;
        RECT 529.950 721.800 532.050 723.900 ;
        RECT 559.950 721.800 562.050 723.900 ;
      LAYER metal3 ;
        RECT 529.950 936.600 532.050 937.050 ;
        RECT 577.950 936.600 580.050 937.050 ;
        RECT 655.950 936.600 658.050 937.050 ;
        RECT 529.950 935.400 658.050 936.600 ;
        RECT 529.950 934.950 532.050 935.400 ;
        RECT 577.950 934.950 580.050 935.400 ;
        RECT 655.950 934.950 658.050 935.400 ;
        RECT 478.950 930.600 481.050 931.050 ;
        RECT 487.950 930.600 490.050 931.050 ;
        RECT 529.950 930.600 532.050 931.050 ;
        RECT 478.950 929.400 532.050 930.600 ;
        RECT 478.950 928.950 481.050 929.400 ;
        RECT 487.950 928.950 490.050 929.400 ;
        RECT 529.950 928.950 532.050 929.400 ;
        RECT 655.950 930.600 658.050 931.050 ;
        RECT 742.950 930.600 745.050 931.050 ;
        RECT 799.950 930.600 802.050 931.050 ;
        RECT 655.950 929.400 802.050 930.600 ;
        RECT 655.950 928.950 658.050 929.400 ;
        RECT 742.950 928.950 745.050 929.400 ;
        RECT 799.950 928.950 802.050 929.400 ;
        RECT 538.950 867.600 541.050 868.050 ;
        RECT 547.950 867.600 550.050 868.050 ;
        RECT 577.950 867.600 580.050 868.050 ;
        RECT 607.950 867.600 610.050 868.050 ;
        RECT 538.950 866.400 610.050 867.600 ;
        RECT 538.950 865.950 541.050 866.400 ;
        RECT 547.950 865.950 550.050 866.400 ;
        RECT 577.950 865.950 580.050 866.400 ;
        RECT 607.950 865.950 610.050 866.400 ;
        RECT 463.950 846.600 466.050 847.050 ;
        RECT 469.950 846.600 472.050 847.050 ;
        RECT 487.950 846.600 490.050 847.050 ;
        RECT 463.950 845.400 490.050 846.600 ;
        RECT 463.950 844.950 466.050 845.400 ;
        RECT 469.950 844.950 472.050 845.400 ;
        RECT 487.950 844.950 490.050 845.400 ;
        RECT 469.950 822.600 472.050 823.050 ;
        RECT 484.950 822.600 487.050 823.050 ;
        RECT 469.950 821.400 487.050 822.600 ;
        RECT 469.950 820.950 472.050 821.400 ;
        RECT 484.950 820.950 487.050 821.400 ;
        RECT 784.950 819.600 787.050 820.050 ;
        RECT 799.950 819.600 802.050 820.050 ;
        RECT 784.950 818.400 802.050 819.600 ;
        RECT 784.950 817.950 787.050 818.400 ;
        RECT 799.950 817.950 802.050 818.400 ;
        RECT 778.950 810.600 781.050 811.050 ;
        RECT 784.950 810.600 787.050 811.050 ;
        RECT 778.950 809.400 787.050 810.600 ;
        RECT 778.950 808.950 781.050 809.400 ;
        RECT 784.950 808.950 787.050 809.400 ;
        RECT 748.950 768.600 751.050 769.050 ;
        RECT 775.950 768.600 778.050 769.050 ;
        RECT 748.950 767.400 778.050 768.600 ;
        RECT 748.950 766.950 751.050 767.400 ;
        RECT 775.950 766.950 778.050 767.400 ;
        RECT 478.950 735.600 481.050 736.050 ;
        RECT 496.950 735.600 499.050 736.050 ;
        RECT 478.950 734.400 499.050 735.600 ;
        RECT 478.950 733.950 481.050 734.400 ;
        RECT 496.950 733.950 499.050 734.400 ;
        RECT 496.950 729.600 499.050 730.200 ;
        RECT 496.950 728.400 528.600 729.600 ;
        RECT 496.950 728.100 499.050 728.400 ;
        RECT 527.400 726.600 528.600 728.400 ;
        RECT 527.400 725.400 531.600 726.600 ;
        RECT 530.400 723.900 531.600 725.400 ;
        RECT 529.950 723.600 532.050 723.900 ;
        RECT 559.950 723.600 562.050 723.900 ;
        RECT 529.950 722.400 562.050 723.600 ;
        RECT 529.950 721.800 532.050 722.400 ;
        RECT 559.950 721.800 562.050 722.400 ;
    END
  END ABCmd_i[5]
  PIN ABCmd_i[4]
    PORT
      LAYER metal1 ;
        RECT 769.950 831.450 772.050 832.050 ;
        RECT 778.950 831.450 781.050 832.050 ;
        RECT 784.950 831.450 787.050 832.050 ;
        RECT 769.950 830.550 787.050 831.450 ;
        RECT 769.950 829.950 772.050 830.550 ;
        RECT 778.950 829.950 781.050 830.550 ;
        RECT 784.950 829.950 787.050 830.550 ;
      LAYER metal2 ;
        RECT 767.400 937.050 768.600 945.600 ;
        RECT 760.950 934.950 763.050 937.050 ;
        RECT 766.950 934.950 769.050 937.050 ;
        RECT 761.400 853.050 762.600 934.950 ;
        RECT 760.950 850.950 763.050 853.050 ;
        RECT 778.950 850.950 781.050 853.050 ;
        RECT 601.950 847.950 604.050 850.050 ;
        RECT 602.400 841.050 603.600 847.950 ;
        RECT 601.950 838.950 604.050 841.050 ;
        RECT 601.950 832.950 604.050 835.050 ;
        RECT 602.400 810.600 603.600 832.950 ;
        RECT 779.400 832.050 780.600 850.950 ;
        RECT 769.950 829.950 772.050 832.050 ;
        RECT 778.950 829.950 781.050 832.050 ;
        RECT 784.950 831.600 789.000 832.050 ;
        RECT 784.950 829.950 789.600 831.600 ;
        RECT 602.400 809.400 606.600 810.600 ;
        RECT 605.400 805.050 606.600 809.400 ;
        RECT 770.400 808.050 771.600 829.950 ;
        RECT 788.400 814.050 789.600 829.950 ;
        RECT 787.950 811.950 790.050 814.050 ;
        RECT 799.800 811.950 801.900 814.050 ;
        RECT 769.950 805.950 772.050 808.050 ;
        RECT 604.950 802.950 607.050 805.050 ;
        RECT 800.400 802.050 801.600 811.950 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 799.950 799.950 802.050 802.050 ;
        RECT 806.400 801.900 807.600 802.950 ;
        RECT 805.950 799.800 808.050 801.900 ;
        RECT 751.950 796.950 754.050 799.050 ;
        RECT 752.400 760.050 753.600 796.950 ;
        RECT 751.950 757.950 754.050 760.050 ;
      LAYER metal3 ;
        RECT 760.950 936.600 763.050 937.050 ;
        RECT 766.950 936.600 769.050 937.050 ;
        RECT 760.950 935.400 769.050 936.600 ;
        RECT 760.950 934.950 763.050 935.400 ;
        RECT 766.950 934.950 769.050 935.400 ;
        RECT 760.950 852.600 763.050 853.050 ;
        RECT 778.950 852.600 781.050 853.050 ;
        RECT 760.950 851.400 781.050 852.600 ;
        RECT 760.950 850.950 763.050 851.400 ;
        RECT 778.950 850.950 781.050 851.400 ;
        RECT 601.950 849.600 604.050 850.050 ;
        RECT 761.400 849.600 762.600 850.950 ;
        RECT 601.950 848.400 762.600 849.600 ;
        RECT 601.950 847.950 604.050 848.400 ;
        RECT 601.950 838.950 604.050 841.050 ;
        RECT 602.400 835.050 603.600 838.950 ;
        RECT 601.950 832.950 604.050 835.050 ;
        RECT 787.950 813.600 790.050 814.050 ;
        RECT 799.800 813.600 801.900 814.050 ;
        RECT 787.950 812.400 801.900 813.600 ;
        RECT 787.950 811.950 790.050 812.400 ;
        RECT 799.800 811.950 801.900 812.400 ;
        RECT 769.950 807.600 772.050 808.050 ;
        RECT 755.400 806.400 772.050 807.600 ;
        RECT 755.400 799.050 756.600 806.400 ;
        RECT 769.950 805.950 772.050 806.400 ;
        RECT 799.950 801.600 802.050 802.050 ;
        RECT 805.950 801.600 808.050 801.900 ;
        RECT 799.950 800.400 808.050 801.600 ;
        RECT 799.950 799.950 802.050 800.400 ;
        RECT 805.950 799.800 808.050 800.400 ;
        RECT 751.950 797.400 756.600 799.050 ;
        RECT 751.950 796.950 756.000 797.400 ;
    END
  END ABCmd_i[4]
  PIN ABCmd_i[3]
    PORT
      LAYER metal1 ;
        RECT 843.000 885.450 847.050 886.050 ;
        RECT 842.550 883.950 847.050 885.450 ;
        RECT 842.550 880.050 843.450 883.950 ;
        RECT 842.550 878.550 847.050 880.050 ;
        RECT 843.000 877.950 847.050 878.550 ;
      LAYER metal2 ;
        RECT 844.950 922.950 847.050 925.050 ;
        RECT 845.400 886.050 846.600 922.950 ;
        RECT 872.400 922.050 873.600 945.600 ;
        RECT 871.950 919.950 874.050 922.050 ;
        RECT 889.950 918.000 892.050 922.050 ;
        RECT 890.400 916.050 891.600 918.000 ;
        RECT 889.950 913.950 892.050 916.050 ;
        RECT 844.950 883.950 847.050 886.050 ;
        RECT 844.950 877.950 847.050 880.050 ;
        RECT 845.400 858.600 846.600 877.950 ;
        RECT 845.400 857.400 849.600 858.600 ;
        RECT 848.400 823.050 849.600 857.400 ;
        RECT 838.950 820.950 841.050 823.050 ;
        RECT 847.950 820.950 850.050 823.050 ;
        RECT 839.400 775.050 840.600 820.950 ;
        RECT 817.950 772.950 820.050 775.050 ;
        RECT 838.950 772.950 841.050 775.050 ;
        RECT 818.400 763.050 819.600 772.950 ;
        RECT 817.950 760.950 820.050 763.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 815.400 756.900 816.600 757.950 ;
        RECT 814.950 754.800 817.050 756.900 ;
      LAYER metal3 ;
        RECT 844.950 924.600 847.050 925.050 ;
        RECT 844.950 923.400 873.600 924.600 ;
        RECT 844.950 922.950 847.050 923.400 ;
        RECT 872.400 922.050 873.600 923.400 ;
        RECT 871.950 921.600 874.050 922.050 ;
        RECT 889.950 921.600 892.050 922.050 ;
        RECT 871.950 920.400 892.050 921.600 ;
        RECT 871.950 919.950 874.050 920.400 ;
        RECT 889.950 919.950 892.050 920.400 ;
        RECT 838.950 822.600 841.050 823.050 ;
        RECT 847.950 822.600 850.050 823.050 ;
        RECT 838.950 821.400 850.050 822.600 ;
        RECT 838.950 820.950 841.050 821.400 ;
        RECT 847.950 820.950 850.050 821.400 ;
        RECT 817.950 774.600 820.050 775.050 ;
        RECT 838.950 774.600 841.050 775.050 ;
        RECT 817.950 773.400 841.050 774.600 ;
        RECT 817.950 772.950 820.050 773.400 ;
        RECT 838.950 772.950 841.050 773.400 ;
        RECT 816.000 762.600 820.050 763.050 ;
        RECT 815.400 760.950 820.050 762.600 ;
        RECT 815.400 756.900 816.600 760.950 ;
        RECT 814.950 754.800 817.050 756.900 ;
    END
  END ABCmd_i[3]
  PIN ABCmd_i[2]
    PORT
      LAYER metal2 ;
        RECT 754.950 884.100 757.050 886.200 ;
        RECT 755.400 883.050 756.600 884.100 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 751.950 877.950 754.050 880.050 ;
        RECT 752.400 826.050 753.600 877.950 ;
        RECT 904.950 835.950 907.050 838.050 ;
        RECT 751.950 823.950 754.050 826.050 ;
        RECT 772.950 823.950 775.050 826.050 ;
        RECT 773.400 817.050 774.600 823.950 ;
        RECT 905.400 817.050 906.600 835.950 ;
        RECT 772.950 814.950 775.050 817.050 ;
        RECT 904.950 814.950 907.050 817.050 ;
        RECT 913.950 814.950 916.050 817.050 ;
        RECT 773.400 805.050 774.600 814.950 ;
        RECT 914.400 805.050 915.600 814.950 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 913.950 802.950 916.050 805.050 ;
      LAYER metal3 ;
        RECT 754.950 884.100 757.050 886.200 ;
        RECT 755.400 880.050 756.600 884.100 ;
        RECT 751.950 878.400 756.600 880.050 ;
        RECT 751.950 877.950 756.000 878.400 ;
        RECT 751.950 825.600 754.050 826.050 ;
        RECT 772.950 825.600 775.050 826.050 ;
        RECT 751.950 824.400 775.050 825.600 ;
        RECT 751.950 823.950 754.050 824.400 ;
        RECT 772.950 823.950 775.050 824.400 ;
        RECT 772.950 816.600 775.050 817.050 ;
        RECT 904.950 816.600 907.050 817.050 ;
        RECT 913.950 816.600 916.050 817.050 ;
        RECT 772.950 815.400 927.600 816.600 ;
        RECT 772.950 814.950 775.050 815.400 ;
        RECT 904.950 814.950 907.050 815.400 ;
        RECT 913.950 814.950 916.050 815.400 ;
    END
  END ABCmd_i[2]
  PIN ABCmd_i[1]
    PORT
      LAYER metal1 ;
        RECT 622.950 732.450 625.050 733.050 ;
        RECT 611.550 731.550 625.050 732.450 ;
        RECT 611.550 724.050 612.450 731.550 ;
        RECT 622.950 730.950 625.050 731.550 ;
        RECT 611.550 722.550 616.050 724.050 ;
        RECT 612.000 721.950 616.050 722.550 ;
      LAYER metal2 ;
        RECT 568.950 839.100 571.050 841.200 ;
        RECT 569.400 838.050 570.600 839.100 ;
        RECT 574.950 838.950 577.050 841.050 ;
        RECT 568.950 835.950 571.050 838.050 ;
        RECT 575.400 808.050 576.600 838.950 ;
        RECT 574.950 805.950 577.050 808.050 ;
        RECT 730.950 806.100 733.050 808.200 ;
        RECT 742.950 806.100 745.050 808.200 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 616.800 799.950 618.900 802.050 ;
        RECT 617.400 772.050 618.600 799.950 ;
        RECT 662.400 793.050 663.600 802.950 ;
        RECT 731.400 796.050 732.600 806.100 ;
        RECT 743.400 805.050 744.600 806.100 ;
        RECT 742.950 802.950 745.050 805.050 ;
        RECT 919.950 802.950 922.050 805.050 ;
        RECT 730.950 793.950 733.050 796.050 ;
        RECT 754.950 793.950 757.050 796.050 ;
        RECT 661.950 790.950 664.050 793.050 ;
        RECT 662.400 772.050 663.600 790.950 ;
        RECT 755.400 778.050 756.600 793.950 ;
        RECT 920.400 793.050 921.600 802.950 ;
        RECT 907.950 790.950 910.050 793.050 ;
        RECT 919.950 790.950 922.050 793.050 ;
        RECT 908.400 784.050 909.600 790.950 ;
        RECT 805.950 781.950 808.050 784.050 ;
        RECT 907.950 781.950 910.050 784.050 ;
        RECT 806.400 778.050 807.600 781.950 ;
        RECT 754.950 775.950 757.050 778.050 ;
        RECT 805.800 775.950 807.900 778.050 ;
        RECT 616.950 769.950 619.050 772.050 ;
        RECT 622.950 769.950 625.050 772.050 ;
        RECT 661.950 769.950 664.050 772.050 ;
        RECT 623.400 733.050 624.600 769.950 ;
        RECT 622.950 730.950 625.050 733.050 ;
        RECT 613.950 721.950 616.050 724.050 ;
        RECT 614.400 700.050 615.600 721.950 ;
        RECT 613.950 697.950 616.050 700.050 ;
        RECT 628.950 697.950 631.050 700.050 ;
        RECT 629.400 678.900 630.600 697.950 ;
        RECT 634.950 679.950 637.050 682.050 ;
        RECT 635.400 678.900 636.600 679.950 ;
        RECT 628.950 676.800 631.050 678.900 ;
        RECT 634.950 676.800 637.050 678.900 ;
      LAYER metal3 ;
        RECT 568.950 840.600 571.050 841.200 ;
        RECT 574.950 840.600 577.050 841.050 ;
        RECT 568.950 839.400 577.050 840.600 ;
        RECT 568.950 839.100 571.050 839.400 ;
        RECT 574.950 838.950 577.050 839.400 ;
        RECT 574.950 807.600 577.050 808.050 ;
        RECT 730.950 807.750 733.050 808.200 ;
        RECT 742.950 807.750 745.050 808.200 ;
        RECT 574.950 806.400 588.600 807.600 ;
        RECT 574.950 805.950 577.050 806.400 ;
        RECT 587.400 804.600 588.600 806.400 ;
        RECT 730.950 806.550 745.050 807.750 ;
        RECT 730.950 806.100 733.050 806.550 ;
        RECT 742.950 806.100 745.050 806.550 ;
        RECT 919.950 804.600 922.050 805.050 ;
        RECT 926.400 804.600 927.600 807.600 ;
        RECT 587.400 804.000 618.450 804.600 ;
        RECT 587.400 803.400 619.050 804.000 ;
        RECT 616.950 802.050 619.050 803.400 ;
        RECT 919.950 803.400 927.600 804.600 ;
        RECT 919.950 802.950 922.050 803.400 ;
        RECT 616.800 801.000 619.050 802.050 ;
        RECT 616.800 799.950 618.900 801.000 ;
        RECT 730.950 795.600 733.050 796.050 ;
        RECT 754.950 795.600 757.050 796.050 ;
        RECT 713.400 794.400 757.050 795.600 ;
        RECT 661.950 792.600 664.050 793.050 ;
        RECT 713.400 792.600 714.600 794.400 ;
        RECT 730.950 793.950 733.050 794.400 ;
        RECT 754.950 793.950 757.050 794.400 ;
        RECT 661.950 791.400 714.600 792.600 ;
        RECT 907.950 792.600 910.050 793.050 ;
        RECT 919.950 792.600 922.050 793.050 ;
        RECT 907.950 791.400 922.050 792.600 ;
        RECT 661.950 790.950 664.050 791.400 ;
        RECT 907.950 790.950 910.050 791.400 ;
        RECT 919.950 790.950 922.050 791.400 ;
        RECT 805.950 783.600 808.050 784.050 ;
        RECT 907.950 783.600 910.050 784.050 ;
        RECT 805.950 782.400 910.050 783.600 ;
        RECT 805.950 781.950 808.050 782.400 ;
        RECT 907.950 781.950 910.050 782.400 ;
        RECT 754.950 777.600 757.050 778.050 ;
        RECT 805.800 777.600 807.900 778.050 ;
        RECT 754.950 776.400 807.900 777.600 ;
        RECT 754.950 775.950 757.050 776.400 ;
        RECT 805.800 775.950 807.900 776.400 ;
        RECT 616.950 771.600 619.050 772.050 ;
        RECT 622.950 771.600 625.050 772.050 ;
        RECT 661.950 771.600 664.050 772.050 ;
        RECT 616.950 770.400 664.050 771.600 ;
        RECT 616.950 769.950 619.050 770.400 ;
        RECT 622.950 769.950 625.050 770.400 ;
        RECT 661.950 769.950 664.050 770.400 ;
        RECT 613.950 699.600 616.050 700.050 ;
        RECT 628.950 699.600 631.050 700.050 ;
        RECT 613.950 698.400 631.050 699.600 ;
        RECT 613.950 697.950 616.050 698.400 ;
        RECT 628.950 697.950 631.050 698.400 ;
        RECT 628.950 678.450 631.050 678.900 ;
        RECT 634.950 678.450 637.050 678.900 ;
        RECT 628.950 677.250 637.050 678.450 ;
        RECT 628.950 676.800 631.050 677.250 ;
        RECT 634.950 676.800 637.050 677.250 ;
    END
  END ABCmd_i[1]
  PIN ABCmd_i[0]
    PORT
      LAYER metal1 ;
        RECT 655.950 840.450 658.050 841.050 ;
        RECT 655.950 839.550 666.450 840.450 ;
        RECT 655.950 838.950 658.050 839.550 ;
        RECT 665.550 835.050 666.450 839.550 ;
        RECT 665.550 833.550 670.050 835.050 ;
        RECT 666.000 832.950 670.050 833.550 ;
        RECT 696.000 762.450 700.050 763.050 ;
        RECT 695.550 760.950 700.050 762.450 ;
        RECT 695.550 757.050 696.450 760.950 ;
        RECT 695.550 755.550 700.050 757.050 ;
        RECT 696.000 754.950 700.050 755.550 ;
        RECT 699.000 729.450 703.050 730.050 ;
        RECT 698.550 727.950 703.050 729.450 ;
        RECT 698.550 724.050 699.450 727.950 ;
        RECT 694.950 722.550 699.450 724.050 ;
        RECT 694.950 721.950 699.000 722.550 ;
      LAYER metal2 ;
        RECT 466.950 913.950 469.050 916.050 ;
        RECT 467.400 897.600 468.600 913.950 ;
        RECT 464.400 896.400 468.600 897.600 ;
        RECT 457.950 880.950 460.050 883.050 ;
        RECT 458.400 865.050 459.600 880.950 ;
        RECT 464.400 865.050 465.600 896.400 ;
        RECT 655.950 868.950 658.050 871.050 ;
        RECT 457.950 862.950 460.050 865.050 ;
        RECT 463.950 862.950 466.050 865.050 ;
        RECT 484.950 862.950 487.050 865.050 ;
        RECT 589.950 862.950 592.050 865.050 ;
        RECT 604.950 862.950 607.050 865.050 ;
        RECT 485.400 853.050 486.600 862.950 ;
        RECT 590.400 853.050 591.600 862.950 ;
        RECT 484.950 850.950 487.050 853.050 ;
        RECT 589.950 850.950 592.050 853.050 ;
        RECT 485.400 838.050 486.600 850.950 ;
        RECT 605.400 847.050 606.600 862.950 ;
        RECT 656.400 847.050 657.600 868.950 ;
        RECT 766.950 865.950 769.050 868.050 ;
        RECT 767.400 847.050 768.600 865.950 ;
        RECT 793.950 859.950 796.050 862.050 ;
        RECT 794.400 847.050 795.600 859.950 ;
        RECT 919.950 853.950 922.050 856.050 ;
        RECT 604.950 844.950 607.050 847.050 ;
        RECT 655.950 844.950 658.050 847.050 ;
        RECT 766.950 844.950 769.050 847.050 ;
        RECT 793.950 844.950 796.050 847.050 ;
        RECT 656.400 841.050 657.600 844.950 ;
        RECT 655.950 838.950 658.050 841.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 667.950 832.950 670.050 835.050 ;
        RECT 668.400 826.050 669.600 832.950 ;
        RECT 680.400 826.050 681.600 835.950 ;
        RECT 667.950 823.950 670.050 826.050 ;
        RECT 679.950 823.950 682.050 826.050 ;
        RECT 680.400 817.050 681.600 823.950 ;
        RECT 679.950 814.950 682.050 817.050 ;
        RECT 706.950 814.950 709.050 817.050 ;
        RECT 707.400 807.600 708.600 814.950 ;
        RECT 920.400 811.050 921.600 853.950 ;
        RECT 919.950 808.950 922.050 811.050 ;
        RECT 707.400 806.400 711.600 807.600 ;
        RECT 710.400 784.050 711.600 806.400 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 755.400 801.600 756.600 802.950 ;
        RECT 755.400 800.400 759.600 801.600 ;
        RECT 758.400 790.050 759.600 800.400 ;
        RECT 745.950 787.950 748.050 790.050 ;
        RECT 757.950 787.950 760.050 790.050 ;
        RECT 746.400 784.050 747.600 787.950 ;
        RECT 697.950 781.950 700.050 784.050 ;
        RECT 709.950 781.950 712.050 784.050 ;
        RECT 745.950 781.950 748.050 784.050 ;
        RECT 698.400 763.050 699.600 781.950 ;
        RECT 697.950 760.950 700.050 763.050 ;
        RECT 697.950 754.950 700.050 757.050 ;
        RECT 698.400 738.600 699.600 754.950 ;
        RECT 698.400 737.400 702.600 738.600 ;
        RECT 701.400 730.050 702.600 737.400 ;
        RECT 700.950 727.950 703.050 730.050 ;
        RECT 694.950 721.950 697.050 724.050 ;
        RECT 695.400 709.050 696.600 721.950 ;
        RECT 676.950 706.950 679.050 709.050 ;
        RECT 694.950 706.950 697.050 709.050 ;
        RECT 677.400 688.050 678.600 706.950 ;
        RECT 676.950 685.950 679.050 688.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 584.400 673.050 585.600 679.950 ;
        RECT 656.400 678.900 657.600 679.950 ;
        RECT 655.950 676.800 658.050 678.900 ;
        RECT 583.950 670.950 586.050 673.050 ;
        RECT 601.950 670.950 604.050 673.050 ;
        RECT 602.400 667.050 603.600 670.950 ;
        RECT 656.400 667.050 657.600 676.800 ;
        RECT 601.950 664.950 604.050 667.050 ;
        RECT 655.950 664.950 658.050 667.050 ;
      LAYER metal3 ;
        RECT 655.950 870.600 658.050 871.050 ;
        RECT 655.950 869.400 738.600 870.600 ;
        RECT 655.950 868.950 658.050 869.400 ;
        RECT 737.400 867.600 738.600 869.400 ;
        RECT 766.950 867.600 769.050 868.050 ;
        RECT 737.400 866.400 769.050 867.600 ;
        RECT 766.950 865.950 769.050 866.400 ;
        RECT 457.950 864.600 460.050 865.050 ;
        RECT 463.950 864.600 466.050 865.050 ;
        RECT 484.950 864.600 487.050 865.050 ;
        RECT 457.950 863.400 487.050 864.600 ;
        RECT 457.950 862.950 460.050 863.400 ;
        RECT 463.950 862.950 466.050 863.400 ;
        RECT 484.950 862.950 487.050 863.400 ;
        RECT 589.950 864.600 592.050 865.050 ;
        RECT 604.950 864.600 607.050 865.050 ;
        RECT 589.950 863.400 607.050 864.600 ;
        RECT 589.950 862.950 592.050 863.400 ;
        RECT 604.950 862.950 607.050 863.400 ;
        RECT 793.950 861.600 796.050 862.050 ;
        RECT 793.950 860.400 834.600 861.600 ;
        RECT 793.950 859.950 796.050 860.400 ;
        RECT 833.400 858.600 834.600 860.400 ;
        RECT 833.400 857.400 918.600 858.600 ;
        RECT 917.400 856.050 918.600 857.400 ;
        RECT 917.400 854.400 922.050 856.050 ;
        RECT 918.000 853.950 922.050 854.400 ;
        RECT 484.950 852.600 487.050 853.050 ;
        RECT 589.950 852.600 592.050 853.050 ;
        RECT 484.950 851.400 592.050 852.600 ;
        RECT 484.950 850.950 487.050 851.400 ;
        RECT 589.950 850.950 592.050 851.400 ;
        RECT 604.950 846.600 607.050 847.050 ;
        RECT 655.950 846.600 658.050 847.050 ;
        RECT 604.950 845.400 658.050 846.600 ;
        RECT 604.950 844.950 607.050 845.400 ;
        RECT 655.950 844.950 658.050 845.400 ;
        RECT 766.950 846.600 769.050 847.050 ;
        RECT 793.950 846.600 796.050 847.050 ;
        RECT 766.950 845.400 796.050 846.600 ;
        RECT 766.950 844.950 769.050 845.400 ;
        RECT 793.950 844.950 796.050 845.400 ;
        RECT 667.950 825.600 670.050 826.050 ;
        RECT 679.950 825.600 682.050 826.050 ;
        RECT 667.950 824.400 682.050 825.600 ;
        RECT 667.950 823.950 670.050 824.400 ;
        RECT 679.950 823.950 682.050 824.400 ;
        RECT 679.950 816.600 682.050 817.050 ;
        RECT 706.950 816.600 709.050 817.050 ;
        RECT 679.950 815.400 709.050 816.600 ;
        RECT 679.950 814.950 682.050 815.400 ;
        RECT 706.950 814.950 709.050 815.400 ;
        RECT 919.950 810.600 922.050 811.050 ;
        RECT 919.950 809.400 930.600 810.600 ;
        RECT 919.950 808.950 922.050 809.400 ;
        RECT 929.400 801.600 930.600 809.400 ;
        RECT 926.400 800.400 930.600 801.600 ;
        RECT 745.950 789.600 748.050 790.050 ;
        RECT 757.950 789.600 760.050 790.050 ;
        RECT 745.950 788.400 760.050 789.600 ;
        RECT 745.950 787.950 748.050 788.400 ;
        RECT 757.950 787.950 760.050 788.400 ;
        RECT 697.950 783.600 700.050 784.050 ;
        RECT 709.950 783.600 712.050 784.050 ;
        RECT 745.950 783.600 748.050 784.050 ;
        RECT 697.950 782.400 748.050 783.600 ;
        RECT 697.950 781.950 700.050 782.400 ;
        RECT 709.950 781.950 712.050 782.400 ;
        RECT 745.950 781.950 748.050 782.400 ;
        RECT 676.950 708.600 679.050 709.050 ;
        RECT 694.950 708.600 697.050 709.050 ;
        RECT 676.950 707.400 697.050 708.600 ;
        RECT 676.950 706.950 679.050 707.400 ;
        RECT 694.950 706.950 697.050 707.400 ;
        RECT 676.950 687.600 679.050 688.050 ;
        RECT 659.400 686.400 679.050 687.600 ;
        RECT 659.400 681.600 660.600 686.400 ;
        RECT 676.950 685.950 679.050 686.400 ;
        RECT 656.400 680.400 660.600 681.600 ;
        RECT 656.400 678.900 657.600 680.400 ;
        RECT 655.950 676.800 658.050 678.900 ;
        RECT 583.950 672.600 586.050 673.050 ;
        RECT 601.950 672.600 604.050 673.050 ;
        RECT 583.950 671.400 604.050 672.600 ;
        RECT 583.950 670.950 586.050 671.400 ;
        RECT 601.950 670.950 604.050 671.400 ;
        RECT 601.950 666.600 604.050 667.050 ;
        RECT 655.950 666.600 658.050 667.050 ;
        RECT 601.950 665.400 658.050 666.600 ;
        RECT 601.950 664.950 604.050 665.400 ;
        RECT 655.950 664.950 658.050 665.400 ;
    END
  END ABCmd_i[0]
  PIN ACC_o[7]
    PORT
      LAYER metal2 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 701.400 -2.400 702.600 22.950 ;
        RECT 698.400 -3.600 702.600 -2.400 ;
    END
  END ACC_o[7]
  PIN ACC_o[6]
    PORT
      LAYER metal2 ;
        RECT 757.950 22.950 760.050 25.050 ;
        RECT 758.400 -2.400 759.600 22.950 ;
        RECT 755.400 -3.600 759.600 -2.400 ;
    END
  END ACC_o[6]
  PIN ACC_o[5]
    PORT
      LAYER metal2 ;
        RECT 811.950 22.950 814.050 25.050 ;
        RECT 812.400 -2.400 813.600 22.950 ;
        RECT 809.400 -3.600 813.600 -2.400 ;
    END
  END ACC_o[5]
  PIN ACC_o[4]
    PORT
      LAYER metal2 ;
        RECT 832.950 22.950 835.050 25.050 ;
        RECT 833.400 -2.400 834.600 22.950 ;
        RECT 830.400 -3.600 834.600 -2.400 ;
    END
  END ACC_o[4]
  PIN ACC_o[3]
    PORT
      LAYER metal2 ;
        RECT 850.950 22.950 853.050 25.050 ;
        RECT 851.400 -3.600 852.600 22.950 ;
    END
  END ACC_o[3]
  PIN ACC_o[2]
    PORT
      LAYER metal2 ;
        RECT 694.950 178.950 697.050 181.050 ;
        RECT 4.950 175.800 7.050 177.900 ;
        RECT 5.400 166.050 6.600 175.800 ;
        RECT 695.400 166.050 696.600 178.950 ;
        RECT 4.950 163.950 7.050 166.050 ;
        RECT 127.950 163.950 130.050 166.050 ;
        RECT 355.950 163.950 358.050 166.050 ;
        RECT 694.950 163.950 697.050 166.050 ;
        RECT 128.400 160.050 129.600 163.950 ;
        RECT 356.400 160.050 357.600 163.950 ;
        RECT 127.950 157.950 130.050 160.050 ;
        RECT 355.950 157.950 358.050 160.050 ;
      LAYER metal3 ;
        RECT 4.950 177.600 7.050 177.900 ;
        RECT -3.600 176.400 7.050 177.600 ;
        RECT 4.950 175.800 7.050 176.400 ;
        RECT 4.950 165.600 7.050 166.050 ;
        RECT 127.950 165.600 130.050 166.050 ;
        RECT 4.950 164.400 130.050 165.600 ;
        RECT 4.950 163.950 7.050 164.400 ;
        RECT 127.950 163.950 130.050 164.400 ;
        RECT 355.950 165.600 358.050 166.050 ;
        RECT 694.950 165.600 697.050 166.050 ;
        RECT 355.950 164.400 697.050 165.600 ;
        RECT 355.950 163.950 358.050 164.400 ;
        RECT 694.950 163.950 697.050 164.400 ;
        RECT 127.950 159.600 130.050 160.050 ;
        RECT 355.950 159.600 358.050 160.050 ;
        RECT 127.950 158.400 358.050 159.600 ;
        RECT 127.950 157.950 130.050 158.400 ;
        RECT 355.950 157.950 358.050 158.400 ;
    END
  END ACC_o[2]
  PIN ACC_o[1]
    PORT
      LAYER metal2 ;
        RECT 394.950 334.950 397.050 337.050 ;
        RECT 395.400 333.900 396.600 334.950 ;
        RECT 394.950 331.800 397.050 333.900 ;
        RECT 10.950 328.950 13.050 331.050 ;
        RECT 331.950 328.950 334.050 331.050 ;
        RECT 11.400 313.050 12.600 328.950 ;
        RECT 332.400 319.050 333.600 328.950 ;
        RECT 283.950 316.950 286.050 319.050 ;
        RECT 331.950 316.950 334.050 319.050 ;
        RECT 10.950 310.950 13.050 313.050 ;
        RECT 208.950 310.950 211.050 313.050 ;
        RECT 209.400 295.050 210.600 310.950 ;
        RECT 208.950 292.950 211.050 295.050 ;
        RECT 284.400 292.050 285.600 316.950 ;
        RECT 283.950 289.950 286.050 292.050 ;
      LAYER metal3 ;
        RECT 394.950 333.600 397.050 333.900 ;
        RECT -3.600 330.600 -2.400 333.600 ;
        RECT 332.400 333.000 397.050 333.600 ;
        RECT 331.950 332.400 397.050 333.000 ;
        RECT 10.950 330.600 13.050 331.050 ;
        RECT -3.600 329.400 13.050 330.600 ;
        RECT 10.950 328.950 13.050 329.400 ;
        RECT 331.950 328.950 334.050 332.400 ;
        RECT 394.950 331.800 397.050 332.400 ;
        RECT 283.950 318.600 286.050 319.050 ;
        RECT 331.950 318.600 334.050 319.050 ;
        RECT 283.950 317.400 334.050 318.600 ;
        RECT 283.950 316.950 286.050 317.400 ;
        RECT 331.950 316.950 334.050 317.400 ;
        RECT 10.950 312.600 13.050 313.050 ;
        RECT 208.950 312.600 211.050 313.050 ;
        RECT 10.950 311.400 211.050 312.600 ;
        RECT 10.950 310.950 13.050 311.400 ;
        RECT 208.950 310.950 211.050 311.400 ;
        RECT 208.950 291.600 211.050 295.050 ;
        RECT 283.950 291.600 286.050 292.050 ;
        RECT 208.950 291.000 286.050 291.600 ;
        RECT 209.400 290.400 286.050 291.000 ;
        RECT 283.950 289.950 286.050 290.400 ;
    END
  END ACC_o[1]
  PIN ACC_o[0]
    PORT
      LAYER metal1 ;
        RECT 322.950 303.450 325.050 304.050 ;
        RECT 331.950 303.450 334.050 304.050 ;
        RECT 322.950 302.550 334.050 303.450 ;
        RECT 322.950 301.950 325.050 302.550 ;
        RECT 331.950 301.950 334.050 302.550 ;
      LAYER metal2 ;
        RECT 4.950 337.950 7.050 340.050 ;
        RECT 5.400 316.050 6.600 337.950 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 497.400 319.050 498.600 334.950 ;
        RECT 241.950 316.800 244.050 318.900 ;
        RECT 376.950 316.950 379.050 319.050 ;
        RECT 496.950 316.950 499.050 319.050 ;
        RECT 4.950 313.950 7.050 316.050 ;
        RECT 242.400 307.050 243.600 316.800 ;
        RECT 304.950 310.950 307.050 313.050 ;
        RECT 313.800 310.950 315.900 313.050 ;
        RECT 305.400 307.050 306.600 310.950 ;
        RECT 314.400 307.050 315.600 310.950 ;
        RECT 377.400 310.050 378.600 316.950 ;
        RECT 367.950 307.050 370.050 310.050 ;
        RECT 376.950 307.950 379.050 310.050 ;
        RECT 241.950 304.950 244.050 307.050 ;
        RECT 304.950 304.950 307.050 307.050 ;
        RECT 313.950 304.950 316.050 307.050 ;
        RECT 322.950 301.950 325.050 307.050 ;
        RECT 331.950 301.950 334.050 307.050 ;
        RECT 364.950 306.000 370.050 307.050 ;
        RECT 364.950 305.400 369.600 306.000 ;
        RECT 364.950 304.950 369.000 305.400 ;
      LAYER metal3 ;
        RECT 4.950 339.600 7.050 340.050 ;
        RECT -3.600 338.400 7.050 339.600 ;
        RECT 4.950 337.950 7.050 338.400 ;
        RECT 241.950 318.600 244.050 318.900 ;
        RECT 215.400 317.400 244.050 318.600 ;
        RECT 4.950 315.600 7.050 316.050 ;
        RECT 215.400 315.600 216.600 317.400 ;
        RECT 241.950 316.800 244.050 317.400 ;
        RECT 376.950 318.600 379.050 319.050 ;
        RECT 496.950 318.600 499.050 319.050 ;
        RECT 376.950 317.400 499.050 318.600 ;
        RECT 376.950 316.950 379.050 317.400 ;
        RECT 496.950 316.950 499.050 317.400 ;
        RECT 4.950 314.400 216.600 315.600 ;
        RECT 4.950 313.950 7.050 314.400 ;
        RECT 304.950 312.600 307.050 313.050 ;
        RECT 313.800 312.600 315.900 313.050 ;
        RECT 304.950 311.400 315.900 312.600 ;
        RECT 304.950 310.950 307.050 311.400 ;
        RECT 313.800 310.950 315.900 311.400 ;
        RECT 367.950 309.600 370.050 310.050 ;
        RECT 376.950 309.600 379.050 310.050 ;
        RECT 367.950 308.400 379.050 309.600 ;
        RECT 367.950 307.950 370.050 308.400 ;
        RECT 376.950 307.950 379.050 308.400 ;
        RECT 241.950 306.600 244.050 307.050 ;
        RECT 304.950 306.600 307.050 307.050 ;
        RECT 241.950 305.400 307.050 306.600 ;
        RECT 241.950 304.950 244.050 305.400 ;
        RECT 304.950 304.950 307.050 305.400 ;
        RECT 313.950 306.600 316.050 307.050 ;
        RECT 322.950 306.600 325.050 307.050 ;
        RECT 313.950 305.400 325.050 306.600 ;
        RECT 313.950 304.950 316.050 305.400 ;
        RECT 322.950 304.950 325.050 305.400 ;
        RECT 331.950 306.600 334.050 307.050 ;
        RECT 364.950 306.600 367.050 307.050 ;
        RECT 331.950 305.400 367.050 306.600 ;
        RECT 331.950 304.950 334.050 305.400 ;
        RECT 364.950 304.950 367.050 305.400 ;
    END
  END ACC_o[0]
  PIN Done_o
    PORT
      LAYER metal2 ;
        RECT 871.950 22.950 874.050 25.050 ;
        RECT 872.400 -2.400 873.600 22.950 ;
        RECT 869.400 -3.600 873.600 -2.400 ;
    END
  END Done_o
  PIN LoadA_i
    PORT
      LAYER metal1 ;
        RECT 844.950 480.450 847.050 480.900 ;
        RECT 850.950 480.450 853.050 481.050 ;
        RECT 844.950 479.550 853.050 480.450 ;
        RECT 844.950 478.800 847.050 479.550 ;
        RECT 850.950 478.950 853.050 479.550 ;
        RECT 849.000 417.450 853.050 418.050 ;
        RECT 848.550 415.950 853.050 417.450 ;
        RECT 848.550 412.050 849.450 415.950 ;
        RECT 848.550 410.550 853.050 412.050 ;
        RECT 849.000 409.950 853.050 410.550 ;
        RECT 850.950 372.450 855.000 373.050 ;
        RECT 850.950 370.950 855.450 372.450 ;
        RECT 854.550 367.050 855.450 370.950 ;
        RECT 854.550 365.550 859.050 367.050 ;
        RECT 855.000 364.950 859.050 365.550 ;
      LAYER metal2 ;
        RECT 890.400 934.050 891.600 945.600 ;
        RECT 883.950 931.950 886.050 934.050 ;
        RECT 889.950 931.950 892.050 934.050 ;
        RECT 884.400 877.050 885.600 931.950 ;
        RECT 883.950 874.950 886.050 877.050 ;
        RECT 892.950 874.950 895.050 877.050 ;
        RECT 893.400 829.050 894.600 874.950 ;
        RECT 880.950 826.950 883.050 829.050 ;
        RECT 892.950 826.950 895.050 829.050 ;
        RECT 881.400 787.050 882.600 826.950 ;
        RECT 865.950 784.950 868.050 787.050 ;
        RECT 880.950 784.950 883.050 787.050 ;
        RECT 866.400 756.600 867.600 784.950 ;
        RECT 863.400 755.400 867.600 756.600 ;
        RECT 863.400 745.050 864.600 755.400 ;
        RECT 853.950 742.950 856.050 745.050 ;
        RECT 862.950 742.950 865.050 745.050 ;
        RECT 854.400 730.050 855.600 742.950 ;
        RECT 853.950 727.950 856.050 730.050 ;
        RECT 853.950 721.950 856.050 724.050 ;
        RECT 854.400 717.600 855.600 721.950 ;
        RECT 851.400 716.400 855.600 717.600 ;
        RECT 851.400 652.050 852.600 716.400 ;
        RECT 850.950 649.950 853.050 652.050 ;
        RECT 850.950 643.950 853.050 646.050 ;
        RECT 851.400 637.050 852.600 643.950 ;
        RECT 838.950 634.950 841.050 637.050 ;
        RECT 850.950 634.950 853.050 637.050 ;
        RECT 839.400 601.050 840.600 634.950 ;
        RECT 838.950 598.950 841.050 601.050 ;
        RECT 853.950 598.950 856.050 601.050 ;
        RECT 854.400 567.600 855.600 598.950 ;
        RECT 851.400 566.400 855.600 567.600 ;
        RECT 851.400 481.050 852.600 566.400 ;
        RECT 844.950 478.800 847.050 480.900 ;
        RECT 850.950 478.950 853.050 481.050 ;
        RECT 845.400 445.050 846.600 478.800 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 844.950 442.950 847.050 445.050 ;
        RECT 857.400 444.900 858.600 445.950 ;
        RECT 856.950 442.800 859.050 444.900 ;
        RECT 857.400 441.600 858.600 442.800 ;
        RECT 854.400 440.400 858.600 441.600 ;
        RECT 854.400 420.600 855.600 440.400 ;
        RECT 851.400 420.000 855.600 420.600 ;
        RECT 850.950 419.400 855.600 420.000 ;
        RECT 850.950 415.950 853.050 419.400 ;
        RECT 850.950 409.950 853.050 412.050 ;
        RECT 851.400 373.050 852.600 409.950 ;
        RECT 850.950 370.950 853.050 373.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 848.400 361.050 849.600 367.950 ;
        RECT 856.950 364.950 859.050 367.050 ;
        RECT 857.400 361.050 858.600 364.950 ;
        RECT 847.950 358.950 850.050 361.050 ;
        RECT 856.950 358.950 859.050 361.050 ;
        RECT 874.950 358.950 877.050 361.050 ;
        RECT 875.400 337.050 876.600 358.950 ;
        RECT 874.950 334.950 877.050 337.050 ;
      LAYER metal3 ;
        RECT 883.950 933.600 886.050 934.050 ;
        RECT 889.950 933.600 892.050 934.050 ;
        RECT 883.950 932.400 892.050 933.600 ;
        RECT 883.950 931.950 886.050 932.400 ;
        RECT 889.950 931.950 892.050 932.400 ;
        RECT 883.950 876.600 886.050 877.050 ;
        RECT 892.950 876.600 895.050 877.050 ;
        RECT 883.950 875.400 895.050 876.600 ;
        RECT 883.950 874.950 886.050 875.400 ;
        RECT 892.950 874.950 895.050 875.400 ;
        RECT 880.950 828.600 883.050 829.050 ;
        RECT 892.950 828.600 895.050 829.050 ;
        RECT 880.950 827.400 895.050 828.600 ;
        RECT 880.950 826.950 883.050 827.400 ;
        RECT 892.950 826.950 895.050 827.400 ;
        RECT 865.950 786.600 868.050 787.050 ;
        RECT 880.950 786.600 883.050 787.050 ;
        RECT 865.950 785.400 883.050 786.600 ;
        RECT 865.950 784.950 868.050 785.400 ;
        RECT 880.950 784.950 883.050 785.400 ;
        RECT 853.950 744.600 856.050 745.050 ;
        RECT 862.950 744.600 865.050 745.050 ;
        RECT 853.950 743.400 865.050 744.600 ;
        RECT 853.950 742.950 856.050 743.400 ;
        RECT 862.950 742.950 865.050 743.400 ;
        RECT 853.950 727.950 856.050 730.050 ;
        RECT 854.400 724.050 855.600 727.950 ;
        RECT 853.950 721.950 856.050 724.050 ;
        RECT 850.950 649.950 853.050 652.050 ;
        RECT 851.400 646.050 852.600 649.950 ;
        RECT 850.950 643.950 853.050 646.050 ;
        RECT 838.950 636.600 841.050 637.050 ;
        RECT 850.950 636.600 853.050 637.050 ;
        RECT 838.950 635.400 853.050 636.600 ;
        RECT 838.950 634.950 841.050 635.400 ;
        RECT 850.950 634.950 853.050 635.400 ;
        RECT 838.950 600.600 841.050 601.050 ;
        RECT 853.950 600.600 856.050 601.050 ;
        RECT 838.950 599.400 856.050 600.600 ;
        RECT 838.950 598.950 841.050 599.400 ;
        RECT 853.950 598.950 856.050 599.400 ;
        RECT 844.950 444.600 847.050 445.050 ;
        RECT 856.950 444.600 859.050 444.900 ;
        RECT 844.950 443.400 859.050 444.600 ;
        RECT 844.950 442.950 847.050 443.400 ;
        RECT 856.950 442.800 859.050 443.400 ;
        RECT 847.950 360.600 850.050 361.050 ;
        RECT 856.950 360.600 859.050 361.050 ;
        RECT 874.950 360.600 877.050 361.050 ;
        RECT 847.950 359.400 877.050 360.600 ;
        RECT 847.950 358.950 850.050 359.400 ;
        RECT 856.950 358.950 859.050 359.400 ;
        RECT 874.950 358.950 877.050 359.400 ;
    END
  END LoadA_i
  PIN LoadB_i
    PORT
      LAYER metal1 ;
        RECT 885.000 918.450 889.050 919.050 ;
        RECT 884.550 916.950 889.050 918.450 ;
        RECT 884.550 913.050 885.450 916.950 ;
        RECT 884.550 911.550 889.050 913.050 ;
        RECT 885.000 910.950 889.050 911.550 ;
      LAYER metal2 ;
        RECT 884.400 944.400 888.600 945.600 ;
        RECT 887.400 919.050 888.600 944.400 ;
        RECT 886.950 916.950 889.050 919.050 ;
        RECT 886.950 910.950 889.050 913.050 ;
        RECT 887.400 834.600 888.600 910.950 ;
        RECT 884.400 833.400 888.600 834.600 ;
        RECT 884.400 796.050 885.600 833.400 ;
        RECT 871.950 793.950 874.050 796.050 ;
        RECT 883.950 793.950 886.050 796.050 ;
        RECT 872.400 745.050 873.600 793.950 ;
        RECT 871.950 742.950 874.050 745.050 ;
        RECT 880.950 742.950 883.050 745.050 ;
        RECT 881.400 676.050 882.600 742.950 ;
        RECT 874.950 673.950 877.050 676.050 ;
        RECT 880.950 673.950 883.050 676.050 ;
        RECT 875.400 645.600 876.600 673.950 ;
        RECT 872.400 644.400 876.600 645.600 ;
        RECT 872.400 640.050 873.600 644.400 ;
        RECT 871.950 637.950 874.050 640.050 ;
        RECT 877.950 637.950 880.050 640.050 ;
        RECT 878.400 577.050 879.600 637.950 ;
        RECT 856.950 574.800 859.050 576.900 ;
        RECT 877.950 574.950 880.050 577.050 ;
        RECT 857.400 564.600 858.600 574.800 ;
        RECT 854.400 563.400 858.600 564.600 ;
        RECT 854.400 529.050 855.600 563.400 ;
        RECT 853.950 526.950 856.050 529.050 ;
        RECT 853.950 520.950 856.050 523.050 ;
        RECT 854.400 487.050 855.600 520.950 ;
        RECT 853.950 484.950 856.050 487.050 ;
        RECT 865.950 484.950 868.050 487.050 ;
        RECT 866.400 451.050 867.600 484.950 ;
        RECT 865.950 448.950 868.050 451.050 ;
        RECT 865.950 442.950 868.050 445.050 ;
        RECT 866.400 421.050 867.600 442.950 ;
        RECT 865.950 418.950 868.050 421.050 ;
        RECT 877.950 416.100 880.050 418.200 ;
        RECT 878.400 415.050 879.600 416.100 ;
        RECT 877.950 412.950 880.050 415.050 ;
        RECT 844.950 409.950 847.050 412.050 ;
        RECT 845.400 376.050 846.600 409.950 ;
        RECT 844.950 372.000 847.050 376.050 ;
        RECT 853.950 373.950 856.050 376.050 ;
        RECT 845.400 370.050 846.600 372.000 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 854.400 364.050 855.600 373.950 ;
        RECT 859.950 372.000 862.050 376.050 ;
        RECT 860.400 370.050 861.600 372.000 ;
        RECT 859.950 367.950 862.050 370.050 ;
        RECT 853.950 361.950 856.050 364.050 ;
        RECT 859.950 361.950 862.050 364.050 ;
        RECT 860.400 342.600 861.600 361.950 ;
        RECT 860.400 341.400 864.600 342.600 ;
        RECT 863.400 337.050 864.600 341.400 ;
        RECT 862.950 334.950 865.050 337.050 ;
      LAYER metal3 ;
        RECT 871.950 795.600 874.050 796.050 ;
        RECT 883.950 795.600 886.050 796.050 ;
        RECT 871.950 794.400 886.050 795.600 ;
        RECT 871.950 793.950 874.050 794.400 ;
        RECT 883.950 793.950 886.050 794.400 ;
        RECT 871.950 744.600 874.050 745.050 ;
        RECT 880.950 744.600 883.050 745.050 ;
        RECT 871.950 743.400 883.050 744.600 ;
        RECT 871.950 742.950 874.050 743.400 ;
        RECT 880.950 742.950 883.050 743.400 ;
        RECT 874.950 675.600 877.050 676.050 ;
        RECT 880.950 675.600 883.050 676.050 ;
        RECT 874.950 674.400 883.050 675.600 ;
        RECT 874.950 673.950 877.050 674.400 ;
        RECT 880.950 673.950 883.050 674.400 ;
        RECT 871.950 639.600 874.050 640.050 ;
        RECT 877.950 639.600 880.050 640.050 ;
        RECT 871.950 638.400 880.050 639.600 ;
        RECT 871.950 637.950 874.050 638.400 ;
        RECT 877.950 637.950 880.050 638.400 ;
        RECT 856.950 576.600 859.050 576.900 ;
        RECT 877.950 576.600 880.050 577.050 ;
        RECT 856.950 575.400 880.050 576.600 ;
        RECT 856.950 574.800 859.050 575.400 ;
        RECT 877.950 574.950 880.050 575.400 ;
        RECT 853.950 526.950 856.050 529.050 ;
        RECT 854.400 523.050 855.600 526.950 ;
        RECT 853.950 520.950 856.050 523.050 ;
        RECT 853.950 486.600 856.050 487.050 ;
        RECT 865.950 486.600 868.050 487.050 ;
        RECT 853.950 485.400 868.050 486.600 ;
        RECT 853.950 484.950 856.050 485.400 ;
        RECT 865.950 484.950 868.050 485.400 ;
        RECT 865.950 448.950 868.050 451.050 ;
        RECT 866.400 445.050 867.600 448.950 ;
        RECT 865.950 442.950 868.050 445.050 ;
        RECT 865.950 417.600 868.050 421.050 ;
        RECT 877.950 417.600 880.050 418.200 ;
        RECT 865.950 417.000 880.050 417.600 ;
        RECT 866.400 416.400 880.050 417.000 ;
        RECT 866.400 414.600 867.600 416.400 ;
        RECT 877.950 416.100 880.050 416.400 ;
        RECT 845.400 414.000 867.600 414.600 ;
        RECT 844.950 413.400 867.600 414.000 ;
        RECT 844.950 409.950 847.050 413.400 ;
        RECT 844.950 375.600 847.050 376.050 ;
        RECT 853.950 375.600 856.050 376.050 ;
        RECT 859.950 375.600 862.050 376.050 ;
        RECT 844.950 374.400 862.050 375.600 ;
        RECT 844.950 373.950 847.050 374.400 ;
        RECT 853.950 373.950 856.050 374.400 ;
        RECT 859.950 373.950 862.050 374.400 ;
        RECT 853.950 363.600 856.050 364.050 ;
        RECT 859.950 363.600 862.050 364.050 ;
        RECT 853.950 362.400 862.050 363.600 ;
        RECT 853.950 361.950 856.050 362.400 ;
        RECT 859.950 361.950 862.050 362.400 ;
    END
  END LoadB_i
  PIN LoadCmd_i
    PORT
      LAYER metal1 ;
        RECT 877.950 723.450 880.050 724.050 ;
        RECT 883.950 723.450 886.050 724.050 ;
        RECT 877.950 722.550 886.050 723.450 ;
        RECT 877.950 721.950 880.050 722.550 ;
        RECT 883.950 721.950 886.050 722.550 ;
      LAYER metal2 ;
        RECT 878.400 940.050 879.600 945.600 ;
        RECT 877.950 937.950 880.050 940.050 ;
        RECT 910.950 937.950 913.050 940.050 ;
        RECT 911.400 835.050 912.600 937.950 ;
        RECT 901.950 832.950 904.050 835.050 ;
        RECT 910.950 832.950 913.050 835.050 ;
        RECT 902.400 793.050 903.600 832.950 ;
        RECT 868.950 790.950 871.050 793.050 ;
        RECT 901.950 790.950 904.050 793.050 ;
        RECT 869.400 742.050 870.600 790.950 ;
        RECT 868.950 739.950 871.050 742.050 ;
        RECT 883.950 739.950 886.050 742.050 ;
        RECT 884.400 724.050 885.600 739.950 ;
        RECT 877.950 721.950 880.050 724.050 ;
        RECT 883.950 721.950 886.050 724.050 ;
        RECT 878.400 642.600 879.600 721.950 ;
        RECT 875.400 641.400 879.600 642.600 ;
        RECT 875.400 592.050 876.600 641.400 ;
        RECT 874.950 589.950 877.050 592.050 ;
        RECT 895.950 589.950 898.050 592.050 ;
        RECT 892.950 420.600 895.050 421.050 ;
        RECT 896.400 420.600 897.600 589.950 ;
        RECT 892.950 419.400 897.600 420.600 ;
        RECT 892.950 418.950 895.050 419.400 ;
        RECT 893.400 411.600 894.600 418.950 ;
        RECT 898.950 417.000 901.050 421.050 ;
        RECT 899.400 415.050 900.600 417.000 ;
        RECT 898.950 412.950 901.050 415.050 ;
        RECT 893.400 410.400 897.600 411.600 ;
        RECT 889.950 367.950 892.050 370.050 ;
        RECT 890.400 366.900 891.600 367.950 ;
        RECT 896.400 367.050 897.600 410.400 ;
        RECT 889.950 364.800 892.050 366.900 ;
        RECT 895.800 364.950 897.900 367.050 ;
      LAYER metal3 ;
        RECT 877.950 939.600 880.050 940.050 ;
        RECT 910.950 939.600 913.050 940.050 ;
        RECT 877.950 938.400 913.050 939.600 ;
        RECT 877.950 937.950 880.050 938.400 ;
        RECT 910.950 937.950 913.050 938.400 ;
        RECT 901.950 834.600 904.050 835.050 ;
        RECT 910.950 834.600 913.050 835.050 ;
        RECT 901.950 833.400 913.050 834.600 ;
        RECT 901.950 832.950 904.050 833.400 ;
        RECT 910.950 832.950 913.050 833.400 ;
        RECT 868.950 792.600 871.050 793.050 ;
        RECT 901.950 792.600 904.050 793.050 ;
        RECT 868.950 791.400 904.050 792.600 ;
        RECT 868.950 790.950 871.050 791.400 ;
        RECT 901.950 790.950 904.050 791.400 ;
        RECT 868.950 741.600 871.050 742.050 ;
        RECT 883.950 741.600 886.050 742.050 ;
        RECT 868.950 740.400 886.050 741.600 ;
        RECT 868.950 739.950 871.050 740.400 ;
        RECT 883.950 739.950 886.050 740.400 ;
        RECT 874.950 591.600 877.050 592.050 ;
        RECT 895.950 591.600 898.050 592.050 ;
        RECT 874.950 590.400 898.050 591.600 ;
        RECT 874.950 589.950 877.050 590.400 ;
        RECT 895.950 589.950 898.050 590.400 ;
        RECT 892.950 420.600 895.050 421.050 ;
        RECT 898.950 420.600 901.050 421.050 ;
        RECT 892.950 419.400 901.050 420.600 ;
        RECT 892.950 418.950 895.050 419.400 ;
        RECT 898.950 418.950 901.050 419.400 ;
        RECT 889.950 366.600 892.050 366.900 ;
        RECT 895.800 366.600 897.900 367.050 ;
        RECT 889.950 365.400 897.900 366.600 ;
        RECT 889.950 364.800 892.050 365.400 ;
        RECT 895.800 364.950 897.900 365.400 ;
    END
  END LoadCmd_i
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 781.950 261.450 786.000 262.050 ;
        RECT 781.950 259.950 786.450 261.450 ;
        RECT 785.550 256.050 786.450 259.950 ;
        RECT 785.550 254.550 790.050 256.050 ;
        RECT 786.000 253.950 790.050 254.550 ;
      LAYER metal2 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 707.400 567.900 708.600 568.950 ;
        RECT 706.950 565.800 709.050 567.900 ;
        RECT 733.950 565.800 736.050 567.900 ;
        RECT 734.400 541.050 735.600 565.800 ;
        RECT 803.400 562.050 804.600 568.950 ;
        RECT 790.950 559.950 793.050 562.050 ;
        RECT 802.950 559.950 805.050 562.050 ;
        RECT 791.400 541.050 792.600 559.950 ;
        RECT 733.950 538.950 736.050 541.050 ;
        RECT 790.950 538.950 793.050 541.050 ;
        RECT 791.400 514.050 792.600 538.950 ;
        RECT 790.950 511.950 793.050 514.050 ;
        RECT 808.950 511.950 811.050 514.050 ;
        RECT 809.400 478.050 810.600 511.950 ;
        RECT 796.950 475.950 799.050 478.050 ;
        RECT 808.950 475.950 811.050 478.050 ;
        RECT 797.400 451.200 798.600 475.950 ;
        RECT 769.950 449.100 772.050 451.200 ;
        RECT 796.950 449.100 799.050 451.200 ;
        RECT 770.400 448.050 771.600 449.100 ;
        RECT 769.950 445.950 772.050 448.050 ;
        RECT 797.400 430.050 798.600 449.100 ;
        RECT 796.950 427.950 799.050 430.050 ;
        RECT 808.950 427.950 811.050 430.050 ;
        RECT 809.400 366.600 810.600 427.950 ;
        RECT 806.400 365.400 810.600 366.600 ;
        RECT 806.400 328.050 807.600 365.400 ;
        RECT 790.950 325.950 793.050 328.050 ;
        RECT 805.950 325.950 808.050 328.050 ;
        RECT 791.400 295.050 792.600 325.950 ;
        RECT 790.800 292.950 792.900 295.050 ;
        RECT 781.950 286.950 784.050 289.050 ;
        RECT 782.400 262.050 783.600 286.950 ;
        RECT 781.950 259.950 784.050 262.050 ;
        RECT 787.950 253.950 790.050 256.050 ;
        RECT 788.400 217.050 789.600 253.950 ;
        RECT 787.950 214.950 790.050 217.050 ;
        RECT 766.950 208.950 769.050 211.050 ;
        RECT 767.400 163.050 768.600 208.950 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 773.400 163.050 774.600 178.950 ;
        RECT 766.950 160.950 769.050 163.050 ;
        RECT 772.950 160.950 775.050 163.050 ;
        RECT 877.950 160.950 880.050 163.050 ;
        RECT 878.400 151.050 879.600 160.950 ;
        RECT 877.950 148.950 880.050 151.050 ;
        RECT 898.950 148.950 901.050 151.050 ;
        RECT 899.400 139.200 900.600 148.950 ;
        RECT 898.950 137.100 901.050 139.200 ;
        RECT 899.400 136.050 900.600 137.100 ;
        RECT 898.950 133.950 901.050 136.050 ;
      LAYER metal3 ;
        RECT 706.950 567.450 709.050 567.900 ;
        RECT 733.950 567.450 736.050 567.900 ;
        RECT 706.950 566.250 736.050 567.450 ;
        RECT 706.950 565.800 709.050 566.250 ;
        RECT 733.950 565.800 736.050 566.250 ;
        RECT 790.950 561.600 793.050 562.050 ;
        RECT 802.950 561.600 805.050 562.050 ;
        RECT 790.950 560.400 805.050 561.600 ;
        RECT 790.950 559.950 793.050 560.400 ;
        RECT 802.950 559.950 805.050 560.400 ;
        RECT 733.950 540.600 736.050 541.050 ;
        RECT 790.950 540.600 793.050 541.050 ;
        RECT 733.950 539.400 793.050 540.600 ;
        RECT 733.950 538.950 736.050 539.400 ;
        RECT 790.950 538.950 793.050 539.400 ;
        RECT 790.950 513.600 793.050 514.050 ;
        RECT 808.950 513.600 811.050 514.050 ;
        RECT 790.950 512.400 811.050 513.600 ;
        RECT 790.950 511.950 793.050 512.400 ;
        RECT 808.950 511.950 811.050 512.400 ;
        RECT 796.950 477.600 799.050 478.050 ;
        RECT 808.950 477.600 811.050 478.050 ;
        RECT 796.950 476.400 811.050 477.600 ;
        RECT 796.950 475.950 799.050 476.400 ;
        RECT 808.950 475.950 811.050 476.400 ;
        RECT 769.950 450.750 772.050 451.200 ;
        RECT 796.950 450.750 799.050 451.200 ;
        RECT 769.950 449.550 799.050 450.750 ;
        RECT 769.950 449.100 772.050 449.550 ;
        RECT 796.950 449.100 799.050 449.550 ;
        RECT 796.950 429.600 799.050 430.050 ;
        RECT 808.950 429.600 811.050 430.050 ;
        RECT 796.950 428.400 811.050 429.600 ;
        RECT 796.950 427.950 799.050 428.400 ;
        RECT 808.950 427.950 811.050 428.400 ;
        RECT 790.950 327.600 793.050 328.050 ;
        RECT 805.950 327.600 808.050 328.050 ;
        RECT 790.950 326.400 808.050 327.600 ;
        RECT 790.950 325.950 793.050 326.400 ;
        RECT 805.950 325.950 808.050 326.400 ;
        RECT 790.800 292.950 792.900 295.050 ;
        RECT 781.950 288.600 784.050 289.050 ;
        RECT 791.250 288.600 792.450 292.950 ;
        RECT 781.950 287.400 792.450 288.600 ;
        RECT 781.950 286.950 784.050 287.400 ;
        RECT 787.950 214.950 790.050 217.050 ;
        RECT 766.950 210.600 769.050 211.050 ;
        RECT 788.400 210.600 789.600 214.950 ;
        RECT 766.950 209.400 789.600 210.600 ;
        RECT 766.950 208.950 769.050 209.400 ;
        RECT 766.950 162.600 769.050 163.050 ;
        RECT 772.950 162.600 775.050 163.050 ;
        RECT 877.950 162.600 880.050 163.050 ;
        RECT 766.950 161.400 880.050 162.600 ;
        RECT 766.950 160.950 769.050 161.400 ;
        RECT 772.950 160.950 775.050 161.400 ;
        RECT 877.950 160.950 880.050 161.400 ;
        RECT 877.950 150.600 880.050 151.050 ;
        RECT 898.950 150.600 901.050 151.050 ;
        RECT 877.950 149.400 901.050 150.600 ;
        RECT 877.950 148.950 880.050 149.400 ;
        RECT 898.950 148.950 901.050 149.400 ;
        RECT 898.950 138.600 901.050 139.200 ;
        RECT 898.950 137.400 927.600 138.600 ;
        RECT 898.950 137.100 901.050 137.400 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal2 ;
        RECT 904.950 211.950 907.050 214.050 ;
        RECT 905.400 210.900 906.600 211.950 ;
        RECT 904.950 208.800 907.050 210.900 ;
      LAYER metal3 ;
        RECT 904.950 210.600 907.050 210.900 ;
        RECT 926.400 210.600 927.600 216.600 ;
        RECT 904.950 209.400 927.600 210.600 ;
        RECT 904.950 208.800 907.050 209.400 ;
    END
  END reset
  OBS
      LAYER metal1 ;
        RECT 13.800 929.400 15.600 935.400 ;
        RECT 35.400 929.400 37.200 935.400 ;
        RECT 56.400 929.400 58.200 935.400 ;
        RECT 76.800 929.400 78.600 935.400 ;
        RECT 94.800 929.400 96.600 935.400 ;
        RECT 14.400 916.050 15.600 929.400 ;
        RECT 17.100 916.050 18.900 917.850 ;
        RECT 35.850 916.050 37.050 929.400 ;
        RECT 41.100 916.050 42.900 917.850 ;
        RECT 56.850 916.050 58.050 929.400 ;
        RECT 62.100 916.050 63.900 917.850 ;
        RECT 77.400 916.050 78.600 929.400 ;
        RECT 95.700 929.100 96.600 929.400 ;
        RECT 100.800 929.400 102.600 935.400 ;
        RECT 116.400 929.400 118.200 935.400 ;
        RECT 100.800 929.100 102.300 929.400 ;
        RECT 95.700 928.200 102.300 929.100 ;
        RECT 116.700 929.100 118.200 929.400 ;
        RECT 122.400 929.400 124.200 935.400 ;
        RECT 140.400 929.400 142.200 935.400 ;
        RECT 160.800 929.400 162.600 935.400 ;
        RECT 122.400 929.100 123.300 929.400 ;
        RECT 116.700 928.200 123.300 929.100 ;
        RECT 80.100 916.050 81.900 917.850 ;
        RECT 95.700 916.050 96.600 928.200 ;
        RECT 101.100 916.050 102.900 917.850 ;
        RECT 116.100 916.050 117.900 917.850 ;
        RECT 122.400 916.050 123.300 928.200 ;
        RECT 140.850 916.050 142.050 929.400 ;
        RECT 161.700 929.100 162.600 929.400 ;
        RECT 166.800 929.400 168.600 935.400 ;
        RECT 184.800 929.400 186.600 935.400 ;
        RECT 203.400 929.400 205.200 935.400 ;
        RECT 224.400 929.400 226.200 935.400 ;
        RECT 166.800 929.100 168.300 929.400 ;
        RECT 161.700 928.200 168.300 929.100 ;
        RECT 146.100 916.050 147.900 917.850 ;
        RECT 161.700 916.050 162.600 928.200 ;
        RECT 167.100 916.050 168.900 917.850 ;
        RECT 185.400 916.050 186.600 929.400 ;
        RECT 188.100 916.050 189.900 917.850 ;
        RECT 203.850 916.050 205.050 929.400 ;
        RECT 224.700 929.100 226.200 929.400 ;
        RECT 230.400 929.400 232.200 935.400 ;
        RECT 230.400 929.100 231.300 929.400 ;
        RECT 224.700 928.200 231.300 929.100 ;
        RECT 209.100 916.050 210.900 917.850 ;
        RECT 224.100 916.050 225.900 917.850 ;
        RECT 230.400 916.050 231.300 928.200 ;
        RECT 244.800 923.400 246.600 935.400 ;
        RECT 247.800 924.300 249.600 935.400 ;
        RECT 253.800 924.300 255.600 935.400 ;
        RECT 269.400 929.400 271.200 935.400 ;
        RECT 269.700 929.100 271.200 929.400 ;
        RECT 275.400 929.400 277.200 935.400 ;
        RECT 295.800 929.400 297.600 935.400 ;
        RECT 314.400 929.400 316.200 935.400 ;
        RECT 275.400 929.100 276.300 929.400 ;
        RECT 269.700 928.200 276.300 929.100 ;
        RECT 247.800 923.400 255.600 924.300 ;
        RECT 245.400 916.050 246.300 923.400 ;
        RECT 251.100 916.050 252.900 917.850 ;
        RECT 269.100 916.050 270.900 917.850 ;
        RECT 275.400 916.050 276.300 928.200 ;
        RECT 296.400 916.050 297.600 929.400 ;
        RECT 314.700 929.100 316.200 929.400 ;
        RECT 320.400 929.400 322.200 935.400 ;
        RECT 337.800 929.400 339.600 935.400 ;
        RECT 353.400 929.400 355.200 935.400 ;
        RECT 320.400 929.100 321.300 929.400 ;
        RECT 314.700 928.200 321.300 929.100 ;
        RECT 314.100 916.050 315.900 917.850 ;
        RECT 320.400 916.050 321.300 928.200 ;
        RECT 338.400 916.050 339.600 929.400 ;
        RECT 353.700 929.100 355.200 929.400 ;
        RECT 359.400 929.400 361.200 935.400 ;
        RECT 376.800 929.400 378.600 935.400 ;
        RECT 359.400 929.100 360.300 929.400 ;
        RECT 353.700 928.200 360.300 929.100 ;
        RECT 340.950 921.450 343.050 922.200 ;
        RECT 349.950 921.450 352.050 922.050 ;
        RECT 340.950 920.550 352.050 921.450 ;
        RECT 340.950 920.100 343.050 920.550 ;
        RECT 349.950 919.950 352.050 920.550 ;
        RECT 353.100 916.050 354.900 917.850 ;
        RECT 359.400 916.050 360.300 928.200 ;
        RECT 377.700 929.100 378.600 929.400 ;
        RECT 382.800 929.400 384.600 935.400 ;
        RECT 382.800 929.100 384.300 929.400 ;
        RECT 377.700 928.200 384.300 929.100 ;
        RECT 377.700 916.050 378.600 928.200 ;
        RECT 402.300 924.900 404.100 935.400 ;
        RECT 401.700 923.400 404.100 924.900 ;
        RECT 409.800 923.400 411.600 935.400 ;
        RECT 379.950 921.450 382.050 922.050 ;
        RECT 397.950 921.450 400.050 922.050 ;
        RECT 379.950 920.550 400.050 921.450 ;
        RECT 379.950 919.950 382.050 920.550 ;
        RECT 397.950 919.950 400.050 920.550 ;
        RECT 383.100 916.050 384.900 917.850 ;
        RECT 401.700 916.050 403.050 923.400 ;
        RECT 410.400 921.900 411.600 923.400 ;
        RECT 13.950 913.950 16.050 916.050 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 31.950 913.950 34.050 916.050 ;
        RECT 34.950 913.950 37.050 916.050 ;
        RECT 37.950 913.950 40.050 916.050 ;
        RECT 40.950 913.950 43.050 916.050 ;
        RECT 52.950 913.950 55.050 916.050 ;
        RECT 55.950 913.950 58.050 916.050 ;
        RECT 58.950 913.950 61.050 916.050 ;
        RECT 61.950 913.950 64.050 916.050 ;
        RECT 76.950 913.950 79.050 916.050 ;
        RECT 79.950 913.950 82.050 916.050 ;
        RECT 94.950 913.950 97.050 916.050 ;
        RECT 97.950 913.950 100.050 916.050 ;
        RECT 100.950 913.950 103.050 916.050 ;
        RECT 103.950 913.950 106.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 115.950 913.950 118.050 916.050 ;
        RECT 118.950 913.950 121.050 916.050 ;
        RECT 121.950 913.950 124.050 916.050 ;
        RECT 136.950 913.950 139.050 916.050 ;
        RECT 139.950 913.950 142.050 916.050 ;
        RECT 142.950 913.950 145.050 916.050 ;
        RECT 145.950 913.950 148.050 916.050 ;
        RECT 160.950 913.950 163.050 916.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 166.950 913.950 169.050 916.050 ;
        RECT 169.950 913.950 172.050 916.050 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 187.950 913.950 190.050 916.050 ;
        RECT 199.950 913.950 202.050 916.050 ;
        RECT 202.950 913.950 205.050 916.050 ;
        RECT 205.950 913.950 208.050 916.050 ;
        RECT 208.950 913.950 211.050 916.050 ;
        RECT 220.950 913.950 223.050 916.050 ;
        RECT 223.950 913.950 226.050 916.050 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 244.950 913.950 247.050 916.050 ;
        RECT 247.950 913.950 250.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 265.950 913.950 268.050 916.050 ;
        RECT 268.950 913.950 271.050 916.050 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 292.950 913.950 295.050 916.050 ;
        RECT 295.950 913.950 298.050 916.050 ;
        RECT 298.950 913.950 301.050 916.050 ;
        RECT 310.950 913.950 313.050 916.050 ;
        RECT 313.950 913.950 316.050 916.050 ;
        RECT 316.950 913.950 319.050 916.050 ;
        RECT 319.950 913.950 322.050 916.050 ;
        RECT 334.950 913.950 337.050 916.050 ;
        RECT 337.950 913.950 340.050 916.050 ;
        RECT 340.950 913.950 343.050 916.050 ;
        RECT 349.950 913.950 352.050 916.050 ;
        RECT 352.950 913.950 355.050 916.050 ;
        RECT 355.950 913.950 358.050 916.050 ;
        RECT 358.950 913.950 361.050 916.050 ;
        RECT 376.950 913.950 379.050 916.050 ;
        RECT 379.950 913.950 382.050 916.050 ;
        RECT 382.950 913.950 385.050 916.050 ;
        RECT 385.950 913.950 388.050 916.050 ;
        RECT 400.950 913.950 403.050 916.050 ;
        RECT 404.400 920.700 411.600 921.900 ;
        RECT 425.400 929.400 427.200 935.400 ;
        RECT 442.800 929.400 444.600 935.400 ;
        RECT 404.400 920.100 406.200 920.700 ;
        RECT 14.400 903.600 15.600 913.950 ;
        RECT 32.100 912.150 33.900 913.950 ;
        RECT 34.950 909.750 36.150 913.950 ;
        RECT 38.100 912.150 39.900 913.950 ;
        RECT 53.100 912.150 54.900 913.950 ;
        RECT 55.950 909.750 57.150 913.950 ;
        RECT 59.100 912.150 60.900 913.950 ;
        RECT 32.400 908.700 36.150 909.750 ;
        RECT 53.400 908.700 57.150 909.750 ;
        RECT 32.400 906.600 33.600 908.700 ;
        RECT 13.800 900.600 15.600 903.600 ;
        RECT 31.800 900.600 33.600 906.600 ;
        RECT 34.800 905.700 42.600 907.050 ;
        RECT 53.400 906.600 54.600 908.700 ;
        RECT 34.800 900.600 36.600 905.700 ;
        RECT 40.800 900.600 42.600 905.700 ;
        RECT 52.800 900.600 54.600 906.600 ;
        RECT 55.800 905.700 63.600 907.050 ;
        RECT 55.800 900.600 57.600 905.700 ;
        RECT 61.800 900.600 63.600 905.700 ;
        RECT 77.400 903.600 78.600 913.950 ;
        RECT 95.700 910.200 96.600 913.950 ;
        RECT 98.100 912.150 99.900 913.950 ;
        RECT 104.100 912.150 105.900 913.950 ;
        RECT 113.100 912.150 114.900 913.950 ;
        RECT 119.100 912.150 120.900 913.950 ;
        RECT 122.400 910.200 123.300 913.950 ;
        RECT 137.100 912.150 138.900 913.950 ;
        RECT 95.700 909.000 99.000 910.200 ;
        RECT 76.800 900.600 78.600 903.600 ;
        RECT 97.200 900.600 99.000 909.000 ;
        RECT 120.000 909.000 123.300 910.200 ;
        RECT 139.950 909.750 141.150 913.950 ;
        RECT 143.100 912.150 144.900 913.950 ;
        RECT 120.000 900.600 121.800 909.000 ;
        RECT 137.400 908.700 141.150 909.750 ;
        RECT 161.700 910.200 162.600 913.950 ;
        RECT 164.100 912.150 165.900 913.950 ;
        RECT 170.100 912.150 171.900 913.950 ;
        RECT 161.700 909.000 165.000 910.200 ;
        RECT 137.400 906.600 138.600 908.700 ;
        RECT 136.800 900.600 138.600 906.600 ;
        RECT 139.800 905.700 147.600 907.050 ;
        RECT 139.800 900.600 141.600 905.700 ;
        RECT 145.800 900.600 147.600 905.700 ;
        RECT 163.200 900.600 165.000 909.000 ;
        RECT 185.400 903.600 186.600 913.950 ;
        RECT 200.100 912.150 201.900 913.950 ;
        RECT 202.950 909.750 204.150 913.950 ;
        RECT 206.100 912.150 207.900 913.950 ;
        RECT 221.100 912.150 222.900 913.950 ;
        RECT 227.100 912.150 228.900 913.950 ;
        RECT 230.400 910.200 231.300 913.950 ;
        RECT 200.400 908.700 204.150 909.750 ;
        RECT 228.000 909.000 231.300 910.200 ;
        RECT 200.400 906.600 201.600 908.700 ;
        RECT 184.800 900.600 186.600 903.600 ;
        RECT 199.800 900.600 201.600 906.600 ;
        RECT 202.800 905.700 210.600 907.050 ;
        RECT 202.800 900.600 204.600 905.700 ;
        RECT 208.800 900.600 210.600 905.700 ;
        RECT 228.000 900.600 229.800 909.000 ;
        RECT 245.400 906.600 246.300 913.950 ;
        RECT 248.100 912.150 249.900 913.950 ;
        RECT 254.100 912.150 255.900 913.950 ;
        RECT 266.100 912.150 267.900 913.950 ;
        RECT 272.100 912.150 273.900 913.950 ;
        RECT 275.400 910.200 276.300 913.950 ;
        RECT 293.100 912.150 294.900 913.950 ;
        RECT 273.000 909.000 276.300 910.200 ;
        RECT 245.400 905.400 250.500 906.600 ;
        RECT 248.700 900.600 250.500 905.400 ;
        RECT 273.000 900.600 274.800 909.000 ;
        RECT 296.400 908.700 297.600 913.950 ;
        RECT 299.100 912.150 300.900 913.950 ;
        RECT 311.100 912.150 312.900 913.950 ;
        RECT 317.100 912.150 318.900 913.950 ;
        RECT 320.400 910.200 321.300 913.950 ;
        RECT 335.100 912.150 336.900 913.950 ;
        RECT 293.400 907.800 297.600 908.700 ;
        RECT 318.000 909.000 321.300 910.200 ;
        RECT 293.400 900.600 295.200 907.800 ;
        RECT 318.000 900.600 319.800 909.000 ;
        RECT 338.400 908.700 339.600 913.950 ;
        RECT 341.100 912.150 342.900 913.950 ;
        RECT 350.100 912.150 351.900 913.950 ;
        RECT 356.100 912.150 357.900 913.950 ;
        RECT 359.400 910.200 360.300 913.950 ;
        RECT 335.400 907.800 339.600 908.700 ;
        RECT 357.000 909.000 360.300 910.200 ;
        RECT 377.700 910.200 378.600 913.950 ;
        RECT 380.100 912.150 381.900 913.950 ;
        RECT 386.100 912.150 387.900 913.950 ;
        RECT 377.700 909.000 381.000 910.200 ;
        RECT 335.400 900.600 337.200 907.800 ;
        RECT 357.000 900.600 358.800 909.000 ;
        RECT 379.200 900.600 381.000 909.000 ;
        RECT 400.950 906.600 402.000 913.950 ;
        RECT 404.400 909.600 405.300 920.100 ;
        RECT 407.100 916.050 408.900 917.850 ;
        RECT 425.400 916.050 426.600 929.400 ;
        RECT 443.400 916.050 444.600 929.400 ;
        RECT 461.700 924.600 463.500 935.400 ;
        RECT 461.700 923.400 465.300 924.600 ;
        RECT 446.100 916.050 447.900 917.850 ;
        RECT 461.100 916.050 462.900 917.850 ;
        RECT 464.400 916.050 465.300 923.400 ;
        RECT 482.400 923.400 484.200 935.400 ;
        RECT 503.400 929.400 505.200 935.400 ;
        RECT 526.800 929.400 528.600 935.400 ;
        RECT 545.400 929.400 547.200 935.400 ;
        RECT 568.800 929.400 570.600 935.400 ;
        RECT 467.100 916.050 468.900 917.850 ;
        RECT 482.400 916.050 483.600 923.400 ;
        RECT 503.850 916.050 505.050 929.400 ;
        RECT 509.100 916.050 510.900 917.850 ;
        RECT 527.400 916.050 528.600 929.400 ;
        RECT 545.850 916.050 547.050 929.400 ;
        RECT 551.100 916.050 552.900 917.850 ;
        RECT 563.100 916.050 564.900 917.850 ;
        RECT 568.950 916.050 570.150 929.400 ;
        RECT 589.800 923.400 591.600 935.400 ;
        RECT 592.800 924.300 594.600 935.400 ;
        RECT 598.800 924.300 600.600 935.400 ;
        RECT 592.800 923.400 600.600 924.300 ;
        RECT 614.400 929.400 616.200 935.400 ;
        RECT 632.400 929.400 634.200 935.400 ;
        RECT 655.800 929.400 657.600 935.400 ;
        RECT 673.800 929.400 675.600 935.400 ;
        RECT 586.950 918.450 589.050 922.050 ;
        RECT 584.550 918.000 589.050 918.450 ;
        RECT 584.550 917.550 588.450 918.000 ;
        RECT 406.950 913.950 409.050 916.050 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 421.950 913.950 424.050 916.050 ;
        RECT 424.950 913.950 427.050 916.050 ;
        RECT 427.950 913.950 430.050 916.050 ;
        RECT 442.950 913.950 445.050 916.050 ;
        RECT 445.950 913.950 448.050 916.050 ;
        RECT 460.950 913.950 463.050 916.050 ;
        RECT 463.950 913.950 466.050 916.050 ;
        RECT 466.950 913.950 469.050 916.050 ;
        RECT 478.950 913.950 481.050 916.050 ;
        RECT 481.950 913.950 484.050 916.050 ;
        RECT 499.950 913.950 502.050 916.050 ;
        RECT 502.950 913.950 505.050 916.050 ;
        RECT 505.950 913.950 508.050 916.050 ;
        RECT 508.950 913.950 511.050 916.050 ;
        RECT 523.950 913.950 526.050 916.050 ;
        RECT 526.950 913.950 529.050 916.050 ;
        RECT 529.950 913.950 532.050 916.050 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 544.950 913.950 547.050 916.050 ;
        RECT 547.950 913.950 550.050 916.050 ;
        RECT 550.950 913.950 553.050 916.050 ;
        RECT 562.950 913.950 565.050 916.050 ;
        RECT 565.950 913.950 568.050 916.050 ;
        RECT 568.950 913.950 571.050 916.050 ;
        RECT 571.950 913.950 574.050 916.050 ;
        RECT 410.100 912.150 411.900 913.950 ;
        RECT 422.100 912.150 423.900 913.950 ;
        RECT 404.400 908.700 406.200 909.600 ;
        RECT 425.400 908.700 426.600 913.950 ;
        RECT 428.100 912.150 429.900 913.950 ;
        RECT 404.400 907.800 407.700 908.700 ;
        RECT 425.400 907.800 429.600 908.700 ;
        RECT 400.800 900.600 402.600 906.600 ;
        RECT 406.800 903.600 407.700 907.800 ;
        RECT 406.800 900.600 408.600 903.600 ;
        RECT 427.800 900.600 429.600 907.800 ;
        RECT 443.400 903.600 444.600 913.950 ;
        RECT 464.400 903.600 465.300 913.950 ;
        RECT 479.100 912.150 480.900 913.950 ;
        RECT 482.400 906.600 483.600 913.950 ;
        RECT 500.100 912.150 501.900 913.950 ;
        RECT 502.950 909.750 504.150 913.950 ;
        RECT 506.100 912.150 507.900 913.950 ;
        RECT 524.100 912.150 525.900 913.950 ;
        RECT 500.400 908.700 504.150 909.750 ;
        RECT 527.400 908.700 528.600 913.950 ;
        RECT 530.100 912.150 531.900 913.950 ;
        RECT 542.100 912.150 543.900 913.950 ;
        RECT 544.950 909.750 546.150 913.950 ;
        RECT 548.100 912.150 549.900 913.950 ;
        RECT 566.100 912.150 567.900 913.950 ;
        RECT 500.400 906.600 501.600 908.700 ;
        RECT 524.400 907.800 528.600 908.700 ;
        RECT 542.400 908.700 546.150 909.750 ;
        RECT 569.850 909.750 571.050 913.950 ;
        RECT 572.100 912.150 573.900 913.950 ;
        RECT 584.550 913.050 585.450 917.550 ;
        RECT 590.400 916.050 591.300 923.400 ;
        RECT 601.950 918.450 606.000 919.050 ;
        RECT 596.100 916.050 597.900 917.850 ;
        RECT 601.950 916.950 606.450 918.450 ;
        RECT 589.950 913.950 592.050 916.050 ;
        RECT 592.950 913.950 595.050 916.050 ;
        RECT 595.950 913.950 598.050 916.050 ;
        RECT 598.950 913.950 601.050 916.050 ;
        RECT 584.550 911.550 589.050 913.050 ;
        RECT 585.000 910.950 589.050 911.550 ;
        RECT 569.850 908.700 573.600 909.750 ;
        RECT 442.800 900.600 444.600 903.600 ;
        RECT 463.800 900.600 465.600 903.600 ;
        RECT 482.400 900.600 484.200 906.600 ;
        RECT 499.800 900.600 501.600 906.600 ;
        RECT 502.800 905.700 510.600 907.050 ;
        RECT 502.800 900.600 504.600 905.700 ;
        RECT 508.800 900.600 510.600 905.700 ;
        RECT 524.400 900.600 526.200 907.800 ;
        RECT 542.400 906.600 543.600 908.700 ;
        RECT 541.800 900.600 543.600 906.600 ;
        RECT 544.800 905.700 552.600 907.050 ;
        RECT 544.800 900.600 546.600 905.700 ;
        RECT 550.800 900.600 552.600 905.700 ;
        RECT 563.400 905.700 571.200 907.050 ;
        RECT 563.400 900.600 565.200 905.700 ;
        RECT 569.400 900.600 571.200 905.700 ;
        RECT 572.400 906.600 573.600 908.700 ;
        RECT 590.400 906.600 591.300 913.950 ;
        RECT 593.100 912.150 594.900 913.950 ;
        RECT 599.100 912.150 600.900 913.950 ;
        RECT 605.550 913.050 606.450 916.950 ;
        RECT 611.100 916.050 612.900 917.850 ;
        RECT 614.400 916.050 615.600 929.400 ;
        RECT 632.850 916.050 634.050 929.400 ;
        RECT 638.100 916.050 639.900 917.850 ;
        RECT 650.100 916.050 651.900 917.850 ;
        RECT 655.950 916.050 657.150 929.400 ;
        RECT 674.400 916.050 675.600 929.400 ;
        RECT 691.800 924.600 693.600 935.400 ;
        RECT 691.800 923.400 696.600 924.600 ;
        RECT 694.500 922.500 696.600 923.400 ;
        RECT 699.300 923.400 701.100 935.400 ;
        RECT 706.800 924.300 708.600 935.400 ;
        RECT 722.400 929.400 724.200 935.400 ;
        RECT 722.700 929.100 724.200 929.400 ;
        RECT 728.400 929.400 730.200 935.400 ;
        RECT 749.400 929.400 751.200 935.400 ;
        RECT 728.400 929.100 729.300 929.400 ;
        RECT 722.700 928.200 729.300 929.100 ;
        RECT 704.100 923.400 708.600 924.300 ;
        RECT 699.300 921.900 700.500 923.400 ;
        RECT 699.000 921.000 700.500 921.900 ;
        RECT 704.100 921.300 706.200 923.400 ;
        RECT 699.000 918.900 699.900 921.000 ;
        RECT 677.100 916.050 678.900 917.850 ;
        RECT 692.100 916.050 693.900 917.850 ;
        RECT 697.800 916.800 699.900 918.900 ;
        RECT 700.800 919.500 702.900 919.800 ;
        RECT 700.800 917.700 704.700 919.500 ;
        RECT 610.950 913.950 613.050 916.050 ;
        RECT 613.950 913.950 616.050 916.050 ;
        RECT 628.950 913.950 631.050 916.050 ;
        RECT 631.950 913.950 634.050 916.050 ;
        RECT 634.950 913.950 637.050 916.050 ;
        RECT 637.950 913.950 640.050 916.050 ;
        RECT 649.950 913.950 652.050 916.050 ;
        RECT 652.950 913.950 655.050 916.050 ;
        RECT 655.950 913.950 658.050 916.050 ;
        RECT 658.950 913.950 661.050 916.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 676.950 913.950 679.050 916.050 ;
        RECT 685.950 915.450 690.000 916.050 ;
        RECT 691.950 915.450 694.050 916.050 ;
        RECT 698.400 915.900 700.800 916.800 ;
        RECT 685.950 914.550 694.050 915.450 ;
        RECT 685.950 913.950 690.000 914.550 ;
        RECT 691.950 913.950 694.050 914.550 ;
        RECT 605.550 911.550 610.050 913.050 ;
        RECT 606.000 910.950 610.050 911.550 ;
        RECT 572.400 900.600 574.200 906.600 ;
        RECT 590.400 905.400 595.500 906.600 ;
        RECT 593.700 900.600 595.500 905.400 ;
        RECT 614.400 903.600 615.600 913.950 ;
        RECT 629.100 912.150 630.900 913.950 ;
        RECT 631.950 909.750 633.150 913.950 ;
        RECT 635.100 912.150 636.900 913.950 ;
        RECT 653.100 912.150 654.900 913.950 ;
        RECT 629.400 908.700 633.150 909.750 ;
        RECT 656.850 909.750 658.050 913.950 ;
        RECT 659.100 912.150 660.900 913.950 ;
        RECT 656.850 908.700 660.600 909.750 ;
        RECT 629.400 906.600 630.600 908.700 ;
        RECT 614.400 900.600 616.200 903.600 ;
        RECT 628.800 900.600 630.600 906.600 ;
        RECT 631.800 905.700 639.600 907.050 ;
        RECT 631.800 900.600 633.600 905.700 ;
        RECT 637.800 900.600 639.600 905.700 ;
        RECT 650.400 905.700 658.200 907.050 ;
        RECT 650.400 900.600 652.200 905.700 ;
        RECT 656.400 900.600 658.200 905.700 ;
        RECT 659.400 906.600 660.600 908.700 ;
        RECT 659.400 900.600 661.200 906.600 ;
        RECT 674.400 903.600 675.600 913.950 ;
        RECT 696.600 913.200 698.400 915.000 ;
        RECT 696.750 911.100 698.850 913.200 ;
        RECT 699.750 910.200 700.800 915.900 ;
        RECT 701.700 915.900 703.500 916.500 ;
        RECT 722.100 916.050 723.900 917.850 ;
        RECT 728.400 916.050 729.300 928.200 ;
        RECT 749.850 916.050 751.050 929.400 ;
        RECT 772.500 924.600 774.300 935.400 ;
        RECT 770.700 923.400 774.300 924.600 ;
        RECT 791.400 929.400 793.200 935.400 ;
        RECT 811.800 929.400 813.600 935.400 ;
        RECT 755.100 916.050 756.900 917.850 ;
        RECT 767.100 916.050 768.900 917.850 ;
        RECT 770.700 916.050 771.600 923.400 ;
        RECT 773.100 916.050 774.900 917.850 ;
        RECT 788.100 916.050 789.900 917.850 ;
        RECT 791.400 916.050 792.600 929.400 ;
        RECT 812.400 916.050 813.600 929.400 ;
        RECT 824.400 928.200 826.200 934.200 ;
        RECT 824.400 923.100 825.300 928.200 ;
        RECT 831.900 924.900 833.700 934.200 ;
        RECT 857.400 929.400 859.200 935.400 ;
        RECT 874.800 929.400 876.600 935.400 ;
        RECT 831.900 924.000 834.000 924.900 ;
        RECT 824.400 922.200 831.750 923.100 ;
        RECT 830.550 917.850 831.750 922.200 ;
        RECT 827.100 916.050 828.900 917.850 ;
        RECT 830.250 916.050 832.050 917.850 ;
        RECT 833.100 916.050 834.000 924.000 ;
        RECT 838.950 921.450 841.050 922.050 ;
        RECT 853.950 921.450 856.050 922.050 ;
        RECT 838.950 920.550 856.050 921.450 ;
        RECT 838.950 919.950 841.050 920.550 ;
        RECT 853.950 919.950 856.050 920.550 ;
        RECT 836.100 916.050 837.900 917.850 ;
        RECT 857.850 916.050 859.050 929.400 ;
        RECT 863.100 916.050 864.900 917.850 ;
        RECT 875.400 916.050 876.600 929.400 ;
        RECT 893.400 923.400 895.200 935.400 ;
        RECT 878.100 916.050 879.900 917.850 ;
        RECT 893.700 916.050 894.750 923.400 ;
        RECT 706.500 915.900 708.600 916.050 ;
        RECT 701.700 914.700 708.600 915.900 ;
        RECT 706.500 913.950 708.600 914.700 ;
        RECT 718.950 913.950 721.050 916.050 ;
        RECT 721.950 913.950 724.050 916.050 ;
        RECT 724.950 913.950 727.050 916.050 ;
        RECT 727.950 913.950 730.050 916.050 ;
        RECT 745.950 913.950 748.050 916.050 ;
        RECT 748.950 913.950 751.050 916.050 ;
        RECT 751.950 913.950 754.050 916.050 ;
        RECT 754.950 913.950 757.050 916.050 ;
        RECT 766.950 913.950 769.050 916.050 ;
        RECT 769.950 913.950 772.050 916.050 ;
        RECT 772.950 913.950 775.050 916.050 ;
        RECT 787.950 913.950 790.050 916.050 ;
        RECT 790.950 913.950 793.050 916.050 ;
        RECT 808.950 913.950 811.050 916.050 ;
        RECT 811.950 913.950 814.050 916.050 ;
        RECT 814.950 913.950 817.050 916.050 ;
        RECT 823.950 913.950 826.050 916.050 ;
        RECT 826.950 913.950 829.050 916.050 ;
        RECT 694.500 907.500 696.600 908.700 ;
        RECT 697.800 908.100 700.800 910.200 ;
        RECT 701.700 911.400 703.500 913.200 ;
        RECT 706.800 913.050 708.600 913.950 ;
        RECT 706.800 912.150 712.050 913.050 ;
        RECT 719.100 912.150 720.900 913.950 ;
        RECT 725.100 912.150 726.900 913.950 ;
        RECT 707.550 911.550 712.050 912.150 ;
        RECT 701.700 909.300 703.800 911.400 ;
        RECT 708.000 910.950 712.050 911.550 ;
        RECT 728.400 910.200 729.300 913.950 ;
        RECT 746.100 912.150 747.900 913.950 ;
        RECT 701.700 908.400 708.000 909.300 ;
        RECT 673.800 900.600 675.600 903.600 ;
        RECT 691.800 906.600 696.600 907.500 ;
        RECT 699.600 906.600 700.800 908.100 ;
        RECT 706.800 906.600 708.000 908.400 ;
        RECT 726.000 909.000 729.300 910.200 ;
        RECT 748.950 909.750 750.150 913.950 ;
        RECT 752.100 912.150 753.900 913.950 ;
        RECT 691.800 900.600 693.600 906.600 ;
        RECT 699.300 900.600 701.100 906.600 ;
        RECT 706.800 900.600 708.600 906.600 ;
        RECT 726.000 900.600 727.800 909.000 ;
        RECT 746.400 908.700 750.150 909.750 ;
        RECT 746.400 906.600 747.600 908.700 ;
        RECT 745.800 900.600 747.600 906.600 ;
        RECT 748.800 905.700 756.600 907.050 ;
        RECT 748.800 900.600 750.600 905.700 ;
        RECT 754.800 900.600 756.600 905.700 ;
        RECT 770.700 903.600 771.600 913.950 ;
        RECT 775.950 909.450 778.050 910.050 ;
        RECT 787.950 909.450 790.050 910.050 ;
        RECT 775.950 908.550 790.050 909.450 ;
        RECT 775.950 907.950 778.050 908.550 ;
        RECT 787.950 907.950 790.050 908.550 ;
        RECT 791.400 903.600 792.600 913.950 ;
        RECT 809.100 912.150 810.900 913.950 ;
        RECT 812.400 908.700 813.600 913.950 ;
        RECT 815.100 912.150 816.900 913.950 ;
        RECT 824.100 912.150 825.900 913.950 ;
        RECT 830.400 909.000 831.600 916.050 ;
        RECT 832.950 913.950 835.050 916.050 ;
        RECT 835.950 913.950 838.050 916.050 ;
        RECT 853.950 913.950 856.050 916.050 ;
        RECT 856.950 913.950 859.050 916.050 ;
        RECT 859.950 913.950 862.050 916.050 ;
        RECT 862.950 913.950 865.050 916.050 ;
        RECT 874.950 913.950 877.050 916.050 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 889.950 913.950 892.050 916.050 ;
        RECT 893.700 913.950 898.050 916.050 ;
        RECT 809.400 907.800 813.600 908.700 ;
        RECT 824.400 908.100 831.600 909.000 ;
        RECT 770.400 900.600 772.200 903.600 ;
        RECT 791.400 900.600 793.200 903.600 ;
        RECT 809.400 900.600 811.200 907.800 ;
        RECT 824.400 904.800 825.300 908.100 ;
        RECT 833.100 907.200 834.000 913.950 ;
        RECT 854.100 912.150 855.900 913.950 ;
        RECT 856.950 909.750 858.150 913.950 ;
        RECT 860.100 912.150 861.900 913.950 ;
        RECT 831.900 906.300 834.000 907.200 ;
        RECT 854.400 908.700 858.150 909.750 ;
        RECT 854.400 906.600 855.600 908.700 ;
        RECT 824.400 901.800 826.200 904.800 ;
        RECT 831.900 901.800 833.700 906.300 ;
        RECT 853.800 900.600 855.600 906.600 ;
        RECT 856.800 905.700 864.600 907.050 ;
        RECT 856.800 900.600 858.600 905.700 ;
        RECT 862.800 900.600 864.600 905.700 ;
        RECT 875.400 903.600 876.600 913.950 ;
        RECT 890.100 912.150 891.900 913.950 ;
        RECT 893.700 906.600 894.750 913.950 ;
        RECT 874.800 900.600 876.600 903.600 ;
        RECT 893.400 900.600 895.200 906.600 ;
        RECT 21.000 890.400 22.800 896.400 ;
        RECT 14.100 883.050 15.900 884.850 ;
        RECT 21.000 883.050 22.050 890.400 ;
        RECT 38.400 889.200 40.200 896.400 ;
        RECT 38.400 888.300 42.600 889.200 ;
        RECT 28.950 885.450 33.000 886.050 ;
        RECT 26.100 883.050 27.900 884.850 ;
        RECT 28.950 883.950 33.450 885.450 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 19.950 880.950 22.050 883.050 ;
        RECT 22.950 880.950 25.050 883.050 ;
        RECT 25.950 880.950 28.050 883.050 ;
        RECT 17.100 879.150 18.900 880.950 ;
        RECT 21.000 875.400 21.900 880.950 ;
        RECT 23.100 879.150 24.900 880.950 ;
        RECT 32.550 880.050 33.450 883.950 ;
        RECT 38.100 883.050 39.900 884.850 ;
        RECT 41.400 883.050 42.600 888.300 ;
        RECT 63.000 888.000 64.800 896.400 ;
        RECT 85.500 891.600 87.300 896.400 ;
        RECT 108.300 892.200 110.100 896.400 ;
        RECT 85.500 890.400 90.600 891.600 ;
        RECT 63.000 886.800 66.300 888.000 ;
        RECT 44.100 883.050 45.900 884.850 ;
        RECT 56.100 883.050 57.900 884.850 ;
        RECT 62.100 883.050 63.900 884.850 ;
        RECT 65.400 883.050 66.300 886.800 ;
        RECT 80.100 883.050 81.900 884.850 ;
        RECT 86.100 883.050 87.900 884.850 ;
        RECT 89.700 883.050 90.600 890.400 ;
        RECT 107.400 890.400 110.100 892.200 ;
        RECT 107.400 883.050 108.300 890.400 ;
        RECT 110.100 888.600 111.900 889.500 ;
        RECT 115.800 888.600 117.600 896.400 ;
        RECT 130.800 890.400 132.600 896.400 ;
        RECT 110.100 887.700 117.600 888.600 ;
        RECT 131.400 888.300 132.600 890.400 ;
        RECT 133.800 891.300 135.600 896.400 ;
        RECT 139.800 891.300 141.600 896.400 ;
        RECT 156.300 892.200 158.100 896.400 ;
        RECT 133.800 889.950 141.600 891.300 ;
        RECT 155.400 890.400 158.100 892.200 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 55.950 880.950 58.050 883.050 ;
        RECT 58.950 880.950 61.050 883.050 ;
        RECT 61.950 880.950 64.050 883.050 ;
        RECT 64.950 880.950 67.050 883.050 ;
        RECT 79.950 880.950 82.050 883.050 ;
        RECT 82.950 880.950 85.050 883.050 ;
        RECT 85.950 880.950 88.050 883.050 ;
        RECT 88.950 880.950 91.050 883.050 ;
        RECT 106.950 880.950 109.050 883.050 ;
        RECT 109.950 880.950 112.050 883.050 ;
        RECT 28.950 878.550 33.450 880.050 ;
        RECT 28.950 877.950 33.000 878.550 ;
        RECT 16.800 874.500 21.900 875.400 ;
        RECT 13.800 862.500 15.600 873.600 ;
        RECT 16.800 863.400 18.600 874.500 ;
        RECT 19.800 872.400 27.600 873.300 ;
        RECT 19.800 862.500 21.600 872.400 ;
        RECT 13.800 861.600 21.600 862.500 ;
        RECT 25.800 861.600 27.600 872.400 ;
        RECT 41.400 867.600 42.600 880.950 ;
        RECT 59.100 879.150 60.900 880.950 ;
        RECT 65.400 868.800 66.300 880.950 ;
        RECT 83.100 879.150 84.900 880.950 ;
        RECT 89.700 873.600 90.600 880.950 ;
        RECT 107.400 873.600 108.300 880.950 ;
        RECT 110.100 879.150 111.900 880.950 ;
        RECT 59.700 867.900 66.300 868.800 ;
        RECT 59.700 867.600 61.200 867.900 ;
        RECT 40.800 861.600 42.600 867.600 ;
        RECT 59.400 861.600 61.200 867.600 ;
        RECT 65.400 867.600 66.300 867.900 ;
        RECT 80.400 872.700 88.200 873.600 ;
        RECT 65.400 861.600 67.200 867.600 ;
        RECT 80.400 861.600 82.200 872.700 ;
        RECT 86.400 861.600 88.200 872.700 ;
        RECT 89.400 861.600 91.200 873.600 ;
        RECT 106.800 861.600 108.600 873.600 ;
        RECT 113.700 867.600 114.600 887.700 ;
        RECT 131.400 887.250 135.150 888.300 ;
        RECT 116.100 883.050 117.900 884.850 ;
        RECT 131.100 883.050 132.900 884.850 ;
        RECT 133.950 883.050 135.150 887.250 ;
        RECT 137.100 883.050 138.900 884.850 ;
        RECT 155.400 883.050 156.300 890.400 ;
        RECT 158.100 888.600 159.900 889.500 ;
        RECT 163.800 888.600 165.600 896.400 ;
        RECT 181.800 893.400 183.600 896.400 ;
        RECT 158.100 887.700 165.600 888.600 ;
        RECT 115.950 880.950 118.050 883.050 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 154.950 880.950 157.050 883.050 ;
        RECT 157.950 880.950 160.050 883.050 ;
        RECT 134.850 867.600 136.050 880.950 ;
        RECT 140.100 879.150 141.900 880.950 ;
        RECT 155.400 873.600 156.300 880.950 ;
        RECT 158.100 879.150 159.900 880.950 ;
        RECT 112.800 861.600 114.600 867.600 ;
        RECT 134.400 861.600 136.200 867.600 ;
        RECT 154.800 861.600 156.600 873.600 ;
        RECT 161.700 867.600 162.600 887.700 ;
        RECT 164.100 883.050 165.900 884.850 ;
        RECT 182.400 883.050 183.300 893.400 ;
        RECT 194.400 891.300 196.200 896.400 ;
        RECT 200.400 891.300 202.200 896.400 ;
        RECT 194.400 889.950 202.200 891.300 ;
        RECT 203.400 890.400 205.200 896.400 ;
        RECT 220.800 893.400 222.600 896.400 ;
        RECT 238.800 893.400 240.600 896.400 ;
        RECT 203.400 888.300 204.600 890.400 ;
        RECT 200.850 887.250 204.600 888.300 ;
        RECT 197.100 883.050 198.900 884.850 ;
        RECT 200.850 883.050 202.050 887.250 ;
        RECT 203.100 883.050 204.900 884.850 ;
        RECT 221.400 883.050 222.600 893.400 ;
        RECT 239.400 883.050 240.600 893.400 ;
        RECT 251.400 891.300 253.200 896.400 ;
        RECT 257.400 891.300 259.200 896.400 ;
        RECT 251.400 889.950 259.200 891.300 ;
        RECT 260.400 890.400 262.200 896.400 ;
        RECT 275.400 893.400 277.200 896.400 ;
        RECT 260.400 888.300 261.600 890.400 ;
        RECT 257.850 887.250 261.600 888.300 ;
        RECT 254.100 883.050 255.900 884.850 ;
        RECT 257.850 883.050 259.050 887.250 ;
        RECT 260.100 883.050 261.900 884.850 ;
        RECT 275.400 883.050 276.600 893.400 ;
        RECT 295.200 888.000 297.000 896.400 ;
        RECT 316.800 893.400 318.600 896.400 ;
        RECT 293.700 886.800 297.000 888.000 ;
        RECT 293.700 883.050 294.600 886.800 ;
        RECT 296.100 883.050 297.900 884.850 ;
        RECT 302.100 883.050 303.900 884.850 ;
        RECT 317.400 883.050 318.600 893.400 ;
        RECT 332.400 891.300 334.200 896.400 ;
        RECT 338.400 891.300 340.200 896.400 ;
        RECT 332.400 889.950 340.200 891.300 ;
        RECT 341.400 890.400 343.200 896.400 ;
        RECT 356.400 893.400 358.200 896.400 ;
        RECT 319.950 888.450 322.050 889.050 ;
        RECT 328.950 888.450 331.050 889.050 ;
        RECT 319.950 887.550 331.050 888.450 ;
        RECT 341.400 888.300 342.600 890.400 ;
        RECT 319.950 886.950 322.050 887.550 ;
        RECT 328.950 886.950 331.050 887.550 ;
        RECT 338.850 887.250 342.600 888.300 ;
        RECT 335.100 883.050 336.900 884.850 ;
        RECT 338.850 883.050 340.050 887.250 ;
        RECT 341.100 883.050 342.900 884.850 ;
        RECT 356.400 883.050 357.600 893.400 ;
        RECT 370.800 890.400 372.600 896.400 ;
        RECT 371.400 888.300 372.600 890.400 ;
        RECT 373.800 891.300 375.600 896.400 ;
        RECT 379.800 891.300 381.600 896.400 ;
        RECT 373.800 889.950 381.600 891.300 ;
        RECT 397.500 891.600 399.300 896.400 ;
        RECT 416.400 893.400 418.200 896.400 ;
        RECT 437.400 893.400 439.200 896.400 ;
        RECT 397.500 890.400 402.600 891.600 ;
        RECT 371.400 887.250 375.150 888.300 ;
        RECT 371.100 883.050 372.900 884.850 ;
        RECT 373.950 883.050 375.150 887.250 ;
        RECT 377.100 883.050 378.900 884.850 ;
        RECT 392.100 883.050 393.900 884.850 ;
        RECT 398.100 883.050 399.900 884.850 ;
        RECT 401.700 883.050 402.600 890.400 ;
        RECT 416.700 883.050 417.600 893.400 ;
        RECT 424.950 891.450 427.050 892.050 ;
        RECT 433.950 891.450 436.050 892.050 ;
        RECT 424.950 890.550 436.050 891.450 ;
        RECT 424.950 889.950 427.050 890.550 ;
        RECT 433.950 889.950 436.050 890.550 ;
        RECT 418.950 888.450 421.050 889.050 ;
        RECT 427.950 888.450 430.050 889.050 ;
        RECT 418.950 887.550 430.050 888.450 ;
        RECT 418.950 886.950 421.050 887.550 ;
        RECT 427.950 886.950 430.050 887.550 ;
        RECT 437.400 883.050 438.600 893.400 ;
        RECT 454.800 890.400 456.600 896.400 ;
        RECT 455.400 883.050 456.600 890.400 ;
        RECT 477.000 888.000 478.800 896.400 ;
        RECT 504.000 890.400 505.800 896.400 ;
        RECT 518.400 891.300 520.200 896.400 ;
        RECT 524.400 891.300 526.200 896.400 ;
        RECT 477.000 886.800 480.300 888.000 ;
        RECT 458.100 883.050 459.900 884.850 ;
        RECT 470.100 883.050 471.900 884.850 ;
        RECT 476.100 883.050 477.900 884.850 ;
        RECT 479.400 883.050 480.300 886.800 ;
        RECT 497.100 883.050 498.900 884.850 ;
        RECT 504.000 883.050 505.050 890.400 ;
        RECT 518.400 889.950 526.200 891.300 ;
        RECT 527.400 890.400 529.200 896.400 ;
        RECT 527.400 888.300 528.600 890.400 ;
        RECT 544.800 889.200 546.600 896.400 ;
        RECT 560.400 891.300 562.200 896.400 ;
        RECT 566.400 891.300 568.200 896.400 ;
        RECT 560.400 889.950 568.200 891.300 ;
        RECT 569.400 890.400 571.200 896.400 ;
        RECT 586.800 890.400 588.600 896.400 ;
        RECT 524.850 887.250 528.600 888.300 ;
        RECT 542.400 888.300 546.600 889.200 ;
        RECT 569.400 888.300 570.600 890.400 ;
        RECT 509.100 883.050 510.900 884.850 ;
        RECT 521.100 883.050 522.900 884.850 ;
        RECT 524.850 883.050 526.050 887.250 ;
        RECT 527.100 883.050 528.900 884.850 ;
        RECT 539.100 883.050 540.900 884.850 ;
        RECT 542.400 883.050 543.600 888.300 ;
        RECT 566.850 887.250 570.600 888.300 ;
        RECT 587.400 888.300 588.600 890.400 ;
        RECT 589.800 891.300 591.600 896.400 ;
        RECT 595.800 891.300 597.600 896.400 ;
        RECT 589.800 889.950 597.600 891.300 ;
        RECT 610.800 890.400 612.600 896.400 ;
        RECT 611.400 888.300 612.600 890.400 ;
        RECT 613.800 891.300 615.600 896.400 ;
        RECT 619.800 891.300 621.600 896.400 ;
        RECT 613.800 889.950 621.600 891.300 ;
        RECT 634.500 891.600 636.300 896.400 ;
        RECT 634.500 890.400 639.600 891.600 ;
        RECT 655.800 890.400 657.600 896.400 ;
        RECT 587.400 887.250 591.150 888.300 ;
        RECT 611.400 887.250 615.150 888.300 ;
        RECT 555.000 885.450 559.050 886.050 ;
        RECT 545.100 883.050 546.900 884.850 ;
        RECT 554.550 883.950 559.050 885.450 ;
        RECT 163.950 880.950 166.050 883.050 ;
        RECT 178.950 880.950 181.050 883.050 ;
        RECT 181.950 880.950 184.050 883.050 ;
        RECT 184.950 880.950 187.050 883.050 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 196.950 880.950 199.050 883.050 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 202.950 880.950 205.050 883.050 ;
        RECT 220.950 880.950 223.050 883.050 ;
        RECT 223.950 880.950 226.050 883.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 241.950 880.950 244.050 883.050 ;
        RECT 250.950 880.950 253.050 883.050 ;
        RECT 253.950 880.950 256.050 883.050 ;
        RECT 256.950 880.950 259.050 883.050 ;
        RECT 259.950 880.950 262.050 883.050 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 274.950 880.950 277.050 883.050 ;
        RECT 292.950 880.950 295.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 298.950 880.950 301.050 883.050 ;
        RECT 301.950 880.950 304.050 883.050 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 331.950 880.950 334.050 883.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 337.950 880.950 340.050 883.050 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 352.950 880.950 355.050 883.050 ;
        RECT 355.950 880.950 358.050 883.050 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 379.950 880.950 382.050 883.050 ;
        RECT 391.950 880.950 394.050 883.050 ;
        RECT 394.950 880.950 397.050 883.050 ;
        RECT 397.950 880.950 400.050 883.050 ;
        RECT 400.950 880.950 403.050 883.050 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 418.950 880.950 421.050 883.050 ;
        RECT 433.950 880.950 436.050 883.050 ;
        RECT 436.950 880.950 439.050 883.050 ;
        RECT 454.950 880.950 457.050 883.050 ;
        RECT 457.950 880.950 460.050 883.050 ;
        RECT 469.950 880.950 472.050 883.050 ;
        RECT 472.950 880.950 475.050 883.050 ;
        RECT 475.950 880.950 478.050 883.050 ;
        RECT 478.950 880.950 481.050 883.050 ;
        RECT 496.950 880.950 499.050 883.050 ;
        RECT 499.950 880.950 502.050 883.050 ;
        RECT 502.950 880.950 505.050 883.050 ;
        RECT 505.950 880.950 508.050 883.050 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 517.950 880.950 520.050 883.050 ;
        RECT 520.950 880.950 523.050 883.050 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 538.950 880.950 541.050 883.050 ;
        RECT 541.950 880.950 544.050 883.050 ;
        RECT 544.950 880.950 547.050 883.050 ;
        RECT 179.100 879.150 180.900 880.950 ;
        RECT 182.400 873.600 183.300 880.950 ;
        RECT 185.100 879.150 186.900 880.950 ;
        RECT 194.100 879.150 195.900 880.950 ;
        RECT 160.800 861.600 162.600 867.600 ;
        RECT 179.700 872.400 183.300 873.600 ;
        RECT 179.700 861.600 181.500 872.400 ;
        RECT 199.950 867.600 201.150 880.950 ;
        RECT 221.400 867.600 222.600 880.950 ;
        RECT 224.100 879.150 225.900 880.950 ;
        RECT 239.400 867.600 240.600 880.950 ;
        RECT 242.100 879.150 243.900 880.950 ;
        RECT 251.100 879.150 252.900 880.950 ;
        RECT 256.950 867.600 258.150 880.950 ;
        RECT 272.100 879.150 273.900 880.950 ;
        RECT 275.400 867.600 276.600 880.950 ;
        RECT 293.700 868.800 294.600 880.950 ;
        RECT 299.100 879.150 300.900 880.950 ;
        RECT 293.700 867.900 300.300 868.800 ;
        RECT 293.700 867.600 294.600 867.900 ;
        RECT 199.800 861.600 201.600 867.600 ;
        RECT 220.800 861.600 222.600 867.600 ;
        RECT 238.800 861.600 240.600 867.600 ;
        RECT 256.800 861.600 258.600 867.600 ;
        RECT 275.400 861.600 277.200 867.600 ;
        RECT 292.800 861.600 294.600 867.600 ;
        RECT 298.800 867.600 300.300 867.900 ;
        RECT 317.400 867.600 318.600 880.950 ;
        RECT 320.100 879.150 321.900 880.950 ;
        RECT 332.100 879.150 333.900 880.950 ;
        RECT 337.950 867.600 339.150 880.950 ;
        RECT 353.100 879.150 354.900 880.950 ;
        RECT 356.400 867.600 357.600 880.950 ;
        RECT 374.850 867.600 376.050 880.950 ;
        RECT 380.100 879.150 381.900 880.950 ;
        RECT 395.100 879.150 396.900 880.950 ;
        RECT 385.950 876.450 388.050 877.050 ;
        RECT 397.950 876.450 400.050 877.050 ;
        RECT 385.950 875.550 400.050 876.450 ;
        RECT 385.950 874.950 388.050 875.550 ;
        RECT 397.950 874.950 400.050 875.550 ;
        RECT 401.700 873.600 402.600 880.950 ;
        RECT 413.100 879.150 414.900 880.950 ;
        RECT 416.700 873.600 417.600 880.950 ;
        RECT 419.100 879.150 420.900 880.950 ;
        RECT 434.100 879.150 435.900 880.950 ;
        RECT 392.400 872.700 400.200 873.600 ;
        RECT 298.800 861.600 300.600 867.600 ;
        RECT 316.800 861.600 318.600 867.600 ;
        RECT 337.800 861.600 339.600 867.600 ;
        RECT 356.400 861.600 358.200 867.600 ;
        RECT 374.400 861.600 376.200 867.600 ;
        RECT 392.400 861.600 394.200 872.700 ;
        RECT 398.400 861.600 400.200 872.700 ;
        RECT 401.400 861.600 403.200 873.600 ;
        RECT 416.700 872.400 420.300 873.600 ;
        RECT 418.500 861.600 420.300 872.400 ;
        RECT 437.400 867.600 438.600 880.950 ;
        RECT 445.950 879.450 448.050 880.050 ;
        RECT 451.950 879.450 454.050 880.050 ;
        RECT 445.950 878.550 454.050 879.450 ;
        RECT 445.950 877.950 448.050 878.550 ;
        RECT 451.950 877.950 454.050 878.550 ;
        RECT 455.400 873.600 456.600 880.950 ;
        RECT 473.100 879.150 474.900 880.950 ;
        RECT 437.400 861.600 439.200 867.600 ;
        RECT 454.800 861.600 456.600 873.600 ;
        RECT 479.400 868.800 480.300 880.950 ;
        RECT 500.100 879.150 501.900 880.950 ;
        RECT 504.000 875.400 504.900 880.950 ;
        RECT 506.100 879.150 507.900 880.950 ;
        RECT 518.100 879.150 519.900 880.950 ;
        RECT 499.800 874.500 504.900 875.400 ;
        RECT 473.700 867.900 480.300 868.800 ;
        RECT 473.700 867.600 475.200 867.900 ;
        RECT 473.400 861.600 475.200 867.600 ;
        RECT 479.400 867.600 480.300 867.900 ;
        RECT 479.400 861.600 481.200 867.600 ;
        RECT 496.800 862.500 498.600 873.600 ;
        RECT 499.800 863.400 501.600 874.500 ;
        RECT 502.800 872.400 510.600 873.300 ;
        RECT 502.800 862.500 504.600 872.400 ;
        RECT 496.800 861.600 504.600 862.500 ;
        RECT 508.800 861.600 510.600 872.400 ;
        RECT 523.950 867.600 525.150 880.950 ;
        RECT 542.400 867.600 543.600 880.950 ;
        RECT 554.550 880.050 555.450 883.950 ;
        RECT 563.100 883.050 564.900 884.850 ;
        RECT 566.850 883.050 568.050 887.250 ;
        RECT 569.100 883.050 570.900 884.850 ;
        RECT 587.100 883.050 588.900 884.850 ;
        RECT 589.950 883.050 591.150 887.250 ;
        RECT 593.100 883.050 594.900 884.850 ;
        RECT 611.100 883.050 612.900 884.850 ;
        RECT 613.950 883.050 615.150 887.250 ;
        RECT 617.100 883.050 618.900 884.850 ;
        RECT 629.100 883.050 630.900 884.850 ;
        RECT 635.100 883.050 636.900 884.850 ;
        RECT 638.700 883.050 639.600 890.400 ;
        RECT 640.950 888.450 643.050 889.050 ;
        RECT 652.950 888.450 655.050 889.050 ;
        RECT 640.950 887.550 655.050 888.450 ;
        RECT 640.950 886.950 643.050 887.550 ;
        RECT 652.950 886.950 655.050 887.550 ;
        RECT 656.400 888.300 657.600 890.400 ;
        RECT 658.800 891.300 660.600 896.400 ;
        RECT 664.800 891.300 666.600 896.400 ;
        RECT 658.800 889.950 666.600 891.300 ;
        RECT 682.200 890.400 684.000 896.400 ;
        RECT 656.400 887.250 660.150 888.300 ;
        RECT 656.100 883.050 657.900 884.850 ;
        RECT 658.950 883.050 660.150 887.250 ;
        RECT 662.100 883.050 663.900 884.850 ;
        RECT 677.100 883.050 678.900 884.850 ;
        RECT 682.950 883.050 684.000 890.400 ;
        RECT 709.800 889.200 711.600 896.400 ;
        RECT 707.400 888.300 711.600 889.200 ;
        RECT 689.100 883.050 690.900 884.850 ;
        RECT 704.100 883.050 705.900 884.850 ;
        RECT 707.400 883.050 708.600 888.300 ;
        RECT 729.000 888.000 730.800 896.400 ;
        RECT 748.800 890.400 750.600 896.400 ;
        RECT 754.800 893.400 756.600 896.400 ;
        RECT 729.000 886.800 732.300 888.000 ;
        RECT 710.100 883.050 711.900 884.850 ;
        RECT 722.100 883.050 723.900 884.850 ;
        RECT 728.100 883.050 729.900 884.850 ;
        RECT 731.400 883.050 732.300 886.800 ;
        RECT 748.800 883.050 750.000 890.400 ;
        RECT 755.400 889.500 756.600 893.400 ;
        RECT 750.900 888.600 756.600 889.500 ;
        RECT 770.400 889.200 772.200 896.400 ;
        RECT 790.800 889.200 792.600 896.400 ;
        RECT 806.400 891.300 808.200 896.400 ;
        RECT 812.400 891.300 814.200 896.400 ;
        RECT 806.400 889.950 814.200 891.300 ;
        RECT 815.400 890.400 817.200 896.400 ;
        RECT 832.800 893.400 834.600 896.400 ;
        RECT 750.900 887.700 752.850 888.600 ;
        RECT 770.400 888.300 774.600 889.200 ;
        RECT 559.950 880.950 562.050 883.050 ;
        RECT 562.950 880.950 565.050 883.050 ;
        RECT 565.950 880.950 568.050 883.050 ;
        RECT 568.950 880.950 571.050 883.050 ;
        RECT 586.950 880.950 589.050 883.050 ;
        RECT 589.950 880.950 592.050 883.050 ;
        RECT 592.950 880.950 595.050 883.050 ;
        RECT 595.950 880.950 598.050 883.050 ;
        RECT 610.950 880.950 613.050 883.050 ;
        RECT 613.950 880.950 616.050 883.050 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 619.950 880.950 622.050 883.050 ;
        RECT 628.950 880.950 631.050 883.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 634.950 880.950 637.050 883.050 ;
        RECT 637.950 880.950 640.050 883.050 ;
        RECT 655.950 880.950 658.050 883.050 ;
        RECT 658.950 880.950 661.050 883.050 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 676.950 880.950 679.050 883.050 ;
        RECT 679.950 880.950 682.050 883.050 ;
        RECT 682.950 880.950 685.050 883.050 ;
        RECT 685.950 880.950 688.050 883.050 ;
        RECT 688.950 880.950 691.050 883.050 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 721.950 880.950 724.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 748.800 880.950 751.050 883.050 ;
        RECT 552.000 879.900 555.450 880.050 ;
        RECT 550.950 878.550 555.450 879.900 ;
        RECT 560.100 879.150 561.900 880.950 ;
        RECT 550.950 877.950 555.000 878.550 ;
        RECT 550.950 877.800 553.050 877.950 ;
        RECT 565.950 867.600 567.150 880.950 ;
        RECT 590.850 867.600 592.050 880.950 ;
        RECT 596.100 879.150 597.900 880.950 ;
        RECT 614.850 867.600 616.050 880.950 ;
        RECT 620.100 879.150 621.900 880.950 ;
        RECT 632.100 879.150 633.900 880.950 ;
        RECT 625.950 876.450 628.050 877.050 ;
        RECT 634.950 876.450 637.050 877.050 ;
        RECT 625.950 875.550 637.050 876.450 ;
        RECT 625.950 874.950 628.050 875.550 ;
        RECT 634.950 874.950 637.050 875.550 ;
        RECT 638.700 873.600 639.600 880.950 ;
        RECT 629.400 872.700 637.200 873.600 ;
        RECT 523.800 861.600 525.600 867.600 ;
        RECT 542.400 861.600 544.200 867.600 ;
        RECT 565.800 861.600 567.600 867.600 ;
        RECT 590.400 861.600 592.200 867.600 ;
        RECT 614.400 861.600 616.200 867.600 ;
        RECT 629.400 861.600 631.200 872.700 ;
        RECT 635.400 861.600 637.200 872.700 ;
        RECT 638.400 861.600 640.200 873.600 ;
        RECT 659.850 867.600 661.050 880.950 ;
        RECT 665.100 879.150 666.900 880.950 ;
        RECT 680.100 879.150 681.900 880.950 ;
        RECT 683.100 875.400 684.000 880.950 ;
        RECT 686.100 879.150 687.900 880.950 ;
        RECT 683.100 874.500 688.200 875.400 ;
        RECT 677.400 872.400 685.200 873.300 ;
        RECT 659.400 861.600 661.200 867.600 ;
        RECT 677.400 861.600 679.200 872.400 ;
        RECT 683.400 862.500 685.200 872.400 ;
        RECT 686.400 863.400 688.200 874.500 ;
        RECT 689.400 862.500 691.200 873.600 ;
        RECT 683.400 861.600 691.200 862.500 ;
        RECT 707.400 867.600 708.600 880.950 ;
        RECT 725.100 879.150 726.900 880.950 ;
        RECT 731.400 868.800 732.300 880.950 ;
        RECT 725.700 867.900 732.300 868.800 ;
        RECT 725.700 867.600 727.200 867.900 ;
        RECT 707.400 861.600 709.200 867.600 ;
        RECT 725.400 861.600 727.200 867.600 ;
        RECT 731.400 867.600 732.300 867.900 ;
        RECT 748.800 873.600 750.000 880.950 ;
        RECT 751.950 876.300 752.850 887.700 ;
        RECT 770.100 883.050 771.900 884.850 ;
        RECT 773.400 883.050 774.600 888.300 ;
        RECT 788.400 888.300 792.600 889.200 ;
        RECT 815.400 888.300 816.600 890.400 ;
        RECT 776.100 883.050 777.900 884.850 ;
        RECT 785.100 883.050 786.900 884.850 ;
        RECT 788.400 883.050 789.600 888.300 ;
        RECT 812.850 887.250 816.600 888.300 ;
        RECT 793.950 885.450 798.000 886.050 ;
        RECT 791.100 883.050 792.900 884.850 ;
        RECT 793.950 883.950 798.450 885.450 ;
        RECT 754.950 880.950 757.050 883.050 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 772.950 880.950 775.050 883.050 ;
        RECT 775.950 880.950 778.050 883.050 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 790.950 880.950 793.050 883.050 ;
        RECT 755.100 879.150 756.900 880.950 ;
        RECT 750.900 875.400 752.850 876.300 ;
        RECT 750.900 874.500 756.600 875.400 ;
        RECT 731.400 861.600 733.200 867.600 ;
        RECT 748.800 861.600 750.600 873.600 ;
        RECT 755.400 867.600 756.600 874.500 ;
        RECT 773.400 867.600 774.600 880.950 ;
        RECT 754.800 861.600 756.600 867.600 ;
        RECT 772.800 861.600 774.600 867.600 ;
        RECT 788.400 867.600 789.600 880.950 ;
        RECT 797.550 880.050 798.450 883.950 ;
        RECT 809.100 883.050 810.900 884.850 ;
        RECT 812.850 883.050 814.050 887.250 ;
        RECT 815.100 883.050 816.900 884.850 ;
        RECT 833.400 883.050 834.300 893.400 ;
        RECT 848.400 891.300 850.200 896.400 ;
        RECT 854.400 891.300 856.200 896.400 ;
        RECT 848.400 889.950 856.200 891.300 ;
        RECT 857.400 890.400 859.200 896.400 ;
        RECT 869.400 891.300 871.200 896.400 ;
        RECT 875.400 891.300 877.200 896.400 ;
        RECT 857.400 888.300 858.600 890.400 ;
        RECT 869.400 889.950 877.200 891.300 ;
        RECT 878.400 890.400 880.200 896.400 ;
        RECT 896.400 893.400 898.200 896.400 ;
        RECT 878.400 888.300 879.600 890.400 ;
        RECT 854.850 887.250 858.600 888.300 ;
        RECT 875.850 887.250 879.600 888.300 ;
        RECT 851.100 883.050 852.900 884.850 ;
        RECT 854.850 883.050 856.050 887.250 ;
        RECT 857.100 883.050 858.900 884.850 ;
        RECT 872.100 883.050 873.900 884.850 ;
        RECT 875.850 883.050 877.050 887.250 ;
        RECT 878.100 883.050 879.900 884.850 ;
        RECT 896.700 883.050 897.600 893.400 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 847.950 880.950 850.050 883.050 ;
        RECT 850.950 880.950 853.050 883.050 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 868.950 880.950 871.050 883.050 ;
        RECT 871.950 880.950 874.050 883.050 ;
        RECT 874.950 880.950 877.050 883.050 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 892.950 880.950 895.050 883.050 ;
        RECT 895.950 880.950 898.050 883.050 ;
        RECT 898.950 880.950 901.050 883.050 ;
        RECT 793.950 878.550 798.450 880.050 ;
        RECT 806.100 879.150 807.900 880.950 ;
        RECT 793.950 877.950 798.000 878.550 ;
        RECT 811.950 867.600 813.150 880.950 ;
        RECT 830.100 879.150 831.900 880.950 ;
        RECT 814.950 876.450 817.050 877.050 ;
        RECT 826.950 876.450 829.050 877.050 ;
        RECT 814.950 875.550 829.050 876.450 ;
        RECT 814.950 874.950 817.050 875.550 ;
        RECT 826.950 874.950 829.050 875.550 ;
        RECT 833.400 873.600 834.300 880.950 ;
        RECT 836.100 879.150 837.900 880.950 ;
        RECT 848.100 879.150 849.900 880.950 ;
        RECT 830.700 872.400 834.300 873.600 ;
        RECT 788.400 861.600 790.200 867.600 ;
        RECT 811.800 861.600 813.600 867.600 ;
        RECT 830.700 861.600 832.500 872.400 ;
        RECT 853.950 867.600 855.150 880.950 ;
        RECT 869.100 879.150 870.900 880.950 ;
        RECT 874.950 867.600 876.150 880.950 ;
        RECT 893.100 879.150 894.900 880.950 ;
        RECT 896.700 873.600 897.600 880.950 ;
        RECT 899.100 879.150 900.900 880.950 ;
        RECT 896.700 872.400 900.300 873.600 ;
        RECT 853.800 861.600 855.600 867.600 ;
        RECT 874.800 861.600 876.600 867.600 ;
        RECT 898.500 861.600 900.300 872.400 ;
        RECT 10.800 851.400 12.600 857.400 ;
        RECT 31.800 851.400 33.600 857.400 ;
        RECT 52.800 851.400 54.600 857.400 ;
        RECT 11.400 838.050 12.600 851.400 ;
        RECT 14.100 838.050 15.900 839.850 ;
        RECT 32.400 838.050 33.600 851.400 ;
        RECT 53.400 838.050 54.600 851.400 ;
        RECT 65.400 846.300 67.200 857.400 ;
        RECT 71.400 846.300 73.200 857.400 ;
        RECT 65.400 845.400 73.200 846.300 ;
        RECT 74.400 845.400 76.200 857.400 ;
        RECT 91.800 851.400 93.600 857.400 ;
        RECT 92.700 851.100 93.600 851.400 ;
        RECT 97.800 851.400 99.600 857.400 ;
        RECT 112.800 851.400 114.600 857.400 ;
        RECT 97.800 851.100 99.300 851.400 ;
        RECT 92.700 850.200 99.300 851.100 ;
        RECT 113.700 851.100 114.600 851.400 ;
        RECT 118.800 851.400 120.600 857.400 ;
        RECT 136.800 851.400 138.600 857.400 ;
        RECT 118.800 851.100 120.300 851.400 ;
        RECT 113.700 850.200 120.300 851.100 ;
        RECT 55.950 843.450 58.050 844.050 ;
        RECT 64.950 843.450 67.050 844.050 ;
        RECT 55.950 842.550 67.050 843.450 ;
        RECT 55.950 841.950 58.050 842.550 ;
        RECT 64.950 841.950 67.050 842.550 ;
        RECT 68.100 838.050 69.900 839.850 ;
        RECT 74.700 838.050 75.600 845.400 ;
        RECT 76.950 840.450 79.050 841.050 ;
        RECT 76.950 839.550 87.450 840.450 ;
        RECT 76.950 838.950 79.050 839.550 ;
        RECT 10.950 835.950 13.050 838.050 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 28.950 835.950 31.050 838.050 ;
        RECT 31.950 835.950 34.050 838.050 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 49.950 835.950 52.050 838.050 ;
        RECT 52.950 835.950 55.050 838.050 ;
        RECT 55.950 835.950 58.050 838.050 ;
        RECT 64.950 835.950 67.050 838.050 ;
        RECT 67.950 835.950 70.050 838.050 ;
        RECT 70.950 835.950 73.050 838.050 ;
        RECT 73.950 835.950 76.050 838.050 ;
        RECT 11.400 825.600 12.600 835.950 ;
        RECT 29.100 834.150 30.900 835.950 ;
        RECT 32.400 830.700 33.600 835.950 ;
        RECT 35.100 834.150 36.900 835.950 ;
        RECT 50.100 834.150 51.900 835.950 ;
        RECT 53.400 830.700 54.600 835.950 ;
        RECT 56.100 834.150 57.900 835.950 ;
        RECT 65.100 834.150 66.900 835.950 ;
        RECT 71.100 834.150 72.900 835.950 ;
        RECT 10.800 822.600 12.600 825.600 ;
        RECT 29.400 829.800 33.600 830.700 ;
        RECT 50.400 829.800 54.600 830.700 ;
        RECT 29.400 822.600 31.200 829.800 ;
        RECT 50.400 822.600 52.200 829.800 ;
        RECT 74.700 828.600 75.600 835.950 ;
        RECT 76.950 834.450 79.050 835.050 ;
        RECT 82.950 834.450 85.050 835.050 ;
        RECT 76.950 833.550 85.050 834.450 ;
        RECT 76.950 832.950 79.050 833.550 ;
        RECT 82.950 832.950 85.050 833.550 ;
        RECT 86.550 832.050 87.450 839.550 ;
        RECT 92.700 838.050 93.600 850.200 ;
        RECT 98.100 838.050 99.900 839.850 ;
        RECT 113.700 838.050 114.600 850.200 ;
        RECT 119.100 838.050 120.900 839.850 ;
        RECT 137.400 838.050 138.600 851.400 ;
        RECT 156.300 846.900 158.100 857.400 ;
        RECT 155.700 845.400 158.100 846.900 ;
        RECT 163.800 845.400 165.600 857.400 ;
        RECT 181.800 851.400 183.600 857.400 ;
        RECT 199.800 851.400 201.600 857.400 ;
        RECT 140.100 838.050 141.900 839.850 ;
        RECT 155.700 838.050 157.050 845.400 ;
        RECT 164.400 843.900 165.600 845.400 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 94.950 835.950 97.050 838.050 ;
        RECT 97.950 835.950 100.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 112.950 835.950 115.050 838.050 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 118.950 835.950 121.050 838.050 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 139.950 835.950 142.050 838.050 ;
        RECT 154.950 835.950 157.050 838.050 ;
        RECT 158.400 842.700 165.600 843.900 ;
        RECT 158.400 842.100 160.200 842.700 ;
        RECT 84.000 831.900 87.450 832.050 ;
        RECT 82.950 830.550 87.450 831.900 ;
        RECT 92.700 832.200 93.600 835.950 ;
        RECT 95.100 834.150 96.900 835.950 ;
        RECT 101.100 834.150 102.900 835.950 ;
        RECT 113.700 832.200 114.600 835.950 ;
        RECT 116.100 834.150 117.900 835.950 ;
        RECT 122.100 834.150 123.900 835.950 ;
        RECT 92.700 831.000 96.000 832.200 ;
        RECT 113.700 831.000 117.000 832.200 ;
        RECT 82.950 829.950 87.000 830.550 ;
        RECT 82.950 829.800 85.050 829.950 ;
        RECT 70.500 827.400 75.600 828.600 ;
        RECT 70.500 822.600 72.300 827.400 ;
        RECT 94.200 822.600 96.000 831.000 ;
        RECT 115.200 822.600 117.000 831.000 ;
        RECT 137.400 825.600 138.600 835.950 ;
        RECT 154.950 828.600 156.000 835.950 ;
        RECT 158.400 831.600 159.300 842.100 ;
        RECT 161.100 838.050 162.900 839.850 ;
        RECT 182.400 838.050 183.600 851.400 ;
        RECT 200.400 838.050 201.600 851.400 ;
        RECT 218.700 846.600 220.500 857.400 ;
        RECT 239.400 851.400 241.200 857.400 ;
        RECT 218.700 845.400 222.300 846.600 ;
        RECT 218.100 838.050 219.900 839.850 ;
        RECT 221.400 838.050 222.300 845.400 ;
        RECT 224.100 838.050 225.900 839.850 ;
        RECT 239.400 838.050 240.600 851.400 ;
        RECT 262.500 846.600 264.300 857.400 ;
        RECT 260.700 845.400 264.300 846.600 ;
        RECT 278.400 851.400 280.200 857.400 ;
        RECT 257.100 838.050 258.900 839.850 ;
        RECT 260.700 838.050 261.600 845.400 ;
        RECT 263.100 838.050 264.900 839.850 ;
        RECT 278.400 838.050 279.600 851.400 ;
        RECT 298.800 845.400 300.600 857.400 ;
        RECT 304.800 851.400 306.600 857.400 ;
        RECT 323.400 851.400 325.200 857.400 ;
        RECT 347.400 851.400 349.200 857.400 ;
        RECT 370.800 851.400 372.600 857.400 ;
        RECT 299.400 838.050 300.300 845.400 ;
        RECT 302.100 838.050 303.900 839.850 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 163.950 835.950 166.050 838.050 ;
        RECT 178.950 835.950 181.050 838.050 ;
        RECT 181.950 835.950 184.050 838.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 196.950 835.950 199.050 838.050 ;
        RECT 199.950 835.950 202.050 838.050 ;
        RECT 202.950 835.950 205.050 838.050 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 220.950 835.950 223.050 838.050 ;
        RECT 223.950 835.950 226.050 838.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 241.950 835.950 244.050 838.050 ;
        RECT 256.950 835.950 259.050 838.050 ;
        RECT 259.950 835.950 262.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 274.950 835.950 277.050 838.050 ;
        RECT 277.950 835.950 280.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 298.950 835.950 301.050 838.050 ;
        RECT 301.950 835.950 304.050 838.050 ;
        RECT 164.100 834.150 165.900 835.950 ;
        RECT 179.100 834.150 180.900 835.950 ;
        RECT 158.400 830.700 160.200 831.600 ;
        RECT 163.950 831.450 166.050 832.050 ;
        RECT 172.950 831.450 175.050 832.050 ;
        RECT 158.400 829.800 161.700 830.700 ;
        RECT 163.950 830.550 175.050 831.450 ;
        RECT 182.400 830.700 183.600 835.950 ;
        RECT 185.100 834.150 186.900 835.950 ;
        RECT 197.100 834.150 198.900 835.950 ;
        RECT 200.400 830.700 201.600 835.950 ;
        RECT 203.100 834.150 204.900 835.950 ;
        RECT 163.950 829.950 166.050 830.550 ;
        RECT 172.950 829.950 175.050 830.550 ;
        RECT 136.800 822.600 138.600 825.600 ;
        RECT 154.800 822.600 156.600 828.600 ;
        RECT 160.800 825.600 161.700 829.800 ;
        RECT 179.400 829.800 183.600 830.700 ;
        RECT 197.400 829.800 201.600 830.700 ;
        RECT 160.800 822.600 162.600 825.600 ;
        RECT 179.400 822.600 181.200 829.800 ;
        RECT 197.400 822.600 199.200 829.800 ;
        RECT 221.400 825.600 222.300 835.950 ;
        RECT 236.100 834.150 237.900 835.950 ;
        RECT 239.400 830.700 240.600 835.950 ;
        RECT 242.100 834.150 243.900 835.950 ;
        RECT 239.400 829.800 243.600 830.700 ;
        RECT 220.800 822.600 222.600 825.600 ;
        RECT 241.800 822.600 243.600 829.800 ;
        RECT 244.950 828.450 247.050 829.050 ;
        RECT 256.950 828.450 259.050 829.050 ;
        RECT 244.950 827.550 259.050 828.450 ;
        RECT 244.950 826.950 247.050 827.550 ;
        RECT 256.950 826.950 259.050 827.550 ;
        RECT 260.700 825.600 261.600 835.950 ;
        RECT 275.100 834.150 276.900 835.950 ;
        RECT 278.400 830.700 279.600 835.950 ;
        RECT 281.100 834.150 282.900 835.950 ;
        RECT 278.400 829.800 282.600 830.700 ;
        RECT 260.400 822.600 262.200 825.600 ;
        RECT 280.800 822.600 282.600 829.800 ;
        RECT 299.400 828.600 300.300 835.950 ;
        RECT 305.700 831.300 306.600 851.400 ;
        RECT 323.850 838.050 325.050 851.400 ;
        RECT 331.950 840.450 334.050 844.050 ;
        RECT 337.950 843.450 340.050 844.050 ;
        RECT 343.950 843.450 346.050 844.050 ;
        RECT 337.950 842.550 346.050 843.450 ;
        RECT 337.950 841.950 340.050 842.550 ;
        RECT 343.950 841.950 346.050 842.550 ;
        RECT 331.950 840.000 336.450 840.450 ;
        RECT 329.100 838.050 330.900 839.850 ;
        RECT 332.550 839.550 336.450 840.000 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 319.950 835.950 322.050 838.050 ;
        RECT 322.950 835.950 325.050 838.050 ;
        RECT 325.950 835.950 328.050 838.050 ;
        RECT 328.950 835.950 331.050 838.050 ;
        RECT 308.100 834.150 309.900 835.950 ;
        RECT 320.100 834.150 321.900 835.950 ;
        RECT 322.950 831.750 324.150 835.950 ;
        RECT 326.100 834.150 327.900 835.950 ;
        RECT 335.550 834.450 336.450 839.550 ;
        RECT 347.850 838.050 349.050 851.400 ;
        RECT 353.100 838.050 354.900 839.850 ;
        RECT 365.100 838.050 366.900 839.850 ;
        RECT 370.950 838.050 372.150 851.400 ;
        RECT 389.400 845.400 391.200 857.400 ;
        RECT 396.900 846.900 398.700 857.400 ;
        RECT 416.400 851.400 418.200 857.400 ;
        RECT 439.800 851.400 441.600 857.400 ;
        RECT 460.800 851.400 462.600 857.400 ;
        RECT 481.800 851.400 483.600 857.400 ;
        RECT 496.800 851.400 498.600 857.400 ;
        RECT 396.900 845.400 399.300 846.900 ;
        RECT 389.400 843.900 390.600 845.400 ;
        RECT 389.400 842.700 396.600 843.900 ;
        RECT 394.800 842.100 396.600 842.700 ;
        RECT 392.100 838.050 393.900 839.850 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 349.950 835.950 352.050 838.050 ;
        RECT 352.950 835.950 355.050 838.050 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 373.950 835.950 376.050 838.050 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 391.950 835.950 394.050 838.050 ;
        RECT 340.950 834.450 343.050 835.050 ;
        RECT 335.550 833.550 343.050 834.450 ;
        RECT 344.100 834.150 345.900 835.950 ;
        RECT 340.950 832.950 343.050 833.550 ;
        RECT 346.950 831.750 348.150 835.950 ;
        RECT 350.100 834.150 351.900 835.950 ;
        RECT 368.100 834.150 369.900 835.950 ;
        RECT 302.100 830.400 309.600 831.300 ;
        RECT 302.100 829.500 303.900 830.400 ;
        RECT 299.400 826.800 302.100 828.600 ;
        RECT 286.950 825.450 289.050 826.050 ;
        RECT 295.950 825.450 298.050 826.050 ;
        RECT 286.950 824.550 298.050 825.450 ;
        RECT 286.950 823.950 289.050 824.550 ;
        RECT 295.950 823.950 298.050 824.550 ;
        RECT 300.300 822.600 302.100 826.800 ;
        RECT 307.800 822.600 309.600 830.400 ;
        RECT 320.400 830.700 324.150 831.750 ;
        RECT 344.400 830.700 348.150 831.750 ;
        RECT 371.850 831.750 373.050 835.950 ;
        RECT 374.100 834.150 375.900 835.950 ;
        RECT 389.100 834.150 390.900 835.950 ;
        RECT 371.850 830.700 375.600 831.750 ;
        RECT 395.700 831.600 396.600 842.100 ;
        RECT 397.950 838.050 399.300 845.400 ;
        RECT 416.400 838.050 417.600 851.400 ;
        RECT 440.400 838.050 441.600 851.400 ;
        RECT 448.950 843.450 451.050 844.050 ;
        RECT 457.950 843.450 460.050 844.050 ;
        RECT 448.950 842.550 460.050 843.450 ;
        RECT 448.950 841.950 451.050 842.550 ;
        RECT 457.950 841.950 460.050 842.550 ;
        RECT 461.400 838.050 462.600 851.400 ;
        RECT 482.400 838.050 483.600 851.400 ;
        RECT 497.700 851.100 498.600 851.400 ;
        RECT 502.800 851.400 504.600 857.400 ;
        RECT 520.800 856.500 528.600 857.400 ;
        RECT 502.800 851.100 504.300 851.400 ;
        RECT 497.700 850.200 504.300 851.100 ;
        RECT 497.700 838.050 498.600 850.200 ;
        RECT 520.800 845.400 522.600 856.500 ;
        RECT 523.800 844.500 525.600 855.600 ;
        RECT 526.800 846.600 528.600 856.500 ;
        RECT 532.800 846.600 534.600 857.400 ;
        RECT 550.800 851.400 552.600 857.400 ;
        RECT 526.800 845.700 534.600 846.600 ;
        RECT 523.800 843.600 528.900 844.500 ;
        RECT 503.100 838.050 504.900 839.850 ;
        RECT 524.100 838.050 525.900 839.850 ;
        RECT 528.000 838.050 528.900 843.600 ;
        RECT 530.100 838.050 531.900 839.850 ;
        RECT 551.400 838.050 552.600 851.400 ;
        RECT 565.800 845.400 567.600 857.400 ;
        RECT 586.800 851.400 588.600 857.400 ;
        RECT 566.400 838.050 567.600 845.400 ;
        RECT 587.400 838.050 588.600 851.400 ;
        RECT 604.800 845.400 606.600 857.400 ;
        RECT 607.800 846.300 609.600 857.400 ;
        RECT 613.800 846.300 615.600 857.400 ;
        RECT 631.800 851.400 633.600 857.400 ;
        RECT 650.400 851.400 652.200 857.400 ;
        RECT 674.400 851.400 676.200 857.400 ;
        RECT 692.400 851.400 694.200 857.400 ;
        RECT 713.400 851.400 715.200 857.400 ;
        RECT 607.800 845.400 615.600 846.300 ;
        RECT 605.400 838.050 606.300 845.400 ;
        RECT 611.100 838.050 612.900 839.850 ;
        RECT 626.100 838.050 627.900 839.850 ;
        RECT 631.950 838.050 633.150 851.400 ;
        RECT 650.400 838.050 651.600 851.400 ;
        RECT 674.850 838.050 676.050 851.400 ;
        RECT 680.100 838.050 681.900 839.850 ;
        RECT 692.400 838.050 693.600 851.400 ;
        RECT 713.700 851.100 715.200 851.400 ;
        RECT 719.400 851.400 721.200 857.400 ;
        RECT 740.400 851.400 742.200 857.400 ;
        RECT 719.400 851.100 720.300 851.400 ;
        RECT 713.700 850.200 720.300 851.100 ;
        RECT 713.100 838.050 714.900 839.850 ;
        RECT 719.400 838.050 720.300 850.200 ;
        RECT 730.950 843.450 733.050 844.050 ;
        RECT 736.950 843.450 739.050 844.200 ;
        RECT 730.950 842.550 739.050 843.450 ;
        RECT 730.950 841.950 733.050 842.550 ;
        RECT 736.950 842.100 739.050 842.550 ;
        RECT 721.950 840.450 724.050 841.050 ;
        RECT 721.950 839.550 732.450 840.450 ;
        RECT 721.950 838.950 724.050 839.550 ;
        RECT 397.950 835.950 400.050 838.050 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 415.950 835.950 418.050 838.050 ;
        RECT 418.950 835.950 421.050 838.050 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 442.950 835.950 445.050 838.050 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 463.950 835.950 466.050 838.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 484.950 835.950 487.050 838.050 ;
        RECT 496.950 835.950 499.050 838.050 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 502.950 835.950 505.050 838.050 ;
        RECT 505.950 835.950 508.050 838.050 ;
        RECT 520.950 835.950 523.050 838.050 ;
        RECT 523.950 835.950 526.050 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 532.950 835.950 535.050 838.050 ;
        RECT 547.950 835.950 550.050 838.050 ;
        RECT 550.950 835.950 553.050 838.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 568.950 835.950 571.050 838.050 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 589.950 835.950 592.050 838.050 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 607.950 835.950 610.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 625.950 835.950 628.050 838.050 ;
        RECT 628.950 835.950 631.050 838.050 ;
        RECT 631.950 835.950 634.050 838.050 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 646.950 835.950 649.050 838.050 ;
        RECT 649.950 835.950 652.050 838.050 ;
        RECT 652.950 835.950 655.050 838.050 ;
        RECT 670.950 835.950 673.050 838.050 ;
        RECT 673.950 835.950 676.050 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 679.950 835.950 682.050 838.050 ;
        RECT 688.950 835.950 691.050 838.050 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 694.950 835.950 697.050 838.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 718.950 835.950 721.050 838.050 ;
        RECT 394.800 830.700 396.600 831.600 ;
        RECT 320.400 828.600 321.600 830.700 ;
        RECT 319.800 822.600 321.600 828.600 ;
        RECT 322.800 827.700 330.600 829.050 ;
        RECT 344.400 828.600 345.600 830.700 ;
        RECT 322.800 822.600 324.600 827.700 ;
        RECT 328.800 822.600 330.600 827.700 ;
        RECT 343.800 822.600 345.600 828.600 ;
        RECT 346.800 827.700 354.600 829.050 ;
        RECT 346.800 822.600 348.600 827.700 ;
        RECT 352.800 822.600 354.600 827.700 ;
        RECT 365.400 827.700 373.200 829.050 ;
        RECT 365.400 822.600 367.200 827.700 ;
        RECT 371.400 822.600 373.200 827.700 ;
        RECT 374.400 828.600 375.600 830.700 ;
        RECT 393.300 829.800 396.600 830.700 ;
        RECT 374.400 822.600 376.200 828.600 ;
        RECT 393.300 825.600 394.200 829.800 ;
        RECT 399.000 828.600 400.050 835.950 ;
        RECT 413.100 834.150 414.900 835.950 ;
        RECT 416.400 830.700 417.600 835.950 ;
        RECT 419.100 834.150 420.900 835.950 ;
        RECT 437.100 834.150 438.900 835.950 ;
        RECT 440.400 830.700 441.600 835.950 ;
        RECT 443.100 834.150 444.900 835.950 ;
        RECT 458.100 834.150 459.900 835.950 ;
        RECT 461.400 830.700 462.600 835.950 ;
        RECT 464.100 834.150 465.900 835.950 ;
        RECT 479.100 834.150 480.900 835.950 ;
        RECT 482.400 830.700 483.600 835.950 ;
        RECT 485.100 834.150 486.900 835.950 ;
        RECT 497.700 832.200 498.600 835.950 ;
        RECT 500.100 834.150 501.900 835.950 ;
        RECT 506.100 834.150 507.900 835.950 ;
        RECT 521.100 834.150 522.900 835.950 ;
        RECT 497.700 831.000 501.000 832.200 ;
        RECT 416.400 829.800 420.600 830.700 ;
        RECT 392.400 822.600 394.200 825.600 ;
        RECT 398.400 822.600 400.200 828.600 ;
        RECT 418.800 822.600 420.600 829.800 ;
        RECT 437.400 829.800 441.600 830.700 ;
        RECT 458.400 829.800 462.600 830.700 ;
        RECT 479.400 829.800 483.600 830.700 ;
        RECT 437.400 822.600 439.200 829.800 ;
        RECT 458.400 822.600 460.200 829.800 ;
        RECT 479.400 822.600 481.200 829.800 ;
        RECT 499.200 822.600 501.000 831.000 ;
        RECT 514.950 831.450 517.050 832.050 ;
        RECT 523.950 831.450 526.050 832.050 ;
        RECT 514.950 830.550 526.050 831.450 ;
        RECT 514.950 829.950 517.050 830.550 ;
        RECT 523.950 829.950 526.050 830.550 ;
        RECT 528.000 828.600 529.050 835.950 ;
        RECT 533.100 834.150 534.900 835.950 ;
        RECT 548.100 834.150 549.900 835.950 ;
        RECT 551.400 830.700 552.600 835.950 ;
        RECT 554.100 834.150 555.900 835.950 ;
        RECT 548.400 829.800 552.600 830.700 ;
        RECT 528.000 822.600 529.800 828.600 ;
        RECT 548.400 822.600 550.200 829.800 ;
        RECT 566.400 828.600 567.600 835.950 ;
        RECT 569.100 834.150 570.900 835.950 ;
        RECT 584.100 834.150 585.900 835.950 ;
        RECT 587.400 830.700 588.600 835.950 ;
        RECT 590.100 834.150 591.900 835.950 ;
        RECT 565.800 822.600 567.600 828.600 ;
        RECT 584.400 829.800 588.600 830.700 ;
        RECT 584.400 822.600 586.200 829.800 ;
        RECT 605.400 828.600 606.300 835.950 ;
        RECT 608.100 834.150 609.900 835.950 ;
        RECT 614.100 834.150 615.900 835.950 ;
        RECT 629.100 834.150 630.900 835.950 ;
        RECT 632.850 831.750 634.050 835.950 ;
        RECT 635.100 834.150 636.900 835.950 ;
        RECT 647.100 834.150 648.900 835.950 ;
        RECT 632.850 830.700 636.600 831.750 ;
        RECT 605.400 827.400 610.500 828.600 ;
        RECT 608.700 822.600 610.500 827.400 ;
        RECT 626.400 827.700 634.200 829.050 ;
        RECT 626.400 822.600 628.200 827.700 ;
        RECT 632.400 822.600 634.200 827.700 ;
        RECT 635.400 828.600 636.600 830.700 ;
        RECT 650.400 830.700 651.600 835.950 ;
        RECT 653.100 834.150 654.900 835.950 ;
        RECT 671.100 834.150 672.900 835.950 ;
        RECT 673.950 831.750 675.150 835.950 ;
        RECT 677.100 834.150 678.900 835.950 ;
        RECT 689.100 834.150 690.900 835.950 ;
        RECT 671.400 830.700 675.150 831.750 ;
        RECT 692.400 830.700 693.600 835.950 ;
        RECT 695.100 834.150 696.900 835.950 ;
        RECT 710.100 834.150 711.900 835.950 ;
        RECT 716.100 834.150 717.900 835.950 ;
        RECT 719.400 832.200 720.300 835.950 ;
        RECT 731.550 835.050 732.450 839.550 ;
        RECT 740.850 838.050 742.050 851.400 ;
        RECT 758.400 846.600 760.200 857.400 ;
        RECT 764.400 856.500 772.200 857.400 ;
        RECT 764.400 846.600 766.200 856.500 ;
        RECT 758.400 845.700 766.200 846.600 ;
        RECT 767.400 844.500 769.200 855.600 ;
        RECT 770.400 845.400 772.200 856.500 ;
        RECT 788.400 851.400 790.200 857.400 ;
        RECT 764.100 843.600 769.200 844.500 ;
        RECT 746.100 838.050 747.900 839.850 ;
        RECT 761.100 838.050 762.900 839.850 ;
        RECT 764.100 838.050 765.000 843.600 ;
        RECT 767.100 838.050 768.900 839.850 ;
        RECT 785.100 838.050 786.900 839.850 ;
        RECT 788.400 838.050 789.600 851.400 ;
        RECT 805.800 846.600 807.600 857.400 ;
        RECT 805.800 845.400 810.600 846.600 ;
        RECT 808.500 844.500 810.600 845.400 ;
        RECT 813.300 845.400 815.100 857.400 ;
        RECT 820.800 846.300 822.600 857.400 ;
        RECT 835.800 851.400 837.600 857.400 ;
        RECT 818.100 845.400 822.600 846.300 ;
        RECT 813.300 843.900 814.500 845.400 ;
        RECT 813.000 843.000 814.500 843.900 ;
        RECT 818.100 843.300 820.200 845.400 ;
        RECT 813.000 840.900 813.900 843.000 ;
        RECT 806.100 838.050 807.900 839.850 ;
        RECT 811.800 838.800 813.900 840.900 ;
        RECT 814.800 841.500 816.900 841.800 ;
        RECT 814.800 839.700 818.700 841.500 ;
        RECT 736.950 835.950 739.050 838.050 ;
        RECT 739.950 835.950 742.050 838.050 ;
        RECT 742.950 835.950 745.050 838.050 ;
        RECT 745.950 835.950 748.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 763.950 835.950 766.050 838.050 ;
        RECT 766.950 835.950 769.050 838.050 ;
        RECT 769.950 835.950 772.050 838.050 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 787.950 835.950 790.050 838.050 ;
        RECT 796.950 837.450 799.050 838.050 ;
        RECT 805.950 837.450 808.050 838.050 ;
        RECT 812.400 837.900 814.800 838.800 ;
        RECT 796.950 836.550 808.050 837.450 ;
        RECT 796.950 835.950 799.050 836.550 ;
        RECT 805.950 835.950 808.050 836.550 ;
        RECT 731.550 833.550 736.050 835.050 ;
        RECT 737.100 834.150 738.900 835.950 ;
        RECT 732.000 832.950 736.050 833.550 ;
        RECT 717.000 831.000 720.300 832.200 ;
        RECT 739.950 831.750 741.150 835.950 ;
        RECT 743.100 834.150 744.900 835.950 ;
        RECT 758.100 834.150 759.900 835.950 ;
        RECT 650.400 829.800 654.600 830.700 ;
        RECT 635.400 822.600 637.200 828.600 ;
        RECT 652.800 822.600 654.600 829.800 ;
        RECT 671.400 828.600 672.600 830.700 ;
        RECT 692.400 829.800 696.600 830.700 ;
        RECT 670.800 822.600 672.600 828.600 ;
        RECT 673.800 827.700 681.600 829.050 ;
        RECT 673.800 822.600 675.600 827.700 ;
        RECT 679.800 822.600 681.600 827.700 ;
        RECT 694.800 822.600 696.600 829.800 ;
        RECT 717.000 822.600 718.800 831.000 ;
        RECT 737.400 830.700 741.150 831.750 ;
        RECT 737.400 828.600 738.600 830.700 ;
        RECT 736.800 822.600 738.600 828.600 ;
        RECT 739.800 827.700 747.600 829.050 ;
        RECT 763.950 828.600 765.000 835.950 ;
        RECT 770.100 834.150 771.900 835.950 ;
        RECT 739.800 822.600 741.600 827.700 ;
        RECT 745.800 822.600 747.600 827.700 ;
        RECT 763.200 822.600 765.000 828.600 ;
        RECT 788.400 825.600 789.600 835.950 ;
        RECT 810.600 835.200 812.400 837.000 ;
        RECT 810.750 833.100 812.850 835.200 ;
        RECT 813.750 832.200 814.800 837.900 ;
        RECT 815.700 837.900 817.500 838.500 ;
        RECT 836.400 838.050 837.600 851.400 ;
        RECT 853.800 845.400 855.600 857.400 ;
        RECT 856.800 846.300 858.600 857.400 ;
        RECT 862.800 846.300 864.600 857.400 ;
        RECT 877.800 851.400 879.600 857.400 ;
        RECT 856.800 845.400 864.600 846.300 ;
        RECT 839.100 838.050 840.900 839.850 ;
        RECT 854.400 838.050 855.300 845.400 ;
        RECT 860.100 838.050 861.900 839.850 ;
        RECT 872.100 838.050 873.900 839.850 ;
        RECT 877.950 838.050 879.150 851.400 ;
        RECT 898.800 845.400 900.600 857.400 ;
        RECT 904.800 851.400 906.600 857.400 ;
        RECT 898.800 838.050 900.000 845.400 ;
        RECT 905.400 844.500 906.600 851.400 ;
        RECT 900.900 843.600 906.600 844.500 ;
        RECT 900.900 842.700 902.850 843.600 ;
        RECT 820.500 837.900 826.050 838.050 ;
        RECT 815.700 836.700 826.050 837.900 ;
        RECT 820.500 835.950 826.050 836.700 ;
        RECT 835.950 835.950 838.050 838.050 ;
        RECT 838.950 835.950 841.050 838.050 ;
        RECT 853.950 835.950 856.050 838.050 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 859.950 835.950 862.050 838.050 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 874.950 835.950 877.050 838.050 ;
        RECT 877.950 835.950 880.050 838.050 ;
        RECT 880.950 835.950 883.050 838.050 ;
        RECT 898.800 835.950 901.050 838.050 ;
        RECT 808.500 829.500 810.600 830.700 ;
        RECT 811.800 830.100 814.800 832.200 ;
        RECT 815.700 833.400 817.500 835.200 ;
        RECT 820.800 834.150 822.600 835.950 ;
        RECT 815.700 831.300 817.800 833.400 ;
        RECT 815.700 830.400 822.000 831.300 ;
        RECT 805.800 828.600 810.600 829.500 ;
        RECT 813.600 828.600 814.800 830.100 ;
        RECT 820.800 828.600 822.000 830.400 ;
        RECT 788.400 822.600 790.200 825.600 ;
        RECT 805.800 822.600 807.600 828.600 ;
        RECT 813.300 822.600 815.100 828.600 ;
        RECT 820.800 822.600 822.600 828.600 ;
        RECT 836.400 825.600 837.600 835.950 ;
        RECT 854.400 828.600 855.300 835.950 ;
        RECT 857.100 834.150 858.900 835.950 ;
        RECT 863.100 834.150 864.900 835.950 ;
        RECT 875.100 834.150 876.900 835.950 ;
        RECT 878.850 831.750 880.050 835.950 ;
        RECT 881.100 834.150 882.900 835.950 ;
        RECT 878.850 830.700 882.600 831.750 ;
        RECT 854.400 827.400 859.500 828.600 ;
        RECT 835.800 822.600 837.600 825.600 ;
        RECT 857.700 822.600 859.500 827.400 ;
        RECT 872.400 827.700 880.200 829.050 ;
        RECT 872.400 822.600 874.200 827.700 ;
        RECT 878.400 822.600 880.200 827.700 ;
        RECT 881.400 828.600 882.600 830.700 ;
        RECT 898.800 828.600 900.000 835.950 ;
        RECT 901.950 831.300 902.850 842.700 ;
        RECT 905.100 838.050 906.900 839.850 ;
        RECT 904.950 835.950 907.050 838.050 ;
        RECT 900.900 830.400 902.850 831.300 ;
        RECT 900.900 829.500 906.600 830.400 ;
        RECT 881.400 822.600 883.200 828.600 ;
        RECT 898.800 822.600 900.600 828.600 ;
        RECT 905.400 825.600 906.600 829.500 ;
        RECT 904.800 822.600 906.600 825.600 ;
        RECT 13.800 812.400 15.600 818.400 ;
        RECT 19.800 815.400 21.600 818.400 ;
        RECT 13.950 805.050 15.000 812.400 ;
        RECT 19.800 811.200 20.700 815.400 ;
        RECT 41.700 813.600 43.500 818.400 ;
        RECT 17.400 810.300 20.700 811.200 ;
        RECT 38.400 812.400 43.500 813.600 ;
        RECT 17.400 809.400 19.200 810.300 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 14.700 795.600 16.050 802.950 ;
        RECT 17.400 798.900 18.300 809.400 ;
        RECT 23.100 805.050 24.900 806.850 ;
        RECT 38.400 805.050 39.300 812.400 ;
        RECT 59.400 811.200 61.200 818.400 ;
        RECT 59.400 810.300 63.600 811.200 ;
        RECT 41.100 805.050 42.900 806.850 ;
        RECT 47.100 805.050 48.900 806.850 ;
        RECT 59.100 805.050 60.900 806.850 ;
        RECT 62.400 805.050 63.600 810.300 ;
        RECT 79.200 810.000 81.000 818.400 ;
        RECT 77.700 808.800 81.000 810.000 ;
        RECT 105.000 810.000 106.800 818.400 ;
        RECT 127.500 813.600 129.300 818.400 ;
        RECT 127.500 812.400 132.600 813.600 ;
        RECT 105.000 808.800 108.300 810.000 ;
        RECT 65.100 805.050 66.900 806.850 ;
        RECT 77.700 805.050 78.600 808.800 ;
        RECT 80.100 805.050 81.900 806.850 ;
        RECT 86.100 805.050 87.900 806.850 ;
        RECT 98.100 805.050 99.900 806.850 ;
        RECT 104.100 805.050 105.900 806.850 ;
        RECT 107.400 805.050 108.300 808.800 ;
        RECT 122.100 805.050 123.900 806.850 ;
        RECT 128.100 805.050 129.900 806.850 ;
        RECT 131.700 805.050 132.600 812.400 ;
        RECT 146.400 813.300 148.200 818.400 ;
        RECT 152.400 813.300 154.200 818.400 ;
        RECT 146.400 811.950 154.200 813.300 ;
        RECT 155.400 812.400 157.200 818.400 ;
        RECT 155.400 810.300 156.600 812.400 ;
        RECT 173.400 811.200 175.200 818.400 ;
        RECT 152.850 809.250 156.600 810.300 ;
        RECT 149.100 805.050 150.900 806.850 ;
        RECT 152.850 805.050 154.050 809.250 ;
        RECT 160.950 808.950 163.050 811.050 ;
        RECT 173.400 810.300 177.600 811.200 ;
        RECT 155.100 805.050 156.900 806.850 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 58.950 802.950 61.050 805.050 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 64.950 802.950 67.050 805.050 ;
        RECT 76.950 802.950 79.050 805.050 ;
        RECT 79.950 802.950 82.050 805.050 ;
        RECT 82.950 802.950 85.050 805.050 ;
        RECT 85.950 802.950 88.050 805.050 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 100.950 802.950 103.050 805.050 ;
        RECT 103.950 802.950 106.050 805.050 ;
        RECT 106.950 802.950 109.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 127.950 802.950 130.050 805.050 ;
        RECT 130.950 802.950 133.050 805.050 ;
        RECT 145.950 802.950 148.050 805.050 ;
        RECT 148.950 802.950 151.050 805.050 ;
        RECT 151.950 802.950 154.050 805.050 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 20.100 801.150 21.900 802.950 ;
        RECT 17.400 798.300 19.200 798.900 ;
        RECT 17.400 797.100 24.600 798.300 ;
        RECT 23.400 795.600 24.600 797.100 ;
        RECT 38.400 795.600 39.300 802.950 ;
        RECT 44.100 801.150 45.900 802.950 ;
        RECT 14.700 794.100 17.100 795.600 ;
        RECT 15.300 783.600 17.100 794.100 ;
        RECT 22.800 783.600 24.600 795.600 ;
        RECT 37.800 783.600 39.600 795.600 ;
        RECT 40.800 794.700 48.600 795.600 ;
        RECT 40.800 783.600 42.600 794.700 ;
        RECT 46.800 783.600 48.600 794.700 ;
        RECT 62.400 789.600 63.600 802.950 ;
        RECT 77.700 790.800 78.600 802.950 ;
        RECT 83.100 801.150 84.900 802.950 ;
        RECT 101.100 801.150 102.900 802.950 ;
        RECT 107.400 790.800 108.300 802.950 ;
        RECT 125.100 801.150 126.900 802.950 ;
        RECT 131.700 795.600 132.600 802.950 ;
        RECT 146.100 801.150 147.900 802.950 ;
        RECT 77.700 789.900 84.300 790.800 ;
        RECT 77.700 789.600 78.600 789.900 ;
        RECT 61.800 783.600 63.600 789.600 ;
        RECT 76.800 783.600 78.600 789.600 ;
        RECT 82.800 789.600 84.300 789.900 ;
        RECT 101.700 789.900 108.300 790.800 ;
        RECT 101.700 789.600 103.200 789.900 ;
        RECT 82.800 783.600 84.600 789.600 ;
        RECT 101.400 783.600 103.200 789.600 ;
        RECT 107.400 789.600 108.300 789.900 ;
        RECT 122.400 794.700 130.200 795.600 ;
        RECT 107.400 783.600 109.200 789.600 ;
        RECT 122.400 783.600 124.200 794.700 ;
        RECT 128.400 783.600 130.200 794.700 ;
        RECT 131.400 783.600 133.200 795.600 ;
        RECT 151.950 789.600 153.150 802.950 ;
        RECT 161.550 801.450 162.450 808.950 ;
        RECT 173.100 805.050 174.900 806.850 ;
        RECT 176.400 805.050 177.600 810.300 ;
        RECT 195.000 810.000 196.800 818.400 ;
        RECT 212.400 812.400 214.200 818.400 ;
        RECT 219.600 813.000 221.400 818.400 ;
        RECT 212.400 811.500 213.900 812.400 ;
        RECT 212.400 810.000 216.750 811.500 ;
        RECT 195.000 808.800 198.300 810.000 ;
        RECT 214.650 809.400 216.750 810.000 ;
        RECT 220.350 810.900 221.400 813.000 ;
        RECT 227.400 812.400 229.200 818.400 ;
        RECT 224.700 811.200 229.200 812.400 ;
        RECT 247.800 811.200 249.600 818.400 ;
        RECT 262.800 817.500 270.600 818.400 ;
        RECT 262.800 812.400 264.600 817.500 ;
        RECT 265.800 812.400 267.600 816.600 ;
        RECT 268.800 813.000 270.600 817.500 ;
        RECT 274.800 813.000 276.600 818.400 ;
        RECT 179.100 805.050 180.900 806.850 ;
        RECT 188.100 805.050 189.900 806.850 ;
        RECT 194.100 805.050 195.900 806.850 ;
        RECT 197.400 805.050 198.300 808.800 ;
        RECT 217.650 807.900 219.450 809.700 ;
        RECT 220.350 808.800 223.500 810.900 ;
        RECT 224.700 809.100 226.800 811.200 ;
        RECT 245.400 810.300 249.600 811.200 ;
        RECT 266.400 810.900 267.300 812.400 ;
        RECT 268.800 812.100 276.600 813.000 ;
        RECT 287.400 813.300 289.200 818.400 ;
        RECT 293.400 813.300 295.200 818.400 ;
        RECT 287.400 811.950 295.200 813.300 ;
        RECT 296.400 812.400 298.200 818.400 ;
        RECT 311.400 815.400 313.200 818.400 ;
        RECT 217.200 807.000 219.300 807.900 ;
        RECT 212.700 805.800 219.300 807.000 ;
        RECT 212.700 805.200 214.500 805.800 ;
        RECT 172.950 802.950 175.050 805.050 ;
        RECT 175.950 802.950 178.050 805.050 ;
        RECT 178.950 802.950 181.050 805.050 ;
        RECT 187.950 802.950 190.050 805.050 ;
        RECT 190.950 802.950 193.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 212.400 803.100 214.500 805.200 ;
        RECT 169.950 801.450 172.050 802.050 ;
        RECT 161.550 800.550 172.050 801.450 ;
        RECT 169.950 799.950 172.050 800.550 ;
        RECT 166.950 798.450 169.050 799.050 ;
        RECT 172.950 798.450 175.050 799.050 ;
        RECT 166.950 797.550 175.050 798.450 ;
        RECT 166.950 796.950 169.050 797.550 ;
        RECT 172.950 796.950 175.050 797.550 ;
        RECT 176.400 789.600 177.600 802.950 ;
        RECT 191.100 801.150 192.900 802.950 ;
        RECT 197.400 790.800 198.300 802.950 ;
        RECT 217.200 802.800 219.300 804.900 ;
        RECT 217.200 801.000 219.000 802.800 ;
        RECT 220.350 802.200 221.250 808.800 ;
        RECT 222.150 804.900 224.250 807.000 ;
        RECT 222.300 803.100 224.100 804.900 ;
        RECT 226.950 803.100 229.050 805.200 ;
        RECT 242.100 805.050 243.900 806.850 ;
        RECT 245.400 805.050 246.600 810.300 ;
        RECT 266.400 809.700 271.050 810.900 ;
        RECT 296.400 810.300 297.600 812.400 ;
        RECT 248.100 805.050 249.900 806.850 ;
        RECT 266.100 805.050 267.900 806.850 ;
        RECT 269.700 805.050 271.050 809.700 ;
        RECT 293.850 809.250 297.600 810.300 ;
        RECT 272.100 805.050 273.900 806.850 ;
        RECT 290.100 805.050 291.900 806.850 ;
        RECT 293.850 805.050 295.050 809.250 ;
        RECT 296.100 805.050 297.900 806.850 ;
        RECT 311.400 805.050 312.600 815.400 ;
        RECT 328.800 812.400 330.600 818.400 ;
        RECT 329.400 810.300 330.600 812.400 ;
        RECT 331.800 813.300 333.600 818.400 ;
        RECT 337.800 813.300 339.600 818.400 ;
        RECT 331.800 811.950 339.600 813.300 ;
        RECT 347.400 813.300 349.200 818.400 ;
        RECT 353.400 813.300 355.200 818.400 ;
        RECT 347.400 811.950 355.200 813.300 ;
        RECT 356.400 812.400 358.200 818.400 ;
        RECT 356.400 810.300 357.600 812.400 ;
        RECT 329.400 809.250 333.150 810.300 ;
        RECT 329.100 805.050 330.900 806.850 ;
        RECT 331.950 805.050 333.150 809.250 ;
        RECT 353.850 809.250 357.600 810.300 ;
        RECT 378.000 810.000 379.800 818.400 ;
        RECT 400.800 811.200 402.600 818.400 ;
        RECT 413.400 813.300 415.200 818.400 ;
        RECT 419.400 813.300 421.200 818.400 ;
        RECT 413.400 811.950 421.200 813.300 ;
        RECT 422.400 812.400 424.200 818.400 ;
        RECT 437.400 815.400 439.200 818.400 ;
        RECT 452.400 815.400 454.200 818.400 ;
        RECT 398.400 810.300 402.600 811.200 ;
        RECT 422.400 810.300 423.600 812.400 ;
        RECT 335.100 805.050 336.900 806.850 ;
        RECT 350.100 805.050 351.900 806.850 ;
        RECT 353.850 805.050 355.050 809.250 ;
        RECT 378.000 808.800 381.300 810.000 ;
        RECT 356.100 805.050 357.900 806.850 ;
        RECT 371.100 805.050 372.900 806.850 ;
        RECT 377.100 805.050 378.900 806.850 ;
        RECT 380.400 805.050 381.300 808.800 ;
        RECT 390.000 807.450 394.050 808.050 ;
        RECT 389.550 805.950 394.050 807.450 ;
        RECT 220.350 800.700 223.500 802.200 ;
        RECT 227.100 801.450 228.900 803.100 ;
        RECT 241.950 802.950 244.050 805.050 ;
        RECT 244.950 802.950 247.050 805.050 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 262.950 802.950 265.050 805.050 ;
        RECT 265.950 802.950 268.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 274.950 802.950 277.050 805.050 ;
        RECT 286.950 802.950 289.050 805.050 ;
        RECT 289.950 802.950 292.050 805.050 ;
        RECT 292.950 802.950 295.050 805.050 ;
        RECT 295.950 802.950 298.050 805.050 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 337.950 802.950 340.050 805.050 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 349.950 802.950 352.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 232.950 801.450 235.050 802.050 ;
        RECT 227.100 801.300 235.050 801.450 ;
        RECT 221.400 800.100 223.500 800.700 ;
        RECT 227.550 800.550 235.050 801.300 ;
        RECT 218.700 797.700 220.500 799.800 ;
        RECT 215.100 796.800 220.500 797.700 ;
        RECT 215.100 795.900 217.200 796.800 ;
        RECT 191.700 789.900 198.300 790.800 ;
        RECT 191.700 789.600 193.200 789.900 ;
        RECT 151.800 783.600 153.600 789.600 ;
        RECT 175.800 783.600 177.600 789.600 ;
        RECT 191.400 783.600 193.200 789.600 ;
        RECT 197.400 789.600 198.300 789.900 ;
        RECT 212.400 794.700 217.200 795.900 ;
        RECT 222.000 795.600 223.200 800.100 ;
        RECT 232.950 799.950 235.050 800.550 ;
        RECT 219.900 794.700 223.200 795.600 ;
        RECT 224.100 795.600 226.200 796.500 ;
        RECT 197.400 783.600 199.200 789.600 ;
        RECT 212.400 783.600 214.200 794.700 ;
        RECT 219.900 783.600 221.700 794.700 ;
        RECT 224.100 794.400 229.200 795.600 ;
        RECT 227.400 783.600 229.200 794.400 ;
        RECT 245.400 789.600 246.600 802.950 ;
        RECT 263.100 801.150 264.900 802.950 ;
        RECT 269.700 795.600 270.900 802.950 ;
        RECT 275.100 801.150 276.900 802.950 ;
        RECT 287.100 801.150 288.900 802.950 ;
        RECT 245.400 783.600 247.200 789.600 ;
        RECT 268.800 783.600 272.100 795.600 ;
        RECT 292.950 789.600 294.150 802.950 ;
        RECT 308.100 801.150 309.900 802.950 ;
        RECT 295.950 798.450 298.050 799.050 ;
        RECT 307.950 798.450 310.050 799.050 ;
        RECT 295.950 797.550 310.050 798.450 ;
        RECT 295.950 796.950 298.050 797.550 ;
        RECT 307.950 796.950 310.050 797.550 ;
        RECT 311.400 789.600 312.600 802.950 ;
        RECT 332.850 789.600 334.050 802.950 ;
        RECT 338.100 801.150 339.900 802.950 ;
        RECT 347.100 801.150 348.900 802.950 ;
        RECT 352.950 789.600 354.150 802.950 ;
        RECT 374.100 801.150 375.900 802.950 ;
        RECT 355.950 798.450 358.050 799.050 ;
        RECT 376.950 798.450 379.050 799.050 ;
        RECT 355.950 797.550 379.050 798.450 ;
        RECT 355.950 796.950 358.050 797.550 ;
        RECT 376.950 796.950 379.050 797.550 ;
        RECT 380.400 790.800 381.300 802.950 ;
        RECT 389.550 802.050 390.450 805.950 ;
        RECT 395.100 805.050 396.900 806.850 ;
        RECT 398.400 805.050 399.600 810.300 ;
        RECT 419.850 809.250 423.600 810.300 ;
        RECT 403.950 807.450 408.000 808.050 ;
        RECT 401.100 805.050 402.900 806.850 ;
        RECT 403.950 805.950 408.450 807.450 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 389.550 800.550 394.050 802.050 ;
        RECT 390.000 799.950 394.050 800.550 ;
        RECT 382.950 795.450 385.050 796.050 ;
        RECT 394.950 795.450 397.050 796.050 ;
        RECT 382.950 794.550 397.050 795.450 ;
        RECT 382.950 793.950 385.050 794.550 ;
        RECT 394.950 793.950 397.050 794.550 ;
        RECT 374.700 789.900 381.300 790.800 ;
        RECT 374.700 789.600 376.200 789.900 ;
        RECT 292.800 783.600 294.600 789.600 ;
        RECT 311.400 783.600 313.200 789.600 ;
        RECT 332.400 783.600 334.200 789.600 ;
        RECT 352.800 783.600 354.600 789.600 ;
        RECT 374.400 783.600 376.200 789.600 ;
        RECT 380.400 789.600 381.300 789.900 ;
        RECT 398.400 789.600 399.600 802.950 ;
        RECT 407.550 802.050 408.450 805.950 ;
        RECT 416.100 805.050 417.900 806.850 ;
        RECT 419.850 805.050 421.050 809.250 ;
        RECT 424.950 807.450 429.000 808.050 ;
        RECT 422.100 805.050 423.900 806.850 ;
        RECT 424.950 805.950 429.450 807.450 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 421.950 802.950 424.050 805.050 ;
        RECT 403.950 800.550 408.450 802.050 ;
        RECT 413.100 801.150 414.900 802.950 ;
        RECT 403.950 799.950 408.000 800.550 ;
        RECT 418.950 789.600 420.150 802.950 ;
        RECT 428.550 802.050 429.450 805.950 ;
        RECT 437.400 805.050 438.600 815.400 ;
        RECT 444.000 807.450 448.050 808.050 ;
        RECT 443.550 805.950 448.050 807.450 ;
        RECT 433.950 802.950 436.050 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 424.950 800.550 429.450 802.050 ;
        RECT 434.100 801.150 435.900 802.950 ;
        RECT 424.950 799.950 429.000 800.550 ;
        RECT 437.400 789.600 438.600 802.950 ;
        RECT 443.550 802.050 444.450 805.950 ;
        RECT 452.400 805.050 453.600 815.400 ;
        RECT 464.400 810.600 466.200 818.400 ;
        RECT 471.900 814.200 473.700 818.400 ;
        RECT 471.900 812.400 474.600 814.200 ;
        RECT 470.100 810.600 471.900 811.500 ;
        RECT 464.400 809.700 471.900 810.600 ;
        RECT 464.100 805.050 465.900 806.850 ;
        RECT 448.950 802.950 451.050 805.050 ;
        RECT 451.950 802.950 454.050 805.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 443.550 800.550 448.050 802.050 ;
        RECT 449.100 801.150 450.900 802.950 ;
        RECT 444.000 799.950 448.050 800.550 ;
        RECT 452.400 789.600 453.600 802.950 ;
        RECT 467.400 789.600 468.300 809.700 ;
        RECT 473.700 805.050 474.600 812.400 ;
        RECT 491.400 811.200 493.200 818.400 ;
        RECT 519.000 812.400 520.800 818.400 ;
        RECT 533.400 813.300 535.200 818.400 ;
        RECT 539.400 813.300 541.200 818.400 ;
        RECT 491.400 810.300 495.600 811.200 ;
        RECT 475.950 807.450 480.000 808.050 ;
        RECT 475.950 805.950 480.450 807.450 ;
        RECT 469.950 802.950 472.050 805.050 ;
        RECT 472.950 802.950 475.050 805.050 ;
        RECT 470.100 801.150 471.900 802.950 ;
        RECT 473.700 795.600 474.600 802.950 ;
        RECT 479.550 802.050 480.450 805.950 ;
        RECT 491.100 805.050 492.900 806.850 ;
        RECT 494.400 805.050 495.600 810.300 ;
        RECT 507.000 807.450 511.050 808.050 ;
        RECT 497.100 805.050 498.900 806.850 ;
        RECT 506.550 805.950 511.050 807.450 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 493.950 802.950 496.050 805.050 ;
        RECT 496.950 802.950 499.050 805.050 ;
        RECT 475.950 800.550 480.450 802.050 ;
        RECT 475.950 799.950 480.000 800.550 ;
        RECT 478.950 798.450 481.050 799.050 ;
        RECT 490.950 798.450 493.050 799.050 ;
        RECT 478.950 797.550 493.050 798.450 ;
        RECT 478.950 796.950 481.050 797.550 ;
        RECT 490.950 796.950 493.050 797.550 ;
        RECT 380.400 783.600 382.200 789.600 ;
        RECT 398.400 783.600 400.200 789.600 ;
        RECT 418.800 783.600 420.600 789.600 ;
        RECT 437.400 783.600 439.200 789.600 ;
        RECT 452.400 783.600 454.200 789.600 ;
        RECT 467.400 783.600 469.200 789.600 ;
        RECT 473.400 783.600 475.200 795.600 ;
        RECT 494.400 789.600 495.600 802.950 ;
        RECT 506.550 802.050 507.450 805.950 ;
        RECT 512.100 805.050 513.900 806.850 ;
        RECT 519.000 805.050 520.050 812.400 ;
        RECT 533.400 811.950 541.200 813.300 ;
        RECT 542.400 812.400 544.200 818.400 ;
        RECT 557.400 813.300 559.200 818.400 ;
        RECT 563.400 813.300 565.200 818.400 ;
        RECT 542.400 810.300 543.600 812.400 ;
        RECT 557.400 811.950 565.200 813.300 ;
        RECT 566.400 812.400 568.200 818.400 ;
        RECT 578.400 813.300 580.200 818.400 ;
        RECT 584.400 813.300 586.200 818.400 ;
        RECT 566.400 810.300 567.600 812.400 ;
        RECT 578.400 811.950 586.200 813.300 ;
        RECT 587.400 812.400 589.200 818.400 ;
        RECT 601.800 815.400 603.600 818.400 ;
        RECT 587.400 810.300 588.600 812.400 ;
        RECT 539.850 809.250 543.600 810.300 ;
        RECT 563.850 809.250 567.600 810.300 ;
        RECT 584.850 809.250 588.600 810.300 ;
        RECT 524.100 805.050 525.900 806.850 ;
        RECT 536.100 805.050 537.900 806.850 ;
        RECT 539.850 805.050 541.050 809.250 ;
        RECT 544.950 807.450 549.000 808.050 ;
        RECT 542.100 805.050 543.900 806.850 ;
        RECT 544.950 805.950 549.450 807.450 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 517.950 802.950 520.050 805.050 ;
        RECT 520.950 802.950 523.050 805.050 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 541.950 802.950 544.050 805.050 ;
        RECT 506.550 800.550 511.050 802.050 ;
        RECT 515.100 801.150 516.900 802.950 ;
        RECT 507.000 799.950 511.050 800.550 ;
        RECT 496.950 798.450 499.050 799.050 ;
        RECT 505.950 798.450 508.050 798.900 ;
        RECT 496.950 797.550 508.050 798.450 ;
        RECT 496.950 796.950 499.050 797.550 ;
        RECT 505.950 796.800 508.050 797.550 ;
        RECT 519.000 797.400 519.900 802.950 ;
        RECT 521.100 801.150 522.900 802.950 ;
        RECT 533.100 801.150 534.900 802.950 ;
        RECT 514.800 796.500 519.900 797.400 ;
        RECT 493.800 783.600 495.600 789.600 ;
        RECT 511.800 784.500 513.600 795.600 ;
        RECT 514.800 785.400 516.600 796.500 ;
        RECT 517.800 794.400 525.600 795.300 ;
        RECT 517.800 784.500 519.600 794.400 ;
        RECT 511.800 783.600 519.600 784.500 ;
        RECT 523.800 783.600 525.600 794.400 ;
        RECT 538.950 789.600 540.150 802.950 ;
        RECT 548.550 802.050 549.450 805.950 ;
        RECT 560.100 805.050 561.900 806.850 ;
        RECT 563.850 805.050 565.050 809.250 ;
        RECT 566.100 805.050 567.900 806.850 ;
        RECT 581.100 805.050 582.900 806.850 ;
        RECT 584.850 805.050 586.050 809.250 ;
        RECT 587.100 805.050 588.900 806.850 ;
        RECT 602.400 805.050 603.600 815.400 ;
        RECT 627.000 812.400 628.800 818.400 ;
        RECT 646.800 815.400 648.600 818.400 ;
        RECT 620.100 805.050 621.900 806.850 ;
        RECT 627.000 805.050 628.050 812.400 ;
        RECT 632.100 805.050 633.900 806.850 ;
        RECT 647.400 805.050 648.600 815.400 ;
        RECT 662.400 811.200 664.200 818.400 ;
        RECT 680.400 811.200 682.200 818.400 ;
        RECT 703.800 811.200 705.600 818.400 ;
        RECT 722.400 815.400 724.200 818.400 ;
        RECT 662.400 810.300 666.600 811.200 ;
        RECT 680.400 810.300 684.600 811.200 ;
        RECT 652.950 807.450 657.000 808.050 ;
        RECT 652.950 805.950 657.450 807.450 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 565.950 802.950 568.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 586.950 802.950 589.050 805.050 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 604.950 802.950 607.050 805.050 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 544.950 800.550 549.450 802.050 ;
        RECT 557.100 801.150 558.900 802.950 ;
        RECT 544.950 799.950 549.000 800.550 ;
        RECT 562.950 789.600 564.150 802.950 ;
        RECT 578.100 801.150 579.900 802.950 ;
        RECT 583.950 789.600 585.150 802.950 ;
        RECT 602.400 789.600 603.600 802.950 ;
        RECT 605.100 801.150 606.900 802.950 ;
        RECT 623.100 801.150 624.900 802.950 ;
        RECT 627.000 797.400 627.900 802.950 ;
        RECT 629.100 801.150 630.900 802.950 ;
        RECT 634.950 801.450 637.050 802.050 ;
        RECT 640.950 801.450 643.050 802.050 ;
        RECT 634.950 800.550 643.050 801.450 ;
        RECT 634.950 799.950 637.050 800.550 ;
        RECT 640.950 799.950 643.050 800.550 ;
        RECT 622.800 796.500 627.900 797.400 ;
        RECT 538.800 783.600 540.600 789.600 ;
        RECT 562.800 783.600 564.600 789.600 ;
        RECT 583.800 783.600 585.600 789.600 ;
        RECT 601.800 783.600 603.600 789.600 ;
        RECT 619.800 784.500 621.600 795.600 ;
        RECT 622.800 785.400 624.600 796.500 ;
        RECT 625.800 794.400 633.600 795.300 ;
        RECT 625.800 784.500 627.600 794.400 ;
        RECT 619.800 783.600 627.600 784.500 ;
        RECT 631.800 783.600 633.600 794.400 ;
        RECT 647.400 789.600 648.600 802.950 ;
        RECT 650.100 801.150 651.900 802.950 ;
        RECT 656.550 802.050 657.450 805.950 ;
        RECT 662.100 805.050 663.900 806.850 ;
        RECT 665.400 805.050 666.600 810.300 ;
        RECT 668.100 805.050 669.900 806.850 ;
        RECT 680.100 805.050 681.900 806.850 ;
        RECT 683.400 805.050 684.600 810.300 ;
        RECT 701.400 810.300 705.600 811.200 ;
        RECT 686.100 805.050 687.900 806.850 ;
        RECT 698.100 805.050 699.900 806.850 ;
        RECT 701.400 805.050 702.600 810.300 ;
        RECT 704.100 805.050 705.900 806.850 ;
        RECT 722.700 805.050 723.600 815.400 ;
        RECT 747.300 812.700 749.100 817.200 ;
        RECT 754.800 814.200 756.600 817.200 ;
        RECT 747.000 811.800 749.100 812.700 ;
        RECT 747.000 805.050 747.900 811.800 ;
        RECT 755.700 810.900 756.600 814.200 ;
        RECT 749.400 810.000 756.600 810.900 ;
        RECT 766.800 812.400 768.600 818.400 ;
        RECT 772.800 815.400 774.600 818.400 ;
        RECT 788.400 815.400 790.200 818.400 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 682.950 802.950 685.050 805.050 ;
        RECT 685.950 802.950 688.050 805.050 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 721.950 802.950 724.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 742.950 802.950 745.050 805.050 ;
        RECT 745.950 802.950 748.050 805.050 ;
        RECT 749.400 802.950 750.600 810.000 ;
        RECT 755.100 805.050 756.900 806.850 ;
        RECT 766.800 805.050 768.000 812.400 ;
        RECT 773.400 811.500 774.600 815.400 ;
        RECT 768.900 810.600 774.600 811.500 ;
        RECT 768.900 809.700 770.850 810.600 ;
        RECT 751.950 802.950 754.050 805.050 ;
        RECT 754.950 802.950 757.050 805.050 ;
        RECT 766.800 802.950 769.050 805.050 ;
        RECT 652.950 800.550 657.450 802.050 ;
        RECT 652.950 799.950 657.000 800.550 ;
        RECT 665.400 789.600 666.600 802.950 ;
        RECT 683.400 789.600 684.600 802.950 ;
        RECT 646.800 783.600 648.600 789.600 ;
        RECT 664.800 783.600 666.600 789.600 ;
        RECT 682.800 783.600 684.600 789.600 ;
        RECT 701.400 789.600 702.600 802.950 ;
        RECT 719.100 801.150 720.900 802.950 ;
        RECT 703.950 798.450 706.050 799.050 ;
        RECT 715.950 798.450 718.050 799.050 ;
        RECT 703.950 797.550 718.050 798.450 ;
        RECT 703.950 796.950 706.050 797.550 ;
        RECT 715.950 796.950 718.050 797.550 ;
        RECT 722.700 795.600 723.600 802.950 ;
        RECT 725.100 801.150 726.900 802.950 ;
        RECT 743.100 801.150 744.900 802.950 ;
        RECT 722.700 794.400 726.300 795.600 ;
        RECT 701.400 783.600 703.200 789.600 ;
        RECT 724.500 783.600 726.300 794.400 ;
        RECT 747.000 795.000 747.900 802.950 ;
        RECT 748.950 801.150 750.750 802.950 ;
        RECT 752.100 801.150 753.900 802.950 ;
        RECT 749.250 796.800 750.450 801.150 ;
        RECT 749.250 795.900 756.600 796.800 ;
        RECT 747.000 794.100 749.100 795.000 ;
        RECT 747.300 784.800 749.100 794.100 ;
        RECT 755.700 790.800 756.600 795.900 ;
        RECT 754.800 784.800 756.600 790.800 ;
        RECT 766.800 795.600 768.000 802.950 ;
        RECT 769.950 798.300 770.850 809.700 ;
        RECT 788.700 805.050 789.600 815.400 ;
        RECT 805.800 812.400 807.600 818.400 ;
        RECT 806.400 810.300 807.600 812.400 ;
        RECT 808.800 813.300 810.600 818.400 ;
        RECT 814.800 813.300 816.600 818.400 ;
        RECT 808.800 811.950 816.600 813.300 ;
        RECT 824.400 813.300 826.200 818.400 ;
        RECT 830.400 813.300 832.200 818.400 ;
        RECT 824.400 811.950 832.200 813.300 ;
        RECT 833.400 812.400 835.200 818.400 ;
        RECT 848.400 813.300 850.200 818.400 ;
        RECT 854.400 813.300 856.200 818.400 ;
        RECT 833.400 810.300 834.600 812.400 ;
        RECT 848.400 811.950 856.200 813.300 ;
        RECT 857.400 812.400 859.200 818.400 ;
        RECT 872.400 815.400 874.200 818.400 ;
        RECT 889.800 815.400 891.600 818.400 ;
        RECT 857.400 810.300 858.600 812.400 ;
        RECT 806.400 809.250 810.150 810.300 ;
        RECT 806.100 805.050 807.900 806.850 ;
        RECT 808.950 805.050 810.150 809.250 ;
        RECT 830.850 809.250 834.600 810.300 ;
        RECT 854.850 809.250 858.600 810.300 ;
        RECT 812.100 805.050 813.900 806.850 ;
        RECT 827.100 805.050 828.900 806.850 ;
        RECT 830.850 805.050 832.050 809.250 ;
        RECT 844.950 807.450 847.050 808.050 ;
        RECT 833.100 805.050 834.900 806.850 ;
        RECT 839.550 806.550 847.050 807.450 ;
        RECT 772.950 802.950 775.050 805.050 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 787.950 802.950 790.050 805.050 ;
        RECT 790.950 802.950 793.050 805.050 ;
        RECT 805.950 802.950 808.050 805.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 829.950 802.950 832.050 805.050 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 773.100 801.150 774.900 802.950 ;
        RECT 785.100 801.150 786.900 802.950 ;
        RECT 768.900 797.400 770.850 798.300 ;
        RECT 768.900 796.500 774.600 797.400 ;
        RECT 766.800 783.600 768.600 795.600 ;
        RECT 773.400 789.600 774.600 796.500 ;
        RECT 788.700 795.600 789.600 802.950 ;
        RECT 791.100 801.150 792.900 802.950 ;
        RECT 788.700 794.400 792.300 795.600 ;
        RECT 772.800 783.600 774.600 789.600 ;
        RECT 790.500 783.600 792.300 794.400 ;
        RECT 809.850 789.600 811.050 802.950 ;
        RECT 815.100 801.150 816.900 802.950 ;
        RECT 824.100 801.150 825.900 802.950 ;
        RECT 829.950 789.600 831.150 802.950 ;
        RECT 839.550 802.050 840.450 806.550 ;
        RECT 844.950 805.950 847.050 806.550 ;
        RECT 851.100 805.050 852.900 806.850 ;
        RECT 854.850 805.050 856.050 809.250 ;
        RECT 857.100 805.050 858.900 806.850 ;
        RECT 872.400 805.050 873.600 815.400 ;
        RECT 890.400 805.050 891.600 815.400 ;
        RECT 907.800 812.400 909.600 818.400 ;
        RECT 913.800 815.400 915.600 818.400 ;
        RECT 907.800 805.050 909.000 812.400 ;
        RECT 914.400 811.500 915.600 815.400 ;
        RECT 909.900 810.600 915.600 811.500 ;
        RECT 909.900 809.700 911.850 810.600 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 856.950 802.950 859.050 805.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 889.950 802.950 892.050 805.050 ;
        RECT 892.950 802.950 895.050 805.050 ;
        RECT 907.800 802.950 910.050 805.050 ;
        RECT 835.950 800.550 840.450 802.050 ;
        RECT 848.100 801.150 849.900 802.950 ;
        RECT 835.950 799.950 840.000 800.550 ;
        RECT 853.950 789.600 855.150 802.950 ;
        RECT 869.100 801.150 870.900 802.950 ;
        RECT 872.400 789.600 873.600 802.950 ;
        RECT 890.400 789.600 891.600 802.950 ;
        RECT 893.100 801.150 894.900 802.950 ;
        RECT 809.400 783.600 811.200 789.600 ;
        RECT 829.800 783.600 831.600 789.600 ;
        RECT 853.800 783.600 855.600 789.600 ;
        RECT 872.400 783.600 874.200 789.600 ;
        RECT 889.800 783.600 891.600 789.600 ;
        RECT 907.800 795.600 909.000 802.950 ;
        RECT 910.950 798.300 911.850 809.700 ;
        RECT 913.950 802.950 916.050 805.050 ;
        RECT 914.100 801.150 915.900 802.950 ;
        RECT 909.900 797.400 911.850 798.300 ;
        RECT 909.900 796.500 915.600 797.400 ;
        RECT 907.800 783.600 909.600 795.600 ;
        RECT 914.400 789.600 915.600 796.500 ;
        RECT 913.800 783.600 915.600 789.600 ;
        RECT 17.400 773.400 19.200 779.400 ;
        RECT 40.800 773.400 42.600 779.400 ;
        RECT 58.800 773.400 60.600 779.400 ;
        RECT 17.850 760.050 19.050 773.400 ;
        RECT 23.100 760.050 24.900 761.850 ;
        RECT 35.100 760.050 36.900 761.850 ;
        RECT 40.950 760.050 42.150 773.400 ;
        RECT 59.700 773.100 60.600 773.400 ;
        RECT 64.800 773.400 66.600 779.400 ;
        RECT 82.800 773.400 84.600 779.400 ;
        RECT 97.800 773.400 99.600 779.400 ;
        RECT 64.800 773.100 66.300 773.400 ;
        RECT 59.700 772.200 66.300 773.100 ;
        RECT 59.700 760.050 60.600 772.200 ;
        RECT 65.100 760.050 66.900 761.850 ;
        RECT 83.400 760.050 84.600 773.400 ;
        RECT 98.700 773.100 99.600 773.400 ;
        RECT 103.800 773.400 105.600 779.400 ;
        RECT 121.800 773.400 123.600 779.400 ;
        RECT 136.800 773.400 138.600 779.400 ;
        RECT 103.800 773.100 105.300 773.400 ;
        RECT 98.700 772.200 105.300 773.100 ;
        RECT 86.100 760.050 87.900 761.850 ;
        RECT 98.700 760.050 99.600 772.200 ;
        RECT 104.100 760.050 105.900 761.850 ;
        RECT 122.400 760.050 123.600 773.400 ;
        RECT 137.700 773.100 138.600 773.400 ;
        RECT 142.800 773.400 144.600 779.400 ;
        RECT 161.400 773.400 163.200 779.400 ;
        RECT 142.800 773.100 144.300 773.400 ;
        RECT 137.700 772.200 144.300 773.100 ;
        RECT 125.100 760.050 126.900 761.850 ;
        RECT 137.700 760.050 138.600 772.200 ;
        RECT 143.100 760.050 144.900 761.850 ;
        RECT 161.850 760.050 163.050 773.400 ;
        RECT 182.700 768.600 184.500 779.400 ;
        RECT 200.400 768.600 202.200 779.400 ;
        RECT 206.400 778.500 214.200 779.400 ;
        RECT 206.400 768.600 208.200 778.500 ;
        RECT 182.700 767.400 186.300 768.600 ;
        RECT 200.400 767.700 208.200 768.600 ;
        RECT 167.100 760.050 168.900 761.850 ;
        RECT 182.100 760.050 183.900 761.850 ;
        RECT 185.400 760.050 186.300 767.400 ;
        RECT 209.400 766.500 211.200 777.600 ;
        RECT 212.400 767.400 214.200 778.500 ;
        RECT 229.800 778.500 237.600 779.400 ;
        RECT 229.800 767.400 231.600 778.500 ;
        RECT 206.100 765.600 211.200 766.500 ;
        RECT 232.800 766.500 234.600 777.600 ;
        RECT 235.800 768.600 237.600 778.500 ;
        RECT 241.800 768.600 243.600 779.400 ;
        RECT 259.800 773.400 261.600 779.400 ;
        RECT 277.800 773.400 279.600 779.400 ;
        RECT 235.800 767.700 243.600 768.600 ;
        RECT 232.800 765.600 237.900 766.500 ;
        RECT 188.100 760.050 189.900 761.850 ;
        RECT 203.100 760.050 204.900 761.850 ;
        RECT 206.100 760.050 207.000 765.600 ;
        RECT 209.100 760.050 210.900 761.850 ;
        RECT 233.100 760.050 234.900 761.850 ;
        RECT 237.000 760.050 237.900 765.600 ;
        RECT 252.000 762.450 256.050 763.050 ;
        RECT 239.100 760.050 240.900 761.850 ;
        RECT 251.550 760.950 256.050 762.450 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 22.950 757.950 25.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 43.950 757.950 46.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 64.950 757.950 67.050 760.050 ;
        RECT 67.950 757.950 70.050 760.050 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 85.950 757.950 88.050 760.050 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 103.950 757.950 106.050 760.050 ;
        RECT 106.950 757.950 109.050 760.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 199.950 757.950 202.050 760.050 ;
        RECT 202.950 757.950 205.050 760.050 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 14.100 756.150 15.900 757.950 ;
        RECT 16.950 753.750 18.150 757.950 ;
        RECT 20.100 756.150 21.900 757.950 ;
        RECT 38.100 756.150 39.900 757.950 ;
        RECT 14.400 752.700 18.150 753.750 ;
        RECT 41.850 753.750 43.050 757.950 ;
        RECT 44.100 756.150 45.900 757.950 ;
        RECT 59.700 754.200 60.600 757.950 ;
        RECT 62.100 756.150 63.900 757.950 ;
        RECT 68.100 756.150 69.900 757.950 ;
        RECT 41.850 752.700 45.600 753.750 ;
        RECT 59.700 753.000 63.000 754.200 ;
        RECT 14.400 750.600 15.600 752.700 ;
        RECT 13.800 744.600 15.600 750.600 ;
        RECT 16.800 749.700 24.600 751.050 ;
        RECT 16.800 744.600 18.600 749.700 ;
        RECT 22.800 744.600 24.600 749.700 ;
        RECT 35.400 749.700 43.200 751.050 ;
        RECT 35.400 744.600 37.200 749.700 ;
        RECT 41.400 744.600 43.200 749.700 ;
        RECT 44.400 750.600 45.600 752.700 ;
        RECT 44.400 744.600 46.200 750.600 ;
        RECT 61.200 744.600 63.000 753.000 ;
        RECT 83.400 747.600 84.600 757.950 ;
        RECT 98.700 754.200 99.600 757.950 ;
        RECT 101.100 756.150 102.900 757.950 ;
        RECT 107.100 756.150 108.900 757.950 ;
        RECT 98.700 753.000 102.000 754.200 ;
        RECT 82.800 744.600 84.600 747.600 ;
        RECT 100.200 744.600 102.000 753.000 ;
        RECT 122.400 747.600 123.600 757.950 ;
        RECT 137.700 754.200 138.600 757.950 ;
        RECT 140.100 756.150 141.900 757.950 ;
        RECT 146.100 756.150 147.900 757.950 ;
        RECT 158.100 756.150 159.900 757.950 ;
        RECT 137.700 753.000 141.000 754.200 ;
        RECT 160.950 753.750 162.150 757.950 ;
        RECT 164.100 756.150 165.900 757.950 ;
        RECT 172.950 756.450 175.050 757.050 ;
        RECT 178.950 756.450 181.050 757.050 ;
        RECT 172.950 755.550 181.050 756.450 ;
        RECT 172.950 754.950 175.050 755.550 ;
        RECT 178.950 754.950 181.050 755.550 ;
        RECT 121.800 744.600 123.600 747.600 ;
        RECT 139.200 744.600 141.000 753.000 ;
        RECT 158.400 752.700 162.150 753.750 ;
        RECT 158.400 750.600 159.600 752.700 ;
        RECT 157.800 744.600 159.600 750.600 ;
        RECT 160.800 749.700 168.600 751.050 ;
        RECT 160.800 744.600 162.600 749.700 ;
        RECT 166.800 744.600 168.600 749.700 ;
        RECT 185.400 747.600 186.300 757.950 ;
        RECT 200.100 756.150 201.900 757.950 ;
        RECT 205.950 750.600 207.000 757.950 ;
        RECT 212.100 756.150 213.900 757.950 ;
        RECT 230.100 756.150 231.900 757.950 ;
        RECT 208.950 753.450 211.050 754.050 ;
        RECT 232.950 753.450 235.050 754.050 ;
        RECT 208.950 752.550 235.050 753.450 ;
        RECT 208.950 751.950 211.050 752.550 ;
        RECT 232.950 751.950 235.050 752.550 ;
        RECT 184.800 744.600 186.600 747.600 ;
        RECT 205.200 744.600 207.000 750.600 ;
        RECT 237.000 750.600 238.050 757.950 ;
        RECT 242.100 756.150 243.900 757.950 ;
        RECT 251.550 757.050 252.450 760.950 ;
        RECT 260.400 760.050 261.600 773.400 ;
        RECT 278.400 760.050 279.600 773.400 ;
        RECT 293.400 767.400 295.200 779.400 ;
        RECT 300.900 768.900 302.700 779.400 ;
        RECT 320.400 773.400 322.200 779.400 ;
        RECT 341.400 773.400 343.200 779.400 ;
        RECT 358.800 773.400 360.600 779.400 ;
        RECT 300.900 767.400 303.300 768.900 ;
        RECT 293.400 765.900 294.600 767.400 ;
        RECT 293.400 764.700 300.600 765.900 ;
        RECT 298.800 764.100 300.600 764.700 ;
        RECT 296.100 760.050 297.900 761.850 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 251.550 755.550 256.050 757.050 ;
        RECT 257.100 756.150 258.900 757.950 ;
        RECT 252.000 754.950 256.050 755.550 ;
        RECT 260.400 752.700 261.600 757.950 ;
        RECT 263.100 756.150 264.900 757.950 ;
        RECT 275.100 756.150 276.900 757.950 ;
        RECT 278.400 752.700 279.600 757.950 ;
        RECT 281.100 756.150 282.900 757.950 ;
        RECT 293.100 756.150 294.900 757.950 ;
        RECT 299.700 753.600 300.600 764.100 ;
        RECT 301.950 760.050 303.300 767.400 ;
        RECT 320.400 760.050 321.600 773.400 ;
        RECT 338.100 760.050 339.900 761.850 ;
        RECT 341.400 760.050 342.600 773.400 ;
        RECT 359.400 760.050 360.600 773.400 ;
        RECT 379.800 767.400 383.100 779.400 ;
        RECT 401.700 768.600 403.500 779.400 ;
        RECT 401.700 767.400 405.300 768.600 ;
        RECT 421.800 767.400 423.600 779.400 ;
        RECT 427.800 773.400 429.600 779.400 ;
        RECT 448.800 773.400 450.600 779.400 ;
        RECT 469.800 773.400 471.600 779.400 ;
        RECT 487.800 778.500 495.600 779.400 ;
        RECT 364.950 762.450 369.000 763.050 ;
        RECT 362.100 760.050 363.900 761.850 ;
        RECT 364.950 760.950 369.450 762.450 ;
        RECT 301.950 757.950 304.050 760.050 ;
        RECT 316.950 757.950 319.050 760.050 ;
        RECT 319.950 757.950 322.050 760.050 ;
        RECT 322.950 757.950 325.050 760.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 340.950 757.950 343.050 760.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 361.950 757.950 364.050 760.050 ;
        RECT 298.800 752.700 300.600 753.600 ;
        RECT 257.400 751.800 261.600 752.700 ;
        RECT 275.400 751.800 279.600 752.700 ;
        RECT 297.300 751.800 300.600 752.700 ;
        RECT 237.000 744.600 238.800 750.600 ;
        RECT 257.400 744.600 259.200 751.800 ;
        RECT 275.400 744.600 277.200 751.800 ;
        RECT 297.300 747.600 298.200 751.800 ;
        RECT 303.000 750.600 304.050 757.950 ;
        RECT 317.100 756.150 318.900 757.950 ;
        RECT 320.400 752.700 321.600 757.950 ;
        RECT 323.100 756.150 324.900 757.950 ;
        RECT 320.400 751.800 324.600 752.700 ;
        RECT 296.400 744.600 298.200 747.600 ;
        RECT 302.400 744.600 304.200 750.600 ;
        RECT 322.800 744.600 324.600 751.800 ;
        RECT 341.400 747.600 342.600 757.950 ;
        RECT 359.400 747.600 360.600 757.950 ;
        RECT 368.550 757.050 369.450 760.950 ;
        RECT 374.100 760.050 375.900 761.850 ;
        RECT 380.700 760.050 381.900 767.400 ;
        RECT 388.950 762.450 391.050 763.050 ;
        RECT 386.100 760.050 387.900 761.850 ;
        RECT 388.950 761.550 396.450 762.450 ;
        RECT 388.950 760.950 391.050 761.550 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 382.950 757.950 385.050 760.050 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 368.550 755.550 373.050 757.050 ;
        RECT 377.100 756.150 378.900 757.950 ;
        RECT 369.000 754.950 373.050 755.550 ;
        RECT 380.700 753.300 382.050 757.950 ;
        RECT 383.100 756.150 384.900 757.950 ;
        RECT 395.550 757.050 396.450 761.550 ;
        RECT 401.100 760.050 402.900 761.850 ;
        RECT 404.400 760.050 405.300 767.400 ;
        RECT 407.100 760.050 408.900 761.850 ;
        RECT 422.400 760.050 423.300 767.400 ;
        RECT 425.100 760.050 426.900 761.850 ;
        RECT 400.950 757.950 403.050 760.050 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 421.950 757.950 424.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 395.550 755.550 400.050 757.050 ;
        RECT 396.000 754.950 400.050 755.550 ;
        RECT 377.400 752.100 382.050 753.300 ;
        RECT 377.400 750.600 378.300 752.100 ;
        RECT 341.400 744.600 343.200 747.600 ;
        RECT 358.800 744.600 360.600 747.600 ;
        RECT 373.800 745.500 375.600 750.600 ;
        RECT 376.800 746.400 378.600 750.600 ;
        RECT 379.800 750.000 387.600 750.900 ;
        RECT 379.800 745.500 381.600 750.000 ;
        RECT 373.800 744.600 381.600 745.500 ;
        RECT 385.800 744.600 387.600 750.000 ;
        RECT 404.400 747.600 405.300 757.950 ;
        RECT 409.950 756.450 412.050 757.050 ;
        RECT 415.950 756.450 418.050 757.050 ;
        RECT 409.950 755.550 418.050 756.450 ;
        RECT 409.950 754.950 412.050 755.550 ;
        RECT 415.950 754.950 418.050 755.550 ;
        RECT 422.400 750.600 423.300 757.950 ;
        RECT 428.700 753.300 429.600 773.400 ;
        RECT 449.400 760.050 450.600 773.400 ;
        RECT 464.100 760.050 465.900 761.850 ;
        RECT 469.950 760.050 471.150 773.400 ;
        RECT 487.800 767.400 489.600 778.500 ;
        RECT 490.800 766.500 492.600 777.600 ;
        RECT 493.800 768.600 495.600 778.500 ;
        RECT 499.800 768.600 501.600 779.400 ;
        RECT 518.400 773.400 520.200 779.400 ;
        RECT 541.800 773.400 543.600 779.400 ;
        RECT 493.800 767.700 501.600 768.600 ;
        RECT 490.800 765.600 495.900 766.500 ;
        RECT 491.100 760.050 492.900 761.850 ;
        RECT 495.000 760.050 495.900 765.600 ;
        RECT 497.100 760.050 498.900 761.850 ;
        RECT 518.850 760.050 520.050 773.400 ;
        RECT 526.950 762.450 529.050 763.050 ;
        RECT 532.950 762.450 535.050 762.900 ;
        RECT 524.100 760.050 525.900 761.850 ;
        RECT 526.950 761.550 535.050 762.450 ;
        RECT 526.950 760.950 529.050 761.550 ;
        RECT 532.950 760.800 535.050 761.550 ;
        RECT 542.400 760.050 543.600 773.400 ;
        RECT 559.800 778.500 567.600 779.400 ;
        RECT 559.800 767.400 561.600 778.500 ;
        RECT 562.800 766.500 564.600 777.600 ;
        RECT 565.800 768.600 567.600 778.500 ;
        RECT 571.800 768.600 573.600 779.400 ;
        RECT 565.800 767.700 573.600 768.600 ;
        RECT 583.800 767.400 585.600 779.400 ;
        RECT 589.800 773.400 591.600 779.400 ;
        RECT 562.800 765.600 567.900 766.500 ;
        RECT 547.950 762.450 552.000 763.050 ;
        RECT 547.950 760.950 552.450 762.450 ;
        RECT 430.950 757.950 433.050 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 463.950 757.950 466.050 760.050 ;
        RECT 466.950 757.950 469.050 760.050 ;
        RECT 469.950 757.950 472.050 760.050 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 487.950 757.950 490.050 760.050 ;
        RECT 490.950 757.950 493.050 760.050 ;
        RECT 493.950 757.950 496.050 760.050 ;
        RECT 496.950 757.950 499.050 760.050 ;
        RECT 499.950 757.950 502.050 760.050 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 517.950 757.950 520.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 538.950 757.950 541.050 760.050 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 431.100 756.150 432.900 757.950 ;
        RECT 446.100 756.150 447.900 757.950 ;
        RECT 425.100 752.400 432.600 753.300 ;
        RECT 449.400 752.700 450.600 757.950 ;
        RECT 452.100 756.150 453.900 757.950 ;
        RECT 467.100 756.150 468.900 757.950 ;
        RECT 470.850 753.750 472.050 757.950 ;
        RECT 473.100 756.150 474.900 757.950 ;
        RECT 488.100 756.150 489.900 757.950 ;
        RECT 470.850 752.700 474.600 753.750 ;
        RECT 425.100 751.500 426.900 752.400 ;
        RECT 422.400 748.800 425.100 750.600 ;
        RECT 403.800 744.600 405.600 747.600 ;
        RECT 423.300 744.600 425.100 748.800 ;
        RECT 430.800 744.600 432.600 752.400 ;
        RECT 446.400 751.800 450.600 752.700 ;
        RECT 446.400 744.600 448.200 751.800 ;
        RECT 464.400 749.700 472.200 751.050 ;
        RECT 464.400 744.600 466.200 749.700 ;
        RECT 470.400 744.600 472.200 749.700 ;
        RECT 473.400 750.600 474.600 752.700 ;
        RECT 481.950 753.450 484.050 754.050 ;
        RECT 487.950 753.450 490.050 754.050 ;
        RECT 481.950 752.550 490.050 753.450 ;
        RECT 481.950 751.950 484.050 752.550 ;
        RECT 487.950 751.950 490.050 752.550 ;
        RECT 495.000 750.600 496.050 757.950 ;
        RECT 500.100 756.150 501.900 757.950 ;
        RECT 515.100 756.150 516.900 757.950 ;
        RECT 517.950 753.750 519.150 757.950 ;
        RECT 521.100 756.150 522.900 757.950 ;
        RECT 539.100 756.150 540.900 757.950 ;
        RECT 515.400 752.700 519.150 753.750 ;
        RECT 542.400 752.700 543.600 757.950 ;
        RECT 545.100 756.150 546.900 757.950 ;
        RECT 551.550 757.050 552.450 760.950 ;
        RECT 563.100 760.050 564.900 761.850 ;
        RECT 567.000 760.050 567.900 765.600 ;
        RECT 569.100 760.050 570.900 761.850 ;
        RECT 584.400 760.050 585.300 767.400 ;
        RECT 587.100 760.050 588.900 761.850 ;
        RECT 559.950 757.950 562.050 760.050 ;
        RECT 562.950 757.950 565.050 760.050 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 586.950 757.950 589.050 760.050 ;
        RECT 547.950 755.550 552.450 757.050 ;
        RECT 560.100 756.150 561.900 757.950 ;
        RECT 547.950 754.950 552.000 755.550 ;
        RECT 515.400 750.600 516.600 752.700 ;
        RECT 539.400 751.800 543.600 752.700 ;
        RECT 473.400 744.600 475.200 750.600 ;
        RECT 495.000 744.600 496.800 750.600 ;
        RECT 514.800 744.600 516.600 750.600 ;
        RECT 517.800 749.700 525.600 751.050 ;
        RECT 517.800 744.600 519.600 749.700 ;
        RECT 523.800 744.600 525.600 749.700 ;
        RECT 539.400 744.600 541.200 751.800 ;
        RECT 567.000 750.600 568.050 757.950 ;
        RECT 572.100 756.150 573.900 757.950 ;
        RECT 584.400 750.600 585.300 757.950 ;
        RECT 590.700 753.300 591.600 773.400 ;
        RECT 605.400 768.600 607.200 779.400 ;
        RECT 611.400 778.500 619.200 779.400 ;
        RECT 611.400 768.600 613.200 778.500 ;
        RECT 605.400 767.700 613.200 768.600 ;
        RECT 614.400 766.500 616.200 777.600 ;
        RECT 617.400 767.400 619.200 778.500 ;
        RECT 622.950 777.450 625.050 778.050 ;
        RECT 628.950 777.450 631.050 778.050 ;
        RECT 622.950 776.550 631.050 777.450 ;
        RECT 622.950 775.950 625.050 776.550 ;
        RECT 628.950 775.950 631.050 776.550 ;
        RECT 632.400 768.600 634.200 779.400 ;
        RECT 638.400 778.500 646.200 779.400 ;
        RECT 638.400 768.600 640.200 778.500 ;
        RECT 632.400 767.700 640.200 768.600 ;
        RECT 641.400 766.500 643.200 777.600 ;
        RECT 644.400 767.400 646.200 778.500 ;
        RECT 659.400 773.400 661.200 779.400 ;
        RECT 680.400 773.400 682.200 779.400 ;
        RECT 607.950 765.450 610.050 766.050 ;
        RECT 599.550 764.550 610.050 765.450 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 593.100 756.150 594.900 757.950 ;
        RECT 599.550 757.050 600.450 764.550 ;
        RECT 607.950 763.950 610.050 764.550 ;
        RECT 611.100 765.600 616.200 766.500 ;
        RECT 638.100 765.600 643.200 766.500 ;
        RECT 608.100 760.050 609.900 761.850 ;
        RECT 611.100 760.050 612.000 765.600 ;
        RECT 627.000 762.450 631.050 763.050 ;
        RECT 614.100 760.050 615.900 761.850 ;
        RECT 626.550 760.950 631.050 762.450 ;
        RECT 604.950 757.950 607.050 760.050 ;
        RECT 607.950 757.950 610.050 760.050 ;
        RECT 610.950 757.950 613.050 760.050 ;
        RECT 613.950 757.950 616.050 760.050 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 595.950 755.550 600.450 757.050 ;
        RECT 605.100 756.150 606.900 757.950 ;
        RECT 595.950 754.950 600.000 755.550 ;
        RECT 587.100 752.400 594.600 753.300 ;
        RECT 587.100 751.500 588.900 752.400 ;
        RECT 567.000 744.600 568.800 750.600 ;
        RECT 584.400 748.800 587.100 750.600 ;
        RECT 585.300 744.600 587.100 748.800 ;
        RECT 592.800 744.600 594.600 752.400 ;
        RECT 610.950 750.600 612.000 757.950 ;
        RECT 617.100 756.150 618.900 757.950 ;
        RECT 626.550 757.050 627.450 760.950 ;
        RECT 635.100 760.050 636.900 761.850 ;
        RECT 638.100 760.050 639.000 765.600 ;
        RECT 641.100 760.050 642.900 761.850 ;
        RECT 659.400 760.050 660.600 773.400 ;
        RECT 631.950 757.950 634.050 760.050 ;
        RECT 634.950 757.950 637.050 760.050 ;
        RECT 637.950 757.950 640.050 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 626.550 755.550 631.050 757.050 ;
        RECT 632.100 756.150 633.900 757.950 ;
        RECT 627.000 754.950 631.050 755.550 ;
        RECT 637.950 750.600 639.000 757.950 ;
        RECT 644.100 756.150 645.900 757.950 ;
        RECT 656.100 756.150 657.900 757.950 ;
        RECT 659.400 752.700 660.600 757.950 ;
        RECT 662.100 756.150 663.900 757.950 ;
        RECT 677.100 756.150 678.900 757.950 ;
        RECT 680.400 753.300 681.300 773.400 ;
        RECT 686.400 767.400 688.200 779.400 ;
        RECT 706.800 773.400 708.600 779.400 ;
        RECT 727.800 773.400 729.600 779.400 ;
        RECT 749.400 773.400 751.200 779.400 ;
        RECT 770.400 773.400 772.200 779.400 ;
        RECT 683.100 760.050 684.900 761.850 ;
        RECT 686.700 760.050 687.600 767.400 ;
        RECT 701.100 760.050 702.900 761.850 ;
        RECT 706.950 760.050 708.150 773.400 ;
        RECT 712.950 762.450 717.000 763.050 ;
        RECT 712.950 760.950 717.450 762.450 ;
        RECT 682.950 757.950 685.050 760.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 659.400 751.800 663.600 752.700 ;
        RECT 610.200 744.600 612.000 750.600 ;
        RECT 637.200 744.600 639.000 750.600 ;
        RECT 661.800 744.600 663.600 751.800 ;
        RECT 677.400 752.400 684.900 753.300 ;
        RECT 677.400 744.600 679.200 752.400 ;
        RECT 683.100 751.500 684.900 752.400 ;
        RECT 686.700 750.600 687.600 757.950 ;
        RECT 704.100 756.150 705.900 757.950 ;
        RECT 707.850 753.750 709.050 757.950 ;
        RECT 710.100 756.150 711.900 757.950 ;
        RECT 716.550 757.050 717.450 760.950 ;
        RECT 722.100 760.050 723.900 761.850 ;
        RECT 727.950 760.050 729.150 773.400 ;
        RECT 749.400 760.050 750.600 773.400 ;
        RECT 766.950 765.450 769.050 766.050 ;
        RECT 758.550 764.550 769.050 765.450 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 745.950 757.950 748.050 760.050 ;
        RECT 748.950 757.950 751.050 760.050 ;
        RECT 751.950 757.950 754.050 760.050 ;
        RECT 716.550 755.550 721.050 757.050 ;
        RECT 725.100 756.150 726.900 757.950 ;
        RECT 717.000 754.950 721.050 755.550 ;
        RECT 728.850 753.750 730.050 757.950 ;
        RECT 731.100 756.150 732.900 757.950 ;
        RECT 746.100 756.150 747.900 757.950 ;
        RECT 707.850 752.700 711.600 753.750 ;
        RECT 728.850 752.700 732.600 753.750 ;
        RECT 684.900 748.800 687.600 750.600 ;
        RECT 701.400 749.700 709.200 751.050 ;
        RECT 684.900 744.600 686.700 748.800 ;
        RECT 701.400 744.600 703.200 749.700 ;
        RECT 707.400 744.600 709.200 749.700 ;
        RECT 710.400 750.600 711.600 752.700 ;
        RECT 710.400 744.600 712.200 750.600 ;
        RECT 722.400 749.700 730.200 751.050 ;
        RECT 722.400 744.600 724.200 749.700 ;
        RECT 728.400 744.600 730.200 749.700 ;
        RECT 731.400 750.600 732.600 752.700 ;
        RECT 749.400 752.700 750.600 757.950 ;
        RECT 752.100 756.150 753.900 757.950 ;
        RECT 758.550 757.050 759.450 764.550 ;
        RECT 766.950 763.950 769.050 764.550 ;
        RECT 770.850 760.050 772.050 773.400 ;
        RECT 788.400 768.300 790.200 779.400 ;
        RECT 794.400 768.300 796.200 779.400 ;
        RECT 788.400 767.400 796.200 768.300 ;
        RECT 797.400 767.400 799.200 779.400 ;
        RECT 811.800 773.400 813.600 779.400 ;
        RECT 778.950 762.450 783.000 763.050 ;
        RECT 776.100 760.050 777.900 761.850 ;
        RECT 778.950 760.950 783.450 762.450 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 769.950 757.950 772.050 760.050 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 775.950 757.950 778.050 760.050 ;
        RECT 754.950 755.550 759.450 757.050 ;
        RECT 767.100 756.150 768.900 757.950 ;
        RECT 754.950 754.950 759.000 755.550 ;
        RECT 769.950 753.750 771.150 757.950 ;
        RECT 773.100 756.150 774.900 757.950 ;
        RECT 767.400 752.700 771.150 753.750 ;
        RECT 782.550 753.450 783.450 760.950 ;
        RECT 791.100 760.050 792.900 761.850 ;
        RECT 797.700 760.050 798.600 767.400 ;
        RECT 807.000 762.450 811.050 763.050 ;
        RECT 806.550 760.950 811.050 762.450 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 793.950 757.950 796.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 788.100 756.150 789.900 757.950 ;
        RECT 794.100 756.150 795.900 757.950 ;
        RECT 787.950 753.450 790.050 754.050 ;
        RECT 749.400 751.800 753.600 752.700 ;
        RECT 731.400 744.600 733.200 750.600 ;
        RECT 751.800 744.600 753.600 751.800 ;
        RECT 767.400 750.600 768.600 752.700 ;
        RECT 782.550 752.550 790.050 753.450 ;
        RECT 787.950 751.950 790.050 752.550 ;
        RECT 766.800 744.600 768.600 750.600 ;
        RECT 769.800 749.700 777.600 751.050 ;
        RECT 797.700 750.600 798.600 757.950 ;
        RECT 799.950 756.450 802.050 757.050 ;
        RECT 806.550 756.450 807.450 760.950 ;
        RECT 812.400 760.050 813.600 773.400 ;
        RECT 827.400 768.300 829.200 779.400 ;
        RECT 833.400 768.300 835.200 779.400 ;
        RECT 827.400 767.400 835.200 768.300 ;
        RECT 836.400 767.400 838.200 779.400 ;
        RECT 851.400 768.300 853.200 779.400 ;
        RECT 857.400 768.300 859.200 779.400 ;
        RECT 851.400 767.400 859.200 768.300 ;
        RECT 860.400 767.400 862.200 779.400 ;
        RECT 881.400 773.400 883.200 779.400 ;
        RECT 901.800 773.400 903.600 779.400 ;
        RECT 815.100 760.050 816.900 761.850 ;
        RECT 830.100 760.050 831.900 761.850 ;
        RECT 836.700 760.050 837.600 767.400 ;
        RECT 854.100 760.050 855.900 761.850 ;
        RECT 860.700 760.050 861.600 767.400 ;
        RECT 881.850 760.050 883.050 773.400 ;
        RECT 887.100 760.050 888.900 761.850 ;
        RECT 896.100 760.050 897.900 761.850 ;
        RECT 901.950 760.050 903.150 773.400 ;
        RECT 811.950 757.950 814.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 826.950 757.950 829.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 832.950 757.950 835.050 760.050 ;
        RECT 835.950 757.950 838.050 760.050 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 856.950 757.950 859.050 760.050 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 877.950 757.950 880.050 760.050 ;
        RECT 880.950 757.950 883.050 760.050 ;
        RECT 883.950 757.950 886.050 760.050 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 895.950 757.950 898.050 760.050 ;
        RECT 898.950 757.950 901.050 760.050 ;
        RECT 901.950 757.950 904.050 760.050 ;
        RECT 904.950 757.950 907.050 760.050 ;
        RECT 799.950 755.550 807.450 756.450 ;
        RECT 799.950 754.950 802.050 755.550 ;
        RECT 769.800 744.600 771.600 749.700 ;
        RECT 775.800 744.600 777.600 749.700 ;
        RECT 793.500 749.400 798.600 750.600 ;
        RECT 793.500 744.600 795.300 749.400 ;
        RECT 812.400 747.600 813.600 757.950 ;
        RECT 827.100 756.150 828.900 757.950 ;
        RECT 833.100 756.150 834.900 757.950 ;
        RECT 836.700 750.600 837.600 757.950 ;
        RECT 851.100 756.150 852.900 757.950 ;
        RECT 857.100 756.150 858.900 757.950 ;
        RECT 860.700 750.600 861.600 757.950 ;
        RECT 878.100 756.150 879.900 757.950 ;
        RECT 880.950 753.750 882.150 757.950 ;
        RECT 884.100 756.150 885.900 757.950 ;
        RECT 899.100 756.150 900.900 757.950 ;
        RECT 878.400 752.700 882.150 753.750 ;
        RECT 902.850 753.750 904.050 757.950 ;
        RECT 905.100 756.150 906.900 757.950 ;
        RECT 902.850 752.700 906.600 753.750 ;
        RECT 878.400 750.600 879.600 752.700 ;
        RECT 811.800 744.600 813.600 747.600 ;
        RECT 832.500 749.400 837.600 750.600 ;
        RECT 856.500 749.400 861.600 750.600 ;
        RECT 832.500 744.600 834.300 749.400 ;
        RECT 856.500 744.600 858.300 749.400 ;
        RECT 877.800 744.600 879.600 750.600 ;
        RECT 880.800 749.700 888.600 751.050 ;
        RECT 880.800 744.600 882.600 749.700 ;
        RECT 886.800 744.600 888.600 749.700 ;
        RECT 896.400 749.700 904.200 751.050 ;
        RECT 896.400 744.600 898.200 749.700 ;
        RECT 902.400 744.600 904.200 749.700 ;
        RECT 905.400 750.600 906.600 752.700 ;
        RECT 905.400 744.600 907.200 750.600 ;
        RECT 14.400 733.200 16.200 740.400 ;
        RECT 37.500 735.600 39.300 740.400 ;
        RECT 37.500 734.400 42.600 735.600 ;
        RECT 14.400 732.300 18.600 733.200 ;
        RECT 14.100 727.050 15.900 728.850 ;
        RECT 17.400 727.050 18.600 732.300 ;
        RECT 20.100 727.050 21.900 728.850 ;
        RECT 32.100 727.050 33.900 728.850 ;
        RECT 38.100 727.050 39.900 728.850 ;
        RECT 41.700 727.050 42.600 734.400 ;
        RECT 56.400 735.300 58.200 740.400 ;
        RECT 62.400 735.300 64.200 740.400 ;
        RECT 56.400 733.950 64.200 735.300 ;
        RECT 65.400 734.400 67.200 740.400 ;
        RECT 65.400 732.300 66.600 734.400 ;
        RECT 62.850 731.250 66.600 732.300 ;
        RECT 87.000 732.000 88.800 740.400 ;
        RECT 106.200 732.000 108.000 740.400 ;
        RECT 130.200 732.000 132.000 740.400 ;
        RECT 151.500 735.600 153.300 740.400 ;
        RECT 173.400 737.400 175.200 740.400 ;
        RECT 151.500 734.400 156.600 735.600 ;
        RECT 59.100 727.050 60.900 728.850 ;
        RECT 62.850 727.050 64.050 731.250 ;
        RECT 87.000 730.800 90.300 732.000 ;
        RECT 65.100 727.050 66.900 728.850 ;
        RECT 80.100 727.050 81.900 728.850 ;
        RECT 86.100 727.050 87.900 728.850 ;
        RECT 89.400 727.050 90.300 730.800 ;
        RECT 104.700 730.800 108.000 732.000 ;
        RECT 128.700 730.800 132.000 732.000 ;
        RECT 104.700 727.050 105.600 730.800 ;
        RECT 107.100 727.050 108.900 728.850 ;
        RECT 113.100 727.050 114.900 728.850 ;
        RECT 128.700 727.050 129.600 730.800 ;
        RECT 131.100 727.050 132.900 728.850 ;
        RECT 137.100 727.050 138.900 728.850 ;
        RECT 146.100 727.050 147.900 728.850 ;
        RECT 152.100 727.050 153.900 728.850 ;
        RECT 155.700 727.050 156.600 734.400 ;
        RECT 173.400 727.050 174.600 737.400 ;
        RECT 188.400 733.200 190.200 740.400 ;
        RECT 210.300 736.200 212.100 740.400 ;
        RECT 209.400 734.400 212.100 736.200 ;
        RECT 188.400 732.300 192.600 733.200 ;
        RECT 188.100 727.050 189.900 728.850 ;
        RECT 191.400 727.050 192.600 732.300 ;
        RECT 194.100 727.050 195.900 728.850 ;
        RECT 209.400 727.050 210.300 734.400 ;
        RECT 212.100 732.600 213.900 733.500 ;
        RECT 217.800 732.600 219.600 740.400 ;
        RECT 212.100 731.700 219.600 732.600 ;
        RECT 233.400 734.400 235.200 740.400 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 19.950 724.950 22.050 727.050 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 37.950 724.950 40.050 727.050 ;
        RECT 40.950 724.950 43.050 727.050 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 58.950 724.950 61.050 727.050 ;
        RECT 61.950 724.950 64.050 727.050 ;
        RECT 64.950 724.950 67.050 727.050 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 130.950 724.950 133.050 727.050 ;
        RECT 133.950 724.950 136.050 727.050 ;
        RECT 136.950 724.950 139.050 727.050 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 154.950 724.950 157.050 727.050 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 187.950 724.950 190.050 727.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 208.950 724.950 211.050 727.050 ;
        RECT 211.950 724.950 214.050 727.050 ;
        RECT 17.400 711.600 18.600 724.950 ;
        RECT 35.100 723.150 36.900 724.950 ;
        RECT 41.700 717.600 42.600 724.950 ;
        RECT 56.100 723.150 57.900 724.950 ;
        RECT 16.800 705.600 18.600 711.600 ;
        RECT 32.400 716.700 40.200 717.600 ;
        RECT 32.400 705.600 34.200 716.700 ;
        RECT 38.400 705.600 40.200 716.700 ;
        RECT 41.400 705.600 43.200 717.600 ;
        RECT 61.950 711.600 63.150 724.950 ;
        RECT 83.100 723.150 84.900 724.950 ;
        RECT 89.400 712.800 90.300 724.950 ;
        RECT 83.700 711.900 90.300 712.800 ;
        RECT 83.700 711.600 85.200 711.900 ;
        RECT 61.800 705.600 63.600 711.600 ;
        RECT 83.400 705.600 85.200 711.600 ;
        RECT 89.400 711.600 90.300 711.900 ;
        RECT 104.700 712.800 105.600 724.950 ;
        RECT 110.100 723.150 111.900 724.950 ;
        RECT 128.700 712.800 129.600 724.950 ;
        RECT 134.100 723.150 135.900 724.950 ;
        RECT 149.100 723.150 150.900 724.950 ;
        RECT 136.950 720.450 139.050 721.050 ;
        RECT 151.950 720.450 154.050 721.050 ;
        RECT 136.950 719.550 154.050 720.450 ;
        RECT 136.950 718.950 139.050 719.550 ;
        RECT 151.950 718.950 154.050 719.550 ;
        RECT 155.700 717.600 156.600 724.950 ;
        RECT 170.100 723.150 171.900 724.950 ;
        RECT 146.400 716.700 154.200 717.600 ;
        RECT 104.700 711.900 111.300 712.800 ;
        RECT 104.700 711.600 105.600 711.900 ;
        RECT 89.400 705.600 91.200 711.600 ;
        RECT 103.800 705.600 105.600 711.600 ;
        RECT 109.800 711.600 111.300 711.900 ;
        RECT 128.700 711.900 135.300 712.800 ;
        RECT 128.700 711.600 129.600 711.900 ;
        RECT 109.800 705.600 111.600 711.600 ;
        RECT 127.800 705.600 129.600 711.600 ;
        RECT 133.800 711.600 135.300 711.900 ;
        RECT 133.800 705.600 135.600 711.600 ;
        RECT 146.400 705.600 148.200 716.700 ;
        RECT 152.400 705.600 154.200 716.700 ;
        RECT 155.400 705.600 157.200 717.600 ;
        RECT 173.400 711.600 174.600 724.950 ;
        RECT 191.400 711.600 192.600 724.950 ;
        RECT 209.400 717.600 210.300 724.950 ;
        RECT 212.100 723.150 213.900 724.950 ;
        RECT 173.400 705.600 175.200 711.600 ;
        RECT 190.800 705.600 192.600 711.600 ;
        RECT 208.800 705.600 210.600 717.600 ;
        RECT 215.700 711.600 216.600 731.700 ;
        RECT 218.100 727.050 219.900 728.850 ;
        RECT 230.100 727.050 231.900 728.850 ;
        RECT 233.400 727.050 234.600 734.400 ;
        RECT 250.800 733.200 252.600 740.400 ;
        RECT 270.300 736.200 272.100 740.400 ;
        RECT 248.400 732.300 252.600 733.200 ;
        RECT 269.400 734.400 272.100 736.200 ;
        RECT 245.100 727.050 246.900 728.850 ;
        RECT 248.400 727.050 249.600 732.300 ;
        RECT 251.100 727.050 252.900 728.850 ;
        RECT 269.400 727.050 270.300 734.400 ;
        RECT 272.100 732.600 273.900 733.500 ;
        RECT 277.800 732.600 279.600 740.400 ;
        RECT 295.800 733.200 297.600 740.400 ;
        RECT 310.800 737.400 312.600 740.400 ;
        RECT 272.100 731.700 279.600 732.600 ;
        RECT 293.400 732.300 297.600 733.200 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 229.950 724.950 232.050 727.050 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 247.950 724.950 250.050 727.050 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 268.950 724.950 271.050 727.050 ;
        RECT 271.950 724.950 274.050 727.050 ;
        RECT 214.800 705.600 216.600 711.600 ;
        RECT 233.400 717.600 234.600 724.950 ;
        RECT 233.400 705.600 235.200 717.600 ;
        RECT 248.400 711.600 249.600 724.950 ;
        RECT 269.400 717.600 270.300 724.950 ;
        RECT 272.100 723.150 273.900 724.950 ;
        RECT 248.400 705.600 250.200 711.600 ;
        RECT 268.800 705.600 270.600 717.600 ;
        RECT 275.700 711.600 276.600 731.700 ;
        RECT 278.100 727.050 279.900 728.850 ;
        RECT 290.100 727.050 291.900 728.850 ;
        RECT 293.400 727.050 294.600 732.300 ;
        RECT 296.100 727.050 297.900 728.850 ;
        RECT 311.400 727.050 312.600 737.400 ;
        RECT 329.400 733.200 331.200 740.400 ;
        RECT 349.800 734.400 351.600 740.400 ;
        RECT 313.950 732.450 316.050 733.050 ;
        RECT 319.950 732.450 322.050 733.050 ;
        RECT 313.950 731.550 322.050 732.450 ;
        RECT 329.400 732.300 333.600 733.200 ;
        RECT 313.950 730.950 316.050 731.550 ;
        RECT 319.950 730.950 322.050 731.550 ;
        RECT 329.100 727.050 330.900 728.850 ;
        RECT 332.400 727.050 333.600 732.300 ;
        RECT 350.400 732.300 351.600 734.400 ;
        RECT 352.800 735.300 354.600 740.400 ;
        RECT 358.800 735.300 360.600 740.400 ;
        RECT 352.800 733.950 360.600 735.300 ;
        RECT 371.400 734.400 373.200 740.400 ;
        RECT 378.600 735.000 380.400 740.400 ;
        RECT 371.400 733.500 372.900 734.400 ;
        RECT 350.400 731.250 354.150 732.300 ;
        RECT 371.400 732.000 375.750 733.500 ;
        RECT 373.650 731.400 375.750 732.000 ;
        RECT 379.350 732.900 380.400 735.000 ;
        RECT 386.400 734.400 388.200 740.400 ;
        RECT 383.700 733.200 388.200 734.400 ;
        RECT 406.800 733.200 408.600 740.400 ;
        RECT 335.100 727.050 336.900 728.850 ;
        RECT 350.100 727.050 351.900 728.850 ;
        RECT 352.950 727.050 354.150 731.250 ;
        RECT 376.650 729.900 378.450 731.700 ;
        RECT 379.350 730.800 382.500 732.900 ;
        RECT 383.700 731.100 385.800 733.200 ;
        RECT 391.950 732.450 394.050 732.900 ;
        RECT 400.950 732.450 403.050 733.050 ;
        RECT 391.950 731.550 403.050 732.450 ;
        RECT 391.950 730.800 394.050 731.550 ;
        RECT 400.950 730.950 403.050 731.550 ;
        RECT 404.400 732.300 408.600 733.200 ;
        RECT 376.200 729.000 378.300 729.900 ;
        RECT 356.100 727.050 357.900 728.850 ;
        RECT 371.700 727.800 378.300 729.000 ;
        RECT 371.700 727.200 373.500 727.800 ;
        RECT 277.950 724.950 280.050 727.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 292.950 724.950 295.050 727.050 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 310.950 724.950 313.050 727.050 ;
        RECT 313.950 724.950 316.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 331.950 724.950 334.050 727.050 ;
        RECT 334.950 724.950 337.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 371.400 725.100 373.500 727.200 ;
        RECT 274.800 705.600 276.600 711.600 ;
        RECT 293.400 711.600 294.600 724.950 ;
        RECT 311.400 711.600 312.600 724.950 ;
        RECT 314.100 723.150 315.900 724.950 ;
        RECT 332.400 711.600 333.600 724.950 ;
        RECT 340.950 720.450 343.050 721.050 ;
        RECT 349.950 720.450 352.050 721.050 ;
        RECT 340.950 719.550 352.050 720.450 ;
        RECT 340.950 718.950 343.050 719.550 ;
        RECT 349.950 718.950 352.050 719.550 ;
        RECT 353.850 711.600 355.050 724.950 ;
        RECT 359.100 723.150 360.900 724.950 ;
        RECT 376.200 724.800 378.300 726.900 ;
        RECT 376.200 723.000 378.000 724.800 ;
        RECT 379.350 724.200 380.250 730.800 ;
        RECT 381.150 726.900 383.250 729.000 ;
        RECT 381.300 725.100 383.100 726.900 ;
        RECT 385.950 725.100 388.050 727.200 ;
        RECT 401.100 727.050 402.900 728.850 ;
        RECT 404.400 727.050 405.600 732.300 ;
        RECT 427.200 732.000 429.000 740.400 ;
        RECT 425.700 730.800 429.000 732.000 ;
        RECT 453.000 732.000 454.800 740.400 ;
        RECT 475.800 733.200 477.600 740.400 ;
        RECT 493.800 737.400 495.600 740.400 ;
        RECT 473.400 732.300 477.600 733.200 ;
        RECT 453.000 730.800 456.300 732.000 ;
        RECT 409.950 729.450 414.000 730.050 ;
        RECT 420.000 729.450 424.050 730.050 ;
        RECT 407.100 727.050 408.900 728.850 ;
        RECT 409.950 727.950 414.450 729.450 ;
        RECT 379.350 722.700 382.500 724.200 ;
        RECT 386.100 723.450 387.900 725.100 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 403.950 724.950 406.050 727.050 ;
        RECT 406.950 724.950 409.050 727.050 ;
        RECT 391.950 723.450 394.050 724.050 ;
        RECT 386.100 723.300 394.050 723.450 ;
        RECT 380.400 722.100 382.500 722.700 ;
        RECT 386.550 722.550 394.050 723.300 ;
        RECT 377.700 719.700 379.500 721.800 ;
        RECT 374.100 718.800 379.500 719.700 ;
        RECT 374.100 717.900 376.200 718.800 ;
        RECT 371.400 716.700 376.200 717.900 ;
        RECT 381.000 717.600 382.200 722.100 ;
        RECT 391.950 721.950 394.050 722.550 ;
        RECT 378.900 716.700 382.200 717.600 ;
        RECT 383.100 717.600 385.200 718.500 ;
        RECT 293.400 705.600 295.200 711.600 ;
        RECT 310.800 705.600 312.600 711.600 ;
        RECT 331.800 705.600 333.600 711.600 ;
        RECT 353.400 705.600 355.200 711.600 ;
        RECT 371.400 705.600 373.200 716.700 ;
        RECT 378.900 705.600 380.700 716.700 ;
        RECT 383.100 716.400 388.200 717.600 ;
        RECT 386.400 705.600 388.200 716.400 ;
        RECT 404.400 711.600 405.600 724.950 ;
        RECT 413.550 724.050 414.450 727.950 ;
        RECT 409.950 722.550 414.450 724.050 ;
        RECT 419.550 727.950 424.050 729.450 ;
        RECT 409.950 721.950 414.000 722.550 ;
        RECT 419.550 720.900 420.450 727.950 ;
        RECT 425.700 727.050 426.600 730.800 ;
        RECT 428.100 727.050 429.900 728.850 ;
        RECT 434.100 727.050 435.900 728.850 ;
        RECT 446.100 727.050 447.900 728.850 ;
        RECT 452.100 727.050 453.900 728.850 ;
        RECT 455.400 727.050 456.300 730.800 ;
        RECT 457.950 729.450 460.050 730.050 ;
        RECT 457.950 728.550 465.450 729.450 ;
        RECT 457.950 727.950 460.050 728.550 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 427.950 724.950 430.050 727.050 ;
        RECT 430.950 724.950 433.050 727.050 ;
        RECT 433.950 724.950 436.050 727.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 451.950 724.950 454.050 727.050 ;
        RECT 454.950 724.950 457.050 727.050 ;
        RECT 418.950 718.800 421.050 720.900 ;
        RECT 425.700 712.800 426.600 724.950 ;
        RECT 431.100 723.150 432.900 724.950 ;
        RECT 449.100 723.150 450.900 724.950 ;
        RECT 455.400 712.800 456.300 724.950 ;
        RECT 464.550 723.450 465.450 728.550 ;
        RECT 470.100 727.050 471.900 728.850 ;
        RECT 473.400 727.050 474.600 732.300 ;
        RECT 476.100 727.050 477.900 728.850 ;
        RECT 494.400 727.050 495.600 737.400 ;
        RECT 509.400 735.300 511.200 740.400 ;
        RECT 515.400 735.300 517.200 740.400 ;
        RECT 509.400 733.950 517.200 735.300 ;
        RECT 518.400 734.400 520.200 740.400 ;
        RECT 518.400 732.300 519.600 734.400 ;
        RECT 535.800 733.200 537.600 740.400 ;
        RECT 515.850 731.250 519.600 732.300 ;
        RECT 533.400 732.300 537.600 733.200 ;
        RECT 554.400 733.200 556.200 740.400 ;
        RECT 569.400 735.300 571.200 740.400 ;
        RECT 575.400 735.300 577.200 740.400 ;
        RECT 569.400 733.950 577.200 735.300 ;
        RECT 578.400 734.400 580.200 740.400 ;
        RECT 595.800 734.400 597.600 740.400 ;
        RECT 554.400 732.300 558.600 733.200 ;
        RECT 578.400 732.300 579.600 734.400 ;
        RECT 504.000 729.450 508.050 730.050 ;
        RECT 503.550 727.950 508.050 729.450 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 475.950 724.950 478.050 727.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 464.550 722.550 468.450 723.450 ;
        RECT 467.550 721.050 468.450 722.550 ;
        RECT 467.550 719.550 472.050 721.050 ;
        RECT 468.000 718.950 472.050 719.550 ;
        RECT 425.700 711.900 432.300 712.800 ;
        RECT 425.700 711.600 426.600 711.900 ;
        RECT 404.400 705.600 406.200 711.600 ;
        RECT 424.800 705.600 426.600 711.600 ;
        RECT 430.800 711.600 432.300 711.900 ;
        RECT 449.700 711.900 456.300 712.800 ;
        RECT 449.700 711.600 451.200 711.900 ;
        RECT 430.800 705.600 432.600 711.600 ;
        RECT 449.400 705.600 451.200 711.600 ;
        RECT 455.400 711.600 456.300 711.900 ;
        RECT 473.400 711.600 474.600 724.950 ;
        RECT 494.400 711.600 495.600 724.950 ;
        RECT 497.100 723.150 498.900 724.950 ;
        RECT 496.950 720.450 499.050 721.050 ;
        RECT 503.550 720.450 504.450 727.950 ;
        RECT 512.100 727.050 513.900 728.850 ;
        RECT 515.850 727.050 517.050 731.250 ;
        RECT 518.100 727.050 519.900 728.850 ;
        RECT 530.100 727.050 531.900 728.850 ;
        RECT 533.400 727.050 534.600 732.300 ;
        RECT 538.950 729.450 543.000 730.050 ;
        RECT 536.100 727.050 537.900 728.850 ;
        RECT 538.950 727.950 543.450 729.450 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 509.100 723.150 510.900 724.950 ;
        RECT 496.950 719.550 504.450 720.450 ;
        RECT 496.950 718.950 499.050 719.550 ;
        RECT 514.950 711.600 516.150 724.950 ;
        RECT 533.400 711.600 534.600 724.950 ;
        RECT 542.550 724.050 543.450 727.950 ;
        RECT 554.100 727.050 555.900 728.850 ;
        RECT 557.400 727.050 558.600 732.300 ;
        RECT 575.850 731.250 579.600 732.300 ;
        RECT 596.400 732.300 597.600 734.400 ;
        RECT 598.800 735.300 600.600 740.400 ;
        RECT 604.800 735.300 606.600 740.400 ;
        RECT 598.800 733.950 606.600 735.300 ;
        RECT 622.500 735.600 624.300 740.400 ;
        RECT 622.500 734.400 627.600 735.600 ;
        RECT 596.400 731.250 600.150 732.300 ;
        RECT 560.100 727.050 561.900 728.850 ;
        RECT 572.100 727.050 573.900 728.850 ;
        RECT 575.850 727.050 577.050 731.250 ;
        RECT 578.100 727.050 579.900 728.850 ;
        RECT 596.100 727.050 597.900 728.850 ;
        RECT 598.950 727.050 600.150 731.250 ;
        RECT 602.100 727.050 603.900 728.850 ;
        RECT 617.100 727.050 618.900 728.850 ;
        RECT 623.100 727.050 624.900 728.850 ;
        RECT 626.700 727.050 627.600 734.400 ;
        RECT 646.800 733.200 648.600 740.400 ;
        RECT 663.300 736.200 665.100 740.400 ;
        RECT 644.400 732.300 648.600 733.200 ;
        RECT 662.400 734.400 665.100 736.200 ;
        RECT 641.100 727.050 642.900 728.850 ;
        RECT 644.400 727.050 645.600 732.300 ;
        RECT 649.950 729.450 654.000 730.050 ;
        RECT 647.100 727.050 648.900 728.850 ;
        RECT 649.950 727.950 654.450 729.450 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 568.950 724.950 571.050 727.050 ;
        RECT 571.950 724.950 574.050 727.050 ;
        RECT 574.950 724.950 577.050 727.050 ;
        RECT 577.950 724.950 580.050 727.050 ;
        RECT 595.950 724.950 598.050 727.050 ;
        RECT 598.950 724.950 601.050 727.050 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 616.950 724.950 619.050 727.050 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 622.950 724.950 625.050 727.050 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 646.950 724.950 649.050 727.050 ;
        RECT 538.950 722.550 543.450 724.050 ;
        RECT 538.950 721.950 543.000 722.550 ;
        RECT 557.400 711.600 558.600 724.950 ;
        RECT 569.100 723.150 570.900 724.950 ;
        RECT 574.950 711.600 576.150 724.950 ;
        RECT 599.850 711.600 601.050 724.950 ;
        RECT 605.100 723.150 606.900 724.950 ;
        RECT 620.100 723.150 621.900 724.950 ;
        RECT 626.700 717.600 627.600 724.950 ;
        RECT 617.400 716.700 625.200 717.600 ;
        RECT 455.400 705.600 457.200 711.600 ;
        RECT 473.400 705.600 475.200 711.600 ;
        RECT 493.800 705.600 495.600 711.600 ;
        RECT 514.800 705.600 516.600 711.600 ;
        RECT 533.400 705.600 535.200 711.600 ;
        RECT 556.800 705.600 558.600 711.600 ;
        RECT 574.800 705.600 576.600 711.600 ;
        RECT 599.400 705.600 601.200 711.600 ;
        RECT 617.400 705.600 619.200 716.700 ;
        RECT 623.400 705.600 625.200 716.700 ;
        RECT 626.400 705.600 628.200 717.600 ;
        RECT 644.400 711.600 645.600 724.950 ;
        RECT 653.550 724.050 654.450 727.950 ;
        RECT 662.400 727.050 663.300 734.400 ;
        RECT 665.100 732.600 666.900 733.500 ;
        RECT 670.800 732.600 672.600 740.400 ;
        RECT 683.400 735.300 685.200 740.400 ;
        RECT 689.400 735.300 691.200 740.400 ;
        RECT 683.400 733.950 691.200 735.300 ;
        RECT 692.400 734.400 694.200 740.400 ;
        RECT 706.800 739.500 714.600 740.400 ;
        RECT 706.800 734.400 708.600 739.500 ;
        RECT 709.800 734.400 711.600 738.600 ;
        RECT 712.800 735.000 714.600 739.500 ;
        RECT 718.800 735.000 720.600 740.400 ;
        RECT 665.100 731.700 672.600 732.600 ;
        RECT 692.400 732.300 693.600 734.400 ;
        RECT 661.950 724.950 664.050 727.050 ;
        RECT 664.950 724.950 667.050 727.050 ;
        RECT 649.950 722.550 654.450 724.050 ;
        RECT 649.950 721.950 654.000 722.550 ;
        RECT 662.400 717.600 663.300 724.950 ;
        RECT 665.100 723.150 666.900 724.950 ;
        RECT 644.400 705.600 646.200 711.600 ;
        RECT 661.800 705.600 663.600 717.600 ;
        RECT 668.700 711.600 669.600 731.700 ;
        RECT 689.850 731.250 693.600 732.300 ;
        RECT 694.950 732.450 697.050 733.050 ;
        RECT 703.950 732.450 706.050 733.050 ;
        RECT 694.950 731.550 706.050 732.450 ;
        RECT 710.400 732.900 711.300 734.400 ;
        RECT 712.800 734.100 720.600 735.000 ;
        RECT 734.400 737.400 736.200 740.400 ;
        RECT 710.400 731.700 715.050 732.900 ;
        RECT 678.000 729.450 682.050 730.050 ;
        RECT 671.100 727.050 672.900 728.850 ;
        RECT 677.550 727.950 682.050 729.450 ;
        RECT 670.950 724.950 673.050 727.050 ;
        RECT 677.550 724.050 678.450 727.950 ;
        RECT 686.100 727.050 687.900 728.850 ;
        RECT 689.850 727.050 691.050 731.250 ;
        RECT 694.950 730.950 697.050 731.550 ;
        RECT 703.950 730.950 706.050 731.550 ;
        RECT 692.100 727.050 693.900 728.850 ;
        RECT 710.100 727.050 711.900 728.850 ;
        RECT 713.700 727.050 715.050 731.700 ;
        RECT 721.950 729.450 726.000 730.050 ;
        RECT 716.100 727.050 717.900 728.850 ;
        RECT 721.950 727.950 726.450 729.450 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 685.950 724.950 688.050 727.050 ;
        RECT 688.950 724.950 691.050 727.050 ;
        RECT 691.950 724.950 694.050 727.050 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 709.950 724.950 712.050 727.050 ;
        RECT 712.950 724.950 715.050 727.050 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 673.950 722.550 678.450 724.050 ;
        RECT 683.100 723.150 684.900 724.950 ;
        RECT 673.950 721.950 678.000 722.550 ;
        RECT 670.950 714.450 673.050 715.050 ;
        RECT 676.950 714.450 679.050 715.050 ;
        RECT 670.950 713.550 679.050 714.450 ;
        RECT 670.950 712.950 673.050 713.550 ;
        RECT 676.950 712.950 679.050 713.550 ;
        RECT 688.950 711.600 690.150 724.950 ;
        RECT 707.100 723.150 708.900 724.950 ;
        RECT 713.700 717.600 714.900 724.950 ;
        RECT 719.100 723.150 720.900 724.950 ;
        RECT 725.550 724.050 726.450 727.950 ;
        RECT 734.400 727.050 735.600 737.400 ;
        RECT 749.400 735.300 751.200 740.400 ;
        RECT 755.400 735.300 757.200 740.400 ;
        RECT 749.400 733.950 757.200 735.300 ;
        RECT 758.400 734.400 760.200 740.400 ;
        RECT 775.800 734.400 777.600 740.400 ;
        RECT 758.400 732.300 759.600 734.400 ;
        RECT 755.850 731.250 759.600 732.300 ;
        RECT 776.400 732.300 777.600 734.400 ;
        RECT 778.800 735.300 780.600 740.400 ;
        RECT 784.800 735.300 786.600 740.400 ;
        RECT 778.800 733.950 786.600 735.300 ;
        RECT 802.500 735.600 804.300 740.400 ;
        RECT 802.500 734.400 807.600 735.600 ;
        RECT 799.950 732.450 802.050 733.050 ;
        RECT 776.400 731.250 780.150 732.300 ;
        RECT 736.950 729.450 739.050 730.050 ;
        RECT 736.950 728.550 744.450 729.450 ;
        RECT 736.950 727.950 739.050 728.550 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 733.950 724.950 736.050 727.050 ;
        RECT 721.950 722.550 726.450 724.050 ;
        RECT 731.100 723.150 732.900 724.950 ;
        RECT 721.950 721.950 726.000 722.550 ;
        RECT 667.800 705.600 669.600 711.600 ;
        RECT 688.800 705.600 690.600 711.600 ;
        RECT 712.800 705.600 716.100 717.600 ;
        RECT 734.400 711.600 735.600 724.950 ;
        RECT 743.550 724.050 744.450 728.550 ;
        RECT 752.100 727.050 753.900 728.850 ;
        RECT 755.850 727.050 757.050 731.250 ;
        RECT 771.000 729.450 775.050 730.050 ;
        RECT 758.100 727.050 759.900 728.850 ;
        RECT 770.550 727.950 775.050 729.450 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 754.950 724.950 757.050 727.050 ;
        RECT 757.950 724.950 760.050 727.050 ;
        RECT 743.550 722.550 748.050 724.050 ;
        RECT 749.100 723.150 750.900 724.950 ;
        RECT 744.000 721.950 748.050 722.550 ;
        RECT 754.950 711.600 756.150 724.950 ;
        RECT 770.550 724.050 771.450 727.950 ;
        RECT 776.100 727.050 777.900 728.850 ;
        RECT 778.950 727.050 780.150 731.250 ;
        RECT 791.550 731.550 802.050 732.450 ;
        RECT 782.100 727.050 783.900 728.850 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 781.950 724.950 784.050 727.050 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 770.550 722.550 775.050 724.050 ;
        RECT 771.000 721.950 775.050 722.550 ;
        RECT 757.950 720.450 760.050 721.050 ;
        RECT 766.950 720.450 769.050 721.050 ;
        RECT 757.950 719.550 769.050 720.450 ;
        RECT 757.950 718.950 760.050 719.550 ;
        RECT 766.950 718.950 769.050 719.550 ;
        RECT 779.850 711.600 781.050 724.950 ;
        RECT 785.100 723.150 786.900 724.950 ;
        RECT 791.550 724.050 792.450 731.550 ;
        RECT 799.950 730.950 802.050 731.550 ;
        RECT 797.100 727.050 798.900 728.850 ;
        RECT 803.100 727.050 804.900 728.850 ;
        RECT 806.700 727.050 807.600 734.400 ;
        RECT 821.400 735.300 823.200 740.400 ;
        RECT 827.400 735.300 829.200 740.400 ;
        RECT 821.400 733.950 829.200 735.300 ;
        RECT 830.400 734.400 832.200 740.400 ;
        RECT 842.400 735.300 844.200 740.400 ;
        RECT 848.400 735.300 850.200 740.400 ;
        RECT 830.400 732.300 831.600 734.400 ;
        RECT 842.400 733.950 850.200 735.300 ;
        RECT 851.400 734.400 853.200 740.400 ;
        RECT 856.950 738.450 859.050 739.050 ;
        RECT 862.950 738.450 865.050 739.050 ;
        RECT 856.950 737.550 865.050 738.450 ;
        RECT 856.950 736.950 859.050 737.550 ;
        RECT 862.950 736.950 865.050 737.550 ;
        RECT 866.400 735.300 868.200 740.400 ;
        RECT 872.400 735.300 874.200 740.400 ;
        RECT 851.400 732.300 852.600 734.400 ;
        RECT 866.400 733.950 874.200 735.300 ;
        RECT 875.400 734.400 877.200 740.400 ;
        RECT 890.400 734.400 892.200 740.400 ;
        RECT 897.900 734.400 899.700 740.400 ;
        RECT 905.400 734.400 907.200 740.400 ;
        RECT 875.400 732.300 876.600 734.400 ;
        RECT 827.850 731.250 831.600 732.300 ;
        RECT 848.850 731.250 852.600 732.300 ;
        RECT 872.850 731.250 876.600 732.300 ;
        RECT 891.000 732.600 892.200 734.400 ;
        RECT 898.200 732.900 899.400 734.400 ;
        RECT 902.400 733.500 907.200 734.400 ;
        RECT 891.000 731.700 897.300 732.600 ;
        RECT 816.000 729.450 820.050 730.050 ;
        RECT 815.550 727.950 820.050 729.450 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 805.950 724.950 808.050 727.050 ;
        RECT 787.950 722.550 792.450 724.050 ;
        RECT 800.100 723.150 801.900 724.950 ;
        RECT 787.950 721.950 792.000 722.550 ;
        RECT 806.700 717.600 807.600 724.950 ;
        RECT 815.550 724.050 816.450 727.950 ;
        RECT 824.100 727.050 825.900 728.850 ;
        RECT 827.850 727.050 829.050 731.250 ;
        RECT 830.100 727.050 831.900 728.850 ;
        RECT 845.100 727.050 846.900 728.850 ;
        RECT 848.850 727.050 850.050 731.250 ;
        RECT 851.100 727.050 852.900 728.850 ;
        RECT 869.100 727.050 870.900 728.850 ;
        RECT 872.850 727.050 874.050 731.250 ;
        RECT 877.950 729.450 880.050 730.050 ;
        RECT 895.200 729.600 897.300 731.700 ;
        RECT 877.950 728.850 891.450 729.450 ;
        RECT 875.100 727.050 876.900 728.850 ;
        RECT 877.950 728.550 892.200 728.850 ;
        RECT 877.950 727.950 880.050 728.550 ;
        RECT 890.400 727.050 892.200 728.550 ;
        RECT 895.500 727.800 897.300 729.600 ;
        RECT 898.200 730.800 901.200 732.900 ;
        RECT 902.400 732.300 904.500 733.500 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 829.950 724.950 832.050 727.050 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 890.400 726.300 892.500 727.050 ;
        RECT 890.400 725.100 897.300 726.300 ;
        RECT 890.400 724.950 892.500 725.100 ;
        RECT 815.550 722.550 820.050 724.050 ;
        RECT 821.100 723.150 822.900 724.950 ;
        RECT 816.000 721.950 820.050 722.550 ;
        RECT 797.400 716.700 805.200 717.600 ;
        RECT 734.400 705.600 736.200 711.600 ;
        RECT 754.800 705.600 756.600 711.600 ;
        RECT 779.400 705.600 781.200 711.600 ;
        RECT 797.400 705.600 799.200 716.700 ;
        RECT 803.400 705.600 805.200 716.700 ;
        RECT 806.400 705.600 808.200 717.600 ;
        RECT 826.950 711.600 828.150 724.950 ;
        RECT 842.100 723.150 843.900 724.950 ;
        RECT 847.950 711.600 849.150 724.950 ;
        RECT 866.100 723.150 867.900 724.950 ;
        RECT 850.950 720.450 853.050 721.050 ;
        RECT 862.950 720.450 865.050 721.050 ;
        RECT 850.950 719.550 865.050 720.450 ;
        RECT 850.950 718.950 853.050 719.550 ;
        RECT 862.950 718.950 865.050 719.550 ;
        RECT 871.950 711.600 873.150 724.950 ;
        RECT 895.500 724.500 897.300 725.100 ;
        RECT 898.200 725.100 899.250 730.800 ;
        RECT 900.150 727.800 902.250 729.900 ;
        RECT 900.600 726.000 902.400 727.800 ;
        RECT 904.950 726.450 907.050 727.050 ;
        RECT 909.000 726.450 913.050 727.050 ;
        RECT 904.950 725.550 913.050 726.450 ;
        RECT 898.200 724.200 900.600 725.100 ;
        RECT 904.950 724.950 907.050 725.550 ;
        RECT 909.000 724.950 913.050 725.550 ;
        RECT 894.300 721.500 898.200 723.300 ;
        RECT 896.100 721.200 898.200 721.500 ;
        RECT 899.100 722.100 901.200 724.200 ;
        RECT 905.100 723.150 906.900 724.950 ;
        RECT 899.100 720.000 900.000 722.100 ;
        RECT 892.800 717.600 894.900 719.700 ;
        RECT 898.500 719.100 900.000 720.000 ;
        RECT 898.500 717.600 899.700 719.100 ;
        RECT 890.400 716.700 894.900 717.600 ;
        RECT 826.800 705.600 828.600 711.600 ;
        RECT 847.800 705.600 849.600 711.600 ;
        RECT 871.800 705.600 873.600 711.600 ;
        RECT 890.400 705.600 892.200 716.700 ;
        RECT 897.900 709.050 899.700 717.600 ;
        RECT 902.400 717.600 904.500 718.500 ;
        RECT 902.400 716.400 907.200 717.600 ;
        RECT 897.900 706.950 901.050 709.050 ;
        RECT 897.900 705.600 899.700 706.950 ;
        RECT 905.400 705.600 907.200 716.400 ;
        RECT 13.800 695.400 15.600 701.400 ;
        RECT 32.400 695.400 34.200 701.400 ;
        RECT 14.400 682.050 15.600 695.400 ;
        RECT 32.700 695.100 34.200 695.400 ;
        RECT 38.400 695.400 40.200 701.400 ;
        RECT 38.400 695.100 39.300 695.400 ;
        RECT 32.700 694.200 39.300 695.100 ;
        RECT 32.100 682.050 33.900 683.850 ;
        RECT 38.400 682.050 39.300 694.200 ;
        RECT 55.800 689.400 57.600 701.400 ;
        RECT 58.800 690.300 60.600 701.400 ;
        RECT 64.800 690.300 66.600 701.400 ;
        RECT 80.400 695.400 82.200 701.400 ;
        RECT 80.700 695.100 82.200 695.400 ;
        RECT 86.400 695.400 88.200 701.400 ;
        RECT 86.400 695.100 87.300 695.400 ;
        RECT 80.700 694.200 87.300 695.100 ;
        RECT 58.800 689.400 66.600 690.300 ;
        RECT 56.400 682.050 57.300 689.400 ;
        RECT 58.950 687.450 61.050 688.200 ;
        RECT 70.950 687.450 73.050 688.050 ;
        RECT 58.950 686.550 73.050 687.450 ;
        RECT 58.950 686.100 61.050 686.550 ;
        RECT 70.950 685.950 73.050 686.550 ;
        RECT 62.100 682.050 63.900 683.850 ;
        RECT 80.100 682.050 81.900 683.850 ;
        RECT 86.400 682.050 87.300 694.200 ;
        RECT 101.400 690.300 103.200 701.400 ;
        RECT 107.400 690.300 109.200 701.400 ;
        RECT 101.400 689.400 109.200 690.300 ;
        RECT 110.400 689.400 112.200 701.400 ;
        RECT 125.400 690.300 127.200 701.400 ;
        RECT 125.400 689.400 129.900 690.300 ;
        RECT 132.900 689.400 134.700 701.400 ;
        RECT 140.400 690.600 142.200 701.400 ;
        RECT 104.100 682.050 105.900 683.850 ;
        RECT 110.700 682.050 111.600 689.400 ;
        RECT 127.800 687.300 129.900 689.400 ;
        RECT 133.500 687.900 134.700 689.400 ;
        RECT 137.400 689.400 142.200 690.600 ;
        RECT 158.700 690.600 160.500 701.400 ;
        RECT 158.700 689.400 162.300 690.600 ;
        RECT 184.800 689.400 188.100 701.400 ;
        RECT 206.400 695.400 208.200 701.400 ;
        RECT 223.800 695.400 225.600 701.400 ;
        RECT 137.400 688.500 139.500 689.400 ;
        RECT 133.500 687.000 135.000 687.900 ;
        RECT 131.100 685.500 133.200 685.800 ;
        RECT 129.300 683.700 133.200 685.500 ;
        RECT 134.100 684.900 135.000 687.000 ;
        RECT 134.100 682.800 136.200 684.900 ;
        RECT 10.950 679.950 13.050 682.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 28.950 679.950 31.050 682.050 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 58.950 679.950 61.050 682.050 ;
        RECT 61.950 679.950 64.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 76.950 679.950 79.050 682.050 ;
        RECT 79.950 679.950 82.050 682.050 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 85.950 679.950 88.050 682.050 ;
        RECT 11.100 678.150 12.900 679.950 ;
        RECT 14.400 674.700 15.600 679.950 ;
        RECT 17.100 678.150 18.900 679.950 ;
        RECT 29.100 678.150 30.900 679.950 ;
        RECT 35.100 678.150 36.900 679.950 ;
        RECT 38.400 676.200 39.300 679.950 ;
        RECT 11.400 673.800 15.600 674.700 ;
        RECT 36.000 675.000 39.300 676.200 ;
        RECT 11.400 666.600 13.200 673.800 ;
        RECT 36.000 666.600 37.800 675.000 ;
        RECT 56.400 672.600 57.300 679.950 ;
        RECT 59.100 678.150 60.900 679.950 ;
        RECT 65.100 678.150 66.900 679.950 ;
        RECT 77.100 678.150 78.900 679.950 ;
        RECT 83.100 678.150 84.900 679.950 ;
        RECT 86.400 676.200 87.300 679.950 ;
        RECT 91.950 678.450 94.050 682.050 ;
        RECT 100.950 679.950 103.050 682.050 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 125.400 681.900 127.500 682.050 ;
        RECT 130.500 681.900 132.300 682.500 ;
        RECT 125.400 680.700 132.300 681.900 ;
        RECT 133.200 681.900 135.600 682.800 ;
        RECT 140.100 682.050 141.900 683.850 ;
        RECT 158.100 682.050 159.900 683.850 ;
        RECT 161.400 682.050 162.300 689.400 ;
        RECT 164.100 682.050 165.900 683.850 ;
        RECT 179.100 682.050 180.900 683.850 ;
        RECT 185.700 682.050 186.900 689.400 ;
        RECT 193.950 684.450 198.000 685.050 ;
        RECT 191.100 682.050 192.900 683.850 ;
        RECT 193.950 682.950 198.450 684.450 ;
        RECT 125.400 679.950 127.500 680.700 ;
        RECT 97.950 678.450 100.050 679.050 ;
        RECT 91.950 678.000 100.050 678.450 ;
        RECT 101.100 678.150 102.900 679.950 ;
        RECT 107.100 678.150 108.900 679.950 ;
        RECT 92.550 677.550 100.050 678.000 ;
        RECT 97.950 676.950 100.050 677.550 ;
        RECT 84.000 675.000 87.300 676.200 ;
        RECT 56.400 671.400 61.500 672.600 ;
        RECT 59.700 666.600 61.500 671.400 ;
        RECT 84.000 666.600 85.800 675.000 ;
        RECT 110.700 672.600 111.600 679.950 ;
        RECT 125.400 679.050 127.200 679.950 ;
        RECT 121.950 678.150 127.200 679.050 ;
        RECT 121.950 677.550 126.450 678.150 ;
        RECT 121.950 676.950 126.000 677.550 ;
        RECT 130.500 677.400 132.300 679.200 ;
        RECT 130.200 675.300 132.300 677.400 ;
        RECT 126.000 674.400 132.300 675.300 ;
        RECT 133.200 676.200 134.250 681.900 ;
        RECT 139.950 681.450 142.050 682.050 ;
        RECT 148.950 681.450 151.050 682.050 ;
        RECT 135.600 679.200 137.400 681.000 ;
        RECT 139.950 680.550 151.050 681.450 ;
        RECT 139.950 679.950 142.050 680.550 ;
        RECT 148.950 679.950 151.050 680.550 ;
        RECT 157.950 679.950 160.050 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 187.950 679.950 190.050 682.050 ;
        RECT 190.950 679.950 193.050 682.050 ;
        RECT 135.150 677.100 137.250 679.200 ;
        RECT 126.000 672.600 127.200 674.400 ;
        RECT 133.200 674.100 136.200 676.200 ;
        RECT 133.200 672.600 134.400 674.100 ;
        RECT 137.400 673.500 139.500 674.700 ;
        RECT 137.400 672.600 142.200 673.500 ;
        RECT 106.500 671.400 111.600 672.600 ;
        RECT 106.500 666.600 108.300 671.400 ;
        RECT 125.400 666.600 127.200 672.600 ;
        RECT 132.900 666.600 134.700 672.600 ;
        RECT 140.400 666.600 142.200 672.600 ;
        RECT 161.400 669.600 162.300 679.950 ;
        RECT 182.100 678.150 183.900 679.950 ;
        RECT 185.700 675.300 187.050 679.950 ;
        RECT 188.100 678.150 189.900 679.950 ;
        RECT 197.550 679.050 198.450 682.950 ;
        RECT 206.400 682.050 207.600 695.400 ;
        RECT 224.700 695.100 225.600 695.400 ;
        RECT 229.800 695.400 231.600 701.400 ;
        RECT 229.800 695.100 231.300 695.400 ;
        RECT 224.700 694.200 231.300 695.100 ;
        RECT 224.700 682.050 225.600 694.200 ;
        RECT 247.800 689.400 249.600 701.400 ;
        RECT 250.800 690.300 252.600 701.400 ;
        RECT 256.800 690.300 258.600 701.400 ;
        RECT 272.400 695.400 274.200 701.400 ;
        RECT 295.800 695.400 297.600 701.400 ;
        RECT 317.400 695.400 319.200 701.400 ;
        RECT 250.800 689.400 258.600 690.300 ;
        RECT 230.100 682.050 231.900 683.850 ;
        RECT 248.400 682.050 249.300 689.400 ;
        RECT 254.100 682.050 255.900 683.850 ;
        RECT 272.850 682.050 274.050 695.400 ;
        RECT 278.100 682.050 279.900 683.850 ;
        RECT 296.400 682.050 297.600 695.400 ;
        RECT 317.850 682.050 319.050 695.400 ;
        RECT 337.800 689.400 339.600 701.400 ;
        RECT 343.800 695.400 345.600 701.400 ;
        RECT 323.100 682.050 324.900 683.850 ;
        RECT 337.800 682.050 339.000 689.400 ;
        RECT 344.400 688.500 345.600 695.400 ;
        RECT 339.900 687.600 345.600 688.500 ;
        RECT 355.800 689.400 357.600 701.400 ;
        RECT 361.800 695.400 363.600 701.400 ;
        RECT 339.900 686.700 341.850 687.600 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 223.950 679.950 226.050 682.050 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 268.950 679.950 271.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 274.950 679.950 277.050 682.050 ;
        RECT 277.950 679.950 280.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 298.950 679.950 301.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 322.950 679.950 325.050 682.050 ;
        RECT 337.800 679.950 340.050 682.050 ;
        RECT 197.550 677.550 202.050 679.050 ;
        RECT 203.100 678.150 204.900 679.950 ;
        RECT 198.000 676.950 202.050 677.550 ;
        RECT 182.400 674.100 187.050 675.300 ;
        RECT 206.400 674.700 207.600 679.950 ;
        RECT 209.100 678.150 210.900 679.950 ;
        RECT 211.950 678.450 214.050 679.050 ;
        RECT 217.950 678.450 220.050 679.050 ;
        RECT 211.950 677.550 220.050 678.450 ;
        RECT 211.950 676.950 214.050 677.550 ;
        RECT 217.950 676.950 220.050 677.550 ;
        RECT 224.700 676.200 225.600 679.950 ;
        RECT 227.100 678.150 228.900 679.950 ;
        RECT 233.100 678.150 234.900 679.950 ;
        RECT 224.700 675.000 228.000 676.200 ;
        RECT 182.400 672.600 183.300 674.100 ;
        RECT 206.400 673.800 210.600 674.700 ;
        RECT 160.800 666.600 162.600 669.600 ;
        RECT 178.800 667.500 180.600 672.600 ;
        RECT 181.800 668.400 183.600 672.600 ;
        RECT 184.800 672.000 192.600 672.900 ;
        RECT 184.800 667.500 186.600 672.000 ;
        RECT 178.800 666.600 186.600 667.500 ;
        RECT 190.800 666.600 192.600 672.000 ;
        RECT 208.800 666.600 210.600 673.800 ;
        RECT 226.200 666.600 228.000 675.000 ;
        RECT 248.400 672.600 249.300 679.950 ;
        RECT 251.100 678.150 252.900 679.950 ;
        RECT 257.100 678.150 258.900 679.950 ;
        RECT 269.100 678.150 270.900 679.950 ;
        RECT 253.950 675.450 256.050 676.050 ;
        RECT 265.950 675.450 268.050 676.050 ;
        RECT 271.950 675.750 273.150 679.950 ;
        RECT 275.100 678.150 276.900 679.950 ;
        RECT 293.100 678.150 294.900 679.950 ;
        RECT 253.950 674.550 268.050 675.450 ;
        RECT 253.950 673.950 256.050 674.550 ;
        RECT 265.950 673.950 268.050 674.550 ;
        RECT 269.400 674.700 273.150 675.750 ;
        RECT 296.400 674.700 297.600 679.950 ;
        RECT 299.100 678.150 300.900 679.950 ;
        RECT 314.100 678.150 315.900 679.950 ;
        RECT 269.400 672.600 270.600 674.700 ;
        RECT 293.400 673.800 297.600 674.700 ;
        RECT 298.950 675.450 301.050 676.050 ;
        RECT 307.950 675.450 310.050 676.050 ;
        RECT 316.950 675.750 318.150 679.950 ;
        RECT 320.100 678.150 321.900 679.950 ;
        RECT 298.950 674.550 310.050 675.450 ;
        RECT 298.950 673.950 301.050 674.550 ;
        RECT 307.950 673.950 310.050 674.550 ;
        RECT 314.400 674.700 318.150 675.750 ;
        RECT 248.400 671.400 253.500 672.600 ;
        RECT 251.700 666.600 253.500 671.400 ;
        RECT 268.800 666.600 270.600 672.600 ;
        RECT 271.800 671.700 279.600 673.050 ;
        RECT 271.800 666.600 273.600 671.700 ;
        RECT 277.800 666.600 279.600 671.700 ;
        RECT 293.400 666.600 295.200 673.800 ;
        RECT 314.400 672.600 315.600 674.700 ;
        RECT 313.800 666.600 315.600 672.600 ;
        RECT 316.800 671.700 324.600 673.050 ;
        RECT 316.800 666.600 318.600 671.700 ;
        RECT 322.800 666.600 324.600 671.700 ;
        RECT 337.800 672.600 339.000 679.950 ;
        RECT 340.950 675.300 341.850 686.700 ;
        RECT 344.100 682.050 345.900 683.850 ;
        RECT 355.800 682.050 357.000 689.400 ;
        RECT 362.400 688.500 363.600 695.400 ;
        RECT 373.800 690.600 375.600 701.400 ;
        RECT 373.800 689.400 378.600 690.600 ;
        RECT 376.500 688.500 378.600 689.400 ;
        RECT 381.300 689.400 383.100 701.400 ;
        RECT 388.800 690.300 390.600 701.400 ;
        RECT 386.100 689.400 390.600 690.300 ;
        RECT 403.800 689.400 405.600 701.400 ;
        RECT 409.800 695.400 411.600 701.400 ;
        RECT 357.900 687.600 363.600 688.500 ;
        RECT 381.300 687.900 382.500 689.400 ;
        RECT 357.900 686.700 359.850 687.600 ;
        RECT 343.950 679.950 346.050 682.050 ;
        RECT 355.800 679.950 358.050 682.050 ;
        RECT 339.900 674.400 341.850 675.300 ;
        RECT 339.900 673.500 345.600 674.400 ;
        RECT 337.800 666.600 339.600 672.600 ;
        RECT 344.400 669.600 345.600 673.500 ;
        RECT 343.800 666.600 345.600 669.600 ;
        RECT 355.800 672.600 357.000 679.950 ;
        RECT 358.950 675.300 359.850 686.700 ;
        RECT 381.000 687.000 382.500 687.900 ;
        RECT 386.100 687.300 388.200 689.400 ;
        RECT 364.950 684.450 369.000 685.050 ;
        RECT 381.000 684.900 381.900 687.000 ;
        RECT 362.100 682.050 363.900 683.850 ;
        RECT 364.950 682.950 369.450 684.450 ;
        RECT 361.950 679.950 364.050 682.050 ;
        RECT 368.550 681.450 369.450 682.950 ;
        RECT 374.100 682.050 375.900 683.850 ;
        RECT 379.800 682.800 381.900 684.900 ;
        RECT 382.800 685.500 384.900 685.800 ;
        RECT 382.800 683.700 386.700 685.500 ;
        RECT 373.950 681.450 376.050 682.050 ;
        RECT 380.400 681.900 382.800 682.800 ;
        RECT 368.550 680.550 376.050 681.450 ;
        RECT 373.950 679.950 376.050 680.550 ;
        RECT 378.600 679.200 380.400 681.000 ;
        RECT 378.750 677.100 380.850 679.200 ;
        RECT 381.750 676.200 382.800 681.900 ;
        RECT 383.700 681.900 385.500 682.500 ;
        RECT 403.800 682.050 405.000 689.400 ;
        RECT 410.400 688.500 411.600 695.400 ;
        RECT 405.900 687.600 411.600 688.500 ;
        RECT 425.400 689.400 427.200 701.400 ;
        RECT 442.800 695.400 444.600 701.400 ;
        RECT 461.400 695.400 463.200 701.400 ;
        RECT 405.900 686.700 407.850 687.600 ;
        RECT 388.500 681.900 394.050 682.050 ;
        RECT 383.700 680.700 394.050 681.900 ;
        RECT 388.500 679.950 394.050 680.700 ;
        RECT 403.800 679.950 406.050 682.050 ;
        RECT 357.900 674.400 359.850 675.300 ;
        RECT 357.900 673.500 363.600 674.400 ;
        RECT 376.500 673.500 378.600 674.700 ;
        RECT 379.800 674.100 382.800 676.200 ;
        RECT 383.700 677.400 385.500 679.200 ;
        RECT 388.800 678.150 390.600 679.950 ;
        RECT 383.700 675.300 385.800 677.400 ;
        RECT 383.700 674.400 390.000 675.300 ;
        RECT 355.800 666.600 357.600 672.600 ;
        RECT 362.400 669.600 363.600 673.500 ;
        RECT 361.800 666.600 363.600 669.600 ;
        RECT 373.800 672.600 378.600 673.500 ;
        RECT 381.600 672.600 382.800 674.100 ;
        RECT 388.800 672.600 390.000 674.400 ;
        RECT 403.800 672.600 405.000 679.950 ;
        RECT 406.950 675.300 407.850 686.700 ;
        RECT 417.000 684.450 421.050 685.050 ;
        RECT 410.100 682.050 411.900 683.850 ;
        RECT 416.550 682.950 421.050 684.450 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 416.550 679.050 417.450 682.950 ;
        RECT 425.400 682.050 426.600 689.400 ;
        RECT 435.000 687.450 439.050 688.050 ;
        RECT 434.550 685.950 439.050 687.450 ;
        RECT 434.550 684.450 435.450 685.950 ;
        RECT 431.550 683.550 435.450 684.450 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 412.950 677.550 417.450 679.050 ;
        RECT 422.100 678.150 423.900 679.950 ;
        RECT 412.950 676.950 417.000 677.550 ;
        RECT 405.900 674.400 407.850 675.300 ;
        RECT 405.900 673.500 411.600 674.400 ;
        RECT 373.800 666.600 375.600 672.600 ;
        RECT 381.300 666.600 383.100 672.600 ;
        RECT 388.800 666.600 390.600 672.600 ;
        RECT 403.800 666.600 405.600 672.600 ;
        RECT 410.400 669.600 411.600 673.500 ;
        RECT 409.800 666.600 411.600 669.600 ;
        RECT 425.400 672.600 426.600 679.950 ;
        RECT 431.550 679.050 432.450 683.550 ;
        RECT 437.100 682.050 438.900 683.850 ;
        RECT 442.950 682.050 444.150 695.400 ;
        RECT 461.400 688.500 462.600 695.400 ;
        RECT 467.400 689.400 469.200 701.400 ;
        RECT 461.400 687.600 467.100 688.500 ;
        RECT 465.150 686.700 467.100 687.600 ;
        RECT 461.100 682.050 462.900 683.850 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 439.950 679.950 442.050 682.050 ;
        RECT 442.950 679.950 445.050 682.050 ;
        RECT 445.950 679.950 448.050 682.050 ;
        RECT 460.950 679.950 463.050 682.050 ;
        RECT 431.550 677.550 436.050 679.050 ;
        RECT 440.100 678.150 441.900 679.950 ;
        RECT 432.000 676.950 436.050 677.550 ;
        RECT 443.850 675.750 445.050 679.950 ;
        RECT 446.100 678.150 447.900 679.950 ;
        RECT 443.850 674.700 447.600 675.750 ;
        RECT 425.400 666.600 427.200 672.600 ;
        RECT 437.400 671.700 445.200 673.050 ;
        RECT 437.400 666.600 439.200 671.700 ;
        RECT 443.400 666.600 445.200 671.700 ;
        RECT 446.400 672.600 447.600 674.700 ;
        RECT 465.150 675.300 466.050 686.700 ;
        RECT 468.000 682.050 469.200 689.400 ;
        RECT 482.400 695.400 484.200 701.400 ;
        RECT 482.400 688.500 483.600 695.400 ;
        RECT 488.400 689.400 490.200 701.400 ;
        RECT 503.400 690.300 505.200 701.400 ;
        RECT 503.400 689.400 507.900 690.300 ;
        RECT 510.900 689.400 512.700 701.400 ;
        RECT 518.400 690.600 520.200 701.400 ;
        RECT 482.400 687.600 488.100 688.500 ;
        RECT 486.150 686.700 488.100 687.600 ;
        RECT 482.100 682.050 483.900 683.850 ;
        RECT 466.950 679.950 469.200 682.050 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 465.150 674.400 467.100 675.300 ;
        RECT 461.400 673.500 467.100 674.400 ;
        RECT 446.400 666.600 448.200 672.600 ;
        RECT 461.400 669.600 462.600 673.500 ;
        RECT 468.000 672.600 469.200 679.950 ;
        RECT 486.150 675.300 487.050 686.700 ;
        RECT 489.000 682.050 490.200 689.400 ;
        RECT 505.800 687.300 507.900 689.400 ;
        RECT 511.500 687.900 512.700 689.400 ;
        RECT 515.400 689.400 520.200 690.600 ;
        RECT 533.400 695.400 535.200 701.400 ;
        RECT 515.400 688.500 517.500 689.400 ;
        RECT 533.400 688.500 534.600 695.400 ;
        RECT 539.400 689.400 541.200 701.400 ;
        RECT 511.500 687.000 513.000 687.900 ;
        RECT 533.400 687.600 539.100 688.500 ;
        RECT 509.100 685.500 511.200 685.800 ;
        RECT 507.300 683.700 511.200 685.500 ;
        RECT 512.100 684.900 513.000 687.000 ;
        RECT 537.150 686.700 539.100 687.600 ;
        RECT 512.100 682.800 514.200 684.900 ;
        RECT 487.950 679.950 490.200 682.050 ;
        RECT 499.950 681.900 505.500 682.050 ;
        RECT 508.500 681.900 510.300 682.500 ;
        RECT 499.950 680.700 510.300 681.900 ;
        RECT 511.200 681.900 513.600 682.800 ;
        RECT 518.100 682.050 519.900 683.850 ;
        RECT 526.950 682.950 529.050 685.050 ;
        RECT 499.950 679.950 505.500 680.700 ;
        RECT 486.150 674.400 488.100 675.300 ;
        RECT 461.400 666.600 463.200 669.600 ;
        RECT 467.400 666.600 469.200 672.600 ;
        RECT 482.400 673.500 488.100 674.400 ;
        RECT 482.400 669.600 483.600 673.500 ;
        RECT 489.000 672.600 490.200 679.950 ;
        RECT 503.400 678.150 505.200 679.950 ;
        RECT 508.500 677.400 510.300 679.200 ;
        RECT 508.200 675.300 510.300 677.400 ;
        RECT 504.000 674.400 510.300 675.300 ;
        RECT 511.200 676.200 512.250 681.900 ;
        RECT 517.950 681.450 520.050 682.050 ;
        RECT 522.000 681.450 526.050 682.050 ;
        RECT 513.600 679.200 515.400 681.000 ;
        RECT 517.950 680.550 526.050 681.450 ;
        RECT 517.950 679.950 520.050 680.550 ;
        RECT 522.000 679.950 526.050 680.550 ;
        RECT 513.150 677.100 515.250 679.200 ;
        RECT 504.000 672.600 505.200 674.400 ;
        RECT 511.200 674.100 514.200 676.200 ;
        RECT 527.550 676.050 528.450 682.950 ;
        RECT 533.100 682.050 534.900 683.850 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 511.200 672.600 512.400 674.100 ;
        RECT 515.400 673.500 517.500 674.700 ;
        RECT 523.950 674.550 528.450 676.050 ;
        RECT 537.150 675.300 538.050 686.700 ;
        RECT 540.000 682.050 541.200 689.400 ;
        RECT 557.400 695.400 559.200 701.400 ;
        RECT 557.400 682.050 558.600 695.400 ;
        RECT 578.700 690.600 580.500 701.400 ;
        RECT 596.400 695.400 598.200 701.400 ;
        RECT 578.700 689.400 582.300 690.600 ;
        RECT 578.100 682.050 579.900 683.850 ;
        RECT 581.400 682.050 582.300 689.400 ;
        RECT 596.400 688.500 597.600 695.400 ;
        RECT 602.400 689.400 604.200 701.400 ;
        RECT 596.400 687.600 602.100 688.500 ;
        RECT 600.150 686.700 602.100 687.600 ;
        RECT 584.100 682.050 585.900 683.850 ;
        RECT 596.100 682.050 597.900 683.850 ;
        RECT 538.950 679.950 541.200 682.050 ;
        RECT 553.950 679.950 556.050 682.050 ;
        RECT 556.950 679.950 559.050 682.050 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 577.950 679.950 580.050 682.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 523.950 673.950 528.000 674.550 ;
        RECT 537.150 674.400 539.100 675.300 ;
        RECT 533.400 673.500 539.100 674.400 ;
        RECT 515.400 672.600 520.200 673.500 ;
        RECT 482.400 666.600 484.200 669.600 ;
        RECT 488.400 666.600 490.200 672.600 ;
        RECT 503.400 666.600 505.200 672.600 ;
        RECT 510.900 666.600 512.700 672.600 ;
        RECT 518.400 666.600 520.200 672.600 ;
        RECT 533.400 669.600 534.600 673.500 ;
        RECT 540.000 672.600 541.200 679.950 ;
        RECT 554.100 678.150 555.900 679.950 ;
        RECT 557.400 674.700 558.600 679.950 ;
        RECT 560.100 678.150 561.900 679.950 ;
        RECT 557.400 673.800 561.600 674.700 ;
        RECT 533.400 666.600 535.200 669.600 ;
        RECT 539.400 666.600 541.200 672.600 ;
        RECT 559.800 666.600 561.600 673.800 ;
        RECT 581.400 669.600 582.300 679.950 ;
        RECT 600.150 675.300 601.050 686.700 ;
        RECT 603.000 682.050 604.200 689.400 ;
        RECT 620.400 695.400 622.200 701.400 ;
        RECT 638.400 695.400 640.200 701.400 ;
        RECT 652.800 695.400 654.600 701.400 ;
        RECT 671.400 695.400 673.200 701.400 ;
        RECT 694.800 695.400 696.600 701.400 ;
        RECT 620.400 682.050 621.600 695.400 ;
        RECT 635.100 682.050 636.900 683.850 ;
        RECT 638.400 682.050 639.600 695.400 ;
        RECT 653.400 682.050 654.600 695.400 ;
        RECT 656.100 682.050 657.900 683.850 ;
        RECT 671.850 682.050 673.050 695.400 ;
        RECT 677.100 682.050 678.900 683.850 ;
        RECT 689.100 682.050 690.900 683.850 ;
        RECT 694.950 682.050 696.150 695.400 ;
        RECT 697.950 693.450 700.050 694.050 ;
        RECT 709.950 693.450 712.050 694.050 ;
        RECT 697.950 692.550 712.050 693.450 ;
        RECT 697.950 691.950 700.050 692.550 ;
        RECT 709.950 691.950 712.050 692.550 ;
        RECT 713.400 690.300 715.200 701.400 ;
        RECT 713.400 689.400 717.900 690.300 ;
        RECT 720.900 689.400 722.700 701.400 ;
        RECT 728.400 690.600 730.200 701.400 ;
        RECT 715.800 687.300 717.900 689.400 ;
        RECT 721.500 687.900 722.700 689.400 ;
        RECT 725.400 689.400 730.200 690.600 ;
        RECT 740.400 690.300 742.200 701.400 ;
        RECT 746.400 690.300 748.200 701.400 ;
        RECT 740.400 689.400 748.200 690.300 ;
        RECT 749.400 689.400 751.200 701.400 ;
        RECT 769.800 695.400 771.600 701.400 ;
        RECT 775.950 699.450 778.050 700.050 ;
        RECT 787.950 699.450 790.050 700.050 ;
        RECT 775.950 698.550 790.050 699.450 ;
        RECT 775.950 697.950 778.050 698.550 ;
        RECT 787.950 697.950 790.050 698.550 ;
        RECT 794.400 695.400 796.200 701.400 ;
        RECT 814.800 695.400 816.600 701.400 ;
        RECT 725.400 688.500 727.500 689.400 ;
        RECT 721.500 687.000 723.000 687.900 ;
        RECT 719.100 685.500 721.200 685.800 ;
        RECT 700.950 684.450 705.000 685.050 ;
        RECT 700.950 682.950 705.450 684.450 ;
        RECT 717.300 683.700 721.200 685.500 ;
        RECT 722.100 684.900 723.000 687.000 ;
        RECT 601.950 679.950 604.200 682.050 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 619.950 679.950 622.050 682.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 634.950 679.950 637.050 682.050 ;
        RECT 637.950 679.950 640.050 682.050 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 667.950 679.950 670.050 682.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 673.950 679.950 676.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 688.950 679.950 691.050 682.050 ;
        RECT 691.950 679.950 694.050 682.050 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 697.950 679.950 700.050 682.050 ;
        RECT 600.150 674.400 602.100 675.300 ;
        RECT 596.400 673.500 602.100 674.400 ;
        RECT 596.400 669.600 597.600 673.500 ;
        RECT 603.000 672.600 604.200 679.950 ;
        RECT 617.100 678.150 618.900 679.950 ;
        RECT 620.400 674.700 621.600 679.950 ;
        RECT 623.100 678.150 624.900 679.950 ;
        RECT 620.400 673.800 624.600 674.700 ;
        RECT 580.800 666.600 582.600 669.600 ;
        RECT 596.400 666.600 598.200 669.600 ;
        RECT 602.400 666.600 604.200 672.600 ;
        RECT 622.800 666.600 624.600 673.800 ;
        RECT 638.400 669.600 639.600 679.950 ;
        RECT 653.400 669.600 654.600 679.950 ;
        RECT 668.100 678.150 669.900 679.950 ;
        RECT 670.950 675.750 672.150 679.950 ;
        RECT 674.100 678.150 675.900 679.950 ;
        RECT 692.100 678.150 693.900 679.950 ;
        RECT 668.400 674.700 672.150 675.750 ;
        RECT 695.850 675.750 697.050 679.950 ;
        RECT 698.100 678.150 699.900 679.950 ;
        RECT 704.550 679.050 705.450 682.950 ;
        RECT 722.100 682.800 724.200 684.900 ;
        RECT 709.950 681.900 715.500 682.050 ;
        RECT 718.500 681.900 720.300 682.500 ;
        RECT 709.950 680.700 720.300 681.900 ;
        RECT 721.200 681.900 723.600 682.800 ;
        RECT 728.100 682.050 729.900 683.850 ;
        RECT 743.100 682.050 744.900 683.850 ;
        RECT 749.700 682.050 750.600 689.400 ;
        RECT 756.000 687.450 760.050 688.050 ;
        RECT 755.550 685.950 760.050 687.450 ;
        RECT 709.950 679.950 715.500 680.700 ;
        RECT 700.950 677.550 705.450 679.050 ;
        RECT 713.400 678.150 715.200 679.950 ;
        RECT 700.950 676.950 705.000 677.550 ;
        RECT 718.500 677.400 720.300 679.200 ;
        RECT 695.850 674.700 699.600 675.750 ;
        RECT 718.200 675.300 720.300 677.400 ;
        RECT 668.400 672.600 669.600 674.700 ;
        RECT 638.400 666.600 640.200 669.600 ;
        RECT 652.800 666.600 654.600 669.600 ;
        RECT 667.800 666.600 669.600 672.600 ;
        RECT 670.800 671.700 678.600 673.050 ;
        RECT 670.800 666.600 672.600 671.700 ;
        RECT 676.800 666.600 678.600 671.700 ;
        RECT 689.400 671.700 697.200 673.050 ;
        RECT 689.400 666.600 691.200 671.700 ;
        RECT 695.400 666.600 697.200 671.700 ;
        RECT 698.400 672.600 699.600 674.700 ;
        RECT 714.000 674.400 720.300 675.300 ;
        RECT 721.200 676.200 722.250 681.900 ;
        RECT 727.950 681.450 730.050 682.050 ;
        RECT 723.600 679.200 725.400 681.000 ;
        RECT 727.950 680.550 735.450 681.450 ;
        RECT 727.950 679.950 730.050 680.550 ;
        RECT 723.150 677.100 725.250 679.200 ;
        RECT 734.550 679.050 735.450 680.550 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 734.550 677.550 739.050 679.050 ;
        RECT 740.100 678.150 741.900 679.950 ;
        RECT 746.100 678.150 747.900 679.950 ;
        RECT 735.000 676.950 739.050 677.550 ;
        RECT 714.000 672.600 715.200 674.400 ;
        RECT 721.200 674.100 724.200 676.200 ;
        RECT 721.200 672.600 722.400 674.100 ;
        RECT 725.400 673.500 727.500 674.700 ;
        RECT 725.400 672.600 730.200 673.500 ;
        RECT 749.700 672.600 750.600 679.950 ;
        RECT 755.550 679.050 756.450 685.950 ;
        RECT 759.000 684.450 763.050 685.050 ;
        RECT 751.950 677.550 756.450 679.050 ;
        RECT 758.550 682.950 763.050 684.450 ;
        RECT 758.550 679.050 759.450 682.950 ;
        RECT 764.100 682.050 765.900 683.850 ;
        RECT 769.950 682.050 771.150 695.400 ;
        RECT 794.850 682.050 796.050 695.400 ;
        RECT 800.100 682.050 801.900 683.850 ;
        RECT 809.100 682.050 810.900 683.850 ;
        RECT 814.950 682.050 816.150 695.400 ;
        RECT 833.400 689.400 835.200 701.400 ;
        RECT 840.900 690.900 842.700 701.400 ;
        RECT 840.900 689.400 843.300 690.900 ;
        RECT 859.800 690.600 861.600 701.400 ;
        RECT 859.800 689.400 864.600 690.600 ;
        RECT 833.400 687.900 834.600 689.400 ;
        RECT 833.400 686.700 840.600 687.900 ;
        RECT 838.800 686.100 840.600 686.700 ;
        RECT 820.950 684.450 823.050 685.050 ;
        RECT 820.950 683.550 828.450 684.450 ;
        RECT 820.950 682.950 823.050 683.550 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 758.550 677.550 763.050 679.050 ;
        RECT 767.100 678.150 768.900 679.950 ;
        RECT 751.950 676.950 756.000 677.550 ;
        RECT 759.000 676.950 763.050 677.550 ;
        RECT 770.850 675.750 772.050 679.950 ;
        RECT 773.100 678.150 774.900 679.950 ;
        RECT 791.100 678.150 792.900 679.950 ;
        RECT 793.950 675.750 795.150 679.950 ;
        RECT 797.100 678.150 798.900 679.950 ;
        RECT 812.100 678.150 813.900 679.950 ;
        RECT 770.850 674.700 774.600 675.750 ;
        RECT 698.400 666.600 700.200 672.600 ;
        RECT 713.400 666.600 715.200 672.600 ;
        RECT 720.900 666.600 722.700 672.600 ;
        RECT 728.400 666.600 730.200 672.600 ;
        RECT 745.500 671.400 750.600 672.600 ;
        RECT 764.400 671.700 772.200 673.050 ;
        RECT 745.500 666.600 747.300 671.400 ;
        RECT 764.400 666.600 766.200 671.700 ;
        RECT 770.400 666.600 772.200 671.700 ;
        RECT 773.400 672.600 774.600 674.700 ;
        RECT 791.400 674.700 795.150 675.750 ;
        RECT 815.850 675.750 817.050 679.950 ;
        RECT 818.100 678.150 819.900 679.950 ;
        RECT 827.550 678.450 828.450 683.550 ;
        RECT 836.100 682.050 837.900 683.850 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 827.550 677.550 831.450 678.450 ;
        RECT 833.100 678.150 834.900 679.950 ;
        RECT 830.550 676.050 831.450 677.550 ;
        RECT 815.850 674.700 819.600 675.750 ;
        RECT 791.400 672.600 792.600 674.700 ;
        RECT 773.400 666.600 775.200 672.600 ;
        RECT 790.800 666.600 792.600 672.600 ;
        RECT 793.800 671.700 801.600 673.050 ;
        RECT 793.800 666.600 795.600 671.700 ;
        RECT 799.800 666.600 801.600 671.700 ;
        RECT 809.400 671.700 817.200 673.050 ;
        RECT 809.400 666.600 811.200 671.700 ;
        RECT 815.400 666.600 817.200 671.700 ;
        RECT 818.400 672.600 819.600 674.700 ;
        RECT 830.550 674.550 835.050 676.050 ;
        RECT 839.700 675.600 840.600 686.100 ;
        RECT 841.950 682.050 843.300 689.400 ;
        RECT 862.500 688.500 864.600 689.400 ;
        RECT 867.300 689.400 869.100 701.400 ;
        RECT 874.800 690.300 876.600 701.400 ;
        RECT 872.100 689.400 876.600 690.300 ;
        RECT 887.700 690.600 889.500 701.400 ;
        RECT 887.700 689.400 891.300 690.600 ;
        RECT 905.400 690.300 907.200 701.400 ;
        RECT 911.400 690.300 913.200 701.400 ;
        RECT 905.400 689.400 913.200 690.300 ;
        RECT 914.400 689.400 916.200 701.400 ;
        RECT 867.300 687.900 868.500 689.400 ;
        RECT 867.000 687.000 868.500 687.900 ;
        RECT 872.100 687.300 874.200 689.400 ;
        RECT 844.950 684.450 847.050 685.050 ;
        RECT 867.000 684.900 867.900 687.000 ;
        RECT 844.950 683.550 855.450 684.450 ;
        RECT 844.950 682.950 847.050 683.550 ;
        RECT 841.950 679.950 844.050 682.050 ;
        RECT 854.550 681.450 855.450 683.550 ;
        RECT 860.100 682.050 861.900 683.850 ;
        RECT 865.800 682.800 867.900 684.900 ;
        RECT 868.800 685.500 870.900 685.800 ;
        RECT 868.800 683.700 872.700 685.500 ;
        RECT 859.950 681.450 862.050 682.050 ;
        RECT 866.400 681.900 868.800 682.800 ;
        RECT 854.550 680.550 862.050 681.450 ;
        RECT 859.950 679.950 862.050 680.550 ;
        RECT 838.800 674.700 840.600 675.600 ;
        RECT 831.000 673.950 835.050 674.550 ;
        RECT 837.300 673.800 840.600 674.700 ;
        RECT 818.400 666.600 820.200 672.600 ;
        RECT 837.300 669.600 838.200 673.800 ;
        RECT 843.000 672.600 844.050 679.950 ;
        RECT 864.600 679.200 866.400 681.000 ;
        RECT 864.750 677.100 866.850 679.200 ;
        RECT 867.750 676.200 868.800 681.900 ;
        RECT 869.700 681.900 871.500 682.500 ;
        RECT 887.100 682.050 888.900 683.850 ;
        RECT 890.400 682.050 891.300 689.400 ;
        RECT 898.950 685.950 901.050 688.050 ;
        RECT 893.100 682.050 894.900 683.850 ;
        RECT 874.500 681.900 876.600 682.050 ;
        RECT 869.700 680.700 876.600 681.900 ;
        RECT 874.500 679.950 876.600 680.700 ;
        RECT 886.950 679.950 889.050 682.050 ;
        RECT 889.950 679.950 892.050 682.050 ;
        RECT 892.950 679.950 895.050 682.050 ;
        RECT 862.500 673.500 864.600 674.700 ;
        RECT 865.800 674.100 868.800 676.200 ;
        RECT 869.700 677.400 871.500 679.200 ;
        RECT 874.800 678.450 876.600 679.950 ;
        RECT 883.950 678.450 886.050 679.050 ;
        RECT 874.800 678.150 886.050 678.450 ;
        RECT 875.550 677.550 886.050 678.150 ;
        RECT 869.700 675.300 871.800 677.400 ;
        RECT 883.950 676.950 886.050 677.550 ;
        RECT 869.700 674.400 876.000 675.300 ;
        RECT 859.800 672.600 864.600 673.500 ;
        RECT 867.600 672.600 868.800 674.100 ;
        RECT 874.800 672.600 876.000 674.400 ;
        RECT 836.400 666.600 838.200 669.600 ;
        RECT 842.400 666.600 844.200 672.600 ;
        RECT 859.800 666.600 861.600 672.600 ;
        RECT 867.300 666.600 869.100 672.600 ;
        RECT 874.800 666.600 876.600 672.600 ;
        RECT 890.400 669.600 891.300 679.950 ;
        RECT 899.550 679.050 900.450 685.950 ;
        RECT 908.100 682.050 909.900 683.850 ;
        RECT 914.700 682.050 915.600 689.400 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 907.950 679.950 910.050 682.050 ;
        RECT 910.950 679.950 913.050 682.050 ;
        RECT 913.950 679.950 916.050 682.050 ;
        RECT 895.950 677.550 900.450 679.050 ;
        RECT 905.100 678.150 906.900 679.950 ;
        RECT 911.100 678.150 912.900 679.950 ;
        RECT 895.950 676.950 900.000 677.550 ;
        RECT 914.700 672.600 915.600 679.950 ;
        RECT 910.500 671.400 915.600 672.600 ;
        RECT 889.800 666.600 891.600 669.600 ;
        RECT 910.500 666.600 912.300 671.400 ;
        RECT 16.800 659.400 18.600 662.400 ;
        RECT 17.400 649.050 18.300 659.400 ;
        RECT 31.800 656.400 33.600 662.400 ;
        RECT 32.400 654.300 33.600 656.400 ;
        RECT 34.800 657.300 36.600 662.400 ;
        RECT 40.800 657.300 42.600 662.400 ;
        RECT 34.800 655.950 42.600 657.300 ;
        RECT 58.500 657.600 60.300 662.400 ;
        RECT 58.500 656.400 63.600 657.600 ;
        RECT 32.400 653.250 36.150 654.300 ;
        RECT 32.100 649.050 33.900 650.850 ;
        RECT 34.950 649.050 36.150 653.250 ;
        RECT 38.100 649.050 39.900 650.850 ;
        RECT 53.100 649.050 54.900 650.850 ;
        RECT 59.100 649.050 60.900 650.850 ;
        RECT 62.700 649.050 63.600 656.400 ;
        RECT 74.400 657.300 76.200 662.400 ;
        RECT 80.400 657.300 82.200 662.400 ;
        RECT 74.400 655.950 82.200 657.300 ;
        RECT 83.400 656.400 85.200 662.400 ;
        RECT 101.400 659.400 103.200 662.400 ;
        RECT 83.400 654.300 84.600 656.400 ;
        RECT 102.300 655.200 103.200 659.400 ;
        RECT 107.400 656.400 109.200 662.400 ;
        RECT 122.400 656.400 124.200 662.400 ;
        RECT 129.600 657.000 131.400 662.400 ;
        RECT 102.300 654.300 105.600 655.200 ;
        RECT 80.850 653.250 84.600 654.300 ;
        RECT 103.800 653.400 105.600 654.300 ;
        RECT 64.950 651.450 69.000 652.050 ;
        RECT 64.950 649.950 69.450 651.450 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 14.100 645.150 15.900 646.950 ;
        RECT 17.400 639.600 18.300 646.950 ;
        RECT 20.100 645.150 21.900 646.950 ;
        RECT 14.700 638.400 18.300 639.600 ;
        RECT 14.700 627.600 16.500 638.400 ;
        RECT 35.850 633.600 37.050 646.950 ;
        RECT 41.100 645.150 42.900 646.950 ;
        RECT 56.100 645.150 57.900 646.950 ;
        RECT 62.700 639.600 63.600 646.950 ;
        RECT 68.550 645.450 69.450 649.950 ;
        RECT 77.100 649.050 78.900 650.850 ;
        RECT 80.850 649.050 82.050 653.250 ;
        RECT 83.100 649.050 84.900 650.850 ;
        RECT 98.100 649.050 99.900 650.850 ;
        RECT 73.950 646.950 76.050 649.050 ;
        RECT 76.950 646.950 79.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 97.950 646.950 100.050 649.050 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 68.550 644.550 72.450 645.450 ;
        RECT 74.100 645.150 75.900 646.950 ;
        RECT 71.550 643.050 72.450 644.550 ;
        RECT 71.550 641.550 76.050 643.050 ;
        RECT 72.000 640.950 76.050 641.550 ;
        RECT 53.400 638.700 61.200 639.600 ;
        RECT 35.400 627.600 37.200 633.600 ;
        RECT 53.400 627.600 55.200 638.700 ;
        RECT 59.400 627.600 61.200 638.700 ;
        RECT 62.400 627.600 64.200 639.600 ;
        RECT 79.950 633.600 81.150 646.950 ;
        RECT 101.100 645.150 102.900 646.950 ;
        RECT 104.700 642.900 105.600 653.400 ;
        RECT 108.000 649.050 109.050 656.400 ;
        RECT 122.400 655.500 123.900 656.400 ;
        RECT 122.400 654.000 126.750 655.500 ;
        RECT 124.650 653.400 126.750 654.000 ;
        RECT 130.350 654.900 131.400 657.000 ;
        RECT 137.400 656.400 139.200 662.400 ;
        RECT 134.700 655.200 139.200 656.400 ;
        RECT 149.400 657.300 151.200 662.400 ;
        RECT 155.400 657.300 157.200 662.400 ;
        RECT 149.400 655.950 157.200 657.300 ;
        RECT 158.400 656.400 160.200 662.400 ;
        RECT 127.650 651.900 129.450 653.700 ;
        RECT 130.350 652.800 133.500 654.900 ;
        RECT 134.700 653.100 136.800 655.200 ;
        RECT 158.400 654.300 159.600 656.400 ;
        RECT 178.800 655.200 180.600 662.400 ;
        RECT 184.950 660.450 187.050 661.050 ;
        RECT 190.950 660.450 193.050 661.050 ;
        RECT 184.950 659.550 193.050 660.450 ;
        RECT 184.950 658.950 187.050 659.550 ;
        RECT 190.950 658.950 193.050 659.550 ;
        RECT 155.850 653.250 159.600 654.300 ;
        RECT 176.400 654.300 180.600 655.200 ;
        RECT 197.400 655.200 199.200 662.400 ;
        RECT 217.800 656.400 219.600 662.400 ;
        RECT 225.600 657.000 227.400 662.400 ;
        RECT 217.800 655.200 222.300 656.400 ;
        RECT 197.400 654.300 201.600 655.200 ;
        RECT 127.200 651.000 129.300 651.900 ;
        RECT 122.700 649.800 129.300 651.000 ;
        RECT 122.700 649.200 124.500 649.800 ;
        RECT 103.800 642.300 105.600 642.900 ;
        RECT 98.400 641.100 105.600 642.300 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 122.400 647.100 124.500 649.200 ;
        RECT 98.400 639.600 99.600 641.100 ;
        RECT 106.950 639.600 108.300 646.950 ;
        RECT 127.200 646.800 129.300 648.900 ;
        RECT 127.200 645.000 129.000 646.800 ;
        RECT 130.350 646.200 131.250 652.800 ;
        RECT 132.150 648.900 134.250 651.000 ;
        RECT 132.300 647.100 134.100 648.900 ;
        RECT 136.950 647.100 139.050 649.200 ;
        RECT 152.100 649.050 153.900 650.850 ;
        RECT 155.850 649.050 157.050 653.250 ;
        RECT 158.100 649.050 159.900 650.850 ;
        RECT 173.100 649.050 174.900 650.850 ;
        RECT 176.400 649.050 177.600 654.300 ;
        RECT 179.100 649.050 180.900 650.850 ;
        RECT 197.100 649.050 198.900 650.850 ;
        RECT 200.400 649.050 201.600 654.300 ;
        RECT 220.200 653.100 222.300 655.200 ;
        RECT 225.600 654.900 226.650 657.000 ;
        RECT 232.800 656.400 234.600 662.400 ;
        RECT 233.100 655.500 234.600 656.400 ;
        RECT 223.500 652.800 226.650 654.900 ;
        RECT 230.250 654.000 234.600 655.500 ;
        RECT 248.400 655.200 250.200 662.400 ;
        RECT 265.800 661.500 273.600 662.400 ;
        RECT 265.800 656.400 267.600 661.500 ;
        RECT 268.800 656.400 270.600 660.600 ;
        RECT 271.800 657.000 273.600 661.500 ;
        RECT 277.800 657.000 279.600 662.400 ;
        RECT 294.300 658.200 296.100 662.400 ;
        RECT 248.400 654.300 252.600 655.200 ;
        RECT 203.100 649.050 204.900 650.850 ;
        RECT 130.350 644.700 133.500 646.200 ;
        RECT 137.100 645.450 138.900 647.100 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 151.950 646.950 154.050 649.050 ;
        RECT 154.950 646.950 157.050 649.050 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 172.950 646.950 175.050 649.050 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 196.950 646.950 199.050 649.050 ;
        RECT 199.950 646.950 202.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 217.950 647.100 220.050 649.200 ;
        RECT 222.750 648.900 224.850 651.000 ;
        RECT 222.900 647.100 224.700 648.900 ;
        RECT 142.950 645.450 145.050 646.050 ;
        RECT 137.100 645.300 145.050 645.450 ;
        RECT 131.400 644.100 133.500 644.700 ;
        RECT 137.550 644.550 145.050 645.300 ;
        RECT 149.100 645.150 150.900 646.950 ;
        RECT 128.700 641.700 130.500 643.800 ;
        RECT 125.100 640.800 130.500 641.700 ;
        RECT 125.100 639.900 127.200 640.800 ;
        RECT 79.800 627.600 81.600 633.600 ;
        RECT 98.400 627.600 100.200 639.600 ;
        RECT 105.900 638.100 108.300 639.600 ;
        RECT 122.400 638.700 127.200 639.900 ;
        RECT 132.000 639.600 133.200 644.100 ;
        RECT 142.950 643.950 145.050 644.550 ;
        RECT 129.900 638.700 133.200 639.600 ;
        RECT 134.100 639.600 136.200 640.500 ;
        RECT 105.900 627.600 107.700 638.100 ;
        RECT 122.400 627.600 124.200 638.700 ;
        RECT 129.900 627.600 131.700 638.700 ;
        RECT 134.100 638.400 139.200 639.600 ;
        RECT 137.400 627.600 139.200 638.400 ;
        RECT 154.950 633.600 156.150 646.950 ;
        RECT 176.400 633.600 177.600 646.950 ;
        RECT 200.400 633.600 201.600 646.950 ;
        RECT 218.100 646.050 219.900 647.100 ;
        RECT 225.750 646.200 226.650 652.800 ;
        RECT 227.550 651.900 229.350 653.700 ;
        RECT 230.250 653.400 232.350 654.000 ;
        RECT 227.700 651.000 229.800 651.900 ;
        RECT 227.700 649.800 234.300 651.000 ;
        RECT 232.500 649.200 234.300 649.800 ;
        RECT 232.500 649.050 234.600 649.200 ;
        RECT 248.100 649.050 249.900 650.850 ;
        RECT 251.400 649.050 252.600 654.300 ;
        RECT 269.400 654.900 270.300 656.400 ;
        RECT 271.800 656.100 279.600 657.000 ;
        RECT 293.400 656.400 296.100 658.200 ;
        RECT 269.400 653.700 274.050 654.900 ;
        RECT 254.100 649.050 255.900 650.850 ;
        RECT 269.100 649.050 270.900 650.850 ;
        RECT 272.700 649.050 274.050 653.700 ;
        RECT 275.100 649.050 276.900 650.850 ;
        RECT 293.400 649.050 294.300 656.400 ;
        RECT 296.100 654.600 297.900 655.500 ;
        RECT 301.800 654.600 303.600 662.400 ;
        RECT 296.100 653.700 303.600 654.600 ;
        RECT 317.400 655.200 319.200 662.400 ;
        RECT 337.800 656.400 339.600 662.400 ;
        RECT 343.800 659.400 345.600 662.400 ;
        RECT 317.400 654.300 321.600 655.200 ;
        RECT 227.700 646.800 229.800 648.900 ;
        RECT 232.500 647.100 238.050 649.050 ;
        RECT 234.000 646.950 238.050 647.100 ;
        RECT 247.950 646.950 250.050 649.050 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 268.950 646.950 271.050 649.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 274.950 646.950 277.050 649.050 ;
        RECT 277.950 646.950 280.050 649.050 ;
        RECT 292.950 646.950 295.050 649.050 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 216.000 645.900 219.900 646.050 ;
        RECT 214.950 645.300 219.900 645.900 ;
        RECT 214.950 644.550 219.450 645.300 ;
        RECT 223.500 644.700 226.650 646.200 ;
        RECT 228.000 645.000 229.800 646.800 ;
        RECT 214.950 643.950 219.000 644.550 ;
        RECT 223.500 644.100 225.600 644.700 ;
        RECT 214.950 643.800 217.050 643.950 ;
        RECT 202.950 642.450 205.050 643.050 ;
        RECT 215.550 642.450 216.450 643.800 ;
        RECT 202.950 641.550 216.450 642.450 ;
        RECT 202.950 640.950 205.050 641.550 ;
        RECT 220.800 639.600 222.900 640.500 ;
        RECT 154.800 627.600 156.600 633.600 ;
        RECT 176.400 627.600 178.200 633.600 ;
        RECT 199.800 627.600 201.600 633.600 ;
        RECT 217.800 638.400 222.900 639.600 ;
        RECT 223.800 639.600 225.000 644.100 ;
        RECT 226.500 641.700 228.300 643.800 ;
        RECT 226.500 640.800 231.900 641.700 ;
        RECT 229.800 639.900 231.900 640.800 ;
        RECT 223.800 638.700 227.100 639.600 ;
        RECT 229.800 638.700 234.600 639.900 ;
        RECT 217.800 627.600 219.600 638.400 ;
        RECT 225.300 627.600 227.100 638.700 ;
        RECT 232.800 627.600 234.600 638.700 ;
        RECT 251.400 633.600 252.600 646.950 ;
        RECT 266.100 645.150 267.900 646.950 ;
        RECT 272.700 639.600 273.900 646.950 ;
        RECT 278.100 645.150 279.900 646.950 ;
        RECT 293.400 639.600 294.300 646.950 ;
        RECT 296.100 645.150 297.900 646.950 ;
        RECT 250.800 627.600 252.600 633.600 ;
        RECT 271.800 627.600 275.100 639.600 ;
        RECT 292.800 627.600 294.600 639.600 ;
        RECT 299.700 633.600 300.600 653.700 ;
        RECT 302.100 649.050 303.900 650.850 ;
        RECT 317.100 649.050 318.900 650.850 ;
        RECT 320.400 649.050 321.600 654.300 ;
        RECT 323.100 649.050 324.900 650.850 ;
        RECT 337.800 649.050 339.000 656.400 ;
        RECT 344.400 655.500 345.600 659.400 ;
        RECT 339.900 654.600 345.600 655.500 ;
        RECT 358.800 656.400 360.600 662.400 ;
        RECT 364.800 659.400 366.600 662.400 ;
        RECT 339.900 653.700 341.850 654.600 ;
        RECT 301.950 646.950 304.050 649.050 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 337.800 646.950 340.050 649.050 ;
        RECT 301.950 642.450 304.050 643.050 ;
        RECT 316.950 642.450 319.050 643.050 ;
        RECT 301.950 641.550 319.050 642.450 ;
        RECT 301.950 640.950 304.050 641.550 ;
        RECT 316.950 640.950 319.050 641.550 ;
        RECT 320.400 633.600 321.600 646.950 ;
        RECT 298.800 627.600 300.600 633.600 ;
        RECT 319.800 627.600 321.600 633.600 ;
        RECT 337.800 639.600 339.000 646.950 ;
        RECT 340.950 642.300 341.850 653.700 ;
        RECT 358.800 649.050 360.000 656.400 ;
        RECT 365.400 655.500 366.600 659.400 ;
        RECT 379.800 656.400 381.600 662.400 ;
        RECT 387.300 656.400 389.100 662.400 ;
        RECT 394.800 656.400 396.600 662.400 ;
        RECT 407.400 657.300 409.200 662.400 ;
        RECT 413.400 657.300 415.200 662.400 ;
        RECT 379.800 655.500 384.600 656.400 ;
        RECT 360.900 654.600 366.600 655.500 ;
        RECT 360.900 653.700 362.850 654.600 ;
        RECT 382.500 654.300 384.600 655.500 ;
        RECT 387.600 654.900 388.800 656.400 ;
        RECT 343.950 646.950 346.050 649.050 ;
        RECT 358.800 646.950 361.050 649.050 ;
        RECT 344.100 645.150 345.900 646.950 ;
        RECT 339.900 641.400 341.850 642.300 ;
        RECT 339.900 640.500 345.600 641.400 ;
        RECT 337.800 627.600 339.600 639.600 ;
        RECT 344.400 633.600 345.600 640.500 ;
        RECT 343.800 627.600 345.600 633.600 ;
        RECT 358.800 639.600 360.000 646.950 ;
        RECT 361.950 642.300 362.850 653.700 ;
        RECT 385.800 652.800 388.800 654.900 ;
        RECT 394.800 654.600 396.000 656.400 ;
        RECT 407.400 655.950 415.200 657.300 ;
        RECT 416.400 656.400 418.200 662.400 ;
        RECT 422.550 656.400 424.350 662.400 ;
        RECT 430.650 659.400 432.450 662.400 ;
        RECT 438.450 659.400 440.250 662.400 ;
        RECT 446.250 660.300 448.050 662.400 ;
        RECT 446.250 659.400 450.000 660.300 ;
        RECT 430.650 658.500 431.700 659.400 ;
        RECT 427.950 657.300 431.700 658.500 ;
        RECT 439.200 658.500 440.250 659.400 ;
        RECT 448.950 658.500 450.000 659.400 ;
        RECT 439.200 657.450 444.150 658.500 ;
        RECT 427.950 656.400 430.050 657.300 ;
        RECT 442.350 656.700 444.150 657.450 ;
        RECT 367.950 651.450 372.000 652.050 ;
        RECT 367.950 649.950 372.450 651.450 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 365.100 645.150 366.900 646.950 ;
        RECT 371.550 645.450 372.450 649.950 ;
        RECT 384.750 649.800 386.850 651.900 ;
        RECT 373.950 648.450 378.000 649.050 ;
        RECT 379.950 648.450 382.050 649.050 ;
        RECT 373.950 647.550 382.050 648.450 ;
        RECT 384.600 648.000 386.400 649.800 ;
        RECT 373.950 646.950 378.000 647.550 ;
        RECT 379.950 646.950 382.050 647.550 ;
        RECT 387.750 647.100 388.800 652.800 ;
        RECT 389.700 653.700 396.000 654.600 ;
        RECT 416.400 654.300 417.600 656.400 ;
        RECT 389.700 651.600 391.800 653.700 ;
        RECT 413.850 653.250 417.600 654.300 ;
        RECT 389.700 649.800 391.500 651.600 ;
        RECT 400.950 651.450 403.050 652.050 ;
        RECT 395.550 650.850 403.050 651.450 ;
        RECT 394.800 650.550 403.050 650.850 ;
        RECT 394.800 649.050 396.600 650.550 ;
        RECT 400.950 649.950 403.050 650.550 ;
        RECT 410.100 649.050 411.900 650.850 ;
        RECT 413.850 649.050 415.050 653.250 ;
        RECT 416.100 649.050 417.900 650.850 ;
        RECT 422.550 649.050 423.750 656.400 ;
        RECT 445.650 655.800 447.450 657.600 ;
        RECT 448.950 656.400 451.050 658.500 ;
        RECT 454.050 656.400 455.850 662.400 ;
        RECT 435.150 654.000 436.950 654.600 ;
        RECT 446.100 654.000 447.150 655.800 ;
        RECT 435.150 652.800 447.150 654.000 ;
        RECT 394.500 648.300 396.600 649.050 ;
        RECT 371.550 644.550 375.450 645.450 ;
        RECT 380.100 645.150 381.900 646.950 ;
        RECT 386.400 646.200 388.800 647.100 ;
        RECT 389.700 647.100 396.600 648.300 ;
        RECT 389.700 646.500 391.500 647.100 ;
        RECT 394.500 646.950 396.600 647.100 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 415.950 646.950 418.050 649.050 ;
        RECT 422.550 647.250 428.850 649.050 ;
        RECT 422.550 646.950 427.050 647.250 ;
        RECT 360.900 641.400 362.850 642.300 ;
        RECT 374.550 643.050 375.450 644.550 ;
        RECT 385.800 644.100 387.900 646.200 ;
        RECT 374.550 641.550 379.050 643.050 ;
        RECT 360.900 640.500 366.600 641.400 ;
        RECT 375.000 640.950 379.050 641.550 ;
        RECT 387.000 642.000 387.900 644.100 ;
        RECT 388.800 643.500 392.700 645.300 ;
        RECT 407.100 645.150 408.900 646.950 ;
        RECT 388.800 643.200 390.900 643.500 ;
        RECT 387.000 641.100 388.500 642.000 ;
        RECT 358.800 627.600 360.600 639.600 ;
        RECT 365.400 633.600 366.600 640.500 ;
        RECT 382.500 639.600 384.600 640.500 ;
        RECT 364.800 627.600 366.600 633.600 ;
        RECT 379.800 638.400 384.600 639.600 ;
        RECT 387.300 639.600 388.500 641.100 ;
        RECT 392.100 639.600 394.200 641.700 ;
        RECT 379.800 627.600 381.600 638.400 ;
        RECT 387.300 631.050 389.100 639.600 ;
        RECT 392.100 638.700 396.600 639.600 ;
        RECT 385.950 628.950 389.100 631.050 ;
        RECT 387.300 627.600 389.100 628.950 ;
        RECT 394.800 627.600 396.600 638.700 ;
        RECT 412.950 633.600 414.150 646.950 ;
        RECT 422.550 639.600 423.750 646.950 ;
        RECT 424.950 641.400 426.750 643.200 ;
        RECT 425.850 640.200 430.050 641.400 ;
        RECT 435.150 640.200 436.050 652.800 ;
        RECT 446.100 651.600 453.000 652.800 ;
        RECT 446.100 651.000 447.900 651.600 ;
        RECT 452.100 650.850 453.000 651.600 ;
        RECT 449.100 649.800 450.900 650.400 ;
        RECT 442.950 648.600 450.900 649.800 ;
        RECT 452.100 649.050 453.900 650.850 ;
        RECT 442.950 646.950 445.050 648.600 ;
        RECT 451.950 646.950 454.050 649.050 ;
        RECT 444.750 641.700 446.550 642.000 ;
        RECT 454.950 641.700 455.850 656.400 ;
        RECT 444.750 641.100 455.850 641.700 ;
        RECT 412.800 627.600 414.600 633.600 ;
        RECT 422.550 627.600 424.350 639.600 ;
        RECT 427.950 639.300 430.050 640.200 ;
        RECT 430.950 639.300 436.050 640.200 ;
        RECT 438.150 640.500 455.850 641.100 ;
        RECT 438.150 640.200 446.550 640.500 ;
        RECT 430.950 638.400 431.850 639.300 ;
        RECT 429.150 636.600 431.850 638.400 ;
        RECT 432.750 638.100 434.550 638.400 ;
        RECT 438.150 638.100 439.050 640.200 ;
        RECT 454.950 639.600 455.850 640.500 ;
        RECT 432.750 637.200 439.050 638.100 ;
        RECT 439.950 638.700 441.750 639.300 ;
        RECT 439.950 637.500 447.450 638.700 ;
        RECT 432.750 636.600 434.550 637.200 ;
        RECT 446.250 636.600 447.450 637.500 ;
        RECT 427.950 633.600 431.850 635.700 ;
        RECT 436.950 635.550 438.750 636.300 ;
        RECT 441.750 635.550 443.550 636.300 ;
        RECT 436.950 634.500 443.550 635.550 ;
        RECT 446.250 634.500 451.050 636.600 ;
        RECT 430.050 627.600 431.850 633.600 ;
        RECT 437.850 627.600 439.650 634.500 ;
        RECT 446.250 633.600 447.450 634.500 ;
        RECT 445.650 627.600 447.450 633.600 ;
        RECT 454.050 627.600 455.850 639.600 ;
        RECT 458.550 656.400 460.350 662.400 ;
        RECT 466.650 659.400 468.450 662.400 ;
        RECT 474.450 659.400 476.250 662.400 ;
        RECT 482.250 660.300 484.050 662.400 ;
        RECT 482.250 659.400 486.000 660.300 ;
        RECT 466.650 658.500 467.700 659.400 ;
        RECT 463.950 657.300 467.700 658.500 ;
        RECT 475.200 658.500 476.250 659.400 ;
        RECT 484.950 658.500 486.000 659.400 ;
        RECT 475.200 657.450 480.150 658.500 ;
        RECT 463.950 656.400 466.050 657.300 ;
        RECT 478.350 656.700 480.150 657.450 ;
        RECT 458.550 649.050 459.750 656.400 ;
        RECT 481.650 655.800 483.450 657.600 ;
        RECT 484.950 656.400 487.050 658.500 ;
        RECT 490.050 656.400 491.850 662.400 ;
        RECT 502.800 656.400 504.600 662.400 ;
        RECT 471.150 654.000 472.950 654.600 ;
        RECT 482.100 654.000 483.150 655.800 ;
        RECT 471.150 652.800 483.150 654.000 ;
        RECT 458.550 647.250 464.850 649.050 ;
        RECT 458.550 646.950 463.050 647.250 ;
        RECT 458.550 639.600 459.750 646.950 ;
        RECT 460.950 641.400 462.750 643.200 ;
        RECT 461.850 640.200 466.050 641.400 ;
        RECT 471.150 640.200 472.050 652.800 ;
        RECT 482.100 651.600 489.000 652.800 ;
        RECT 482.100 651.000 483.900 651.600 ;
        RECT 488.100 650.850 489.000 651.600 ;
        RECT 485.100 649.800 486.900 650.400 ;
        RECT 478.950 648.600 486.900 649.800 ;
        RECT 488.100 649.050 489.900 650.850 ;
        RECT 478.950 646.950 481.050 648.600 ;
        RECT 487.950 646.950 490.050 649.050 ;
        RECT 480.750 641.700 482.550 642.000 ;
        RECT 490.950 641.700 491.850 656.400 ;
        RECT 503.400 654.300 504.600 656.400 ;
        RECT 505.800 657.300 507.600 662.400 ;
        RECT 511.800 657.300 513.600 662.400 ;
        RECT 505.800 655.950 513.600 657.300 ;
        RECT 524.400 657.300 526.200 662.400 ;
        RECT 530.400 657.300 532.200 662.400 ;
        RECT 524.400 655.950 532.200 657.300 ;
        RECT 533.400 656.400 535.200 662.400 ;
        RECT 550.800 659.400 552.600 662.400 ;
        RECT 533.400 654.300 534.600 656.400 ;
        RECT 503.400 653.250 507.150 654.300 ;
        RECT 503.100 649.050 504.900 650.850 ;
        RECT 505.950 649.050 507.150 653.250 ;
        RECT 530.850 653.250 534.600 654.300 ;
        RECT 509.100 649.050 510.900 650.850 ;
        RECT 527.100 649.050 528.900 650.850 ;
        RECT 530.850 649.050 532.050 653.250 ;
        RECT 533.100 649.050 534.900 650.850 ;
        RECT 551.400 649.050 552.600 659.400 ;
        RECT 557.550 656.400 559.350 662.400 ;
        RECT 565.650 659.400 567.450 662.400 ;
        RECT 573.450 659.400 575.250 662.400 ;
        RECT 581.250 660.300 583.050 662.400 ;
        RECT 581.250 659.400 585.000 660.300 ;
        RECT 565.650 658.500 566.700 659.400 ;
        RECT 562.950 657.300 566.700 658.500 ;
        RECT 574.200 658.500 575.250 659.400 ;
        RECT 583.950 658.500 585.000 659.400 ;
        RECT 574.200 657.450 579.150 658.500 ;
        RECT 562.950 656.400 565.050 657.300 ;
        RECT 577.350 656.700 579.150 657.450 ;
        RECT 557.550 649.050 558.750 656.400 ;
        RECT 580.650 655.800 582.450 657.600 ;
        RECT 583.950 656.400 586.050 658.500 ;
        RECT 589.050 656.400 590.850 662.400 ;
        RECT 604.800 656.400 606.600 662.400 ;
        RECT 570.150 654.000 571.950 654.600 ;
        RECT 581.100 654.000 582.150 655.800 ;
        RECT 570.150 652.800 582.150 654.000 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 508.950 646.950 511.050 649.050 ;
        RECT 511.950 646.950 514.050 649.050 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 526.950 646.950 529.050 649.050 ;
        RECT 529.950 646.950 532.050 649.050 ;
        RECT 532.950 646.950 535.050 649.050 ;
        RECT 550.950 646.950 553.050 649.050 ;
        RECT 553.950 646.950 556.050 649.050 ;
        RECT 557.550 647.250 563.850 649.050 ;
        RECT 557.550 646.950 562.050 647.250 ;
        RECT 480.750 641.100 491.850 641.700 ;
        RECT 458.550 627.600 460.350 639.600 ;
        RECT 463.950 639.300 466.050 640.200 ;
        RECT 466.950 639.300 472.050 640.200 ;
        RECT 474.150 640.500 491.850 641.100 ;
        RECT 474.150 640.200 482.550 640.500 ;
        RECT 466.950 638.400 467.850 639.300 ;
        RECT 465.150 636.600 467.850 638.400 ;
        RECT 468.750 638.100 470.550 638.400 ;
        RECT 474.150 638.100 475.050 640.200 ;
        RECT 490.950 639.600 491.850 640.500 ;
        RECT 468.750 637.200 475.050 638.100 ;
        RECT 475.950 638.700 477.750 639.300 ;
        RECT 475.950 637.500 483.450 638.700 ;
        RECT 468.750 636.600 470.550 637.200 ;
        RECT 482.250 636.600 483.450 637.500 ;
        RECT 463.950 633.600 467.850 635.700 ;
        RECT 472.950 635.550 474.750 636.300 ;
        RECT 477.750 635.550 479.550 636.300 ;
        RECT 472.950 634.500 479.550 635.550 ;
        RECT 482.250 634.500 487.050 636.600 ;
        RECT 466.050 627.600 467.850 633.600 ;
        RECT 473.850 627.600 475.650 634.500 ;
        RECT 482.250 633.600 483.450 634.500 ;
        RECT 481.650 627.600 483.450 633.600 ;
        RECT 490.050 627.600 491.850 639.600 ;
        RECT 506.850 633.600 508.050 646.950 ;
        RECT 512.100 645.150 513.900 646.950 ;
        RECT 524.100 645.150 525.900 646.950 ;
        RECT 529.950 633.600 531.150 646.950 ;
        RECT 551.400 633.600 552.600 646.950 ;
        RECT 554.100 645.150 555.900 646.950 ;
        RECT 506.400 627.600 508.200 633.600 ;
        RECT 529.800 627.600 531.600 633.600 ;
        RECT 550.800 627.600 552.600 633.600 ;
        RECT 557.550 639.600 558.750 646.950 ;
        RECT 559.950 641.400 561.750 643.200 ;
        RECT 560.850 640.200 565.050 641.400 ;
        RECT 570.150 640.200 571.050 652.800 ;
        RECT 581.100 651.600 588.000 652.800 ;
        RECT 581.100 651.000 582.900 651.600 ;
        RECT 587.100 650.850 588.000 651.600 ;
        RECT 584.100 649.800 585.900 650.400 ;
        RECT 577.950 648.600 585.900 649.800 ;
        RECT 587.100 649.050 588.900 650.850 ;
        RECT 577.950 646.950 580.050 648.600 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 579.750 641.700 581.550 642.000 ;
        RECT 589.950 641.700 590.850 656.400 ;
        RECT 605.400 654.300 606.600 656.400 ;
        RECT 607.800 657.300 609.600 662.400 ;
        RECT 613.800 657.300 615.600 662.400 ;
        RECT 607.800 655.950 615.600 657.300 ;
        RECT 626.400 659.400 628.200 662.400 ;
        RECT 605.400 653.250 609.150 654.300 ;
        RECT 605.100 649.050 606.900 650.850 ;
        RECT 607.950 649.050 609.150 653.250 ;
        RECT 611.100 649.050 612.900 650.850 ;
        RECT 626.400 649.050 627.600 659.400 ;
        RECT 638.400 656.400 640.200 662.400 ;
        RECT 645.600 657.000 647.400 662.400 ;
        RECT 638.400 655.500 639.900 656.400 ;
        RECT 638.400 654.000 642.750 655.500 ;
        RECT 640.650 653.400 642.750 654.000 ;
        RECT 646.350 654.900 647.400 657.000 ;
        RECT 653.400 656.400 655.200 662.400 ;
        RECT 650.700 655.200 655.200 656.400 ;
        RECT 668.400 657.300 670.200 662.400 ;
        RECT 674.400 657.300 676.200 662.400 ;
        RECT 668.400 655.950 676.200 657.300 ;
        RECT 677.400 656.400 679.200 662.400 ;
        RECT 643.650 651.900 645.450 653.700 ;
        RECT 646.350 652.800 649.500 654.900 ;
        RECT 650.700 653.100 652.800 655.200 ;
        RECT 677.400 654.300 678.600 656.400 ;
        RECT 688.950 655.950 691.050 658.050 ;
        RECT 698.700 657.600 700.500 662.400 ;
        RECT 722.700 657.600 724.500 662.400 ;
        RECT 695.400 656.400 700.500 657.600 ;
        RECT 719.400 656.400 724.500 657.600 ;
        RECT 740.400 659.400 742.200 662.400 ;
        RECT 674.850 653.250 678.600 654.300 ;
        RECT 643.200 651.000 645.300 651.900 ;
        RECT 638.700 649.800 645.300 651.000 ;
        RECT 638.700 649.200 640.500 649.800 ;
        RECT 604.950 646.950 607.050 649.050 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 610.950 646.950 613.050 649.050 ;
        RECT 613.950 646.950 616.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 638.400 647.100 640.500 649.200 ;
        RECT 579.750 641.100 590.850 641.700 ;
        RECT 557.550 627.600 559.350 639.600 ;
        RECT 562.950 639.300 565.050 640.200 ;
        RECT 565.950 639.300 571.050 640.200 ;
        RECT 573.150 640.500 590.850 641.100 ;
        RECT 573.150 640.200 581.550 640.500 ;
        RECT 565.950 638.400 566.850 639.300 ;
        RECT 564.150 636.600 566.850 638.400 ;
        RECT 567.750 638.100 569.550 638.400 ;
        RECT 573.150 638.100 574.050 640.200 ;
        RECT 589.950 639.600 590.850 640.500 ;
        RECT 567.750 637.200 574.050 638.100 ;
        RECT 574.950 638.700 576.750 639.300 ;
        RECT 574.950 637.500 582.450 638.700 ;
        RECT 567.750 636.600 569.550 637.200 ;
        RECT 581.250 636.600 582.450 637.500 ;
        RECT 562.950 633.600 566.850 635.700 ;
        RECT 571.950 635.550 573.750 636.300 ;
        RECT 576.750 635.550 578.550 636.300 ;
        RECT 571.950 634.500 578.550 635.550 ;
        RECT 581.250 634.500 586.050 636.600 ;
        RECT 565.050 627.600 566.850 633.600 ;
        RECT 572.850 627.600 574.650 634.500 ;
        RECT 581.250 633.600 582.450 634.500 ;
        RECT 580.650 627.600 582.450 633.600 ;
        RECT 589.050 627.600 590.850 639.600 ;
        RECT 608.850 633.600 610.050 646.950 ;
        RECT 614.100 645.150 615.900 646.950 ;
        RECT 623.100 645.150 624.900 646.950 ;
        RECT 626.400 633.600 627.600 646.950 ;
        RECT 643.200 646.800 645.300 648.900 ;
        RECT 643.200 645.000 645.000 646.800 ;
        RECT 646.350 646.200 647.250 652.800 ;
        RECT 664.950 651.450 667.050 652.050 ;
        RECT 648.150 648.900 650.250 651.000 ;
        RECT 659.550 650.550 667.050 651.450 ;
        RECT 648.300 647.100 650.100 648.900 ;
        RECT 652.950 647.100 655.050 649.200 ;
        RECT 646.350 644.700 649.500 646.200 ;
        RECT 653.100 645.450 654.900 647.100 ;
        RECT 659.550 645.450 660.450 650.550 ;
        RECT 664.950 649.950 667.050 650.550 ;
        RECT 671.100 649.050 672.900 650.850 ;
        RECT 674.850 649.050 676.050 653.250 ;
        RECT 682.950 651.450 685.050 651.900 ;
        RECT 689.550 651.450 690.450 655.950 ;
        RECT 677.100 649.050 678.900 650.850 ;
        RECT 682.950 650.550 690.450 651.450 ;
        RECT 682.950 649.800 685.050 650.550 ;
        RECT 695.400 649.050 696.300 656.400 ;
        RECT 700.950 654.450 703.050 655.050 ;
        RECT 715.950 654.450 718.050 655.050 ;
        RECT 700.950 653.550 718.050 654.450 ;
        RECT 700.950 652.950 703.050 653.550 ;
        RECT 715.950 652.950 718.050 653.550 ;
        RECT 706.950 651.450 709.050 652.050 ;
        RECT 698.100 649.050 699.900 650.850 ;
        RECT 704.100 649.050 705.900 650.850 ;
        RECT 706.950 650.550 714.450 651.450 ;
        RECT 706.950 649.950 709.050 650.550 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 670.950 646.950 673.050 649.050 ;
        RECT 673.950 646.950 676.050 649.050 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 694.950 646.950 697.050 649.050 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 703.950 646.950 706.050 649.050 ;
        RECT 653.100 645.300 660.450 645.450 ;
        RECT 647.400 644.100 649.500 644.700 ;
        RECT 653.550 644.550 660.450 645.300 ;
        RECT 668.100 645.150 669.900 646.950 ;
        RECT 644.700 641.700 646.500 643.800 ;
        RECT 641.100 640.800 646.500 641.700 ;
        RECT 641.100 639.900 643.200 640.800 ;
        RECT 638.400 638.700 643.200 639.900 ;
        RECT 648.000 639.600 649.200 644.100 ;
        RECT 645.900 638.700 649.200 639.600 ;
        RECT 650.100 639.600 652.200 640.500 ;
        RECT 608.400 627.600 610.200 633.600 ;
        RECT 626.400 627.600 628.200 633.600 ;
        RECT 638.400 627.600 640.200 638.700 ;
        RECT 645.900 627.600 647.700 638.700 ;
        RECT 650.100 638.400 655.200 639.600 ;
        RECT 653.400 627.600 655.200 638.400 ;
        RECT 673.950 633.600 675.150 646.950 ;
        RECT 676.950 642.450 679.050 643.050 ;
        RECT 688.950 642.450 691.050 643.050 ;
        RECT 676.950 641.550 691.050 642.450 ;
        RECT 676.950 640.950 679.050 641.550 ;
        RECT 688.950 640.950 691.050 641.550 ;
        RECT 695.400 639.600 696.300 646.950 ;
        RECT 701.100 645.150 702.900 646.950 ;
        RECT 713.550 646.050 714.450 650.550 ;
        RECT 719.400 649.050 720.300 656.400 ;
        RECT 722.100 649.050 723.900 650.850 ;
        RECT 728.100 649.050 729.900 650.850 ;
        RECT 740.400 649.050 741.600 659.400 ;
        RECT 754.800 656.400 756.600 662.400 ;
        RECT 755.400 654.300 756.600 656.400 ;
        RECT 757.800 657.300 759.600 662.400 ;
        RECT 763.800 657.300 765.600 662.400 ;
        RECT 778.800 659.400 780.600 662.400 ;
        RECT 796.800 659.400 798.600 662.400 ;
        RECT 757.800 655.950 765.600 657.300 ;
        RECT 755.400 653.250 759.150 654.300 ;
        RECT 751.950 651.450 754.050 652.050 ;
        RECT 746.550 650.550 754.050 651.450 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 739.950 646.950 742.050 649.050 ;
        RECT 713.550 644.550 718.050 646.050 ;
        RECT 714.000 643.950 718.050 644.550 ;
        RECT 697.950 642.450 700.050 643.050 ;
        RECT 712.950 642.450 715.050 643.050 ;
        RECT 697.950 641.550 715.050 642.450 ;
        RECT 697.950 640.950 700.050 641.550 ;
        RECT 712.950 640.950 715.050 641.550 ;
        RECT 719.400 639.600 720.300 646.950 ;
        RECT 725.100 645.150 726.900 646.950 ;
        RECT 737.100 645.150 738.900 646.950 ;
        RECT 673.800 627.600 675.600 633.600 ;
        RECT 694.800 627.600 696.600 639.600 ;
        RECT 697.800 638.700 705.600 639.600 ;
        RECT 697.800 627.600 699.600 638.700 ;
        RECT 703.800 627.600 705.600 638.700 ;
        RECT 718.800 627.600 720.600 639.600 ;
        RECT 721.800 638.700 729.600 639.600 ;
        RECT 721.800 627.600 723.600 638.700 ;
        RECT 727.800 627.600 729.600 638.700 ;
        RECT 740.400 633.600 741.600 646.950 ;
        RECT 746.550 646.050 747.450 650.550 ;
        RECT 751.950 649.950 754.050 650.550 ;
        RECT 755.100 649.050 756.900 650.850 ;
        RECT 757.950 649.050 759.150 653.250 ;
        RECT 766.950 651.450 769.050 652.050 ;
        RECT 761.100 649.050 762.900 650.850 ;
        RECT 766.950 650.550 774.450 651.450 ;
        RECT 766.950 649.950 769.050 650.550 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 757.950 646.950 760.050 649.050 ;
        RECT 760.950 646.950 763.050 649.050 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 742.950 644.550 747.450 646.050 ;
        RECT 742.950 643.950 747.000 644.550 ;
        RECT 758.850 633.600 760.050 646.950 ;
        RECT 764.100 645.150 765.900 646.950 ;
        RECT 773.550 646.050 774.450 650.550 ;
        RECT 779.400 649.050 780.600 659.400 ;
        RECT 781.950 654.450 784.050 655.050 ;
        RECT 793.950 654.450 796.050 655.050 ;
        RECT 781.950 653.550 796.050 654.450 ;
        RECT 781.950 652.950 784.050 653.550 ;
        RECT 793.950 652.950 796.050 653.550 ;
        RECT 797.400 649.050 798.600 659.400 ;
        RECT 812.400 657.300 814.200 662.400 ;
        RECT 818.400 657.300 820.200 662.400 ;
        RECT 812.400 655.950 820.200 657.300 ;
        RECT 821.400 656.400 823.200 662.400 ;
        RECT 841.200 656.400 843.000 662.400 ;
        RECT 821.400 654.300 822.600 656.400 ;
        RECT 818.850 653.250 822.600 654.300 ;
        RECT 802.950 651.450 807.000 652.050 ;
        RECT 802.950 649.950 807.450 651.450 ;
        RECT 778.950 646.950 781.050 649.050 ;
        RECT 781.950 646.950 784.050 649.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 799.950 646.950 802.050 649.050 ;
        RECT 773.550 644.550 778.050 646.050 ;
        RECT 774.000 643.950 778.050 644.550 ;
        RECT 779.400 633.600 780.600 646.950 ;
        RECT 782.100 645.150 783.900 646.950 ;
        RECT 797.400 633.600 798.600 646.950 ;
        RECT 800.100 645.150 801.900 646.950 ;
        RECT 806.550 646.050 807.450 649.950 ;
        RECT 815.100 649.050 816.900 650.850 ;
        RECT 818.850 649.050 820.050 653.250 ;
        RECT 826.950 651.450 829.050 652.050 ;
        RECT 832.950 651.450 835.050 652.050 ;
        RECT 821.100 649.050 822.900 650.850 ;
        RECT 826.950 650.550 835.050 651.450 ;
        RECT 826.950 649.950 829.050 650.550 ;
        RECT 832.950 649.950 835.050 650.550 ;
        RECT 836.100 649.050 837.900 650.850 ;
        RECT 841.950 649.050 843.000 656.400 ;
        RECT 860.400 657.300 862.200 662.400 ;
        RECT 866.400 657.300 868.200 662.400 ;
        RECT 860.400 655.950 868.200 657.300 ;
        RECT 869.400 656.400 871.200 662.400 ;
        RECT 869.400 654.300 870.600 656.400 ;
        RECT 887.400 655.200 889.200 662.400 ;
        RECT 905.400 659.400 907.200 662.400 ;
        RECT 887.400 654.300 891.600 655.200 ;
        RECT 866.850 653.250 870.600 654.300 ;
        RECT 855.000 651.450 859.050 652.050 ;
        RECT 848.100 649.050 849.900 650.850 ;
        RECT 854.550 649.950 859.050 651.450 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 838.950 646.950 841.050 649.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 844.950 646.950 847.050 649.050 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 802.950 644.550 807.450 646.050 ;
        RECT 812.100 645.150 813.900 646.950 ;
        RECT 802.950 643.950 807.000 644.550 ;
        RECT 817.950 633.600 819.150 646.950 ;
        RECT 839.100 645.150 840.900 646.950 ;
        RECT 842.100 641.400 843.000 646.950 ;
        RECT 845.100 645.150 846.900 646.950 ;
        RECT 854.550 645.450 855.450 649.950 ;
        RECT 863.100 649.050 864.900 650.850 ;
        RECT 866.850 649.050 868.050 653.250 ;
        RECT 871.950 651.450 876.000 652.050 ;
        RECT 869.100 649.050 870.900 650.850 ;
        RECT 871.950 649.950 876.450 651.450 ;
        RECT 859.950 646.950 862.050 649.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 854.550 644.550 858.450 645.450 ;
        RECT 860.100 645.150 861.900 646.950 ;
        RECT 857.550 643.050 858.450 644.550 ;
        RECT 857.550 641.550 862.050 643.050 ;
        RECT 842.100 640.500 847.200 641.400 ;
        RECT 858.000 640.950 862.050 641.550 ;
        RECT 836.400 638.400 844.200 639.300 ;
        RECT 740.400 627.600 742.200 633.600 ;
        RECT 758.400 627.600 760.200 633.600 ;
        RECT 778.800 627.600 780.600 633.600 ;
        RECT 796.800 627.600 798.600 633.600 ;
        RECT 817.800 627.600 819.600 633.600 ;
        RECT 836.400 627.600 838.200 638.400 ;
        RECT 842.400 628.500 844.200 638.400 ;
        RECT 845.400 629.400 847.200 640.500 ;
        RECT 848.400 628.500 850.200 639.600 ;
        RECT 865.950 633.600 867.150 646.950 ;
        RECT 875.550 645.450 876.450 649.950 ;
        RECT 887.100 649.050 888.900 650.850 ;
        RECT 890.400 649.050 891.600 654.300 ;
        RECT 893.100 649.050 894.900 650.850 ;
        RECT 905.400 649.050 906.600 659.400 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 901.950 646.950 904.050 649.050 ;
        RECT 904.950 646.950 907.050 649.050 ;
        RECT 872.550 644.550 876.450 645.450 ;
        RECT 872.550 643.050 873.450 644.550 ;
        RECT 868.950 641.550 873.450 643.050 ;
        RECT 868.950 640.950 873.000 641.550 ;
        RECT 890.400 633.600 891.600 646.950 ;
        RECT 902.100 645.150 903.900 646.950 ;
        RECT 842.400 627.600 850.200 628.500 ;
        RECT 865.800 627.600 867.600 633.600 ;
        RECT 889.800 627.600 891.600 633.600 ;
        RECT 905.400 633.600 906.600 646.950 ;
        RECT 905.400 627.600 907.200 633.600 ;
        RECT 13.800 611.400 15.600 623.400 ;
        RECT 16.800 612.300 18.600 623.400 ;
        RECT 22.800 612.300 24.600 623.400 ;
        RECT 38.400 617.400 40.200 623.400 ;
        RECT 38.700 617.100 40.200 617.400 ;
        RECT 44.400 617.400 46.200 623.400 ;
        RECT 44.400 617.100 45.300 617.400 ;
        RECT 38.700 616.200 45.300 617.100 ;
        RECT 16.800 611.400 24.600 612.300 ;
        RECT 14.400 604.050 15.300 611.400 ;
        RECT 28.950 609.450 31.050 610.050 ;
        RECT 40.950 609.450 43.050 610.050 ;
        RECT 28.950 608.550 43.050 609.450 ;
        RECT 28.950 607.950 31.050 608.550 ;
        RECT 40.950 607.950 43.050 608.550 ;
        RECT 20.100 604.050 21.900 605.850 ;
        RECT 38.100 604.050 39.900 605.850 ;
        RECT 44.400 604.050 45.300 616.200 ;
        RECT 61.500 612.600 63.300 623.400 ;
        RECT 83.400 617.400 85.200 623.400 ;
        RECT 59.700 611.400 63.300 612.600 ;
        RECT 56.100 604.050 57.900 605.850 ;
        RECT 59.700 604.050 60.600 611.400 ;
        RECT 62.100 604.050 63.900 605.850 ;
        RECT 83.850 604.050 85.050 617.400 ;
        RECT 103.500 612.600 105.300 623.400 ;
        RECT 101.700 611.400 105.300 612.600 ;
        RECT 116.400 612.300 118.200 623.400 ;
        RECT 123.900 612.300 125.700 623.400 ;
        RECT 131.400 612.600 133.200 623.400 ;
        RECT 89.100 604.050 90.900 605.850 ;
        RECT 98.100 604.050 99.900 605.850 ;
        RECT 101.700 604.050 102.600 611.400 ;
        RECT 116.400 611.100 121.200 612.300 ;
        RECT 123.900 611.400 127.200 612.300 ;
        RECT 119.100 610.200 121.200 611.100 ;
        RECT 119.100 609.300 124.500 610.200 ;
        RECT 122.700 607.200 124.500 609.300 ;
        RECT 126.000 606.900 127.200 611.400 ;
        RECT 128.100 611.400 133.200 612.600 ;
        RECT 143.400 612.300 145.200 623.400 ;
        RECT 143.400 611.400 147.900 612.300 ;
        RECT 150.900 611.400 152.700 623.400 ;
        RECT 158.400 612.600 160.200 623.400 ;
        RECT 176.400 617.400 178.200 623.400 ;
        RECT 176.700 617.100 178.200 617.400 ;
        RECT 182.400 617.400 184.200 623.400 ;
        RECT 202.800 617.400 204.600 623.400 ;
        RECT 182.400 617.100 183.300 617.400 ;
        RECT 176.700 616.200 183.300 617.100 ;
        RECT 128.100 610.500 130.200 611.400 ;
        RECT 145.800 609.300 147.900 611.400 ;
        RECT 151.500 609.900 152.700 611.400 ;
        RECT 155.400 611.400 160.200 612.600 ;
        RECT 155.400 610.500 157.500 611.400 ;
        RECT 151.500 609.000 153.000 609.900 ;
        RECT 149.100 607.500 151.200 607.800 ;
        RECT 125.400 606.300 127.500 606.900 ;
        RECT 132.000 606.450 136.050 607.050 ;
        RECT 104.100 604.050 105.900 605.850 ;
        RECT 121.200 604.200 123.000 606.000 ;
        RECT 124.350 604.800 127.500 606.300 ;
        RECT 131.550 605.700 136.050 606.450 ;
        RECT 147.300 605.700 151.200 607.500 ;
        RECT 152.100 606.900 153.000 609.000 ;
        RECT 131.100 604.950 136.050 605.700 ;
        RECT 13.950 601.950 16.050 604.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 19.950 601.950 22.050 604.050 ;
        RECT 22.950 601.950 25.050 604.050 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 43.950 601.950 46.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 58.950 601.950 61.050 604.050 ;
        RECT 61.950 601.950 64.050 604.050 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 85.950 601.950 88.050 604.050 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 100.950 601.950 103.050 604.050 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 14.400 594.600 15.300 601.950 ;
        RECT 17.100 600.150 18.900 601.950 ;
        RECT 23.100 600.150 24.900 601.950 ;
        RECT 35.100 600.150 36.900 601.950 ;
        RECT 41.100 600.150 42.900 601.950 ;
        RECT 44.400 598.200 45.300 601.950 ;
        RECT 42.000 597.000 45.300 598.200 ;
        RECT 14.400 593.400 19.500 594.600 ;
        RECT 17.700 588.600 19.500 593.400 ;
        RECT 42.000 588.600 43.800 597.000 ;
        RECT 59.700 591.600 60.600 601.950 ;
        RECT 67.950 600.450 70.050 601.050 ;
        RECT 76.950 600.450 79.050 601.050 ;
        RECT 67.950 599.550 79.050 600.450 ;
        RECT 80.100 600.150 81.900 601.950 ;
        RECT 67.950 598.950 70.050 599.550 ;
        RECT 76.950 598.950 79.050 599.550 ;
        RECT 82.950 597.750 84.150 601.950 ;
        RECT 86.100 600.150 87.900 601.950 ;
        RECT 80.400 596.700 84.150 597.750 ;
        RECT 80.400 594.600 81.600 596.700 ;
        RECT 59.400 588.600 61.200 591.600 ;
        RECT 79.800 588.600 81.600 594.600 ;
        RECT 82.800 593.700 90.600 595.050 ;
        RECT 82.800 588.600 84.600 593.700 ;
        RECT 88.800 588.600 90.600 593.700 ;
        RECT 101.700 591.600 102.600 601.950 ;
        RECT 116.400 601.800 118.500 603.900 ;
        RECT 121.200 602.100 123.300 604.200 ;
        RECT 116.700 601.200 118.500 601.800 ;
        RECT 116.700 600.000 123.300 601.200 ;
        RECT 121.200 599.100 123.300 600.000 ;
        RECT 118.650 597.000 120.750 597.600 ;
        RECT 121.650 597.300 123.450 599.100 ;
        RECT 124.350 598.200 125.250 604.800 ;
        RECT 131.100 603.900 132.900 604.950 ;
        RECT 152.100 604.800 154.200 606.900 ;
        RECT 143.400 603.900 145.500 604.050 ;
        RECT 148.500 603.900 150.300 604.500 ;
        RECT 126.300 602.100 128.100 603.900 ;
        RECT 126.150 600.000 128.250 602.100 ;
        RECT 130.950 601.800 133.050 603.900 ;
        RECT 143.400 602.700 150.300 603.900 ;
        RECT 151.200 603.900 153.600 604.800 ;
        RECT 158.100 604.050 159.900 605.850 ;
        RECT 176.100 604.050 177.900 605.850 ;
        RECT 182.400 604.050 183.300 616.200 ;
        RECT 203.400 604.050 204.600 617.400 ;
        RECT 220.800 611.400 222.600 623.400 ;
        RECT 226.800 617.400 228.600 623.400 ;
        RECT 221.400 604.050 222.300 611.400 ;
        RECT 224.100 604.050 225.900 605.850 ;
        RECT 143.400 601.950 145.500 602.700 ;
        RECT 143.400 600.150 145.200 601.950 ;
        RECT 148.500 599.400 150.300 601.200 ;
        RECT 116.400 595.500 120.750 597.000 ;
        RECT 124.350 596.100 127.500 598.200 ;
        RECT 116.400 594.600 117.900 595.500 ;
        RECT 101.400 588.600 103.200 591.600 ;
        RECT 116.400 588.600 118.200 594.600 ;
        RECT 124.350 594.000 125.400 596.100 ;
        RECT 128.700 595.800 130.800 597.900 ;
        RECT 148.200 597.300 150.300 599.400 ;
        RECT 144.000 596.400 150.300 597.300 ;
        RECT 151.200 598.200 152.250 603.900 ;
        RECT 157.950 603.450 160.050 604.050 ;
        RECT 162.000 603.450 166.050 604.050 ;
        RECT 153.600 601.200 155.400 603.000 ;
        RECT 157.950 602.550 166.050 603.450 ;
        RECT 157.950 601.950 160.050 602.550 ;
        RECT 162.000 601.950 166.050 602.550 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 175.950 601.950 178.050 604.050 ;
        RECT 178.950 601.950 181.050 604.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 202.950 601.950 205.050 604.050 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 153.150 599.100 155.250 601.200 ;
        RECT 173.100 600.150 174.900 601.950 ;
        RECT 179.100 600.150 180.900 601.950 ;
        RECT 182.400 598.200 183.300 601.950 ;
        RECT 200.100 600.150 201.900 601.950 ;
        RECT 128.700 594.600 133.200 595.800 ;
        RECT 144.000 594.600 145.200 596.400 ;
        RECT 151.200 596.100 154.200 598.200 ;
        RECT 180.000 597.000 183.300 598.200 ;
        RECT 151.200 594.600 152.400 596.100 ;
        RECT 155.400 595.500 157.500 596.700 ;
        RECT 155.400 594.600 160.200 595.500 ;
        RECT 123.600 588.600 125.400 594.000 ;
        RECT 131.400 588.600 133.200 594.600 ;
        RECT 143.400 588.600 145.200 594.600 ;
        RECT 150.900 588.600 152.700 594.600 ;
        RECT 158.400 588.600 160.200 594.600 ;
        RECT 180.000 588.600 181.800 597.000 ;
        RECT 203.400 596.700 204.600 601.950 ;
        RECT 206.100 600.150 207.900 601.950 ;
        RECT 200.400 595.800 204.600 596.700 ;
        RECT 200.400 588.600 202.200 595.800 ;
        RECT 221.400 594.600 222.300 601.950 ;
        RECT 227.700 597.300 228.600 617.400 ;
        RECT 245.400 617.400 247.200 623.400 ;
        RECT 262.800 617.400 264.600 623.400 ;
        RECT 237.000 606.450 241.050 607.050 ;
        RECT 236.550 604.950 241.050 606.450 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 230.100 600.150 231.900 601.950 ;
        RECT 236.550 601.050 237.450 604.950 ;
        RECT 242.100 604.050 243.900 605.850 ;
        RECT 245.400 604.050 246.600 617.400 ;
        RECT 263.700 617.100 264.600 617.400 ;
        RECT 268.800 617.400 270.600 623.400 ;
        RECT 287.400 617.400 289.200 623.400 ;
        RECT 305.400 617.400 307.200 623.400 ;
        RECT 268.800 617.100 270.300 617.400 ;
        RECT 263.700 616.200 270.300 617.100 ;
        RECT 247.950 606.450 252.000 607.050 ;
        RECT 247.950 604.950 252.450 606.450 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 236.550 599.550 241.050 601.050 ;
        RECT 237.000 598.950 241.050 599.550 ;
        RECT 224.100 596.400 231.600 597.300 ;
        RECT 224.100 595.500 225.900 596.400 ;
        RECT 221.400 592.800 224.100 594.600 ;
        RECT 222.300 588.600 224.100 592.800 ;
        RECT 229.800 588.600 231.600 596.400 ;
        RECT 245.400 591.600 246.600 601.950 ;
        RECT 251.550 600.450 252.450 604.950 ;
        RECT 263.700 604.050 264.600 616.200 ;
        RECT 265.950 609.450 268.050 610.050 ;
        RECT 277.950 609.450 280.050 610.050 ;
        RECT 265.950 608.550 280.050 609.450 ;
        RECT 265.950 607.950 268.050 608.550 ;
        RECT 277.950 607.950 280.050 608.550 ;
        RECT 279.000 606.450 283.050 607.050 ;
        RECT 269.100 604.050 270.900 605.850 ;
        RECT 278.550 604.950 283.050 606.450 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 259.950 600.450 262.050 601.050 ;
        RECT 251.550 599.550 262.050 600.450 ;
        RECT 259.950 598.950 262.050 599.550 ;
        RECT 263.700 598.200 264.600 601.950 ;
        RECT 266.100 600.150 267.900 601.950 ;
        RECT 272.100 600.150 273.900 601.950 ;
        RECT 278.550 601.050 279.450 604.950 ;
        RECT 284.100 604.050 285.900 605.850 ;
        RECT 287.400 604.050 288.600 617.400 ;
        RECT 292.950 609.450 295.050 610.050 ;
        RECT 301.950 609.450 304.050 610.050 ;
        RECT 292.950 608.550 304.050 609.450 ;
        RECT 292.950 607.950 295.050 608.550 ;
        RECT 301.950 607.950 304.050 608.550 ;
        RECT 297.000 606.450 301.050 607.050 ;
        RECT 296.550 604.950 301.050 606.450 ;
        RECT 283.950 601.950 286.050 604.050 ;
        RECT 286.950 601.950 289.050 604.050 ;
        RECT 274.950 599.550 279.450 601.050 ;
        RECT 274.950 598.950 279.000 599.550 ;
        RECT 263.700 597.000 267.000 598.200 ;
        RECT 245.400 588.600 247.200 591.600 ;
        RECT 265.200 588.600 267.000 597.000 ;
        RECT 287.400 591.600 288.600 601.950 ;
        RECT 296.550 598.050 297.450 604.950 ;
        RECT 305.400 604.050 306.600 617.400 ;
        RECT 326.400 611.400 328.200 623.400 ;
        RECT 338.400 612.600 340.200 623.400 ;
        RECT 344.400 622.500 352.200 623.400 ;
        RECT 344.400 612.600 346.200 622.500 ;
        RECT 338.400 611.700 346.200 612.600 ;
        RECT 319.950 606.450 322.050 607.050 ;
        RECT 314.550 605.550 322.050 606.450 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 304.950 601.950 307.050 604.050 ;
        RECT 307.950 601.950 310.050 604.050 ;
        RECT 302.100 600.150 303.900 601.950 ;
        RECT 292.950 596.550 297.450 598.050 ;
        RECT 305.400 596.700 306.600 601.950 ;
        RECT 308.100 600.150 309.900 601.950 ;
        RECT 314.550 601.050 315.450 605.550 ;
        RECT 319.950 604.950 322.050 605.550 ;
        RECT 326.400 604.050 327.600 611.400 ;
        RECT 347.400 610.500 349.200 621.600 ;
        RECT 350.400 611.400 352.200 622.500 ;
        RECT 368.400 617.400 370.200 623.400 ;
        RECT 386.400 617.400 388.200 623.400 ;
        RECT 344.100 609.600 349.200 610.500 ;
        RECT 341.100 604.050 342.900 605.850 ;
        RECT 344.100 604.050 345.000 609.600 ;
        RECT 352.950 609.450 355.050 610.050 ;
        RECT 358.950 609.450 361.050 610.050 ;
        RECT 352.950 608.550 361.050 609.450 ;
        RECT 352.950 607.950 355.050 608.550 ;
        RECT 358.950 607.950 361.050 608.550 ;
        RECT 347.100 604.050 348.900 605.850 ;
        RECT 368.400 604.050 369.600 617.400 ;
        RECT 386.400 610.500 387.600 617.400 ;
        RECT 392.400 611.400 394.200 623.400 ;
        RECT 409.800 617.400 411.600 623.400 ;
        RECT 397.950 613.950 403.050 616.050 ;
        RECT 386.400 609.600 392.100 610.500 ;
        RECT 390.150 608.700 392.100 609.600 ;
        RECT 386.100 604.050 387.900 605.850 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 337.950 601.950 340.050 604.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 310.950 599.550 315.450 601.050 ;
        RECT 323.100 600.150 324.900 601.950 ;
        RECT 310.950 598.950 315.000 599.550 ;
        RECT 292.950 595.950 297.000 596.550 ;
        RECT 305.400 595.800 309.600 596.700 ;
        RECT 287.400 588.600 289.200 591.600 ;
        RECT 307.800 588.600 309.600 595.800 ;
        RECT 326.400 594.600 327.600 601.950 ;
        RECT 338.100 600.150 339.900 601.950 ;
        RECT 343.950 594.600 345.000 601.950 ;
        RECT 350.100 600.150 351.900 601.950 ;
        RECT 365.100 600.150 366.900 601.950 ;
        RECT 349.950 597.450 352.050 598.050 ;
        RECT 355.950 597.450 358.050 598.050 ;
        RECT 349.950 596.550 358.050 597.450 ;
        RECT 349.950 595.950 352.050 596.550 ;
        RECT 355.950 595.950 358.050 596.550 ;
        RECT 368.400 596.700 369.600 601.950 ;
        RECT 371.100 600.150 372.900 601.950 ;
        RECT 390.150 597.300 391.050 608.700 ;
        RECT 393.000 604.050 394.200 611.400 ;
        RECT 410.400 604.050 411.600 617.400 ;
        RECT 428.400 617.400 430.200 623.400 ;
        RECT 415.950 606.450 420.000 607.050 ;
        RECT 415.950 604.950 420.450 606.450 ;
        RECT 391.950 601.950 394.200 604.050 ;
        RECT 406.950 601.950 409.050 604.050 ;
        RECT 409.950 601.950 412.050 604.050 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 368.400 595.800 372.600 596.700 ;
        RECT 390.150 596.400 392.100 597.300 ;
        RECT 326.400 588.600 328.200 594.600 ;
        RECT 343.200 588.600 345.000 594.600 ;
        RECT 370.800 588.600 372.600 595.800 ;
        RECT 386.400 595.500 392.100 596.400 ;
        RECT 386.400 591.600 387.600 595.500 ;
        RECT 393.000 594.600 394.200 601.950 ;
        RECT 407.100 600.150 408.900 601.950 ;
        RECT 410.400 596.700 411.600 601.950 ;
        RECT 413.100 600.150 414.900 601.950 ;
        RECT 419.550 601.050 420.450 604.950 ;
        RECT 425.100 604.050 426.900 605.850 ;
        RECT 428.400 604.050 429.600 617.400 ;
        RECT 448.800 611.400 450.600 623.400 ;
        RECT 455.550 611.400 457.350 623.400 ;
        RECT 463.050 617.400 464.850 623.400 ;
        RECT 460.950 615.300 464.850 617.400 ;
        RECT 470.850 616.500 472.650 623.400 ;
        RECT 478.650 617.400 480.450 623.400 ;
        RECT 479.250 616.500 480.450 617.400 ;
        RECT 469.950 615.450 476.550 616.500 ;
        RECT 469.950 614.700 471.750 615.450 ;
        RECT 474.750 614.700 476.550 615.450 ;
        RECT 479.250 614.400 484.050 616.500 ;
        RECT 462.150 612.600 464.850 614.400 ;
        RECT 465.750 613.800 467.550 614.400 ;
        RECT 465.750 612.900 472.050 613.800 ;
        RECT 479.250 613.500 480.450 614.400 ;
        RECT 465.750 612.600 467.550 612.900 ;
        RECT 463.950 611.700 464.850 612.600 ;
        RECT 441.000 606.450 445.050 607.050 ;
        RECT 440.550 604.950 445.050 606.450 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 415.950 599.550 420.450 601.050 ;
        RECT 415.950 598.950 420.000 599.550 ;
        RECT 386.400 588.600 388.200 591.600 ;
        RECT 392.400 588.600 394.200 594.600 ;
        RECT 407.400 595.800 411.600 596.700 ;
        RECT 407.400 588.600 409.200 595.800 ;
        RECT 428.400 591.600 429.600 601.950 ;
        RECT 440.550 601.050 441.450 604.950 ;
        RECT 449.250 604.050 450.300 611.400 ;
        RECT 455.550 604.050 456.750 611.400 ;
        RECT 460.950 610.800 463.050 611.700 ;
        RECT 463.950 610.800 469.050 611.700 ;
        RECT 458.850 609.600 463.050 610.800 ;
        RECT 457.950 607.800 459.750 609.600 ;
        RECT 445.950 601.950 450.300 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 455.550 603.750 460.050 604.050 ;
        RECT 455.550 601.950 461.850 603.750 ;
        RECT 440.550 599.550 445.050 601.050 ;
        RECT 441.000 598.950 445.050 599.550 ;
        RECT 449.250 594.600 450.300 601.950 ;
        RECT 452.100 600.150 453.900 601.950 ;
        RECT 455.550 594.600 456.750 601.950 ;
        RECT 468.150 598.200 469.050 610.800 ;
        RECT 471.150 610.800 472.050 612.900 ;
        RECT 472.950 612.300 480.450 613.500 ;
        RECT 472.950 611.700 474.750 612.300 ;
        RECT 487.050 611.400 488.850 623.400 ;
        RECT 471.150 610.500 479.550 610.800 ;
        RECT 487.950 610.500 488.850 611.400 ;
        RECT 471.150 609.900 488.850 610.500 ;
        RECT 477.750 609.300 488.850 609.900 ;
        RECT 477.750 609.000 479.550 609.300 ;
        RECT 475.950 602.400 478.050 604.050 ;
        RECT 475.950 601.200 483.900 602.400 ;
        RECT 484.950 601.950 487.050 604.050 ;
        RECT 482.100 600.600 483.900 601.200 ;
        RECT 485.100 600.150 486.900 601.950 ;
        RECT 479.100 599.400 480.900 600.000 ;
        RECT 485.100 599.400 486.000 600.150 ;
        RECT 479.100 598.200 486.000 599.400 ;
        RECT 468.150 597.000 480.150 598.200 ;
        RECT 468.150 596.400 469.950 597.000 ;
        RECT 479.100 595.200 480.150 597.000 ;
        RECT 428.400 588.600 430.200 591.600 ;
        RECT 448.800 588.600 450.600 594.600 ;
        RECT 455.550 588.600 457.350 594.600 ;
        RECT 460.950 593.700 463.050 594.600 ;
        RECT 460.950 592.500 464.700 593.700 ;
        RECT 475.350 593.550 477.150 594.300 ;
        RECT 463.650 591.600 464.700 592.500 ;
        RECT 472.200 592.500 477.150 593.550 ;
        RECT 478.650 593.400 480.450 595.200 ;
        RECT 487.950 594.600 488.850 609.300 ;
        RECT 503.400 617.400 505.200 623.400 ;
        RECT 503.400 604.050 504.600 617.400 ;
        RECT 512.550 611.400 514.350 623.400 ;
        RECT 520.050 617.400 521.850 623.400 ;
        RECT 517.950 615.300 521.850 617.400 ;
        RECT 527.850 616.500 529.650 623.400 ;
        RECT 535.650 617.400 537.450 623.400 ;
        RECT 536.250 616.500 537.450 617.400 ;
        RECT 526.950 615.450 533.550 616.500 ;
        RECT 526.950 614.700 528.750 615.450 ;
        RECT 531.750 614.700 533.550 615.450 ;
        RECT 536.250 614.400 541.050 616.500 ;
        RECT 519.150 612.600 521.850 614.400 ;
        RECT 522.750 613.800 524.550 614.400 ;
        RECT 522.750 612.900 529.050 613.800 ;
        RECT 536.250 613.500 537.450 614.400 ;
        RECT 522.750 612.600 524.550 612.900 ;
        RECT 520.950 611.700 521.850 612.600 ;
        RECT 512.550 604.050 513.750 611.400 ;
        RECT 517.950 610.800 520.050 611.700 ;
        RECT 520.950 610.800 526.050 611.700 ;
        RECT 515.850 609.600 520.050 610.800 ;
        RECT 514.950 607.800 516.750 609.600 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 502.950 601.950 505.050 604.050 ;
        RECT 505.950 601.950 508.050 604.050 ;
        RECT 512.550 603.750 517.050 604.050 ;
        RECT 512.550 601.950 518.850 603.750 ;
        RECT 500.100 600.150 501.900 601.950 ;
        RECT 503.400 596.700 504.600 601.950 ;
        RECT 506.100 600.150 507.900 601.950 ;
        RECT 503.400 595.800 507.600 596.700 ;
        RECT 481.950 592.500 484.050 594.600 ;
        RECT 472.200 591.600 473.250 592.500 ;
        RECT 481.950 591.600 483.000 592.500 ;
        RECT 463.650 588.600 465.450 591.600 ;
        RECT 471.450 588.600 473.250 591.600 ;
        RECT 479.250 590.700 483.000 591.600 ;
        RECT 479.250 588.600 481.050 590.700 ;
        RECT 487.050 588.600 488.850 594.600 ;
        RECT 505.800 588.600 507.600 595.800 ;
        RECT 512.550 594.600 513.750 601.950 ;
        RECT 525.150 598.200 526.050 610.800 ;
        RECT 528.150 610.800 529.050 612.900 ;
        RECT 529.950 612.300 537.450 613.500 ;
        RECT 529.950 611.700 531.750 612.300 ;
        RECT 544.050 611.400 545.850 623.400 ;
        RECT 528.150 610.500 536.550 610.800 ;
        RECT 544.950 610.500 545.850 611.400 ;
        RECT 528.150 609.900 545.850 610.500 ;
        RECT 534.750 609.300 545.850 609.900 ;
        RECT 534.750 609.000 536.550 609.300 ;
        RECT 532.950 602.400 535.050 604.050 ;
        RECT 532.950 601.200 540.900 602.400 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 539.100 600.600 540.900 601.200 ;
        RECT 542.100 600.150 543.900 601.950 ;
        RECT 536.100 599.400 537.900 600.000 ;
        RECT 542.100 599.400 543.000 600.150 ;
        RECT 536.100 598.200 543.000 599.400 ;
        RECT 525.150 597.000 537.150 598.200 ;
        RECT 525.150 596.400 526.950 597.000 ;
        RECT 536.100 595.200 537.150 597.000 ;
        RECT 512.550 588.600 514.350 594.600 ;
        RECT 517.950 593.700 520.050 594.600 ;
        RECT 517.950 592.500 521.700 593.700 ;
        RECT 532.350 593.550 534.150 594.300 ;
        RECT 520.650 591.600 521.700 592.500 ;
        RECT 529.200 592.500 534.150 593.550 ;
        RECT 535.650 593.400 537.450 595.200 ;
        RECT 544.950 594.600 545.850 609.300 ;
        RECT 560.400 617.400 562.200 623.400 ;
        RECT 584.400 617.400 586.200 623.400 ;
        RECT 605.400 617.400 607.200 623.400 ;
        RECT 626.400 617.400 628.200 623.400 ;
        RECT 643.800 617.400 645.600 623.400 ;
        RECT 665.400 617.400 667.200 623.400 ;
        RECT 686.400 617.400 688.200 623.400 ;
        RECT 560.400 604.050 561.600 617.400 ;
        RECT 584.850 604.050 586.050 617.400 ;
        RECT 590.100 604.050 591.900 605.850 ;
        RECT 605.400 604.050 606.600 617.400 ;
        RECT 610.950 609.450 613.050 610.050 ;
        RECT 622.950 609.450 625.050 610.050 ;
        RECT 610.950 608.550 625.050 609.450 ;
        RECT 610.950 607.950 613.050 608.550 ;
        RECT 622.950 607.950 625.050 608.550 ;
        RECT 626.850 604.050 628.050 617.400 ;
        RECT 634.950 606.450 639.000 607.050 ;
        RECT 632.100 604.050 633.900 605.850 ;
        RECT 634.950 604.950 639.450 606.450 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 580.950 601.950 583.050 604.050 ;
        RECT 583.950 601.950 586.050 604.050 ;
        RECT 586.950 601.950 589.050 604.050 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 604.950 601.950 607.050 604.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 625.950 601.950 628.050 604.050 ;
        RECT 628.950 601.950 631.050 604.050 ;
        RECT 631.950 601.950 634.050 604.050 ;
        RECT 557.100 600.150 558.900 601.950 ;
        RECT 560.400 596.700 561.600 601.950 ;
        RECT 563.100 600.150 564.900 601.950 ;
        RECT 581.100 600.150 582.900 601.950 ;
        RECT 583.950 597.750 585.150 601.950 ;
        RECT 587.100 600.150 588.900 601.950 ;
        RECT 602.100 600.150 603.900 601.950 ;
        RECT 581.400 596.700 585.150 597.750 ;
        RECT 605.400 596.700 606.600 601.950 ;
        RECT 608.100 600.150 609.900 601.950 ;
        RECT 623.100 600.150 624.900 601.950 ;
        RECT 625.950 597.750 627.150 601.950 ;
        RECT 629.100 600.150 630.900 601.950 ;
        RECT 638.550 598.050 639.450 604.950 ;
        RECT 644.400 604.050 645.600 617.400 ;
        RECT 646.950 609.450 649.050 610.050 ;
        RECT 661.950 609.450 664.050 609.900 ;
        RECT 646.950 608.550 664.050 609.450 ;
        RECT 646.950 607.950 649.050 608.550 ;
        RECT 661.950 607.800 664.050 608.550 ;
        RECT 647.100 604.050 648.900 605.850 ;
        RECT 665.850 604.050 667.050 617.400 ;
        RECT 671.100 604.050 672.900 605.850 ;
        RECT 686.400 604.050 687.600 617.400 ;
        RECT 706.500 612.600 708.300 623.400 ;
        RECT 727.800 617.400 729.600 623.400 ;
        RECT 704.700 611.400 708.300 612.600 ;
        RECT 691.950 606.450 696.000 607.050 ;
        RECT 691.950 604.950 696.450 606.450 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 646.950 601.950 649.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 623.400 596.700 627.150 597.750 ;
        RECT 560.400 595.800 564.600 596.700 ;
        RECT 538.950 592.500 541.050 594.600 ;
        RECT 529.200 591.600 530.250 592.500 ;
        RECT 538.950 591.600 540.000 592.500 ;
        RECT 520.650 588.600 522.450 591.600 ;
        RECT 528.450 588.600 530.250 591.600 ;
        RECT 536.250 590.700 540.000 591.600 ;
        RECT 536.250 588.600 538.050 590.700 ;
        RECT 544.050 588.600 545.850 594.600 ;
        RECT 562.800 588.600 564.600 595.800 ;
        RECT 581.400 594.600 582.600 596.700 ;
        RECT 605.400 595.800 609.600 596.700 ;
        RECT 580.800 588.600 582.600 594.600 ;
        RECT 583.800 593.700 591.600 595.050 ;
        RECT 583.800 588.600 585.600 593.700 ;
        RECT 589.800 588.600 591.600 593.700 ;
        RECT 607.800 588.600 609.600 595.800 ;
        RECT 623.400 594.600 624.600 596.700 ;
        RECT 637.950 595.950 640.050 598.050 ;
        RECT 622.800 588.600 624.600 594.600 ;
        RECT 625.800 593.700 633.600 595.050 ;
        RECT 625.800 588.600 627.600 593.700 ;
        RECT 631.800 588.600 633.600 593.700 ;
        RECT 644.400 591.600 645.600 601.950 ;
        RECT 662.100 600.150 663.900 601.950 ;
        RECT 664.950 597.750 666.150 601.950 ;
        RECT 668.100 600.150 669.900 601.950 ;
        RECT 683.100 600.150 684.900 601.950 ;
        RECT 662.400 596.700 666.150 597.750 ;
        RECT 673.950 597.450 676.050 598.050 ;
        RECT 682.950 597.450 685.050 598.050 ;
        RECT 662.400 594.600 663.600 596.700 ;
        RECT 673.950 596.550 685.050 597.450 ;
        RECT 673.950 595.950 676.050 596.550 ;
        RECT 682.950 595.950 685.050 596.550 ;
        RECT 686.400 596.700 687.600 601.950 ;
        RECT 689.100 600.150 690.900 601.950 ;
        RECT 686.400 595.800 690.600 596.700 ;
        RECT 643.800 588.600 645.600 591.600 ;
        RECT 661.800 588.600 663.600 594.600 ;
        RECT 664.800 593.700 672.600 595.050 ;
        RECT 664.800 588.600 666.600 593.700 ;
        RECT 670.800 588.600 672.600 593.700 ;
        RECT 688.800 588.600 690.600 595.800 ;
        RECT 695.550 594.900 696.450 604.950 ;
        RECT 701.100 604.050 702.900 605.850 ;
        RECT 704.700 604.050 705.600 611.400 ;
        RECT 707.100 604.050 708.900 605.850 ;
        RECT 728.400 604.050 729.600 617.400 ;
        RECT 740.400 612.300 742.200 623.400 ;
        RECT 740.400 611.400 744.900 612.300 ;
        RECT 747.900 611.400 749.700 623.400 ;
        RECT 755.400 612.600 757.200 623.400 ;
        RECT 742.800 609.300 744.900 611.400 ;
        RECT 748.500 609.900 749.700 611.400 ;
        RECT 752.400 611.400 757.200 612.600 ;
        RECT 773.400 617.400 775.200 623.400 ;
        RECT 752.400 610.500 754.500 611.400 ;
        RECT 748.500 609.000 750.000 609.900 ;
        RECT 746.100 607.500 748.200 607.800 ;
        RECT 744.300 605.700 748.200 607.500 ;
        RECT 749.100 606.900 750.000 609.000 ;
        RECT 749.100 604.800 751.200 606.900 ;
        RECT 765.000 606.450 769.050 607.050 ;
        RECT 700.950 601.950 703.050 604.050 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 740.400 603.900 742.500 604.050 ;
        RECT 745.500 603.900 747.300 604.500 ;
        RECT 740.400 602.700 747.300 603.900 ;
        RECT 748.200 603.900 750.600 604.800 ;
        RECT 755.100 604.050 756.900 605.850 ;
        RECT 764.550 604.950 769.050 606.450 ;
        RECT 740.400 601.950 742.500 602.700 ;
        RECT 694.950 592.800 697.050 594.900 ;
        RECT 704.700 591.600 705.600 601.950 ;
        RECT 725.100 600.150 726.900 601.950 ;
        RECT 728.400 596.700 729.600 601.950 ;
        RECT 731.100 600.150 732.900 601.950 ;
        RECT 740.400 601.050 742.200 601.950 ;
        RECT 736.950 600.150 742.200 601.050 ;
        RECT 736.950 599.550 741.450 600.150 ;
        RECT 736.950 598.950 741.000 599.550 ;
        RECT 745.500 599.400 747.300 601.200 ;
        RECT 745.200 597.300 747.300 599.400 ;
        RECT 725.400 595.800 729.600 596.700 ;
        RECT 741.000 596.400 747.300 597.300 ;
        RECT 748.200 598.200 749.250 603.900 ;
        RECT 754.950 603.450 757.050 604.050 ;
        RECT 764.550 603.450 765.450 604.950 ;
        RECT 770.100 604.050 771.900 605.850 ;
        RECT 773.400 604.050 774.600 617.400 ;
        RECT 788.400 612.300 790.200 623.400 ;
        RECT 794.400 612.300 796.200 623.400 ;
        RECT 788.400 611.400 796.200 612.300 ;
        RECT 797.400 611.400 799.200 623.400 ;
        RECT 812.400 612.300 814.200 623.400 ;
        RECT 812.400 611.400 816.900 612.300 ;
        RECT 819.900 611.400 821.700 623.400 ;
        RECT 827.400 612.600 829.200 623.400 ;
        RECT 847.800 617.400 849.600 623.400 ;
        RECT 778.950 609.450 781.050 610.050 ;
        RECT 793.950 609.450 796.050 610.050 ;
        RECT 778.950 608.550 796.050 609.450 ;
        RECT 778.950 607.950 781.050 608.550 ;
        RECT 793.950 607.950 796.050 608.550 ;
        RECT 791.100 604.050 792.900 605.850 ;
        RECT 797.700 604.050 798.600 611.400 ;
        RECT 814.800 609.300 816.900 611.400 ;
        RECT 820.500 609.900 821.700 611.400 ;
        RECT 824.400 611.400 829.200 612.600 ;
        RECT 824.400 610.500 826.500 611.400 ;
        RECT 820.500 609.000 822.000 609.900 ;
        RECT 818.100 607.500 820.200 607.800 ;
        RECT 808.950 606.450 813.000 607.050 ;
        RECT 808.950 604.950 814.050 606.450 ;
        RECT 816.300 605.700 820.200 607.500 ;
        RECT 821.100 606.900 822.000 609.000 ;
        RECT 811.950 604.050 814.050 604.950 ;
        RECT 821.100 604.800 823.200 606.900 ;
        RECT 750.600 601.200 752.400 603.000 ;
        RECT 754.950 602.550 765.450 603.450 ;
        RECT 754.950 601.950 757.050 602.550 ;
        RECT 750.150 599.100 752.250 601.200 ;
        RECT 764.550 601.050 765.450 602.550 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 787.950 601.950 790.050 604.050 ;
        RECT 790.950 601.950 793.050 604.050 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 812.400 603.900 814.500 604.050 ;
        RECT 817.500 603.900 819.300 604.500 ;
        RECT 812.400 602.700 819.300 603.900 ;
        RECT 820.200 603.900 822.600 604.800 ;
        RECT 827.100 604.050 828.900 605.850 ;
        RECT 848.400 604.050 849.600 617.400 ;
        RECT 866.400 617.400 868.200 623.400 ;
        RECT 883.800 617.400 885.600 623.400 ;
        RECT 853.950 609.450 856.050 610.050 ;
        RECT 862.950 609.450 865.050 609.900 ;
        RECT 853.950 608.550 865.050 609.450 ;
        RECT 853.950 607.950 856.050 608.550 ;
        RECT 862.950 607.800 865.050 608.550 ;
        RECT 866.400 604.050 867.600 617.400 ;
        RECT 884.700 617.100 885.600 617.400 ;
        RECT 889.800 617.400 891.600 623.400 ;
        RECT 908.400 617.400 910.200 623.400 ;
        RECT 889.800 617.100 891.300 617.400 ;
        RECT 884.700 616.200 891.300 617.100 ;
        RECT 908.700 617.100 910.200 617.400 ;
        RECT 914.400 617.400 916.200 623.400 ;
        RECT 914.400 617.100 915.300 617.400 ;
        RECT 908.700 616.200 915.300 617.100 ;
        RECT 884.700 604.050 885.600 616.200 ;
        RECT 886.950 609.450 889.050 610.200 ;
        RECT 898.950 609.450 901.050 610.050 ;
        RECT 910.950 609.450 913.050 610.200 ;
        RECT 886.950 608.550 901.050 609.450 ;
        RECT 886.950 608.100 889.050 608.550 ;
        RECT 898.950 607.950 901.050 608.550 ;
        RECT 902.550 608.550 913.050 609.450 ;
        RECT 902.550 606.450 903.450 608.550 ;
        RECT 910.950 608.100 913.050 608.550 ;
        RECT 890.100 604.050 891.900 605.850 ;
        RECT 899.550 605.550 903.450 606.450 ;
        RECT 812.400 601.950 814.500 602.700 ;
        RECT 764.550 599.550 769.050 601.050 ;
        RECT 765.000 598.950 769.050 599.550 ;
        RECT 704.400 588.600 706.200 591.600 ;
        RECT 725.400 588.600 727.200 595.800 ;
        RECT 741.000 594.600 742.200 596.400 ;
        RECT 748.200 596.100 751.200 598.200 ;
        RECT 748.200 594.600 749.400 596.100 ;
        RECT 752.400 595.500 754.500 596.700 ;
        RECT 752.400 594.600 757.200 595.500 ;
        RECT 740.400 588.600 742.200 594.600 ;
        RECT 747.900 588.600 749.700 594.600 ;
        RECT 755.400 588.600 757.200 594.600 ;
        RECT 773.400 591.600 774.600 601.950 ;
        RECT 788.100 600.150 789.900 601.950 ;
        RECT 794.100 600.150 795.900 601.950 ;
        RECT 797.700 594.600 798.600 601.950 ;
        RECT 799.950 600.450 802.050 601.050 ;
        RECT 812.400 600.450 814.200 601.950 ;
        RECT 799.950 600.150 814.200 600.450 ;
        RECT 799.950 599.550 813.450 600.150 ;
        RECT 799.950 598.950 802.050 599.550 ;
        RECT 817.500 599.400 819.300 601.200 ;
        RECT 817.200 597.300 819.300 599.400 ;
        RECT 813.000 596.400 819.300 597.300 ;
        RECT 820.200 598.200 821.250 603.900 ;
        RECT 826.950 603.450 829.050 604.050 ;
        RECT 831.000 603.450 835.050 604.050 ;
        RECT 822.600 601.200 824.400 603.000 ;
        RECT 826.950 602.550 835.050 603.450 ;
        RECT 826.950 601.950 829.050 602.550 ;
        RECT 831.000 601.950 835.050 602.550 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 850.950 601.950 853.050 604.050 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 886.950 601.950 889.050 604.050 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 892.950 601.950 895.050 604.050 ;
        RECT 822.150 599.100 824.250 601.200 ;
        RECT 845.100 600.150 846.900 601.950 ;
        RECT 813.000 594.600 814.200 596.400 ;
        RECT 820.200 596.100 823.200 598.200 ;
        RECT 848.400 596.700 849.600 601.950 ;
        RECT 851.100 600.150 852.900 601.950 ;
        RECT 863.100 600.150 864.900 601.950 ;
        RECT 820.200 594.600 821.400 596.100 ;
        RECT 824.400 595.500 826.500 596.700 ;
        RECT 845.400 595.800 849.600 596.700 ;
        RECT 866.400 596.700 867.600 601.950 ;
        RECT 869.100 600.150 870.900 601.950 ;
        RECT 884.700 598.200 885.600 601.950 ;
        RECT 887.100 600.150 888.900 601.950 ;
        RECT 893.100 600.150 894.900 601.950 ;
        RECT 899.550 601.050 900.450 605.550 ;
        RECT 908.100 604.050 909.900 605.850 ;
        RECT 914.400 604.050 915.300 616.200 ;
        RECT 904.950 601.950 907.050 604.050 ;
        RECT 907.950 601.950 910.050 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 913.950 601.950 916.050 604.050 ;
        RECT 899.550 599.550 904.050 601.050 ;
        RECT 905.100 600.150 906.900 601.950 ;
        RECT 911.100 600.150 912.900 601.950 ;
        RECT 900.000 598.950 904.050 599.550 ;
        RECT 914.400 598.200 915.300 601.950 ;
        RECT 884.700 597.000 888.000 598.200 ;
        RECT 866.400 595.800 870.600 596.700 ;
        RECT 824.400 594.600 829.200 595.500 ;
        RECT 793.500 593.400 798.600 594.600 ;
        RECT 773.400 588.600 775.200 591.600 ;
        RECT 793.500 588.600 795.300 593.400 ;
        RECT 812.400 588.600 814.200 594.600 ;
        RECT 819.900 588.600 821.700 594.600 ;
        RECT 827.400 588.600 829.200 594.600 ;
        RECT 845.400 588.600 847.200 595.800 ;
        RECT 868.800 588.600 870.600 595.800 ;
        RECT 886.200 588.600 888.000 597.000 ;
        RECT 912.000 597.000 915.300 598.200 ;
        RECT 912.000 588.600 913.800 597.000 ;
        RECT 21.000 578.400 22.800 584.400 ;
        RECT 39.300 580.200 41.100 584.400 ;
        RECT 38.400 578.400 41.100 580.200 ;
        RECT 14.100 571.050 15.900 572.850 ;
        RECT 21.000 571.050 22.050 578.400 ;
        RECT 26.100 571.050 27.900 572.850 ;
        RECT 38.400 571.050 39.300 578.400 ;
        RECT 41.100 576.600 42.900 577.500 ;
        RECT 46.800 576.600 48.600 584.400 ;
        RECT 64.800 577.200 66.600 584.400 ;
        RECT 41.100 575.700 48.600 576.600 ;
        RECT 62.400 576.300 66.600 577.200 ;
        RECT 83.400 577.200 85.200 584.400 ;
        RECT 106.800 577.200 108.600 584.400 ;
        RECT 124.800 577.200 126.600 584.400 ;
        RECT 83.400 576.300 87.600 577.200 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 22.950 568.950 25.050 571.050 ;
        RECT 25.950 568.950 28.050 571.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 40.950 568.950 43.050 571.050 ;
        RECT 17.100 567.150 18.900 568.950 ;
        RECT 21.000 563.400 21.900 568.950 ;
        RECT 23.100 567.150 24.900 568.950 ;
        RECT 16.800 562.500 21.900 563.400 ;
        RECT 13.800 550.500 15.600 561.600 ;
        RECT 16.800 551.400 18.600 562.500 ;
        RECT 38.400 561.600 39.300 568.950 ;
        RECT 41.100 567.150 42.900 568.950 ;
        RECT 19.800 560.400 27.600 561.300 ;
        RECT 19.800 550.500 21.600 560.400 ;
        RECT 13.800 549.600 21.600 550.500 ;
        RECT 25.800 549.600 27.600 560.400 ;
        RECT 37.800 549.600 39.600 561.600 ;
        RECT 44.700 555.600 45.600 575.700 ;
        RECT 47.100 571.050 48.900 572.850 ;
        RECT 59.100 571.050 60.900 572.850 ;
        RECT 62.400 571.050 63.600 576.300 ;
        RECT 65.100 571.050 66.900 572.850 ;
        RECT 83.100 571.050 84.900 572.850 ;
        RECT 86.400 571.050 87.600 576.300 ;
        RECT 104.400 576.300 108.600 577.200 ;
        RECT 122.400 576.300 126.600 577.200 ;
        RECT 89.100 571.050 90.900 572.850 ;
        RECT 101.100 571.050 102.900 572.850 ;
        RECT 104.400 571.050 105.600 576.300 ;
        RECT 114.000 573.450 118.050 574.050 ;
        RECT 107.100 571.050 108.900 572.850 ;
        RECT 113.550 571.950 118.050 573.450 ;
        RECT 46.950 568.950 49.050 571.050 ;
        RECT 58.950 568.950 61.050 571.050 ;
        RECT 61.950 568.950 64.050 571.050 ;
        RECT 64.950 568.950 67.050 571.050 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 85.950 568.950 88.050 571.050 ;
        RECT 88.950 568.950 91.050 571.050 ;
        RECT 100.950 568.950 103.050 571.050 ;
        RECT 103.950 568.950 106.050 571.050 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 43.800 549.600 45.600 555.600 ;
        RECT 62.400 555.600 63.600 568.950 ;
        RECT 86.400 555.600 87.600 568.950 ;
        RECT 62.400 549.600 64.200 555.600 ;
        RECT 85.800 549.600 87.600 555.600 ;
        RECT 104.400 555.600 105.600 568.950 ;
        RECT 113.550 568.050 114.450 571.950 ;
        RECT 119.100 571.050 120.900 572.850 ;
        RECT 122.400 571.050 123.600 576.300 ;
        RECT 147.000 576.000 148.800 584.400 ;
        RECT 166.500 579.600 168.300 584.400 ;
        RECT 166.500 578.400 171.600 579.600 ;
        RECT 187.800 578.400 189.600 584.400 ;
        RECT 147.000 574.800 150.300 576.000 ;
        RECT 127.950 573.450 130.050 574.050 ;
        RECT 133.950 573.450 136.050 574.050 ;
        RECT 125.100 571.050 126.900 572.850 ;
        RECT 127.950 572.550 136.050 573.450 ;
        RECT 127.950 571.950 130.050 572.550 ;
        RECT 133.950 571.950 136.050 572.550 ;
        RECT 140.100 571.050 141.900 572.850 ;
        RECT 146.100 571.050 147.900 572.850 ;
        RECT 149.400 571.050 150.300 574.800 ;
        RECT 161.100 571.050 162.900 572.850 ;
        RECT 167.100 571.050 168.900 572.850 ;
        RECT 170.700 571.050 171.600 578.400 ;
        RECT 188.400 576.300 189.600 578.400 ;
        RECT 190.800 579.300 192.600 584.400 ;
        RECT 196.800 579.300 198.600 584.400 ;
        RECT 190.800 577.950 198.600 579.300 ;
        RECT 188.400 575.250 192.150 576.300 ;
        RECT 183.000 573.450 187.050 574.050 ;
        RECT 182.550 571.950 187.050 573.450 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 121.950 568.950 124.050 571.050 ;
        RECT 124.950 568.950 127.050 571.050 ;
        RECT 139.950 568.950 142.050 571.050 ;
        RECT 142.950 568.950 145.050 571.050 ;
        RECT 145.950 568.950 148.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 163.950 568.950 166.050 571.050 ;
        RECT 166.950 568.950 169.050 571.050 ;
        RECT 169.950 568.950 172.050 571.050 ;
        RECT 113.550 566.550 118.050 568.050 ;
        RECT 114.000 565.950 118.050 566.550 ;
        RECT 122.400 555.600 123.600 568.950 ;
        RECT 143.100 567.150 144.900 568.950 ;
        RECT 136.950 564.450 139.050 565.050 ;
        RECT 145.950 564.450 148.050 565.050 ;
        RECT 136.950 563.550 148.050 564.450 ;
        RECT 136.950 562.950 139.050 563.550 ;
        RECT 145.950 562.950 148.050 563.550 ;
        RECT 149.400 556.800 150.300 568.950 ;
        RECT 164.100 567.150 165.900 568.950 ;
        RECT 170.700 561.600 171.600 568.950 ;
        RECT 182.550 568.050 183.450 571.950 ;
        RECT 188.100 571.050 189.900 572.850 ;
        RECT 190.950 571.050 192.150 575.250 ;
        RECT 216.000 576.000 217.800 584.400 ;
        RECT 236.400 577.200 238.200 584.400 ;
        RECT 223.950 576.450 226.050 577.050 ;
        RECT 216.000 574.800 219.300 576.000 ;
        RECT 223.950 575.550 231.450 576.450 ;
        RECT 236.400 576.300 240.600 577.200 ;
        RECT 223.950 574.950 226.050 575.550 ;
        RECT 194.100 571.050 195.900 572.850 ;
        RECT 202.950 571.950 205.050 574.050 ;
        RECT 187.950 568.950 190.050 571.050 ;
        RECT 190.950 568.950 193.050 571.050 ;
        RECT 193.950 568.950 196.050 571.050 ;
        RECT 196.950 568.950 199.050 571.050 ;
        RECT 182.550 566.550 187.050 568.050 ;
        RECT 183.000 565.950 187.050 566.550 ;
        RECT 143.700 555.900 150.300 556.800 ;
        RECT 143.700 555.600 145.200 555.900 ;
        RECT 104.400 549.600 106.200 555.600 ;
        RECT 122.400 549.600 124.200 555.600 ;
        RECT 143.400 549.600 145.200 555.600 ;
        RECT 149.400 555.600 150.300 555.900 ;
        RECT 161.400 560.700 169.200 561.600 ;
        RECT 149.400 549.600 151.200 555.600 ;
        RECT 161.400 549.600 163.200 560.700 ;
        RECT 167.400 549.600 169.200 560.700 ;
        RECT 170.400 549.600 172.200 561.600 ;
        RECT 191.850 555.600 193.050 568.950 ;
        RECT 197.100 567.150 198.900 568.950 ;
        RECT 203.550 568.050 204.450 571.950 ;
        RECT 209.100 571.050 210.900 572.850 ;
        RECT 215.100 571.050 216.900 572.850 ;
        RECT 218.400 571.050 219.300 574.800 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 217.950 568.950 220.050 571.050 ;
        RECT 203.550 566.550 208.050 568.050 ;
        RECT 212.100 567.150 213.900 568.950 ;
        RECT 204.000 565.950 208.050 566.550 ;
        RECT 218.400 556.800 219.300 568.950 ;
        RECT 230.550 568.050 231.450 575.550 ;
        RECT 236.100 571.050 237.900 572.850 ;
        RECT 239.400 571.050 240.600 576.300 ;
        RECT 241.950 576.450 244.050 577.050 ;
        RECT 241.950 575.550 249.450 576.450 ;
        RECT 256.200 576.000 258.000 584.400 ;
        RECT 272.400 579.300 274.200 584.400 ;
        RECT 278.400 579.300 280.200 584.400 ;
        RECT 272.400 577.950 280.200 579.300 ;
        RECT 281.400 578.400 283.200 584.400 ;
        RECT 296.400 579.300 298.200 584.400 ;
        RECT 302.400 579.300 304.200 584.400 ;
        RECT 281.400 576.300 282.600 578.400 ;
        RECT 296.400 577.950 304.200 579.300 ;
        RECT 305.400 578.400 307.200 584.400 ;
        RECT 324.300 580.200 326.100 584.400 ;
        RECT 323.400 578.400 326.100 580.200 ;
        RECT 288.000 576.450 292.050 577.050 ;
        RECT 241.950 574.950 244.050 575.550 ;
        RECT 242.100 571.050 243.900 572.850 ;
        RECT 235.950 568.950 238.050 571.050 ;
        RECT 238.950 568.950 241.050 571.050 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 230.550 566.550 235.050 568.050 ;
        RECT 231.000 565.950 235.050 566.550 ;
        RECT 212.700 555.900 219.300 556.800 ;
        RECT 212.700 555.600 214.200 555.900 ;
        RECT 191.400 549.600 193.200 555.600 ;
        RECT 212.400 549.600 214.200 555.600 ;
        RECT 218.400 555.600 219.300 555.900 ;
        RECT 239.400 555.600 240.600 568.950 ;
        RECT 248.550 568.050 249.450 575.550 ;
        RECT 254.700 574.800 258.000 576.000 ;
        RECT 278.850 575.250 282.600 576.300 ;
        RECT 254.700 571.050 255.600 574.800 ;
        RECT 257.100 571.050 258.900 572.850 ;
        RECT 263.100 571.050 264.900 572.850 ;
        RECT 275.100 571.050 276.900 572.850 ;
        RECT 278.850 571.050 280.050 575.250 ;
        RECT 287.550 574.950 292.050 576.450 ;
        RECT 305.400 576.300 306.600 578.400 ;
        RECT 302.850 575.250 306.600 576.300 ;
        RECT 281.100 571.050 282.900 572.850 ;
        RECT 253.950 568.950 256.050 571.050 ;
        RECT 256.950 568.950 259.050 571.050 ;
        RECT 259.950 568.950 262.050 571.050 ;
        RECT 262.950 568.950 265.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 277.950 568.950 280.050 571.050 ;
        RECT 280.950 568.950 283.050 571.050 ;
        RECT 244.950 566.550 249.450 568.050 ;
        RECT 244.950 565.950 249.000 566.550 ;
        RECT 254.700 556.800 255.600 568.950 ;
        RECT 260.100 567.150 261.900 568.950 ;
        RECT 272.100 567.150 273.900 568.950 ;
        RECT 256.950 564.450 259.050 564.750 ;
        RECT 262.950 564.450 265.050 565.050 ;
        RECT 256.950 563.550 265.050 564.450 ;
        RECT 256.950 562.650 259.050 563.550 ;
        RECT 262.950 562.950 265.050 563.550 ;
        RECT 254.700 555.900 261.300 556.800 ;
        RECT 254.700 555.600 255.600 555.900 ;
        RECT 218.400 549.600 220.200 555.600 ;
        RECT 238.800 549.600 240.600 555.600 ;
        RECT 253.800 549.600 255.600 555.600 ;
        RECT 259.800 555.600 261.300 555.900 ;
        RECT 277.950 555.600 279.150 568.950 ;
        RECT 287.550 568.050 288.450 574.950 ;
        RECT 291.000 573.450 295.050 574.050 ;
        RECT 283.950 566.550 288.450 568.050 ;
        RECT 290.550 571.950 295.050 573.450 ;
        RECT 290.550 568.050 291.450 571.950 ;
        RECT 299.100 571.050 300.900 572.850 ;
        RECT 302.850 571.050 304.050 575.250 ;
        RECT 319.950 573.450 322.050 574.050 ;
        RECT 305.100 571.050 306.900 572.850 ;
        RECT 311.550 572.550 322.050 573.450 ;
        RECT 295.950 568.950 298.050 571.050 ;
        RECT 298.950 568.950 301.050 571.050 ;
        RECT 301.950 568.950 304.050 571.050 ;
        RECT 304.950 568.950 307.050 571.050 ;
        RECT 290.550 566.550 295.050 568.050 ;
        RECT 296.100 567.150 297.900 568.950 ;
        RECT 283.950 565.950 288.000 566.550 ;
        RECT 291.000 565.950 295.050 566.550 ;
        RECT 301.950 555.600 303.150 568.950 ;
        RECT 311.550 568.050 312.450 572.550 ;
        RECT 319.950 571.950 322.050 572.550 ;
        RECT 323.400 571.050 324.300 578.400 ;
        RECT 326.100 576.600 327.900 577.500 ;
        RECT 331.800 576.600 333.600 584.400 ;
        RECT 326.100 575.700 333.600 576.600 ;
        RECT 346.800 578.400 348.600 584.400 ;
        RECT 352.800 581.400 354.600 584.400 ;
        RECT 322.950 568.950 325.050 571.050 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 307.950 566.550 312.450 568.050 ;
        RECT 307.950 565.950 312.000 566.550 ;
        RECT 310.950 564.450 313.050 565.050 ;
        RECT 319.950 564.450 322.050 565.050 ;
        RECT 310.950 563.550 322.050 564.450 ;
        RECT 310.950 562.950 313.050 563.550 ;
        RECT 319.950 562.950 322.050 563.550 ;
        RECT 323.400 561.600 324.300 568.950 ;
        RECT 326.100 567.150 327.900 568.950 ;
        RECT 259.800 549.600 261.600 555.600 ;
        RECT 277.800 549.600 279.600 555.600 ;
        RECT 301.800 549.600 303.600 555.600 ;
        RECT 322.800 549.600 324.600 561.600 ;
        RECT 329.700 555.600 330.600 575.700 ;
        RECT 332.100 571.050 333.900 572.850 ;
        RECT 346.800 571.050 348.000 578.400 ;
        RECT 353.400 577.500 354.600 581.400 ;
        RECT 348.900 576.600 354.600 577.500 ;
        RECT 364.800 578.400 366.600 584.400 ;
        RECT 370.800 581.400 372.600 584.400 ;
        RECT 348.900 575.700 350.850 576.600 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 346.800 568.950 349.050 571.050 ;
        RECT 328.800 549.600 330.600 555.600 ;
        RECT 346.800 561.600 348.000 568.950 ;
        RECT 349.950 564.300 350.850 575.700 ;
        RECT 364.800 571.050 366.000 578.400 ;
        RECT 371.400 577.500 372.600 581.400 ;
        RECT 366.900 576.600 372.600 577.500 ;
        RECT 366.900 575.700 368.850 576.600 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 364.800 568.950 367.050 571.050 ;
        RECT 353.100 567.150 354.900 568.950 ;
        RECT 348.900 563.400 350.850 564.300 ;
        RECT 348.900 562.500 354.600 563.400 ;
        RECT 346.800 549.600 348.600 561.600 ;
        RECT 353.400 555.600 354.600 562.500 ;
        RECT 352.800 549.600 354.600 555.600 ;
        RECT 364.800 561.600 366.000 568.950 ;
        RECT 367.950 564.300 368.850 575.700 ;
        RECT 387.000 576.000 388.800 584.400 ;
        RECT 391.950 582.450 394.050 583.050 ;
        RECT 397.950 582.450 400.050 582.900 ;
        RECT 391.950 581.550 400.050 582.450 ;
        RECT 391.950 580.950 394.050 581.550 ;
        RECT 397.950 580.800 400.050 581.550 ;
        RECT 409.800 581.400 411.600 584.400 ;
        RECT 394.950 579.450 397.050 579.900 ;
        RECT 406.950 579.450 409.050 580.050 ;
        RECT 394.950 578.550 409.050 579.450 ;
        RECT 394.950 577.800 397.050 578.550 ;
        RECT 406.950 577.950 409.050 578.550 ;
        RECT 387.000 574.800 390.300 576.000 ;
        RECT 380.100 571.050 381.900 572.850 ;
        RECT 386.100 571.050 387.900 572.850 ;
        RECT 389.400 571.050 390.300 574.800 ;
        RECT 410.400 571.050 411.300 581.400 ;
        RECT 424.800 578.400 426.600 584.400 ;
        RECT 425.400 576.300 426.600 578.400 ;
        RECT 427.800 579.300 429.600 584.400 ;
        RECT 433.800 579.300 435.600 584.400 ;
        RECT 427.800 577.950 435.600 579.300 ;
        RECT 451.800 577.200 453.600 584.400 ;
        RECT 469.800 578.400 471.600 584.400 ;
        RECT 449.400 576.300 453.600 577.200 ;
        RECT 470.400 576.300 471.600 578.400 ;
        RECT 472.800 579.300 474.600 584.400 ;
        RECT 478.800 579.300 480.600 584.400 ;
        RECT 472.800 577.950 480.600 579.300 ;
        RECT 482.550 578.400 484.350 584.400 ;
        RECT 490.650 581.400 492.450 584.400 ;
        RECT 498.450 581.400 500.250 584.400 ;
        RECT 506.250 582.300 508.050 584.400 ;
        RECT 506.250 581.400 510.000 582.300 ;
        RECT 490.650 580.500 491.700 581.400 ;
        RECT 487.950 579.300 491.700 580.500 ;
        RECT 499.200 580.500 500.250 581.400 ;
        RECT 508.950 580.500 510.000 581.400 ;
        RECT 499.200 579.450 504.150 580.500 ;
        RECT 487.950 578.400 490.050 579.300 ;
        RECT 502.350 578.700 504.150 579.450 ;
        RECT 425.400 575.250 429.150 576.300 ;
        RECT 420.000 573.450 424.050 574.050 ;
        RECT 419.550 571.950 424.050 573.450 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 379.950 568.950 382.050 571.050 ;
        RECT 382.950 568.950 385.050 571.050 ;
        RECT 385.950 568.950 388.050 571.050 ;
        RECT 388.950 568.950 391.050 571.050 ;
        RECT 406.950 568.950 409.050 571.050 ;
        RECT 409.950 568.950 412.050 571.050 ;
        RECT 412.950 568.950 415.050 571.050 ;
        RECT 371.100 567.150 372.900 568.950 ;
        RECT 383.100 567.150 384.900 568.950 ;
        RECT 366.900 563.400 368.850 564.300 ;
        RECT 366.900 562.500 372.600 563.400 ;
        RECT 364.800 549.600 366.600 561.600 ;
        RECT 371.400 555.600 372.600 562.500 ;
        RECT 389.400 556.800 390.300 568.950 ;
        RECT 407.100 567.150 408.900 568.950 ;
        RECT 410.400 561.600 411.300 568.950 ;
        RECT 413.100 567.150 414.900 568.950 ;
        RECT 419.550 564.900 420.450 571.950 ;
        RECT 425.100 571.050 426.900 572.850 ;
        RECT 427.950 571.050 429.150 575.250 ;
        RECT 431.100 571.050 432.900 572.850 ;
        RECT 446.100 571.050 447.900 572.850 ;
        RECT 449.400 571.050 450.600 576.300 ;
        RECT 470.400 575.250 474.150 576.300 ;
        RECT 452.100 571.050 453.900 572.850 ;
        RECT 470.100 571.050 471.900 572.850 ;
        RECT 472.950 571.050 474.150 575.250 ;
        RECT 476.100 571.050 477.900 572.850 ;
        RECT 482.550 571.050 483.750 578.400 ;
        RECT 505.650 577.800 507.450 579.600 ;
        RECT 508.950 578.400 511.050 580.500 ;
        RECT 514.050 578.400 515.850 584.400 ;
        RECT 495.150 576.000 496.950 576.600 ;
        RECT 506.100 576.000 507.150 577.800 ;
        RECT 495.150 574.800 507.150 576.000 ;
        RECT 424.950 568.950 427.050 571.050 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 445.950 568.950 448.050 571.050 ;
        RECT 448.950 568.950 451.050 571.050 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 469.950 568.950 472.050 571.050 ;
        RECT 472.950 568.950 475.050 571.050 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 478.950 568.950 481.050 571.050 ;
        RECT 482.550 569.250 488.850 571.050 ;
        RECT 482.550 568.950 487.050 569.250 ;
        RECT 418.950 562.800 421.050 564.900 ;
        RECT 383.700 555.900 390.300 556.800 ;
        RECT 383.700 555.600 385.200 555.900 ;
        RECT 370.800 549.600 372.600 555.600 ;
        RECT 383.400 549.600 385.200 555.600 ;
        RECT 389.400 555.600 390.300 555.900 ;
        RECT 407.700 560.400 411.300 561.600 ;
        RECT 389.400 549.600 391.200 555.600 ;
        RECT 407.700 549.600 409.500 560.400 ;
        RECT 428.850 555.600 430.050 568.950 ;
        RECT 434.100 567.150 435.900 568.950 ;
        RECT 449.400 555.600 450.600 568.950 ;
        RECT 457.950 564.450 460.050 565.050 ;
        RECT 469.950 564.450 472.050 565.050 ;
        RECT 457.950 563.550 472.050 564.450 ;
        RECT 457.950 562.950 460.050 563.550 ;
        RECT 469.950 562.950 472.050 563.550 ;
        RECT 473.850 555.600 475.050 568.950 ;
        RECT 479.100 567.150 480.900 568.950 ;
        RECT 482.550 561.600 483.750 568.950 ;
        RECT 484.950 563.400 486.750 565.200 ;
        RECT 485.850 562.200 490.050 563.400 ;
        RECT 495.150 562.200 496.050 574.800 ;
        RECT 506.100 573.600 513.000 574.800 ;
        RECT 506.100 573.000 507.900 573.600 ;
        RECT 512.100 572.850 513.000 573.600 ;
        RECT 509.100 571.800 510.900 572.400 ;
        RECT 502.950 570.600 510.900 571.800 ;
        RECT 512.100 571.050 513.900 572.850 ;
        RECT 502.950 568.950 505.050 570.600 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 504.750 563.700 506.550 564.000 ;
        RECT 514.950 563.700 515.850 578.400 ;
        RECT 527.400 579.300 529.200 584.400 ;
        RECT 533.400 579.300 535.200 584.400 ;
        RECT 527.400 577.950 535.200 579.300 ;
        RECT 536.400 578.400 538.200 584.400 ;
        RECT 536.400 576.300 537.600 578.400 ;
        RECT 553.800 577.200 555.600 584.400 ;
        RECT 533.850 575.250 537.600 576.300 ;
        RECT 551.400 576.300 555.600 577.200 ;
        RECT 568.800 578.400 570.600 584.400 ;
        RECT 574.800 581.400 576.600 584.400 ;
        RECT 530.100 571.050 531.900 572.850 ;
        RECT 533.850 571.050 535.050 575.250 ;
        RECT 536.100 571.050 537.900 572.850 ;
        RECT 548.100 571.050 549.900 572.850 ;
        RECT 551.400 571.050 552.600 576.300 ;
        RECT 554.100 571.050 555.900 572.850 ;
        RECT 568.800 571.050 570.000 578.400 ;
        RECT 575.400 577.500 576.600 581.400 ;
        RECT 570.900 576.600 576.600 577.500 ;
        RECT 587.400 577.200 589.200 584.400 ;
        RECT 607.800 578.400 609.600 584.400 ;
        RECT 570.900 575.700 572.850 576.600 ;
        RECT 587.400 576.300 591.600 577.200 ;
        RECT 526.950 568.950 529.050 571.050 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 553.950 568.950 556.050 571.050 ;
        RECT 568.800 568.950 571.050 571.050 ;
        RECT 527.100 567.150 528.900 568.950 ;
        RECT 504.750 563.100 515.850 563.700 ;
        RECT 428.400 549.600 430.200 555.600 ;
        RECT 449.400 549.600 451.200 555.600 ;
        RECT 473.400 549.600 475.200 555.600 ;
        RECT 482.550 549.600 484.350 561.600 ;
        RECT 487.950 561.300 490.050 562.200 ;
        RECT 490.950 561.300 496.050 562.200 ;
        RECT 498.150 562.500 515.850 563.100 ;
        RECT 498.150 562.200 506.550 562.500 ;
        RECT 490.950 560.400 491.850 561.300 ;
        RECT 489.150 558.600 491.850 560.400 ;
        RECT 492.750 560.100 494.550 560.400 ;
        RECT 498.150 560.100 499.050 562.200 ;
        RECT 514.950 561.600 515.850 562.500 ;
        RECT 492.750 559.200 499.050 560.100 ;
        RECT 499.950 560.700 501.750 561.300 ;
        RECT 499.950 559.500 507.450 560.700 ;
        RECT 492.750 558.600 494.550 559.200 ;
        RECT 506.250 558.600 507.450 559.500 ;
        RECT 487.950 555.600 491.850 557.700 ;
        RECT 496.950 557.550 498.750 558.300 ;
        RECT 501.750 557.550 503.550 558.300 ;
        RECT 496.950 556.500 503.550 557.550 ;
        RECT 506.250 556.500 511.050 558.600 ;
        RECT 490.050 549.600 491.850 555.600 ;
        RECT 497.850 549.600 499.650 556.500 ;
        RECT 506.250 555.600 507.450 556.500 ;
        RECT 505.650 549.600 507.450 555.600 ;
        RECT 514.050 549.600 515.850 561.600 ;
        RECT 532.950 555.600 534.150 568.950 ;
        RECT 551.400 555.600 552.600 568.950 ;
        RECT 568.800 561.600 570.000 568.950 ;
        RECT 571.950 564.300 572.850 575.700 ;
        RECT 587.100 571.050 588.900 572.850 ;
        RECT 590.400 571.050 591.600 576.300 ;
        RECT 608.400 576.300 609.600 578.400 ;
        RECT 610.800 579.300 612.600 584.400 ;
        RECT 616.800 579.300 618.600 584.400 ;
        RECT 610.800 577.950 618.600 579.300 ;
        RECT 620.550 578.400 622.350 584.400 ;
        RECT 628.650 581.400 630.450 584.400 ;
        RECT 636.450 581.400 638.250 584.400 ;
        RECT 644.250 582.300 646.050 584.400 ;
        RECT 644.250 581.400 648.000 582.300 ;
        RECT 628.650 580.500 629.700 581.400 ;
        RECT 625.950 579.300 629.700 580.500 ;
        RECT 637.200 580.500 638.250 581.400 ;
        RECT 646.950 580.500 648.000 581.400 ;
        RECT 637.200 579.450 642.150 580.500 ;
        RECT 625.950 578.400 628.050 579.300 ;
        RECT 640.350 578.700 642.150 579.450 ;
        RECT 608.400 575.250 612.150 576.300 ;
        RECT 595.950 573.450 600.000 574.050 ;
        RECT 593.100 571.050 594.900 572.850 ;
        RECT 595.950 571.950 600.450 573.450 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 575.100 567.150 576.900 568.950 ;
        RECT 570.900 563.400 572.850 564.300 ;
        RECT 570.900 562.500 576.600 563.400 ;
        RECT 532.800 549.600 534.600 555.600 ;
        RECT 551.400 549.600 553.200 555.600 ;
        RECT 568.800 549.600 570.600 561.600 ;
        RECT 575.400 555.600 576.600 562.500 ;
        RECT 590.400 555.600 591.600 568.950 ;
        RECT 599.550 567.900 600.450 571.950 ;
        RECT 608.100 571.050 609.900 572.850 ;
        RECT 610.950 571.050 612.150 575.250 ;
        RECT 614.100 571.050 615.900 572.850 ;
        RECT 620.550 571.050 621.750 578.400 ;
        RECT 643.650 577.800 645.450 579.600 ;
        RECT 646.950 578.400 649.050 580.500 ;
        RECT 652.050 578.400 653.850 584.400 ;
        RECT 633.150 576.000 634.950 576.600 ;
        RECT 644.100 576.000 645.150 577.800 ;
        RECT 633.150 574.800 645.150 576.000 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 616.950 568.950 619.050 571.050 ;
        RECT 620.550 569.250 626.850 571.050 ;
        RECT 620.550 568.950 625.050 569.250 ;
        RECT 598.950 565.800 601.050 567.900 ;
        RECT 611.850 555.600 613.050 568.950 ;
        RECT 617.100 567.150 618.900 568.950 ;
        RECT 620.550 561.600 621.750 568.950 ;
        RECT 622.950 563.400 624.750 565.200 ;
        RECT 623.850 562.200 628.050 563.400 ;
        RECT 633.150 562.200 634.050 574.800 ;
        RECT 644.100 573.600 651.000 574.800 ;
        RECT 644.100 573.000 645.900 573.600 ;
        RECT 650.100 572.850 651.000 573.600 ;
        RECT 647.100 571.800 648.900 572.400 ;
        RECT 640.950 570.600 648.900 571.800 ;
        RECT 650.100 571.050 651.900 572.850 ;
        RECT 640.950 568.950 643.050 570.600 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 642.750 563.700 644.550 564.000 ;
        RECT 652.950 563.700 653.850 578.400 ;
        RECT 642.750 563.100 653.850 563.700 ;
        RECT 574.800 549.600 576.600 555.600 ;
        RECT 589.800 549.600 591.600 555.600 ;
        RECT 611.400 549.600 613.200 555.600 ;
        RECT 620.550 549.600 622.350 561.600 ;
        RECT 625.950 561.300 628.050 562.200 ;
        RECT 628.950 561.300 634.050 562.200 ;
        RECT 636.150 562.500 653.850 563.100 ;
        RECT 636.150 562.200 644.550 562.500 ;
        RECT 628.950 560.400 629.850 561.300 ;
        RECT 627.150 558.600 629.850 560.400 ;
        RECT 630.750 560.100 632.550 560.400 ;
        RECT 636.150 560.100 637.050 562.200 ;
        RECT 652.950 561.600 653.850 562.500 ;
        RECT 630.750 559.200 637.050 560.100 ;
        RECT 637.950 560.700 639.750 561.300 ;
        RECT 637.950 559.500 645.450 560.700 ;
        RECT 630.750 558.600 632.550 559.200 ;
        RECT 644.250 558.600 645.450 559.500 ;
        RECT 625.950 555.600 629.850 557.700 ;
        RECT 634.950 557.550 636.750 558.300 ;
        RECT 639.750 557.550 641.550 558.300 ;
        RECT 634.950 556.500 641.550 557.550 ;
        RECT 644.250 556.500 649.050 558.600 ;
        RECT 628.050 549.600 629.850 555.600 ;
        RECT 635.850 549.600 637.650 556.500 ;
        RECT 644.250 555.600 645.450 556.500 ;
        RECT 643.650 549.600 645.450 555.600 ;
        RECT 652.050 549.600 653.850 561.600 ;
        RECT 667.800 578.400 669.600 584.400 ;
        RECT 673.800 581.400 675.600 584.400 ;
        RECT 667.800 571.050 669.000 578.400 ;
        RECT 674.400 577.500 675.600 581.400 ;
        RECT 688.800 577.500 690.600 584.400 ;
        RECT 694.800 577.500 696.600 584.400 ;
        RECT 700.800 577.500 702.600 584.400 ;
        RECT 706.800 577.500 708.600 584.400 ;
        RECT 721.800 581.400 723.600 584.400 ;
        RECT 740.400 581.400 742.200 584.400 ;
        RECT 669.900 576.600 675.600 577.500 ;
        RECT 669.900 575.700 671.850 576.600 ;
        RECT 667.800 568.950 670.050 571.050 ;
        RECT 667.800 561.600 669.000 568.950 ;
        RECT 670.950 564.300 671.850 575.700 ;
        RECT 687.900 576.300 690.600 577.500 ;
        RECT 692.700 576.300 696.600 577.500 ;
        RECT 698.700 576.300 702.600 577.500 ;
        RECT 704.700 576.300 708.600 577.500 ;
        RECT 687.900 571.050 688.800 576.300 ;
        RECT 692.700 575.400 693.900 576.300 ;
        RECT 698.700 575.400 699.900 576.300 ;
        RECT 704.700 575.400 705.900 576.300 ;
        RECT 689.700 574.200 693.900 575.400 ;
        RECT 689.700 573.600 691.500 574.200 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 685.950 568.950 688.800 571.050 ;
        RECT 674.100 567.150 675.900 568.950 ;
        RECT 669.900 563.400 671.850 564.300 ;
        RECT 687.900 563.700 688.800 568.950 ;
        RECT 692.700 563.700 693.900 574.200 ;
        RECT 695.700 574.200 699.900 575.400 ;
        RECT 695.700 573.600 697.500 574.200 ;
        RECT 698.700 563.700 699.900 574.200 ;
        RECT 701.700 574.200 705.900 575.400 ;
        RECT 701.700 573.600 703.500 574.200 ;
        RECT 704.700 563.700 705.900 574.200 ;
        RECT 707.100 571.050 708.900 572.850 ;
        RECT 722.400 571.050 723.600 581.400 ;
        RECT 740.700 571.050 741.600 581.400 ;
        RECT 762.300 580.200 764.100 584.400 ;
        RECT 761.400 578.400 764.100 580.200 ;
        RECT 742.950 576.450 745.050 577.050 ;
        RECT 748.950 576.450 751.050 577.050 ;
        RECT 754.950 576.450 757.050 577.050 ;
        RECT 742.950 575.550 757.050 576.450 ;
        RECT 742.950 574.950 745.050 575.550 ;
        RECT 748.950 574.950 751.050 575.550 ;
        RECT 754.950 574.950 757.050 575.550 ;
        RECT 761.400 571.050 762.300 578.400 ;
        RECT 764.100 576.600 765.900 577.500 ;
        RECT 769.800 576.600 771.600 584.400 ;
        RECT 784.800 577.500 786.600 584.400 ;
        RECT 790.800 577.500 792.600 584.400 ;
        RECT 796.800 577.500 798.600 584.400 ;
        RECT 802.800 577.500 804.600 584.400 ;
        RECT 821.400 581.400 823.200 584.400 ;
        RECT 764.100 575.700 771.600 576.600 ;
        RECT 783.900 576.300 786.600 577.500 ;
        RECT 788.700 576.300 792.600 577.500 ;
        RECT 794.700 576.300 798.600 577.500 ;
        RECT 800.700 576.300 804.600 577.500 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 724.950 568.950 727.050 571.050 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 739.950 568.950 742.050 571.050 ;
        RECT 742.950 568.950 745.050 571.050 ;
        RECT 760.950 568.950 763.050 571.050 ;
        RECT 763.950 568.950 766.050 571.050 ;
        RECT 669.900 562.500 675.600 563.400 ;
        RECT 687.900 562.500 690.600 563.700 ;
        RECT 692.700 562.500 696.600 563.700 ;
        RECT 698.700 562.500 702.600 563.700 ;
        RECT 704.700 562.500 708.600 563.700 ;
        RECT 667.800 549.600 669.600 561.600 ;
        RECT 674.400 555.600 675.600 562.500 ;
        RECT 673.800 549.600 675.600 555.600 ;
        RECT 688.800 549.600 690.600 562.500 ;
        RECT 694.800 549.600 696.600 562.500 ;
        RECT 700.800 549.600 702.600 562.500 ;
        RECT 706.800 549.600 708.600 562.500 ;
        RECT 722.400 555.600 723.600 568.950 ;
        RECT 725.100 567.150 726.900 568.950 ;
        RECT 737.100 567.150 738.900 568.950 ;
        RECT 740.700 561.600 741.600 568.950 ;
        RECT 743.100 567.150 744.900 568.950 ;
        RECT 761.400 561.600 762.300 568.950 ;
        RECT 764.100 567.150 765.900 568.950 ;
        RECT 740.700 560.400 744.300 561.600 ;
        RECT 721.800 549.600 723.600 555.600 ;
        RECT 742.500 549.600 744.300 560.400 ;
        RECT 760.800 549.600 762.600 561.600 ;
        RECT 767.700 555.600 768.600 575.700 ;
        RECT 770.100 571.050 771.900 572.850 ;
        RECT 783.900 571.050 784.800 576.300 ;
        RECT 788.700 575.400 789.900 576.300 ;
        RECT 794.700 575.400 795.900 576.300 ;
        RECT 800.700 575.400 801.900 576.300 ;
        RECT 785.700 574.200 789.900 575.400 ;
        RECT 785.700 573.600 787.500 574.200 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 781.950 568.950 784.800 571.050 ;
        RECT 783.900 563.700 784.800 568.950 ;
        RECT 788.700 563.700 789.900 574.200 ;
        RECT 791.700 574.200 795.900 575.400 ;
        RECT 791.700 573.600 793.500 574.200 ;
        RECT 794.700 563.700 795.900 574.200 ;
        RECT 797.700 574.200 801.900 575.400 ;
        RECT 797.700 573.600 799.500 574.200 ;
        RECT 800.700 563.700 801.900 574.200 ;
        RECT 803.100 571.050 804.900 572.850 ;
        RECT 821.700 571.050 822.600 581.400 ;
        RECT 841.200 576.000 843.000 584.400 ;
        RECT 850.950 579.450 853.050 580.050 ;
        RECT 856.950 579.450 859.050 580.050 ;
        RECT 850.950 578.550 859.050 579.450 ;
        RECT 850.950 577.950 853.050 578.550 ;
        RECT 856.950 577.950 859.050 578.550 ;
        RECT 863.400 577.200 865.200 584.400 ;
        RECT 886.800 577.200 888.600 584.400 ;
        RECT 863.400 576.300 867.600 577.200 ;
        RECT 839.700 574.800 843.000 576.000 ;
        RECT 839.700 571.050 840.600 574.800 ;
        RECT 850.950 573.450 853.050 574.050 ;
        RECT 842.100 571.050 843.900 572.850 ;
        RECT 848.100 571.050 849.900 572.850 ;
        RECT 850.950 572.550 858.450 573.450 ;
        RECT 850.950 571.950 853.050 572.550 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 847.950 568.950 850.050 571.050 ;
        RECT 818.100 567.150 819.900 568.950 ;
        RECT 783.900 562.500 786.600 563.700 ;
        RECT 788.700 562.500 792.600 563.700 ;
        RECT 794.700 562.500 798.600 563.700 ;
        RECT 800.700 562.500 804.600 563.700 ;
        RECT 766.800 549.600 768.600 555.600 ;
        RECT 784.800 549.600 786.600 562.500 ;
        RECT 790.800 549.600 792.600 562.500 ;
        RECT 796.800 549.600 798.600 562.500 ;
        RECT 802.800 549.600 804.600 562.500 ;
        RECT 821.700 561.600 822.600 568.950 ;
        RECT 824.100 567.150 825.900 568.950 ;
        RECT 821.700 560.400 825.300 561.600 ;
        RECT 823.500 549.600 825.300 560.400 ;
        RECT 839.700 556.800 840.600 568.950 ;
        RECT 845.100 567.150 846.900 568.950 ;
        RECT 857.550 568.050 858.450 572.550 ;
        RECT 863.100 571.050 864.900 572.850 ;
        RECT 866.400 571.050 867.600 576.300 ;
        RECT 868.950 576.450 871.050 577.050 ;
        RECT 880.950 576.450 883.050 577.050 ;
        RECT 868.950 575.550 883.050 576.450 ;
        RECT 868.950 574.950 871.050 575.550 ;
        RECT 880.950 574.950 883.050 575.550 ;
        RECT 884.400 576.300 888.600 577.200 ;
        RECT 905.400 581.400 907.200 584.400 ;
        RECT 871.950 573.450 876.000 574.050 ;
        RECT 869.100 571.050 870.900 572.850 ;
        RECT 871.950 571.950 876.450 573.450 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 857.550 566.550 862.050 568.050 ;
        RECT 858.000 565.950 862.050 566.550 ;
        RECT 841.950 564.450 844.050 565.050 ;
        RECT 862.950 564.450 865.050 565.050 ;
        RECT 841.950 563.550 865.050 564.450 ;
        RECT 841.950 562.950 844.050 563.550 ;
        RECT 862.950 562.950 865.050 563.550 ;
        RECT 839.700 555.900 846.300 556.800 ;
        RECT 839.700 555.600 840.600 555.900 ;
        RECT 838.800 549.600 840.600 555.600 ;
        RECT 844.800 555.600 846.300 555.900 ;
        RECT 866.400 555.600 867.600 568.950 ;
        RECT 875.550 568.050 876.450 571.950 ;
        RECT 881.100 571.050 882.900 572.850 ;
        RECT 884.400 571.050 885.600 576.300 ;
        RECT 889.950 573.450 894.000 574.050 ;
        RECT 887.100 571.050 888.900 572.850 ;
        RECT 889.950 571.950 894.450 573.450 ;
        RECT 880.950 568.950 883.050 571.050 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 875.550 566.550 880.050 568.050 ;
        RECT 876.000 565.950 880.050 566.550 ;
        RECT 868.950 564.450 871.050 564.750 ;
        RECT 880.950 564.450 883.050 565.050 ;
        RECT 868.950 563.550 883.050 564.450 ;
        RECT 868.950 562.650 871.050 563.550 ;
        RECT 880.950 562.950 883.050 563.550 ;
        RECT 844.800 549.600 846.600 555.600 ;
        RECT 865.800 549.600 867.600 555.600 ;
        RECT 884.400 555.600 885.600 568.950 ;
        RECT 893.550 568.050 894.450 571.950 ;
        RECT 905.400 571.050 906.600 581.400 ;
        RECT 901.950 568.950 904.050 571.050 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 889.950 566.550 894.450 568.050 ;
        RECT 902.100 567.150 903.900 568.950 ;
        RECT 889.950 565.950 894.000 566.550 ;
        RECT 905.400 555.600 906.600 568.950 ;
        RECT 884.400 549.600 886.200 555.600 ;
        RECT 905.400 549.600 907.200 555.600 ;
        RECT 11.400 535.500 13.200 545.400 ;
        RECT 17.400 544.500 25.200 545.400 ;
        RECT 17.400 535.500 19.200 544.500 ;
        RECT 11.400 534.600 19.200 535.500 ;
        RECT 20.400 535.800 22.200 543.600 ;
        RECT 23.400 536.700 25.200 544.500 ;
        RECT 27.000 544.500 34.800 545.400 ;
        RECT 27.000 535.800 28.800 544.500 ;
        RECT 20.400 534.900 28.800 535.800 ;
        RECT 30.000 535.800 31.800 543.600 ;
        RECT 30.000 533.400 31.200 535.800 ;
        RECT 33.000 535.200 34.800 544.500 ;
        RECT 52.800 539.400 54.600 545.400 ;
        RECT 70.800 539.400 72.600 545.400 ;
        RECT 27.750 532.200 31.200 533.400 ;
        RECT 7.950 531.450 10.050 532.050 ;
        RECT 19.950 531.450 22.050 532.050 ;
        RECT 7.950 530.550 22.050 531.450 ;
        RECT 7.950 529.950 10.050 530.550 ;
        RECT 19.950 529.950 22.050 530.550 ;
        RECT 14.100 525.900 15.900 527.700 ;
        RECT 23.100 525.900 24.900 527.700 ;
        RECT 27.750 525.900 28.950 532.200 ;
        RECT 53.400 526.050 54.600 539.400 ;
        RECT 71.700 539.100 72.600 539.400 ;
        RECT 76.800 539.400 78.600 545.400 ;
        RECT 76.800 539.100 78.300 539.400 ;
        RECT 71.700 538.200 78.300 539.100 ;
        RECT 71.700 526.050 72.600 538.200 ;
        RECT 89.400 534.300 91.200 545.400 ;
        RECT 95.400 534.300 97.200 545.400 ;
        RECT 89.400 533.400 97.200 534.300 ;
        RECT 98.400 533.400 100.200 545.400 ;
        RECT 110.400 534.300 112.200 545.400 ;
        RECT 116.400 534.300 118.200 545.400 ;
        RECT 110.400 533.400 118.200 534.300 ;
        RECT 119.400 533.400 121.200 545.400 ;
        RECT 140.400 539.400 142.200 545.400 ;
        RECT 163.800 539.400 165.600 545.400 ;
        RECT 184.800 539.400 186.600 545.400 ;
        RECT 73.950 531.450 76.050 532.050 ;
        RECT 88.950 531.450 91.050 532.050 ;
        RECT 73.950 530.550 91.050 531.450 ;
        RECT 73.950 529.950 76.050 530.550 ;
        RECT 88.950 529.950 91.050 530.550 ;
        RECT 77.100 526.050 78.900 527.850 ;
        RECT 92.100 526.050 93.900 527.850 ;
        RECT 98.700 526.050 99.600 533.400 ;
        RECT 113.100 526.050 114.900 527.850 ;
        RECT 119.700 526.050 120.600 533.400 ;
        RECT 140.850 526.050 142.050 539.400 ;
        RECT 146.100 526.050 147.900 527.850 ;
        RECT 158.100 526.050 159.900 527.850 ;
        RECT 163.950 526.050 165.150 539.400 ;
        RECT 185.700 539.100 186.600 539.400 ;
        RECT 190.800 539.400 192.600 545.400 ;
        RECT 205.800 539.400 207.600 545.400 ;
        RECT 190.800 539.100 192.300 539.400 ;
        RECT 185.700 538.200 192.300 539.100 ;
        RECT 206.700 539.100 207.600 539.400 ;
        RECT 211.800 539.400 213.600 545.400 ;
        RECT 226.800 539.400 228.600 545.400 ;
        RECT 211.800 539.100 213.300 539.400 ;
        RECT 206.700 538.200 213.300 539.100 ;
        RECT 227.700 539.100 228.600 539.400 ;
        RECT 232.800 539.400 234.600 545.400 ;
        RECT 251.400 539.400 253.200 545.400 ;
        RECT 269.400 539.400 271.200 545.400 ;
        RECT 232.800 539.100 234.300 539.400 ;
        RECT 227.700 538.200 234.300 539.100 ;
        RECT 185.700 526.050 186.600 538.200 ;
        RECT 191.100 526.050 192.900 527.850 ;
        RECT 206.700 526.050 207.600 538.200 ;
        RECT 212.100 526.050 213.900 527.850 ;
        RECT 227.700 526.050 228.600 538.200 ;
        RECT 232.950 534.450 235.050 535.050 ;
        RECT 247.950 534.450 250.050 535.050 ;
        RECT 232.950 533.550 250.050 534.450 ;
        RECT 232.950 532.950 235.050 533.550 ;
        RECT 247.950 532.950 250.050 533.550 ;
        RECT 243.000 528.450 247.050 529.050 ;
        RECT 233.100 526.050 234.900 527.850 ;
        RECT 242.550 526.950 247.050 528.450 ;
        RECT 13.950 523.800 16.050 525.900 ;
        RECT 19.950 523.800 22.050 525.900 ;
        RECT 22.950 523.800 25.050 525.900 ;
        RECT 27.750 523.800 31.050 525.900 ;
        RECT 49.950 523.950 52.050 526.050 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 70.950 523.950 73.050 526.050 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 166.950 523.950 169.050 526.050 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 190.950 523.950 193.050 526.050 ;
        RECT 193.950 523.950 196.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 211.950 523.950 214.050 526.050 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 226.950 523.950 229.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 20.100 522.000 21.900 523.800 ;
        RECT 27.750 515.400 28.950 523.800 ;
        RECT 50.100 522.150 51.900 523.950 ;
        RECT 53.400 518.700 54.600 523.950 ;
        RECT 56.100 522.150 57.900 523.950 ;
        RECT 71.700 520.200 72.600 523.950 ;
        RECT 74.100 522.150 75.900 523.950 ;
        RECT 80.100 522.150 81.900 523.950 ;
        RECT 89.100 522.150 90.900 523.950 ;
        RECT 95.100 522.150 96.900 523.950 ;
        RECT 71.700 519.000 75.000 520.200 ;
        RECT 18.150 514.500 28.950 515.400 ;
        RECT 50.400 517.800 54.600 518.700 ;
        RECT 18.150 513.600 19.200 514.500 ;
        RECT 24.150 513.600 25.200 514.500 ;
        RECT 17.400 510.600 19.200 513.600 ;
        RECT 23.400 510.600 25.200 513.600 ;
        RECT 50.400 510.600 52.200 517.800 ;
        RECT 73.200 510.600 75.000 519.000 ;
        RECT 98.700 516.600 99.600 523.950 ;
        RECT 110.100 522.150 111.900 523.950 ;
        RECT 116.100 522.150 117.900 523.950 ;
        RECT 119.700 516.600 120.600 523.950 ;
        RECT 137.100 522.150 138.900 523.950 ;
        RECT 139.950 519.750 141.150 523.950 ;
        RECT 143.100 522.150 144.900 523.950 ;
        RECT 161.100 522.150 162.900 523.950 ;
        RECT 137.400 518.700 141.150 519.750 ;
        RECT 164.850 519.750 166.050 523.950 ;
        RECT 167.100 522.150 168.900 523.950 ;
        RECT 185.700 520.200 186.600 523.950 ;
        RECT 188.100 522.150 189.900 523.950 ;
        RECT 194.100 522.150 195.900 523.950 ;
        RECT 206.700 520.200 207.600 523.950 ;
        RECT 209.100 522.150 210.900 523.950 ;
        RECT 215.100 522.150 216.900 523.950 ;
        RECT 227.700 520.200 228.600 523.950 ;
        RECT 230.100 522.150 231.900 523.950 ;
        RECT 236.100 522.150 237.900 523.950 ;
        RECT 242.550 523.050 243.450 526.950 ;
        RECT 248.100 526.050 249.900 527.850 ;
        RECT 251.400 526.050 252.600 539.400 ;
        RECT 269.700 539.100 271.200 539.400 ;
        RECT 275.400 539.400 277.200 545.400 ;
        RECT 293.400 539.400 295.200 545.400 ;
        RECT 275.400 539.100 276.300 539.400 ;
        RECT 269.700 538.200 276.300 539.100 ;
        RECT 293.700 539.100 295.200 539.400 ;
        RECT 299.400 539.400 301.200 545.400 ;
        RECT 299.400 539.100 300.300 539.400 ;
        RECT 293.700 538.200 300.300 539.100 ;
        RECT 269.100 526.050 270.900 527.850 ;
        RECT 275.400 526.050 276.300 538.200 ;
        RECT 277.950 537.450 280.050 538.050 ;
        RECT 289.950 537.450 292.050 538.050 ;
        RECT 277.950 536.550 292.050 537.450 ;
        RECT 277.950 535.950 280.050 536.550 ;
        RECT 289.950 535.950 292.050 536.550 ;
        RECT 292.950 531.450 295.050 532.050 ;
        RECT 287.550 530.550 295.050 531.450 ;
        RECT 287.550 528.450 288.450 530.550 ;
        RECT 292.950 529.950 295.050 530.550 ;
        RECT 284.550 528.000 288.450 528.450 ;
        RECT 283.950 527.550 288.450 528.000 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 250.950 523.950 253.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 271.950 523.950 274.050 526.050 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 242.550 521.550 247.050 523.050 ;
        RECT 243.000 520.950 247.050 521.550 ;
        RECT 164.850 518.700 168.600 519.750 ;
        RECT 185.700 519.000 189.000 520.200 ;
        RECT 206.700 519.000 210.000 520.200 ;
        RECT 227.700 519.000 231.000 520.200 ;
        RECT 137.400 516.600 138.600 518.700 ;
        RECT 94.500 515.400 99.600 516.600 ;
        RECT 115.500 515.400 120.600 516.600 ;
        RECT 94.500 510.600 96.300 515.400 ;
        RECT 115.500 510.600 117.300 515.400 ;
        RECT 136.800 510.600 138.600 516.600 ;
        RECT 139.800 515.700 147.600 517.050 ;
        RECT 139.800 510.600 141.600 515.700 ;
        RECT 145.800 510.600 147.600 515.700 ;
        RECT 158.400 515.700 166.200 517.050 ;
        RECT 158.400 510.600 160.200 515.700 ;
        RECT 164.400 510.600 166.200 515.700 ;
        RECT 167.400 516.600 168.600 518.700 ;
        RECT 167.400 510.600 169.200 516.600 ;
        RECT 187.200 510.600 189.000 519.000 ;
        RECT 208.200 510.600 210.000 519.000 ;
        RECT 229.200 510.600 231.000 519.000 ;
        RECT 251.400 513.600 252.600 523.950 ;
        RECT 266.100 522.150 267.900 523.950 ;
        RECT 272.100 522.150 273.900 523.950 ;
        RECT 275.400 520.200 276.300 523.950 ;
        RECT 283.950 523.800 286.050 527.550 ;
        RECT 293.100 526.050 294.900 527.850 ;
        RECT 299.400 526.050 300.300 538.200 ;
        RECT 316.500 534.600 318.300 545.400 ;
        RECT 314.700 533.400 318.300 534.600 ;
        RECT 329.400 534.600 331.200 545.400 ;
        RECT 335.400 544.500 343.200 545.400 ;
        RECT 335.400 534.600 337.200 544.500 ;
        RECT 329.400 533.700 337.200 534.600 ;
        RECT 306.000 528.450 310.050 529.050 ;
        RECT 305.550 526.950 310.050 528.450 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 292.950 523.950 295.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 290.100 522.150 291.900 523.950 ;
        RECT 296.100 522.150 297.900 523.950 ;
        RECT 299.400 520.200 300.300 523.950 ;
        RECT 305.550 523.050 306.450 526.950 ;
        RECT 311.100 526.050 312.900 527.850 ;
        RECT 314.700 526.050 315.600 533.400 ;
        RECT 338.400 532.500 340.200 543.600 ;
        RECT 341.400 533.400 343.200 544.500 ;
        RECT 359.400 533.400 361.200 545.400 ;
        RECT 376.800 539.400 378.600 545.400 ;
        RECT 335.100 531.600 340.200 532.500 ;
        RECT 317.100 526.050 318.900 527.850 ;
        RECT 332.100 526.050 333.900 527.850 ;
        RECT 335.100 526.050 336.000 531.600 ;
        RECT 338.100 526.050 339.900 527.850 ;
        RECT 359.400 526.050 360.600 533.400 ;
        RECT 377.400 526.050 378.600 539.400 ;
        RECT 395.400 539.400 397.200 545.400 ;
        RECT 400.950 543.450 403.050 544.050 ;
        RECT 406.950 543.450 409.050 544.050 ;
        RECT 400.950 542.550 409.050 543.450 ;
        RECT 400.950 541.950 403.050 542.550 ;
        RECT 406.950 541.950 409.050 542.550 ;
        RECT 415.800 539.400 417.600 545.400 ;
        RECT 392.100 526.050 393.900 527.850 ;
        RECT 395.400 526.050 396.600 539.400 ;
        RECT 416.400 526.050 417.600 539.400 ;
        RECT 431.400 534.600 433.200 545.400 ;
        RECT 437.400 544.500 445.200 545.400 ;
        RECT 437.400 534.600 439.200 544.500 ;
        RECT 431.400 533.700 439.200 534.600 ;
        RECT 440.400 532.500 442.200 543.600 ;
        RECT 443.400 533.400 445.200 544.500 ;
        RECT 464.400 539.400 466.200 545.400 ;
        RECT 482.400 539.400 484.200 545.400 ;
        RECT 502.800 539.400 504.600 545.400 ;
        RECT 526.800 539.400 528.600 545.400 ;
        RECT 544.800 539.400 546.600 545.400 ;
        RECT 418.950 531.450 421.050 532.050 ;
        RECT 427.950 531.450 430.050 532.050 ;
        RECT 418.950 530.550 430.050 531.450 ;
        RECT 418.950 529.950 421.050 530.550 ;
        RECT 427.950 529.950 430.050 530.550 ;
        RECT 437.100 531.600 442.200 532.500 ;
        RECT 434.100 526.050 435.900 527.850 ;
        RECT 437.100 526.050 438.000 531.600 ;
        RECT 440.100 526.050 441.900 527.850 ;
        RECT 464.850 526.050 466.050 539.400 ;
        RECT 470.100 526.050 471.900 527.850 ;
        RECT 482.400 526.050 483.600 539.400 ;
        RECT 497.100 526.050 498.900 527.850 ;
        RECT 502.950 526.050 504.150 539.400 ;
        RECT 521.100 526.050 522.900 527.850 ;
        RECT 526.950 526.050 528.150 539.400 ;
        RECT 545.400 526.050 546.600 539.400 ;
        RECT 563.400 539.400 565.200 545.400 ;
        RECT 548.100 526.050 549.900 527.850 ;
        RECT 560.100 526.050 561.900 527.850 ;
        RECT 563.400 526.050 564.600 539.400 ;
        RECT 580.800 533.400 582.600 545.400 ;
        RECT 586.800 539.400 588.600 545.400 ;
        RECT 565.950 528.450 568.050 529.050 ;
        RECT 571.950 528.450 574.050 529.050 ;
        RECT 565.950 527.550 574.050 528.450 ;
        RECT 565.950 526.950 568.050 527.550 ;
        RECT 571.950 526.950 574.050 527.550 ;
        RECT 580.800 526.050 582.000 533.400 ;
        RECT 587.400 532.500 588.600 539.400 ;
        RECT 582.900 531.600 588.600 532.500 ;
        RECT 590.550 533.400 592.350 545.400 ;
        RECT 598.050 539.400 599.850 545.400 ;
        RECT 595.950 537.300 599.850 539.400 ;
        RECT 605.850 538.500 607.650 545.400 ;
        RECT 613.650 539.400 615.450 545.400 ;
        RECT 614.250 538.500 615.450 539.400 ;
        RECT 604.950 537.450 611.550 538.500 ;
        RECT 604.950 536.700 606.750 537.450 ;
        RECT 609.750 536.700 611.550 537.450 ;
        RECT 614.250 536.400 619.050 538.500 ;
        RECT 597.150 534.600 599.850 536.400 ;
        RECT 600.750 535.800 602.550 536.400 ;
        RECT 600.750 534.900 607.050 535.800 ;
        RECT 614.250 535.500 615.450 536.400 ;
        RECT 600.750 534.600 602.550 534.900 ;
        RECT 598.950 533.700 599.850 534.600 ;
        RECT 582.900 530.700 584.850 531.600 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 328.950 523.950 331.050 526.050 ;
        RECT 331.950 523.950 334.050 526.050 ;
        RECT 334.950 523.950 337.050 526.050 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 355.950 523.950 358.050 526.050 ;
        RECT 358.950 523.950 361.050 526.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 379.950 523.950 382.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 433.950 523.950 436.050 526.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 439.950 523.950 442.050 526.050 ;
        RECT 442.950 523.950 445.050 526.050 ;
        RECT 460.950 523.950 463.050 526.050 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 478.950 523.950 481.050 526.050 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 499.950 523.950 502.050 526.050 ;
        RECT 502.950 523.950 505.050 526.050 ;
        RECT 505.950 523.950 508.050 526.050 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 523.950 523.950 526.050 526.050 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 529.950 523.950 532.050 526.050 ;
        RECT 544.950 523.950 547.050 526.050 ;
        RECT 547.950 523.950 550.050 526.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 580.800 523.950 583.050 526.050 ;
        RECT 305.550 521.550 310.050 523.050 ;
        RECT 306.000 520.950 310.050 521.550 ;
        RECT 273.000 519.000 276.300 520.200 ;
        RECT 297.000 519.000 300.300 520.200 ;
        RECT 251.400 510.600 253.200 513.600 ;
        RECT 273.000 510.600 274.800 519.000 ;
        RECT 297.000 510.600 298.800 519.000 ;
        RECT 314.700 513.600 315.600 523.950 ;
        RECT 329.100 522.150 330.900 523.950 ;
        RECT 334.950 516.600 336.000 523.950 ;
        RECT 341.100 522.150 342.900 523.950 ;
        RECT 356.100 522.150 357.900 523.950 ;
        RECT 337.950 519.450 340.050 520.050 ;
        RECT 352.950 519.450 355.050 520.050 ;
        RECT 337.950 518.550 355.050 519.450 ;
        RECT 337.950 517.950 340.050 518.550 ;
        RECT 352.950 517.950 355.050 518.550 ;
        RECT 314.400 510.600 316.200 513.600 ;
        RECT 334.200 510.600 336.000 516.600 ;
        RECT 359.400 516.600 360.600 523.950 ;
        RECT 374.100 522.150 375.900 523.950 ;
        RECT 377.400 518.700 378.600 523.950 ;
        RECT 380.100 522.150 381.900 523.950 ;
        RECT 374.400 517.800 378.600 518.700 ;
        RECT 359.400 510.600 361.200 516.600 ;
        RECT 374.400 510.600 376.200 517.800 ;
        RECT 395.400 513.600 396.600 523.950 ;
        RECT 413.100 522.150 414.900 523.950 ;
        RECT 416.400 518.700 417.600 523.950 ;
        RECT 419.100 522.150 420.900 523.950 ;
        RECT 431.100 522.150 432.900 523.950 ;
        RECT 413.400 517.800 417.600 518.700 ;
        RECT 395.400 510.600 397.200 513.600 ;
        RECT 413.400 510.600 415.200 517.800 ;
        RECT 436.950 516.600 438.000 523.950 ;
        RECT 443.100 522.150 444.900 523.950 ;
        RECT 461.100 522.150 462.900 523.950 ;
        RECT 463.950 519.750 465.150 523.950 ;
        RECT 467.100 522.150 468.900 523.950 ;
        RECT 479.100 522.150 480.900 523.950 ;
        RECT 461.400 518.700 465.150 519.750 ;
        RECT 482.400 518.700 483.600 523.950 ;
        RECT 485.100 522.150 486.900 523.950 ;
        RECT 500.100 522.150 501.900 523.950 ;
        RECT 503.850 519.750 505.050 523.950 ;
        RECT 506.100 522.150 507.900 523.950 ;
        RECT 524.100 522.150 525.900 523.950 ;
        RECT 527.850 519.750 529.050 523.950 ;
        RECT 530.100 522.150 531.900 523.950 ;
        RECT 503.850 518.700 507.600 519.750 ;
        RECT 527.850 518.700 531.600 519.750 ;
        RECT 461.400 516.600 462.600 518.700 ;
        RECT 482.400 517.800 486.600 518.700 ;
        RECT 436.200 510.600 438.000 516.600 ;
        RECT 460.800 510.600 462.600 516.600 ;
        RECT 463.800 515.700 471.600 517.050 ;
        RECT 463.800 510.600 465.600 515.700 ;
        RECT 469.800 510.600 471.600 515.700 ;
        RECT 484.800 510.600 486.600 517.800 ;
        RECT 497.400 515.700 505.200 517.050 ;
        RECT 497.400 510.600 499.200 515.700 ;
        RECT 503.400 510.600 505.200 515.700 ;
        RECT 506.400 516.600 507.600 518.700 ;
        RECT 506.400 510.600 508.200 516.600 ;
        RECT 521.400 515.700 529.200 517.050 ;
        RECT 521.400 510.600 523.200 515.700 ;
        RECT 527.400 510.600 529.200 515.700 ;
        RECT 530.400 516.600 531.600 518.700 ;
        RECT 530.400 510.600 532.200 516.600 ;
        RECT 545.400 513.600 546.600 523.950 ;
        RECT 544.800 510.600 546.600 513.600 ;
        RECT 563.400 513.600 564.600 523.950 ;
        RECT 580.800 516.600 582.000 523.950 ;
        RECT 583.950 519.300 584.850 530.700 ;
        RECT 587.100 526.050 588.900 527.850 ;
        RECT 590.550 526.050 591.750 533.400 ;
        RECT 595.950 532.800 598.050 533.700 ;
        RECT 598.950 532.800 604.050 533.700 ;
        RECT 593.850 531.600 598.050 532.800 ;
        RECT 592.950 529.800 594.750 531.600 ;
        RECT 586.950 523.950 589.050 526.050 ;
        RECT 590.550 525.750 595.050 526.050 ;
        RECT 590.550 523.950 596.850 525.750 ;
        RECT 582.900 518.400 584.850 519.300 ;
        RECT 582.900 517.500 588.600 518.400 ;
        RECT 563.400 510.600 565.200 513.600 ;
        RECT 580.800 510.600 582.600 516.600 ;
        RECT 587.400 513.600 588.600 517.500 ;
        RECT 586.800 510.600 588.600 513.600 ;
        RECT 590.550 516.600 591.750 523.950 ;
        RECT 603.150 520.200 604.050 532.800 ;
        RECT 606.150 532.800 607.050 534.900 ;
        RECT 607.950 534.300 615.450 535.500 ;
        RECT 607.950 533.700 609.750 534.300 ;
        RECT 622.050 533.400 623.850 545.400 ;
        RECT 606.150 532.500 614.550 532.800 ;
        RECT 622.950 532.500 623.850 533.400 ;
        RECT 606.150 531.900 623.850 532.500 ;
        RECT 612.750 531.300 623.850 531.900 ;
        RECT 612.750 531.000 614.550 531.300 ;
        RECT 610.950 524.400 613.050 526.050 ;
        RECT 610.950 523.200 618.900 524.400 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 617.100 522.600 618.900 523.200 ;
        RECT 620.100 522.150 621.900 523.950 ;
        RECT 614.100 521.400 615.900 522.000 ;
        RECT 620.100 521.400 621.000 522.150 ;
        RECT 614.100 520.200 621.000 521.400 ;
        RECT 603.150 519.000 615.150 520.200 ;
        RECT 603.150 518.400 604.950 519.000 ;
        RECT 614.100 517.200 615.150 519.000 ;
        RECT 590.550 510.600 592.350 516.600 ;
        RECT 595.950 515.700 598.050 516.600 ;
        RECT 595.950 514.500 599.700 515.700 ;
        RECT 610.350 515.550 612.150 516.300 ;
        RECT 598.650 513.600 599.700 514.500 ;
        RECT 607.200 514.500 612.150 515.550 ;
        RECT 613.650 515.400 615.450 517.200 ;
        RECT 622.950 516.600 623.850 531.300 ;
        RECT 616.950 514.500 619.050 516.600 ;
        RECT 607.200 513.600 608.250 514.500 ;
        RECT 616.950 513.600 618.000 514.500 ;
        RECT 598.650 510.600 600.450 513.600 ;
        RECT 606.450 510.600 608.250 513.600 ;
        RECT 614.250 512.700 618.000 513.600 ;
        RECT 614.250 510.600 616.050 512.700 ;
        RECT 622.050 510.600 623.850 516.600 ;
        RECT 637.800 533.400 639.600 545.400 ;
        RECT 643.800 539.400 645.600 545.400 ;
        RECT 637.800 526.050 639.000 533.400 ;
        RECT 644.400 532.500 645.600 539.400 ;
        RECT 639.900 531.600 645.600 532.500 ;
        RECT 655.800 533.400 657.600 545.400 ;
        RECT 661.800 539.400 663.600 545.400 ;
        RECT 676.800 539.400 678.600 545.400 ;
        RECT 639.900 530.700 641.850 531.600 ;
        RECT 637.800 523.950 640.050 526.050 ;
        RECT 637.800 516.600 639.000 523.950 ;
        RECT 640.950 519.300 641.850 530.700 ;
        RECT 644.100 526.050 645.900 527.850 ;
        RECT 655.800 526.050 657.000 533.400 ;
        RECT 662.400 532.500 663.600 539.400 ;
        RECT 657.900 531.600 663.600 532.500 ;
        RECT 657.900 530.700 659.850 531.600 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 655.800 523.950 658.050 526.050 ;
        RECT 639.900 518.400 641.850 519.300 ;
        RECT 639.900 517.500 645.600 518.400 ;
        RECT 637.800 510.600 639.600 516.600 ;
        RECT 644.400 513.600 645.600 517.500 ;
        RECT 643.800 510.600 645.600 513.600 ;
        RECT 655.800 516.600 657.000 523.950 ;
        RECT 658.950 519.300 659.850 530.700 ;
        RECT 669.000 528.450 673.050 529.050 ;
        RECT 662.100 526.050 663.900 527.850 ;
        RECT 668.550 526.950 673.050 528.450 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 668.550 523.050 669.450 526.950 ;
        RECT 677.400 526.050 678.600 539.400 ;
        RECT 683.550 533.400 685.350 545.400 ;
        RECT 691.050 539.400 692.850 545.400 ;
        RECT 688.950 537.300 692.850 539.400 ;
        RECT 698.850 538.500 700.650 545.400 ;
        RECT 706.650 539.400 708.450 545.400 ;
        RECT 707.250 538.500 708.450 539.400 ;
        RECT 697.950 537.450 704.550 538.500 ;
        RECT 697.950 536.700 699.750 537.450 ;
        RECT 702.750 536.700 704.550 537.450 ;
        RECT 707.250 536.400 712.050 538.500 ;
        RECT 690.150 534.600 692.850 536.400 ;
        RECT 693.750 535.800 695.550 536.400 ;
        RECT 693.750 534.900 700.050 535.800 ;
        RECT 707.250 535.500 708.450 536.400 ;
        RECT 693.750 534.600 695.550 534.900 ;
        RECT 691.950 533.700 692.850 534.600 ;
        RECT 683.550 526.050 684.750 533.400 ;
        RECT 688.950 532.800 691.050 533.700 ;
        RECT 691.950 532.800 697.050 533.700 ;
        RECT 686.850 531.600 691.050 532.800 ;
        RECT 685.950 529.800 687.750 531.600 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 683.550 525.750 688.050 526.050 ;
        RECT 683.550 523.950 689.850 525.750 ;
        RECT 664.950 521.550 669.450 523.050 ;
        RECT 674.100 522.150 675.900 523.950 ;
        RECT 664.950 520.950 669.000 521.550 ;
        RECT 657.900 518.400 659.850 519.300 ;
        RECT 677.400 518.700 678.600 523.950 ;
        RECT 680.100 522.150 681.900 523.950 ;
        RECT 657.900 517.500 663.600 518.400 ;
        RECT 655.800 510.600 657.600 516.600 ;
        RECT 662.400 513.600 663.600 517.500 ;
        RECT 661.800 510.600 663.600 513.600 ;
        RECT 674.400 517.800 678.600 518.700 ;
        RECT 674.400 510.600 676.200 517.800 ;
        RECT 683.550 516.600 684.750 523.950 ;
        RECT 696.150 520.200 697.050 532.800 ;
        RECT 699.150 532.800 700.050 534.900 ;
        RECT 700.950 534.300 708.450 535.500 ;
        RECT 700.950 533.700 702.750 534.300 ;
        RECT 715.050 533.400 716.850 545.400 ;
        RECT 699.150 532.500 707.550 532.800 ;
        RECT 715.950 532.500 716.850 533.400 ;
        RECT 699.150 531.900 716.850 532.500 ;
        RECT 705.750 531.300 716.850 531.900 ;
        RECT 705.750 531.000 707.550 531.300 ;
        RECT 703.950 524.400 706.050 526.050 ;
        RECT 703.950 523.200 711.900 524.400 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 710.100 522.600 711.900 523.200 ;
        RECT 713.100 522.150 714.900 523.950 ;
        RECT 707.100 521.400 708.900 522.000 ;
        RECT 713.100 521.400 714.000 522.150 ;
        RECT 707.100 520.200 714.000 521.400 ;
        RECT 696.150 519.000 708.150 520.200 ;
        RECT 696.150 518.400 697.950 519.000 ;
        RECT 707.100 517.200 708.150 519.000 ;
        RECT 683.550 510.600 685.350 516.600 ;
        RECT 688.950 515.700 691.050 516.600 ;
        RECT 688.950 514.500 692.700 515.700 ;
        RECT 703.350 515.550 705.150 516.300 ;
        RECT 691.650 513.600 692.700 514.500 ;
        RECT 700.200 514.500 705.150 515.550 ;
        RECT 706.650 515.400 708.450 517.200 ;
        RECT 715.950 516.600 716.850 531.300 ;
        RECT 709.950 514.500 712.050 516.600 ;
        RECT 700.200 513.600 701.250 514.500 ;
        RECT 709.950 513.600 711.000 514.500 ;
        RECT 691.650 510.600 693.450 513.600 ;
        RECT 699.450 510.600 701.250 513.600 ;
        RECT 707.250 512.700 711.000 513.600 ;
        RECT 707.250 510.600 709.050 512.700 ;
        RECT 715.050 510.600 716.850 516.600 ;
        RECT 719.550 533.400 721.350 545.400 ;
        RECT 727.050 539.400 728.850 545.400 ;
        RECT 724.950 537.300 728.850 539.400 ;
        RECT 734.850 538.500 736.650 545.400 ;
        RECT 742.650 539.400 744.450 545.400 ;
        RECT 743.250 538.500 744.450 539.400 ;
        RECT 733.950 537.450 740.550 538.500 ;
        RECT 733.950 536.700 735.750 537.450 ;
        RECT 738.750 536.700 740.550 537.450 ;
        RECT 743.250 536.400 748.050 538.500 ;
        RECT 726.150 534.600 728.850 536.400 ;
        RECT 729.750 535.800 731.550 536.400 ;
        RECT 729.750 534.900 736.050 535.800 ;
        RECT 743.250 535.500 744.450 536.400 ;
        RECT 729.750 534.600 731.550 534.900 ;
        RECT 727.950 533.700 728.850 534.600 ;
        RECT 719.550 526.050 720.750 533.400 ;
        RECT 724.950 532.800 727.050 533.700 ;
        RECT 727.950 532.800 733.050 533.700 ;
        RECT 722.850 531.600 727.050 532.800 ;
        RECT 721.950 529.800 723.750 531.600 ;
        RECT 719.550 525.750 724.050 526.050 ;
        RECT 719.550 523.950 725.850 525.750 ;
        RECT 719.550 516.600 720.750 523.950 ;
        RECT 732.150 520.200 733.050 532.800 ;
        RECT 735.150 532.800 736.050 534.900 ;
        RECT 736.950 534.300 744.450 535.500 ;
        RECT 736.950 533.700 738.750 534.300 ;
        RECT 751.050 533.400 752.850 545.400 ;
        RECT 735.150 532.500 743.550 532.800 ;
        RECT 751.950 532.500 752.850 533.400 ;
        RECT 735.150 531.900 752.850 532.500 ;
        RECT 741.750 531.300 752.850 531.900 ;
        RECT 741.750 531.000 743.550 531.300 ;
        RECT 739.950 524.400 742.050 526.050 ;
        RECT 739.950 523.200 747.900 524.400 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 746.100 522.600 747.900 523.200 ;
        RECT 749.100 522.150 750.900 523.950 ;
        RECT 743.100 521.400 744.900 522.000 ;
        RECT 749.100 521.400 750.000 522.150 ;
        RECT 743.100 520.200 750.000 521.400 ;
        RECT 732.150 519.000 744.150 520.200 ;
        RECT 732.150 518.400 733.950 519.000 ;
        RECT 743.100 517.200 744.150 519.000 ;
        RECT 719.550 510.600 721.350 516.600 ;
        RECT 724.950 515.700 727.050 516.600 ;
        RECT 724.950 514.500 728.700 515.700 ;
        RECT 739.350 515.550 741.150 516.300 ;
        RECT 727.650 513.600 728.700 514.500 ;
        RECT 736.200 514.500 741.150 515.550 ;
        RECT 742.650 515.400 744.450 517.200 ;
        RECT 751.950 516.600 752.850 531.300 ;
        RECT 745.950 514.500 748.050 516.600 ;
        RECT 736.200 513.600 737.250 514.500 ;
        RECT 745.950 513.600 747.000 514.500 ;
        RECT 727.650 510.600 729.450 513.600 ;
        RECT 735.450 510.600 737.250 513.600 ;
        RECT 743.250 512.700 747.000 513.600 ;
        RECT 743.250 510.600 745.050 512.700 ;
        RECT 751.050 510.600 752.850 516.600 ;
        RECT 755.550 533.400 757.350 545.400 ;
        RECT 763.050 539.400 764.850 545.400 ;
        RECT 760.950 537.300 764.850 539.400 ;
        RECT 770.850 538.500 772.650 545.400 ;
        RECT 778.650 539.400 780.450 545.400 ;
        RECT 779.250 538.500 780.450 539.400 ;
        RECT 769.950 537.450 776.550 538.500 ;
        RECT 769.950 536.700 771.750 537.450 ;
        RECT 774.750 536.700 776.550 537.450 ;
        RECT 779.250 536.400 784.050 538.500 ;
        RECT 762.150 534.600 764.850 536.400 ;
        RECT 765.750 535.800 767.550 536.400 ;
        RECT 765.750 534.900 772.050 535.800 ;
        RECT 779.250 535.500 780.450 536.400 ;
        RECT 765.750 534.600 767.550 534.900 ;
        RECT 763.950 533.700 764.850 534.600 ;
        RECT 755.550 526.050 756.750 533.400 ;
        RECT 760.950 532.800 763.050 533.700 ;
        RECT 763.950 532.800 769.050 533.700 ;
        RECT 758.850 531.600 763.050 532.800 ;
        RECT 757.950 529.800 759.750 531.600 ;
        RECT 755.550 525.750 760.050 526.050 ;
        RECT 755.550 523.950 761.850 525.750 ;
        RECT 755.550 516.600 756.750 523.950 ;
        RECT 768.150 520.200 769.050 532.800 ;
        RECT 771.150 532.800 772.050 534.900 ;
        RECT 772.950 534.300 780.450 535.500 ;
        RECT 772.950 533.700 774.750 534.300 ;
        RECT 787.050 533.400 788.850 545.400 ;
        RECT 802.800 539.400 804.600 545.400 ;
        RECT 771.150 532.500 779.550 532.800 ;
        RECT 787.950 532.500 788.850 533.400 ;
        RECT 771.150 531.900 788.850 532.500 ;
        RECT 777.750 531.300 788.850 531.900 ;
        RECT 777.750 531.000 779.550 531.300 ;
        RECT 775.950 524.400 778.050 526.050 ;
        RECT 775.950 523.200 783.900 524.400 ;
        RECT 784.950 523.950 787.050 526.050 ;
        RECT 782.100 522.600 783.900 523.200 ;
        RECT 785.100 522.150 786.900 523.950 ;
        RECT 779.100 521.400 780.900 522.000 ;
        RECT 785.100 521.400 786.000 522.150 ;
        RECT 779.100 520.200 786.000 521.400 ;
        RECT 768.150 519.000 780.150 520.200 ;
        RECT 768.150 518.400 769.950 519.000 ;
        RECT 779.100 517.200 780.150 519.000 ;
        RECT 755.550 510.600 757.350 516.600 ;
        RECT 760.950 515.700 763.050 516.600 ;
        RECT 760.950 514.500 764.700 515.700 ;
        RECT 775.350 515.550 777.150 516.300 ;
        RECT 763.650 513.600 764.700 514.500 ;
        RECT 772.200 514.500 777.150 515.550 ;
        RECT 778.650 515.400 780.450 517.200 ;
        RECT 787.950 516.600 788.850 531.300 ;
        RECT 798.000 528.450 802.050 529.050 ;
        RECT 797.550 526.950 802.050 528.450 ;
        RECT 797.550 523.050 798.450 526.950 ;
        RECT 803.400 526.050 804.600 539.400 ;
        RECT 818.400 539.400 820.200 545.400 ;
        RECT 836.400 539.400 838.200 545.400 ;
        RECT 806.100 526.050 807.900 527.850 ;
        RECT 818.400 526.050 819.600 539.400 ;
        RECT 836.700 539.100 838.200 539.400 ;
        RECT 842.400 539.400 844.200 545.400 ;
        RECT 862.800 539.400 864.600 545.400 ;
        RECT 886.800 539.400 888.600 545.400 ;
        RECT 904.800 539.400 906.600 545.400 ;
        RECT 842.400 539.100 843.300 539.400 ;
        RECT 836.700 538.200 843.300 539.100 ;
        RECT 820.950 531.450 823.050 532.050 ;
        RECT 829.950 531.450 832.050 532.050 ;
        RECT 820.950 530.550 832.050 531.450 ;
        RECT 820.950 529.950 823.050 530.550 ;
        RECT 829.950 529.950 832.050 530.550 ;
        RECT 836.100 526.050 837.900 527.850 ;
        RECT 842.400 526.050 843.300 538.200 ;
        RECT 856.950 531.450 859.050 532.050 ;
        RECT 848.550 530.550 859.050 531.450 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 805.950 523.950 808.050 526.050 ;
        RECT 814.950 523.950 817.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 832.950 523.950 835.050 526.050 ;
        RECT 835.950 523.950 838.050 526.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 797.550 521.550 802.050 523.050 ;
        RECT 798.000 520.950 802.050 521.550 ;
        RECT 781.950 514.500 784.050 516.600 ;
        RECT 772.200 513.600 773.250 514.500 ;
        RECT 781.950 513.600 783.000 514.500 ;
        RECT 763.650 510.600 765.450 513.600 ;
        RECT 771.450 510.600 773.250 513.600 ;
        RECT 779.250 512.700 783.000 513.600 ;
        RECT 779.250 510.600 781.050 512.700 ;
        RECT 787.050 510.600 788.850 516.600 ;
        RECT 803.400 513.600 804.600 523.950 ;
        RECT 815.100 522.150 816.900 523.950 ;
        RECT 818.400 518.700 819.600 523.950 ;
        RECT 821.100 522.150 822.900 523.950 ;
        RECT 833.100 522.150 834.900 523.950 ;
        RECT 839.100 522.150 840.900 523.950 ;
        RECT 842.400 520.200 843.300 523.950 ;
        RECT 848.550 523.050 849.450 530.550 ;
        RECT 856.950 529.950 859.050 530.550 ;
        RECT 857.100 526.050 858.900 527.850 ;
        RECT 862.950 526.050 864.150 539.400 ;
        RECT 887.400 526.050 888.600 539.400 ;
        RECT 905.700 539.100 906.600 539.400 ;
        RECT 910.800 539.400 912.600 545.400 ;
        RECT 910.800 539.100 912.300 539.400 ;
        RECT 905.700 538.200 912.300 539.100 ;
        RECT 901.950 528.450 904.050 529.050 ;
        RECT 896.550 527.550 904.050 528.450 ;
        RECT 856.950 523.950 859.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 883.950 523.950 886.050 526.050 ;
        RECT 886.950 523.950 889.050 526.050 ;
        RECT 889.950 523.950 892.050 526.050 ;
        RECT 844.950 521.550 849.450 523.050 ;
        RECT 860.100 522.150 861.900 523.950 ;
        RECT 844.950 520.950 849.000 521.550 ;
        RECT 840.000 519.000 843.300 520.200 ;
        RECT 863.850 519.750 865.050 523.950 ;
        RECT 866.100 522.150 867.900 523.950 ;
        RECT 884.100 522.150 885.900 523.950 ;
        RECT 818.400 517.800 822.600 518.700 ;
        RECT 802.800 510.600 804.600 513.600 ;
        RECT 820.800 510.600 822.600 517.800 ;
        RECT 840.000 510.600 841.800 519.000 ;
        RECT 863.850 518.700 867.600 519.750 ;
        RECT 887.400 518.700 888.600 523.950 ;
        RECT 890.100 522.150 891.900 523.950 ;
        RECT 896.550 523.050 897.450 527.550 ;
        RECT 901.950 526.950 904.050 527.550 ;
        RECT 905.700 526.050 906.600 538.200 ;
        RECT 911.100 526.050 912.900 527.850 ;
        RECT 904.950 523.950 907.050 526.050 ;
        RECT 907.950 523.950 910.050 526.050 ;
        RECT 910.950 523.950 913.050 526.050 ;
        RECT 913.950 523.950 916.050 526.050 ;
        RECT 892.950 521.550 897.450 523.050 ;
        RECT 892.950 520.950 897.000 521.550 ;
        RECT 905.700 520.200 906.600 523.950 ;
        RECT 908.100 522.150 909.900 523.950 ;
        RECT 914.100 522.150 915.900 523.950 ;
        RECT 905.700 519.000 909.000 520.200 ;
        RECT 857.400 515.700 865.200 517.050 ;
        RECT 857.400 510.600 859.200 515.700 ;
        RECT 863.400 510.600 865.200 515.700 ;
        RECT 866.400 516.600 867.600 518.700 ;
        RECT 884.400 517.800 888.600 518.700 ;
        RECT 866.400 510.600 868.200 516.600 ;
        RECT 884.400 510.600 886.200 517.800 ;
        RECT 907.200 510.600 909.000 519.000 ;
        RECT 11.400 501.300 13.200 506.400 ;
        RECT 17.400 501.300 19.200 506.400 ;
        RECT 11.400 499.950 19.200 501.300 ;
        RECT 20.400 500.400 22.200 506.400 ;
        RECT 20.400 498.300 21.600 500.400 ;
        RECT 17.850 497.250 21.600 498.300 ;
        RECT 37.200 498.000 39.000 506.400 ;
        RECT 58.500 501.600 60.300 506.400 ;
        RECT 58.500 500.400 63.600 501.600 ;
        RECT 14.100 493.050 15.900 494.850 ;
        RECT 17.850 493.050 19.050 497.250 ;
        RECT 35.700 496.800 39.000 498.000 ;
        RECT 20.100 493.050 21.900 494.850 ;
        RECT 35.700 493.050 36.600 496.800 ;
        RECT 38.100 493.050 39.900 494.850 ;
        RECT 44.100 493.050 45.900 494.850 ;
        RECT 53.100 493.050 54.900 494.850 ;
        RECT 59.100 493.050 60.900 494.850 ;
        RECT 62.700 493.050 63.600 500.400 ;
        RECT 84.000 498.000 85.800 506.400 ;
        RECT 103.200 498.000 105.000 506.400 ;
        RECT 122.400 501.300 124.200 506.400 ;
        RECT 128.400 501.300 130.200 506.400 ;
        RECT 122.400 499.950 130.200 501.300 ;
        RECT 131.400 500.400 133.200 506.400 ;
        RECT 153.000 500.400 154.800 506.400 ;
        RECT 171.300 502.200 173.100 506.400 ;
        RECT 170.400 500.400 173.100 502.200 ;
        RECT 131.400 498.300 132.600 500.400 ;
        RECT 84.000 496.800 87.300 498.000 ;
        RECT 77.100 493.050 78.900 494.850 ;
        RECT 83.100 493.050 84.900 494.850 ;
        RECT 86.400 493.050 87.300 496.800 ;
        RECT 101.700 496.800 105.000 498.000 ;
        RECT 128.850 497.250 132.600 498.300 ;
        RECT 88.950 495.450 93.000 496.050 ;
        RECT 96.000 495.450 100.050 496.050 ;
        RECT 88.950 493.950 93.450 495.450 ;
        RECT 10.950 490.950 13.050 493.050 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 19.950 490.950 22.050 493.050 ;
        RECT 34.950 490.950 37.050 493.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 55.950 490.950 58.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 61.950 490.950 64.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 11.100 489.150 12.900 490.950 ;
        RECT 16.950 477.600 18.150 490.950 ;
        RECT 35.700 478.800 36.600 490.950 ;
        RECT 41.100 489.150 42.900 490.950 ;
        RECT 56.100 489.150 57.900 490.950 ;
        RECT 62.700 483.600 63.600 490.950 ;
        RECT 80.100 489.150 81.900 490.950 ;
        RECT 67.950 486.450 70.050 487.050 ;
        RECT 76.950 486.450 79.050 487.050 ;
        RECT 67.950 485.550 79.050 486.450 ;
        RECT 67.950 484.950 70.050 485.550 ;
        RECT 76.950 484.950 79.050 485.550 ;
        RECT 53.400 482.700 61.200 483.600 ;
        RECT 35.700 477.900 42.300 478.800 ;
        RECT 35.700 477.600 36.600 477.900 ;
        RECT 16.800 471.600 18.600 477.600 ;
        RECT 34.800 471.600 36.600 477.600 ;
        RECT 40.800 477.600 42.300 477.900 ;
        RECT 40.800 471.600 42.600 477.600 ;
        RECT 53.400 471.600 55.200 482.700 ;
        RECT 59.400 471.600 61.200 482.700 ;
        RECT 62.400 471.600 64.200 483.600 ;
        RECT 86.400 478.800 87.300 490.950 ;
        RECT 92.550 490.050 93.450 493.950 ;
        RECT 88.950 488.550 93.450 490.050 ;
        RECT 95.550 493.950 100.050 495.450 ;
        RECT 88.950 487.950 93.000 488.550 ;
        RECT 95.550 487.050 96.450 493.950 ;
        RECT 101.700 493.050 102.600 496.800 ;
        RECT 112.950 495.450 117.000 496.050 ;
        RECT 104.100 493.050 105.900 494.850 ;
        RECT 110.100 493.050 111.900 494.850 ;
        RECT 112.950 493.950 117.450 495.450 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 94.950 484.950 97.050 487.050 ;
        RECT 80.700 477.900 87.300 478.800 ;
        RECT 80.700 477.600 82.200 477.900 ;
        RECT 80.400 471.600 82.200 477.600 ;
        RECT 86.400 477.600 87.300 477.900 ;
        RECT 101.700 478.800 102.600 490.950 ;
        RECT 107.100 489.150 108.900 490.950 ;
        RECT 116.550 490.050 117.450 493.950 ;
        RECT 125.100 493.050 126.900 494.850 ;
        RECT 128.850 493.050 130.050 497.250 ;
        RECT 131.100 493.050 132.900 494.850 ;
        RECT 146.100 493.050 147.900 494.850 ;
        RECT 153.000 493.050 154.050 500.400 ;
        RECT 158.100 493.050 159.900 494.850 ;
        RECT 170.400 493.050 171.300 500.400 ;
        RECT 173.100 498.600 174.900 499.500 ;
        RECT 178.800 498.600 180.600 506.400 ;
        RECT 196.800 499.200 198.600 506.400 ;
        RECT 173.100 497.700 180.600 498.600 ;
        RECT 194.400 498.300 198.600 499.200 ;
        RECT 121.950 490.950 124.050 493.050 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 127.950 490.950 130.050 493.050 ;
        RECT 130.950 490.950 133.050 493.050 ;
        RECT 145.950 490.950 148.050 493.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 157.950 490.950 160.050 493.050 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 112.950 488.550 117.450 490.050 ;
        RECT 122.100 489.150 123.900 490.950 ;
        RECT 112.950 487.950 117.000 488.550 ;
        RECT 101.700 477.900 108.300 478.800 ;
        RECT 101.700 477.600 102.600 477.900 ;
        RECT 86.400 471.600 88.200 477.600 ;
        RECT 100.800 471.600 102.600 477.600 ;
        RECT 106.800 477.600 108.300 477.900 ;
        RECT 127.950 477.600 129.150 490.950 ;
        RECT 149.100 489.150 150.900 490.950 ;
        RECT 153.000 485.400 153.900 490.950 ;
        RECT 155.100 489.150 156.900 490.950 ;
        RECT 148.800 484.500 153.900 485.400 ;
        RECT 106.800 471.600 108.600 477.600 ;
        RECT 127.800 471.600 129.600 477.600 ;
        RECT 145.800 472.500 147.600 483.600 ;
        RECT 148.800 473.400 150.600 484.500 ;
        RECT 170.400 483.600 171.300 490.950 ;
        RECT 173.100 489.150 174.900 490.950 ;
        RECT 151.800 482.400 159.600 483.300 ;
        RECT 151.800 472.500 153.600 482.400 ;
        RECT 145.800 471.600 153.600 472.500 ;
        RECT 157.800 471.600 159.600 482.400 ;
        RECT 169.800 471.600 171.600 483.600 ;
        RECT 176.700 477.600 177.600 497.700 ;
        RECT 179.100 493.050 180.900 494.850 ;
        RECT 191.100 493.050 192.900 494.850 ;
        RECT 194.400 493.050 195.600 498.300 ;
        RECT 217.200 498.000 219.000 506.400 ;
        RECT 235.800 503.400 237.600 506.400 ;
        RECT 215.700 496.800 219.000 498.000 ;
        RECT 197.100 493.050 198.900 494.850 ;
        RECT 215.700 493.050 216.600 496.800 ;
        RECT 231.000 495.450 235.050 496.050 ;
        RECT 218.100 493.050 219.900 494.850 ;
        RECT 224.100 493.050 225.900 494.850 ;
        RECT 230.550 493.950 235.050 495.450 ;
        RECT 178.950 490.950 181.050 493.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 178.950 486.450 181.050 487.050 ;
        RECT 190.950 486.450 193.050 487.050 ;
        RECT 178.950 485.550 193.050 486.450 ;
        RECT 178.950 484.950 181.050 485.550 ;
        RECT 190.950 484.950 193.050 485.550 ;
        RECT 175.800 471.600 177.600 477.600 ;
        RECT 194.400 477.600 195.600 490.950 ;
        RECT 215.700 478.800 216.600 490.950 ;
        RECT 221.100 489.150 222.900 490.950 ;
        RECT 230.550 490.050 231.450 493.950 ;
        RECT 236.400 493.050 237.600 503.400 ;
        RECT 253.800 500.400 255.600 506.400 ;
        RECT 254.400 498.300 255.600 500.400 ;
        RECT 256.800 501.300 258.600 506.400 ;
        RECT 262.800 501.300 264.600 506.400 ;
        RECT 256.800 499.950 264.600 501.300 ;
        RECT 277.800 500.400 279.600 506.400 ;
        RECT 278.400 498.300 279.600 500.400 ;
        RECT 280.800 501.300 282.600 506.400 ;
        RECT 286.800 501.300 288.600 506.400 ;
        RECT 300.300 502.200 302.100 506.400 ;
        RECT 280.800 499.950 288.600 501.300 ;
        RECT 299.400 500.400 302.100 502.200 ;
        RECT 254.400 497.250 258.150 498.300 ;
        RECT 278.400 497.250 282.150 498.300 ;
        RECT 241.950 495.450 246.000 496.050 ;
        RECT 241.950 493.950 246.450 495.450 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 230.550 488.550 235.050 490.050 ;
        RECT 231.000 487.950 235.050 488.550 ;
        RECT 215.700 477.900 222.300 478.800 ;
        RECT 215.700 477.600 216.600 477.900 ;
        RECT 194.400 471.600 196.200 477.600 ;
        RECT 214.800 471.600 216.600 477.600 ;
        RECT 220.800 477.600 222.300 477.900 ;
        RECT 236.400 477.600 237.600 490.950 ;
        RECT 239.100 489.150 240.900 490.950 ;
        RECT 245.550 486.450 246.450 493.950 ;
        RECT 254.100 493.050 255.900 494.850 ;
        RECT 256.950 493.050 258.150 497.250 ;
        RECT 260.100 493.050 261.900 494.850 ;
        RECT 278.100 493.050 279.900 494.850 ;
        RECT 280.950 493.050 282.150 497.250 ;
        RECT 289.950 495.450 294.000 496.050 ;
        RECT 284.100 493.050 285.900 494.850 ;
        RECT 289.950 493.950 294.450 495.450 ;
        RECT 253.950 490.950 256.050 493.050 ;
        RECT 256.950 490.950 259.050 493.050 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 277.950 490.950 280.050 493.050 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 286.950 490.950 289.050 493.050 ;
        RECT 253.950 486.450 256.050 487.050 ;
        RECT 245.550 485.550 256.050 486.450 ;
        RECT 253.950 484.950 256.050 485.550 ;
        RECT 257.850 477.600 259.050 490.950 ;
        RECT 263.100 489.150 264.900 490.950 ;
        RECT 281.850 477.600 283.050 490.950 ;
        RECT 287.100 489.150 288.900 490.950 ;
        RECT 293.550 490.050 294.450 493.950 ;
        RECT 299.400 493.050 300.300 500.400 ;
        RECT 302.100 498.600 303.900 499.500 ;
        RECT 307.800 498.600 309.600 506.400 ;
        RECT 322.800 499.200 324.600 506.400 ;
        RECT 341.400 503.400 343.200 506.400 ;
        RECT 302.100 497.700 309.600 498.600 ;
        RECT 320.400 498.300 324.600 499.200 ;
        RECT 342.300 499.200 343.200 503.400 ;
        RECT 347.400 500.400 349.200 506.400 ;
        RECT 342.300 498.300 345.600 499.200 ;
        RECT 298.950 490.950 301.050 493.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 289.950 488.550 294.450 490.050 ;
        RECT 289.950 487.950 294.000 488.550 ;
        RECT 299.400 483.600 300.300 490.950 ;
        RECT 302.100 489.150 303.900 490.950 ;
        RECT 220.800 471.600 222.600 477.600 ;
        RECT 235.800 471.600 237.600 477.600 ;
        RECT 257.400 471.600 259.200 477.600 ;
        RECT 281.400 471.600 283.200 477.600 ;
        RECT 298.800 471.600 300.600 483.600 ;
        RECT 305.700 477.600 306.600 497.700 ;
        RECT 308.100 493.050 309.900 494.850 ;
        RECT 317.100 493.050 318.900 494.850 ;
        RECT 320.400 493.050 321.600 498.300 ;
        RECT 343.800 497.400 345.600 498.300 ;
        RECT 323.100 493.050 324.900 494.850 ;
        RECT 338.100 493.050 339.900 494.850 ;
        RECT 307.950 490.950 310.050 493.050 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 304.800 471.600 306.600 477.600 ;
        RECT 320.400 477.600 321.600 490.950 ;
        RECT 341.100 489.150 342.900 490.950 ;
        RECT 344.700 486.900 345.600 497.400 ;
        RECT 348.000 493.050 349.050 500.400 ;
        RECT 367.800 499.200 369.600 506.400 ;
        RECT 373.950 504.450 376.050 505.050 ;
        RECT 382.950 504.450 385.050 505.050 ;
        RECT 373.950 503.550 385.050 504.450 ;
        RECT 373.950 502.950 376.050 503.550 ;
        RECT 382.950 502.950 385.050 503.550 ;
        RECT 354.000 498.450 358.050 499.050 ;
        RECT 343.800 486.300 345.600 486.900 ;
        RECT 338.400 485.100 345.600 486.300 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 353.550 496.950 358.050 498.450 ;
        RECT 365.400 498.300 369.600 499.200 ;
        RECT 386.400 499.200 388.200 506.400 ;
        RECT 407.400 503.400 409.200 506.400 ;
        RECT 386.400 498.300 390.600 499.200 ;
        RECT 338.400 483.600 339.600 485.100 ;
        RECT 346.950 483.600 348.300 490.950 ;
        RECT 353.550 489.450 354.450 496.950 ;
        RECT 357.000 495.450 361.050 496.050 ;
        RECT 350.550 488.550 354.450 489.450 ;
        RECT 356.550 493.950 361.050 495.450 ;
        RECT 356.550 490.050 357.450 493.950 ;
        RECT 362.100 493.050 363.900 494.850 ;
        RECT 365.400 493.050 366.600 498.300 ;
        RECT 368.100 493.050 369.900 494.850 ;
        RECT 386.100 493.050 387.900 494.850 ;
        RECT 389.400 493.050 390.600 498.300 ;
        RECT 394.950 495.450 399.000 496.050 ;
        RECT 392.100 493.050 393.900 494.850 ;
        RECT 394.950 493.950 399.450 495.450 ;
        RECT 361.950 490.950 364.050 493.050 ;
        RECT 364.950 490.950 367.050 493.050 ;
        RECT 367.950 490.950 370.050 493.050 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 388.950 490.950 391.050 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 356.550 488.550 361.050 490.050 ;
        RECT 350.550 487.050 351.450 488.550 ;
        RECT 357.000 487.950 361.050 488.550 ;
        RECT 349.950 486.450 352.050 487.050 ;
        RECT 361.950 486.450 364.050 487.050 ;
        RECT 349.950 485.550 364.050 486.450 ;
        RECT 349.950 484.950 352.050 485.550 ;
        RECT 361.950 484.950 364.050 485.550 ;
        RECT 320.400 471.600 322.200 477.600 ;
        RECT 338.400 471.600 340.200 483.600 ;
        RECT 345.900 482.100 348.300 483.600 ;
        RECT 345.900 471.600 347.700 482.100 ;
        RECT 365.400 477.600 366.600 490.950 ;
        RECT 373.950 486.450 376.050 487.050 ;
        RECT 382.950 486.450 385.050 486.750 ;
        RECT 373.950 485.550 385.050 486.450 ;
        RECT 373.950 484.950 376.050 485.550 ;
        RECT 382.950 484.650 385.050 485.550 ;
        RECT 389.400 477.600 390.600 490.950 ;
        RECT 398.550 490.050 399.450 493.950 ;
        RECT 407.400 493.050 408.600 503.400 ;
        RECT 427.800 499.200 429.600 506.400 ;
        RECT 448.800 499.200 450.600 506.400 ;
        RECT 454.950 502.950 457.050 505.050 ;
        RECT 425.400 498.300 429.600 499.200 ;
        RECT 446.400 498.300 450.600 499.200 ;
        RECT 455.550 499.050 456.450 502.950 ;
        RECT 461.400 501.300 463.200 506.400 ;
        RECT 467.400 501.300 469.200 506.400 ;
        RECT 461.400 499.950 469.200 501.300 ;
        RECT 470.400 500.400 472.200 506.400 ;
        RECT 491.700 501.600 493.500 506.400 ;
        RECT 488.400 500.400 493.500 501.600 ;
        RECT 514.500 501.600 516.300 506.400 ;
        RECT 536.400 503.400 538.200 506.400 ;
        RECT 514.500 500.400 519.600 501.600 ;
        RECT 422.100 493.050 423.900 494.850 ;
        RECT 425.400 493.050 426.600 498.300 ;
        RECT 430.950 495.450 435.000 496.050 ;
        RECT 428.100 493.050 429.900 494.850 ;
        RECT 430.950 493.950 435.450 495.450 ;
        RECT 403.950 490.950 406.050 493.050 ;
        RECT 406.950 490.950 409.050 493.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 434.550 492.450 435.450 493.950 ;
        RECT 443.100 493.050 444.900 494.850 ;
        RECT 446.400 493.050 447.600 498.300 ;
        RECT 454.950 496.950 457.050 499.050 ;
        RECT 470.400 498.300 471.600 500.400 ;
        RECT 467.850 497.250 471.600 498.300 ;
        RECT 449.100 493.050 450.900 494.850 ;
        RECT 464.100 493.050 465.900 494.850 ;
        RECT 467.850 493.050 469.050 497.250 ;
        RECT 470.100 493.050 471.900 494.850 ;
        RECT 488.400 493.050 489.300 500.400 ;
        RECT 491.100 493.050 492.900 494.850 ;
        RECT 497.100 493.050 498.900 494.850 ;
        RECT 509.100 493.050 510.900 494.850 ;
        RECT 515.100 493.050 516.900 494.850 ;
        RECT 518.700 493.050 519.600 500.400 ;
        RECT 536.400 493.050 537.600 503.400 ;
        RECT 558.000 498.000 559.800 506.400 ;
        RECT 578.700 501.600 580.500 506.400 ;
        RECT 575.400 500.400 580.500 501.600 ;
        RECT 558.000 496.800 561.300 498.000 ;
        RECT 551.100 493.050 552.900 494.850 ;
        RECT 557.100 493.050 558.900 494.850 ;
        RECT 560.400 493.050 561.300 496.800 ;
        RECT 575.400 493.050 576.300 500.400 ;
        RECT 603.000 498.000 604.800 506.400 ;
        RECT 627.000 498.000 628.800 506.400 ;
        RECT 644.400 503.400 646.200 506.400 ;
        RECT 644.400 499.500 645.600 503.400 ;
        RECT 650.400 500.400 652.200 506.400 ;
        RECT 644.400 498.600 650.100 499.500 ;
        RECT 603.000 496.800 606.300 498.000 ;
        RECT 627.000 496.800 630.300 498.000 ;
        RECT 578.100 493.050 579.900 494.850 ;
        RECT 584.100 493.050 585.900 494.850 ;
        RECT 596.100 493.050 597.900 494.850 ;
        RECT 602.100 493.050 603.900 494.850 ;
        RECT 605.400 493.050 606.300 496.800 ;
        RECT 607.950 495.450 612.000 496.050 ;
        RECT 607.950 493.950 612.450 495.450 ;
        RECT 434.550 491.550 438.450 492.450 ;
        RECT 394.950 488.550 399.450 490.050 ;
        RECT 404.100 489.150 405.900 490.950 ;
        RECT 394.950 487.950 399.000 488.550 ;
        RECT 365.400 471.600 367.200 477.600 ;
        RECT 388.800 471.600 390.600 477.600 ;
        RECT 407.400 477.600 408.600 490.950 ;
        RECT 425.400 477.600 426.600 490.950 ;
        RECT 437.550 490.050 438.450 491.550 ;
        RECT 442.950 490.950 445.050 493.050 ;
        RECT 445.950 490.950 448.050 493.050 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 466.950 490.950 469.050 493.050 ;
        RECT 469.950 490.950 472.050 493.050 ;
        RECT 487.950 490.950 490.050 493.050 ;
        RECT 490.950 490.950 493.050 493.050 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 508.950 490.950 511.050 493.050 ;
        RECT 511.950 490.950 514.050 493.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 556.950 490.950 559.050 493.050 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 574.950 490.950 577.050 493.050 ;
        RECT 577.950 490.950 580.050 493.050 ;
        RECT 580.950 490.950 583.050 493.050 ;
        RECT 583.950 490.950 586.050 493.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 598.950 490.950 601.050 493.050 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 604.950 490.950 607.050 493.050 ;
        RECT 437.550 488.550 442.050 490.050 ;
        RECT 438.000 487.950 442.050 488.550 ;
        RECT 446.400 477.600 447.600 490.950 ;
        RECT 461.100 489.150 462.900 490.950 ;
        RECT 466.950 477.600 468.150 490.950 ;
        RECT 488.400 483.600 489.300 490.950 ;
        RECT 494.100 489.150 495.900 490.950 ;
        RECT 512.100 489.150 513.900 490.950 ;
        RECT 518.700 483.600 519.600 490.950 ;
        RECT 533.100 489.150 534.900 490.950 ;
        RECT 407.400 471.600 409.200 477.600 ;
        RECT 425.400 471.600 427.200 477.600 ;
        RECT 446.400 471.600 448.200 477.600 ;
        RECT 466.800 471.600 468.600 477.600 ;
        RECT 487.800 471.600 489.600 483.600 ;
        RECT 490.800 482.700 498.600 483.600 ;
        RECT 490.800 471.600 492.600 482.700 ;
        RECT 496.800 471.600 498.600 482.700 ;
        RECT 509.400 482.700 517.200 483.600 ;
        RECT 509.400 471.600 511.200 482.700 ;
        RECT 515.400 471.600 517.200 482.700 ;
        RECT 518.400 471.600 520.200 483.600 ;
        RECT 536.400 477.600 537.600 490.950 ;
        RECT 554.100 489.150 555.900 490.950 ;
        RECT 560.400 478.800 561.300 490.950 ;
        RECT 575.400 483.600 576.300 490.950 ;
        RECT 581.100 489.150 582.900 490.950 ;
        RECT 599.100 489.150 600.900 490.950 ;
        RECT 580.950 486.450 583.050 487.050 ;
        RECT 598.950 486.450 601.050 487.050 ;
        RECT 580.950 485.550 601.050 486.450 ;
        RECT 580.950 484.950 583.050 485.550 ;
        RECT 598.950 484.950 601.050 485.550 ;
        RECT 554.700 477.900 561.300 478.800 ;
        RECT 554.700 477.600 556.200 477.900 ;
        RECT 536.400 471.600 538.200 477.600 ;
        RECT 554.400 471.600 556.200 477.600 ;
        RECT 560.400 477.600 561.300 477.900 ;
        RECT 560.400 471.600 562.200 477.600 ;
        RECT 574.800 471.600 576.600 483.600 ;
        RECT 577.800 482.700 585.600 483.600 ;
        RECT 577.800 471.600 579.600 482.700 ;
        RECT 583.800 471.600 585.600 482.700 ;
        RECT 605.400 478.800 606.300 490.950 ;
        RECT 611.550 490.050 612.450 493.950 ;
        RECT 620.100 493.050 621.900 494.850 ;
        RECT 626.100 493.050 627.900 494.850 ;
        RECT 629.400 493.050 630.300 496.800 ;
        RECT 648.150 497.700 650.100 498.600 ;
        RECT 619.950 490.950 622.050 493.050 ;
        RECT 622.950 490.950 625.050 493.050 ;
        RECT 625.950 490.950 628.050 493.050 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 643.950 490.950 646.050 493.050 ;
        RECT 607.950 488.550 612.450 490.050 ;
        RECT 623.100 489.150 624.900 490.950 ;
        RECT 607.950 487.950 612.000 488.550 ;
        RECT 629.400 478.800 630.300 490.950 ;
        RECT 644.100 489.150 645.900 490.950 ;
        RECT 648.150 486.300 649.050 497.700 ;
        RECT 651.000 493.050 652.200 500.400 ;
        RECT 668.400 499.200 670.200 506.400 ;
        RECT 686.400 501.300 688.200 506.400 ;
        RECT 692.400 501.300 694.200 506.400 ;
        RECT 686.400 499.950 694.200 501.300 ;
        RECT 695.400 500.400 697.200 506.400 ;
        RECT 710.400 501.300 712.200 506.400 ;
        RECT 716.400 501.300 718.200 506.400 ;
        RECT 668.400 498.300 672.600 499.200 ;
        RECT 695.400 498.300 696.600 500.400 ;
        RECT 710.400 499.950 718.200 501.300 ;
        RECT 719.400 500.400 721.200 506.400 ;
        RECT 719.400 498.300 720.600 500.400 ;
        RECT 739.800 499.200 741.600 506.400 ;
        RECT 758.400 503.400 760.200 506.400 ;
        RECT 668.100 493.050 669.900 494.850 ;
        RECT 671.400 493.050 672.600 498.300 ;
        RECT 692.850 497.250 696.600 498.300 ;
        RECT 716.850 497.250 720.600 498.300 ;
        RECT 737.400 498.300 741.600 499.200 ;
        RECT 674.100 493.050 675.900 494.850 ;
        RECT 689.100 493.050 690.900 494.850 ;
        RECT 692.850 493.050 694.050 497.250 ;
        RECT 695.100 493.050 696.900 494.850 ;
        RECT 713.100 493.050 714.900 494.850 ;
        RECT 716.850 493.050 718.050 497.250 ;
        RECT 730.950 495.450 733.050 496.050 ;
        RECT 719.100 493.050 720.900 494.850 ;
        RECT 725.550 494.550 733.050 495.450 ;
        RECT 649.950 490.950 652.200 493.050 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 673.950 490.950 676.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 691.950 490.950 694.050 493.050 ;
        RECT 694.950 490.950 697.050 493.050 ;
        RECT 709.950 490.950 712.050 493.050 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 715.950 490.950 718.050 493.050 ;
        RECT 718.950 490.950 721.050 493.050 ;
        RECT 648.150 485.400 650.100 486.300 ;
        RECT 599.700 477.900 606.300 478.800 ;
        RECT 599.700 477.600 601.200 477.900 ;
        RECT 599.400 471.600 601.200 477.600 ;
        RECT 605.400 477.600 606.300 477.900 ;
        RECT 623.700 477.900 630.300 478.800 ;
        RECT 623.700 477.600 625.200 477.900 ;
        RECT 605.400 471.600 607.200 477.600 ;
        RECT 623.400 471.600 625.200 477.600 ;
        RECT 629.400 477.600 630.300 477.900 ;
        RECT 644.400 484.500 650.100 485.400 ;
        RECT 644.400 477.600 645.600 484.500 ;
        RECT 651.000 483.600 652.200 490.950 ;
        RECT 660.000 489.450 664.050 490.050 ;
        RECT 659.550 487.950 664.050 489.450 ;
        RECT 659.550 483.900 660.450 487.950 ;
        RECT 661.950 486.450 664.050 486.900 ;
        RECT 667.950 486.450 670.050 487.050 ;
        RECT 661.950 485.550 670.050 486.450 ;
        RECT 661.950 484.800 664.050 485.550 ;
        RECT 667.950 484.950 670.050 485.550 ;
        RECT 629.400 471.600 631.200 477.600 ;
        RECT 644.400 471.600 646.200 477.600 ;
        RECT 650.400 471.600 652.200 483.600 ;
        RECT 658.950 481.800 661.050 483.900 ;
        RECT 671.400 477.600 672.600 490.950 ;
        RECT 686.100 489.150 687.900 490.950 ;
        RECT 691.950 477.600 693.150 490.950 ;
        RECT 710.100 489.150 711.900 490.950 ;
        RECT 715.950 477.600 717.150 490.950 ;
        RECT 725.550 490.050 726.450 494.550 ;
        RECT 730.950 493.950 733.050 494.550 ;
        RECT 734.100 493.050 735.900 494.850 ;
        RECT 737.400 493.050 738.600 498.300 ;
        RECT 740.100 493.050 741.900 494.850 ;
        RECT 758.700 493.050 759.600 503.400 ;
        RECT 778.800 500.400 780.600 506.400 ;
        RECT 772.950 496.950 775.050 499.050 ;
        RECT 779.400 498.300 780.600 500.400 ;
        RECT 781.800 501.300 783.600 506.400 ;
        RECT 787.800 501.300 789.600 506.400 ;
        RECT 781.800 499.950 789.600 501.300 ;
        RECT 797.400 503.400 799.200 506.400 ;
        RECT 797.400 499.500 798.600 503.400 ;
        RECT 803.400 500.400 805.200 506.400 ;
        RECT 797.400 498.600 803.100 499.500 ;
        RECT 779.400 497.250 783.150 498.300 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 754.950 490.950 757.050 493.050 ;
        RECT 757.950 490.950 760.050 493.050 ;
        RECT 760.950 490.950 763.050 493.050 ;
        RECT 721.950 488.550 726.450 490.050 ;
        RECT 721.950 487.950 726.000 488.550 ;
        RECT 737.400 477.600 738.600 490.950 ;
        RECT 755.100 489.150 756.900 490.950 ;
        RECT 739.950 486.450 742.050 487.050 ;
        RECT 751.950 486.450 754.050 487.050 ;
        RECT 739.950 485.550 754.050 486.450 ;
        RECT 739.950 484.950 742.050 485.550 ;
        RECT 751.950 484.950 754.050 485.550 ;
        RECT 758.700 483.600 759.600 490.950 ;
        RECT 761.100 489.150 762.900 490.950 ;
        RECT 763.950 489.450 766.050 490.050 ;
        RECT 773.550 489.450 774.450 496.950 ;
        RECT 779.100 493.050 780.900 494.850 ;
        RECT 781.950 493.050 783.150 497.250 ;
        RECT 801.150 497.700 803.100 498.600 ;
        RECT 785.100 493.050 786.900 494.850 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 763.950 488.550 774.450 489.450 ;
        RECT 763.950 487.950 766.050 488.550 ;
        RECT 758.700 482.400 762.300 483.600 ;
        RECT 670.800 471.600 672.600 477.600 ;
        RECT 691.800 471.600 693.600 477.600 ;
        RECT 715.800 471.600 717.600 477.600 ;
        RECT 737.400 471.600 739.200 477.600 ;
        RECT 760.500 471.600 762.300 482.400 ;
        RECT 782.850 477.600 784.050 490.950 ;
        RECT 788.100 489.150 789.900 490.950 ;
        RECT 797.100 489.150 798.900 490.950 ;
        RECT 801.150 486.300 802.050 497.700 ;
        RECT 804.000 493.050 805.200 500.400 ;
        RECT 818.400 501.300 820.200 506.400 ;
        RECT 824.400 501.300 826.200 506.400 ;
        RECT 818.400 499.950 826.200 501.300 ;
        RECT 827.400 500.400 829.200 506.400 ;
        RECT 827.400 498.300 828.600 500.400 ;
        RECT 844.800 499.200 846.600 506.400 ;
        RECT 863.400 503.400 865.200 506.400 ;
        RECT 824.850 497.250 828.600 498.300 ;
        RECT 842.400 498.300 846.600 499.200 ;
        RECT 821.100 493.050 822.900 494.850 ;
        RECT 824.850 493.050 826.050 497.250 ;
        RECT 829.950 495.450 834.000 496.050 ;
        RECT 827.100 493.050 828.900 494.850 ;
        RECT 829.950 493.950 834.450 495.450 ;
        RECT 802.950 490.950 805.200 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 823.950 490.950 826.050 493.050 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 801.150 485.400 803.100 486.300 ;
        RECT 797.400 484.500 803.100 485.400 ;
        RECT 797.400 477.600 798.600 484.500 ;
        RECT 804.000 483.600 805.200 490.950 ;
        RECT 818.100 489.150 819.900 490.950 ;
        RECT 782.400 471.600 784.200 477.600 ;
        RECT 797.400 471.600 799.200 477.600 ;
        RECT 803.400 471.600 805.200 483.600 ;
        RECT 823.950 477.600 825.150 490.950 ;
        RECT 833.550 490.050 834.450 493.950 ;
        RECT 839.100 493.050 840.900 494.850 ;
        RECT 842.400 493.050 843.600 498.300 ;
        RECT 845.100 493.050 846.900 494.850 ;
        RECT 863.700 493.050 864.600 503.400 ;
        RECT 888.000 498.000 889.800 506.400 ;
        RECT 905.400 499.200 907.200 506.400 ;
        RECT 905.400 498.300 909.600 499.200 ;
        RECT 888.000 496.800 891.300 498.000 ;
        RECT 881.100 493.050 882.900 494.850 ;
        RECT 887.100 493.050 888.900 494.850 ;
        RECT 890.400 493.050 891.300 496.800 ;
        RECT 892.950 495.450 895.050 495.900 ;
        RECT 892.950 494.550 900.450 495.450 ;
        RECT 892.950 493.800 895.050 494.550 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 844.950 490.950 847.050 493.050 ;
        RECT 859.950 490.950 862.050 493.050 ;
        RECT 862.950 490.950 865.050 493.050 ;
        RECT 865.950 490.950 868.050 493.050 ;
        RECT 880.950 490.950 883.050 493.050 ;
        RECT 883.950 490.950 886.050 493.050 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 889.950 490.950 892.050 493.050 ;
        RECT 829.950 488.550 834.450 490.050 ;
        RECT 829.950 487.950 834.000 488.550 ;
        RECT 842.400 477.600 843.600 490.950 ;
        RECT 860.100 489.150 861.900 490.950 ;
        RECT 863.700 483.600 864.600 490.950 ;
        RECT 866.100 489.150 867.900 490.950 ;
        RECT 884.100 489.150 885.900 490.950 ;
        RECT 863.700 482.400 867.300 483.600 ;
        RECT 823.800 471.600 825.600 477.600 ;
        RECT 842.400 471.600 844.200 477.600 ;
        RECT 865.500 471.600 867.300 482.400 ;
        RECT 890.400 478.800 891.300 490.950 ;
        RECT 899.550 489.450 900.450 494.550 ;
        RECT 905.100 493.050 906.900 494.850 ;
        RECT 908.400 493.050 909.600 498.300 ;
        RECT 911.100 493.050 912.900 494.850 ;
        RECT 904.950 490.950 907.050 493.050 ;
        RECT 907.950 490.950 910.050 493.050 ;
        RECT 910.950 490.950 913.050 493.050 ;
        RECT 899.550 488.550 903.450 489.450 ;
        RECT 902.550 486.450 903.450 488.550 ;
        RECT 902.550 486.000 906.450 486.450 ;
        RECT 902.550 485.550 907.050 486.000 ;
        RECT 904.950 481.800 907.050 485.550 ;
        RECT 884.700 477.900 891.300 478.800 ;
        RECT 884.700 477.600 886.200 477.900 ;
        RECT 884.400 471.600 886.200 477.600 ;
        RECT 890.400 477.600 891.300 477.900 ;
        RECT 908.400 477.600 909.600 490.950 ;
        RECT 890.400 471.600 892.200 477.600 ;
        RECT 907.800 471.600 909.600 477.600 ;
        RECT 16.800 461.400 18.600 467.400 ;
        RECT 37.800 461.400 39.600 467.400 ;
        RECT 11.100 448.050 12.900 449.850 ;
        RECT 16.950 448.050 18.150 461.400 ;
        RECT 38.700 461.100 39.600 461.400 ;
        RECT 43.800 461.400 45.600 467.400 ;
        RECT 43.800 461.100 45.300 461.400 ;
        RECT 38.700 460.200 45.300 461.100 ;
        RECT 38.700 448.050 39.600 460.200 ;
        RECT 59.400 456.300 61.200 467.400 ;
        RECT 65.400 456.300 67.200 467.400 ;
        RECT 59.400 455.400 67.200 456.300 ;
        RECT 68.400 455.400 70.200 467.400 ;
        RECT 83.400 456.300 85.200 467.400 ;
        RECT 89.400 456.300 91.200 467.400 ;
        RECT 83.400 455.400 91.200 456.300 ;
        RECT 92.400 455.400 94.200 467.400 ;
        RECT 110.400 461.400 112.200 467.400 ;
        RECT 134.400 461.400 136.200 467.400 ;
        RECT 154.800 461.400 156.600 467.400 ;
        RECT 40.950 453.450 43.050 454.050 ;
        RECT 58.950 453.450 61.050 454.050 ;
        RECT 40.950 452.550 61.050 453.450 ;
        RECT 40.950 451.950 43.050 452.550 ;
        RECT 58.950 451.950 61.050 452.550 ;
        RECT 44.100 448.050 45.900 449.850 ;
        RECT 62.100 448.050 63.900 449.850 ;
        RECT 68.700 448.050 69.600 455.400 ;
        RECT 86.100 448.050 87.900 449.850 ;
        RECT 92.700 448.050 93.600 455.400 ;
        RECT 110.850 448.050 112.050 461.400 ;
        RECT 116.100 448.050 117.900 449.850 ;
        RECT 134.850 448.050 136.050 461.400 ;
        RECT 140.100 448.050 141.900 449.850 ;
        RECT 149.100 448.050 150.900 449.850 ;
        RECT 154.950 448.050 156.150 461.400 ;
        RECT 170.400 456.300 172.200 467.400 ;
        RECT 176.400 456.300 178.200 467.400 ;
        RECT 170.400 455.400 178.200 456.300 ;
        RECT 179.400 455.400 181.200 467.400 ;
        RECT 197.400 461.400 199.200 467.400 ;
        RECT 214.800 461.400 216.600 467.400 ;
        RECT 160.950 450.450 165.000 451.050 ;
        RECT 160.950 448.950 165.450 450.450 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 37.950 445.950 40.050 448.050 ;
        RECT 40.950 445.950 43.050 448.050 ;
        RECT 43.950 445.950 46.050 448.050 ;
        RECT 46.950 445.950 49.050 448.050 ;
        RECT 58.950 445.950 61.050 448.050 ;
        RECT 61.950 445.950 64.050 448.050 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 67.950 445.950 70.050 448.050 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 91.950 445.950 94.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 133.950 445.950 136.050 448.050 ;
        RECT 136.950 445.950 139.050 448.050 ;
        RECT 139.950 445.950 142.050 448.050 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 151.950 445.950 154.050 448.050 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 14.100 444.150 15.900 445.950 ;
        RECT 17.850 441.750 19.050 445.950 ;
        RECT 20.100 444.150 21.900 445.950 ;
        RECT 38.700 442.200 39.600 445.950 ;
        RECT 41.100 444.150 42.900 445.950 ;
        RECT 47.100 444.150 48.900 445.950 ;
        RECT 59.100 444.150 60.900 445.950 ;
        RECT 65.100 444.150 66.900 445.950 ;
        RECT 17.850 440.700 21.600 441.750 ;
        RECT 38.700 441.000 42.000 442.200 ;
        RECT 11.400 437.700 19.200 439.050 ;
        RECT 11.400 432.600 13.200 437.700 ;
        RECT 17.400 432.600 19.200 437.700 ;
        RECT 20.400 438.600 21.600 440.700 ;
        RECT 20.400 432.600 22.200 438.600 ;
        RECT 40.200 432.600 42.000 441.000 ;
        RECT 68.700 438.600 69.600 445.950 ;
        RECT 83.100 444.150 84.900 445.950 ;
        RECT 89.100 444.150 90.900 445.950 ;
        RECT 92.700 438.600 93.600 445.950 ;
        RECT 107.100 444.150 108.900 445.950 ;
        RECT 109.950 441.750 111.150 445.950 ;
        RECT 113.100 444.150 114.900 445.950 ;
        RECT 118.950 444.450 121.050 445.050 ;
        RECT 127.950 444.450 130.050 445.050 ;
        RECT 118.950 443.550 130.050 444.450 ;
        RECT 131.100 444.150 132.900 445.950 ;
        RECT 118.950 442.950 121.050 443.550 ;
        RECT 127.950 442.950 130.050 443.550 ;
        RECT 133.950 441.750 135.150 445.950 ;
        RECT 137.100 444.150 138.900 445.950 ;
        RECT 152.100 444.150 153.900 445.950 ;
        RECT 107.400 440.700 111.150 441.750 ;
        RECT 131.400 440.700 135.150 441.750 ;
        RECT 155.850 441.750 157.050 445.950 ;
        RECT 158.100 444.150 159.900 445.950 ;
        RECT 164.550 445.050 165.450 448.950 ;
        RECT 173.100 448.050 174.900 449.850 ;
        RECT 179.700 448.050 180.600 455.400 ;
        RECT 194.100 448.050 195.900 449.850 ;
        RECT 197.400 448.050 198.600 461.400 ;
        RECT 215.700 461.100 216.600 461.400 ;
        RECT 220.800 461.400 222.600 467.400 ;
        RECT 220.800 461.100 222.300 461.400 ;
        RECT 215.700 460.200 222.300 461.100 ;
        RECT 211.950 450.450 214.050 451.050 ;
        RECT 203.550 449.550 214.050 450.450 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 172.950 445.950 175.050 448.050 ;
        RECT 175.950 445.950 178.050 448.050 ;
        RECT 178.950 445.950 181.050 448.050 ;
        RECT 193.950 445.950 196.050 448.050 ;
        RECT 196.950 445.950 199.050 448.050 ;
        RECT 160.950 443.550 165.450 445.050 ;
        RECT 170.100 444.150 171.900 445.950 ;
        RECT 176.100 444.150 177.900 445.950 ;
        RECT 160.950 442.950 165.000 443.550 ;
        RECT 155.850 440.700 159.600 441.750 ;
        RECT 107.400 438.600 108.600 440.700 ;
        RECT 64.500 437.400 69.600 438.600 ;
        RECT 88.500 437.400 93.600 438.600 ;
        RECT 64.500 432.600 66.300 437.400 ;
        RECT 88.500 432.600 90.300 437.400 ;
        RECT 106.800 432.600 108.600 438.600 ;
        RECT 109.800 437.700 117.600 439.050 ;
        RECT 131.400 438.600 132.600 440.700 ;
        RECT 109.800 432.600 111.600 437.700 ;
        RECT 115.800 432.600 117.600 437.700 ;
        RECT 130.800 432.600 132.600 438.600 ;
        RECT 133.800 437.700 141.600 439.050 ;
        RECT 133.800 432.600 135.600 437.700 ;
        RECT 139.800 432.600 141.600 437.700 ;
        RECT 149.400 437.700 157.200 439.050 ;
        RECT 149.400 432.600 151.200 437.700 ;
        RECT 155.400 432.600 157.200 437.700 ;
        RECT 158.400 438.600 159.600 440.700 ;
        RECT 179.700 438.600 180.600 445.950 ;
        RECT 158.400 432.600 160.200 438.600 ;
        RECT 175.500 437.400 180.600 438.600 ;
        RECT 175.500 432.600 177.300 437.400 ;
        RECT 197.400 435.600 198.600 445.950 ;
        RECT 203.550 445.050 204.450 449.550 ;
        RECT 211.950 448.950 214.050 449.550 ;
        RECT 215.700 448.050 216.600 460.200 ;
        RECT 238.800 455.400 240.600 467.400 ;
        RECT 241.800 456.300 243.600 467.400 ;
        RECT 247.800 456.300 249.600 467.400 ;
        RECT 260.400 461.400 262.200 467.400 ;
        RECT 260.700 461.100 262.200 461.400 ;
        RECT 266.400 461.400 268.200 467.400 ;
        RECT 286.800 461.400 288.600 467.400 ;
        RECT 266.400 461.100 267.300 461.400 ;
        RECT 260.700 460.200 267.300 461.100 ;
        RECT 241.800 455.400 249.600 456.300 ;
        RECT 221.100 448.050 222.900 449.850 ;
        RECT 239.400 448.050 240.300 455.400 ;
        RECT 247.950 453.450 250.050 454.050 ;
        RECT 256.950 453.450 259.050 454.050 ;
        RECT 247.950 452.550 259.050 453.450 ;
        RECT 247.950 451.950 250.050 452.550 ;
        RECT 256.950 451.950 259.050 452.550 ;
        RECT 245.100 448.050 246.900 449.850 ;
        RECT 260.100 448.050 261.900 449.850 ;
        RECT 266.400 448.050 267.300 460.200 ;
        RECT 271.950 450.450 274.050 450.900 ;
        RECT 277.950 450.450 280.050 451.050 ;
        RECT 271.950 449.550 280.050 450.450 ;
        RECT 271.950 448.800 274.050 449.550 ;
        RECT 277.950 448.950 280.050 449.550 ;
        RECT 281.100 448.050 282.900 449.850 ;
        RECT 286.950 448.050 288.150 461.400 ;
        RECT 310.500 456.600 312.300 467.400 ;
        RECT 313.950 465.450 316.050 466.050 ;
        RECT 322.950 465.450 325.050 466.050 ;
        RECT 313.950 464.550 325.050 465.450 ;
        RECT 313.950 463.950 316.050 464.550 ;
        RECT 322.950 463.950 325.050 464.550 ;
        RECT 331.800 461.400 333.600 467.400 ;
        RECT 308.700 455.400 312.300 456.600 ;
        RECT 289.950 453.450 292.050 453.900 ;
        RECT 304.950 453.450 307.050 454.050 ;
        RECT 289.950 452.550 307.050 453.450 ;
        RECT 289.950 451.800 292.050 452.550 ;
        RECT 304.950 451.950 307.050 452.550 ;
        RECT 292.950 450.450 297.000 451.050 ;
        RECT 292.950 448.950 297.450 450.450 ;
        RECT 214.950 445.950 217.050 448.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 220.950 445.950 223.050 448.050 ;
        RECT 223.950 445.950 226.050 448.050 ;
        RECT 238.950 445.950 241.050 448.050 ;
        RECT 241.950 445.950 244.050 448.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 280.950 445.950 283.050 448.050 ;
        RECT 283.950 445.950 286.050 448.050 ;
        RECT 286.950 445.950 289.050 448.050 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 199.950 443.550 204.450 445.050 ;
        RECT 199.950 442.950 204.000 443.550 ;
        RECT 215.700 442.200 216.600 445.950 ;
        RECT 218.100 444.150 219.900 445.950 ;
        RECT 224.100 444.150 225.900 445.950 ;
        RECT 215.700 441.000 219.000 442.200 ;
        RECT 197.400 432.600 199.200 435.600 ;
        RECT 217.200 432.600 219.000 441.000 ;
        RECT 239.400 438.600 240.300 445.950 ;
        RECT 242.100 444.150 243.900 445.950 ;
        RECT 248.100 444.150 249.900 445.950 ;
        RECT 257.100 444.150 258.900 445.950 ;
        RECT 263.100 444.150 264.900 445.950 ;
        RECT 266.400 442.200 267.300 445.950 ;
        RECT 284.100 444.150 285.900 445.950 ;
        RECT 264.000 441.000 267.300 442.200 ;
        RECT 287.850 441.750 289.050 445.950 ;
        RECT 290.100 444.150 291.900 445.950 ;
        RECT 296.550 442.050 297.450 448.950 ;
        RECT 305.100 448.050 306.900 449.850 ;
        RECT 308.700 448.050 309.600 455.400 ;
        RECT 324.000 450.450 328.050 451.050 ;
        RECT 311.100 448.050 312.900 449.850 ;
        RECT 323.550 448.950 328.050 450.450 ;
        RECT 304.950 445.950 307.050 448.050 ;
        RECT 307.950 445.950 310.050 448.050 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 239.400 437.400 244.500 438.600 ;
        RECT 242.700 432.600 244.500 437.400 ;
        RECT 264.000 432.600 265.800 441.000 ;
        RECT 287.850 440.700 291.600 441.750 ;
        RECT 281.400 437.700 289.200 439.050 ;
        RECT 281.400 432.600 283.200 437.700 ;
        RECT 287.400 432.600 289.200 437.700 ;
        RECT 290.400 438.600 291.600 440.700 ;
        RECT 295.950 439.950 298.050 442.050 ;
        RECT 290.400 432.600 292.200 438.600 ;
        RECT 308.700 435.600 309.600 445.950 ;
        RECT 323.550 445.050 324.450 448.950 ;
        RECT 332.400 448.050 333.600 461.400 ;
        RECT 344.400 456.300 346.200 467.400 ;
        RECT 350.400 456.300 352.200 467.400 ;
        RECT 344.400 455.400 352.200 456.300 ;
        RECT 353.400 455.400 355.200 467.400 ;
        RECT 370.800 455.400 372.600 467.400 ;
        RECT 376.800 461.400 378.600 467.400 ;
        RECT 347.100 448.050 348.900 449.850 ;
        RECT 353.700 448.050 354.600 455.400 ;
        RECT 370.800 448.050 372.000 455.400 ;
        RECT 377.400 454.500 378.600 461.400 ;
        RECT 389.400 456.300 391.200 467.400 ;
        RECT 395.400 456.300 397.200 467.400 ;
        RECT 389.400 455.400 397.200 456.300 ;
        RECT 398.400 455.400 400.200 467.400 ;
        RECT 418.800 461.400 420.600 467.400 ;
        RECT 372.900 453.600 378.600 454.500 ;
        RECT 372.900 452.700 374.850 453.600 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 331.950 445.950 334.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 343.950 445.950 346.050 448.050 ;
        RECT 346.950 445.950 349.050 448.050 ;
        RECT 349.950 445.950 352.050 448.050 ;
        RECT 352.950 445.950 355.050 448.050 ;
        RECT 370.800 445.950 373.050 448.050 ;
        RECT 323.550 443.550 328.050 445.050 ;
        RECT 329.100 444.150 330.900 445.950 ;
        RECT 324.000 442.950 328.050 443.550 ;
        RECT 332.400 440.700 333.600 445.950 ;
        RECT 335.100 444.150 336.900 445.950 ;
        RECT 344.100 444.150 345.900 445.950 ;
        RECT 350.100 444.150 351.900 445.950 ;
        RECT 329.400 439.800 333.600 440.700 ;
        RECT 334.950 441.450 337.050 442.050 ;
        RECT 349.950 441.450 352.050 442.050 ;
        RECT 334.950 440.550 352.050 441.450 ;
        RECT 334.950 439.950 337.050 440.550 ;
        RECT 349.950 439.950 352.050 440.550 ;
        RECT 308.400 432.600 310.200 435.600 ;
        RECT 329.400 432.600 331.200 439.800 ;
        RECT 353.700 438.600 354.600 445.950 ;
        RECT 349.500 437.400 354.600 438.600 ;
        RECT 370.800 438.600 372.000 445.950 ;
        RECT 373.950 441.300 374.850 452.700 ;
        RECT 384.000 450.450 388.050 451.050 ;
        RECT 377.100 448.050 378.900 449.850 ;
        RECT 383.550 448.950 388.050 450.450 ;
        RECT 376.950 445.950 379.050 448.050 ;
        RECT 372.900 440.400 374.850 441.300 ;
        RECT 383.550 441.450 384.450 448.950 ;
        RECT 392.100 448.050 393.900 449.850 ;
        RECT 398.700 448.050 399.600 455.400 ;
        RECT 406.950 453.450 409.050 454.050 ;
        RECT 412.950 453.450 415.050 454.050 ;
        RECT 406.950 452.550 415.050 453.450 ;
        RECT 406.950 451.950 409.050 452.550 ;
        RECT 412.950 451.950 415.050 452.550 ;
        RECT 413.100 448.050 414.900 449.850 ;
        RECT 418.950 448.050 420.150 461.400 ;
        RECT 434.400 456.600 436.200 467.400 ;
        RECT 440.400 466.500 448.200 467.400 ;
        RECT 440.400 456.600 442.200 466.500 ;
        RECT 434.400 455.700 442.200 456.600 ;
        RECT 443.400 454.500 445.200 465.600 ;
        RECT 446.400 455.400 448.200 466.500 ;
        RECT 461.700 456.600 463.500 467.400 ;
        RECT 482.400 461.400 484.200 467.400 ;
        RECT 482.700 461.100 484.200 461.400 ;
        RECT 488.400 461.400 490.200 467.400 ;
        RECT 488.400 461.100 489.300 461.400 ;
        RECT 482.700 460.200 489.300 461.100 ;
        RECT 461.700 455.400 465.300 456.600 ;
        RECT 421.950 453.450 424.050 454.200 ;
        RECT 433.950 453.450 436.050 453.900 ;
        RECT 421.950 452.550 436.050 453.450 ;
        RECT 421.950 452.100 424.050 452.550 ;
        RECT 433.950 451.800 436.050 452.550 ;
        RECT 440.100 453.600 445.200 454.500 ;
        RECT 437.100 448.050 438.900 449.850 ;
        RECT 440.100 448.050 441.000 453.600 ;
        RECT 456.000 450.450 460.050 451.050 ;
        RECT 443.100 448.050 444.900 449.850 ;
        RECT 455.550 448.950 460.050 450.450 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 433.950 445.950 436.050 448.050 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 389.100 444.150 390.900 445.950 ;
        RECT 395.100 444.150 396.900 445.950 ;
        RECT 388.950 441.450 391.050 442.050 ;
        RECT 383.550 440.550 391.050 441.450 ;
        RECT 372.900 439.500 378.600 440.400 ;
        RECT 388.950 439.950 391.050 440.550 ;
        RECT 349.500 432.600 351.300 437.400 ;
        RECT 370.800 432.600 372.600 438.600 ;
        RECT 377.400 435.600 378.600 439.500 ;
        RECT 398.700 438.600 399.600 445.950 ;
        RECT 416.100 444.150 417.900 445.950 ;
        RECT 419.850 441.750 421.050 445.950 ;
        RECT 422.100 444.150 423.900 445.950 ;
        RECT 434.100 444.150 435.900 445.950 ;
        RECT 419.850 440.700 423.600 441.750 ;
        RECT 376.800 432.600 378.600 435.600 ;
        RECT 394.500 437.400 399.600 438.600 ;
        RECT 413.400 437.700 421.200 439.050 ;
        RECT 394.500 432.600 396.300 437.400 ;
        RECT 413.400 432.600 415.200 437.700 ;
        RECT 419.400 432.600 421.200 437.700 ;
        RECT 422.400 438.600 423.600 440.700 ;
        RECT 439.950 438.600 441.000 445.950 ;
        RECT 446.100 444.150 447.900 445.950 ;
        RECT 455.550 441.900 456.450 448.950 ;
        RECT 461.100 448.050 462.900 449.850 ;
        RECT 464.400 448.050 465.300 455.400 ;
        RECT 474.000 450.450 478.050 451.050 ;
        RECT 467.100 448.050 468.900 449.850 ;
        RECT 473.550 448.950 478.050 450.450 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 463.950 445.950 466.050 448.050 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 454.950 439.800 457.050 441.900 ;
        RECT 422.400 432.600 424.200 438.600 ;
        RECT 439.200 432.600 441.000 438.600 ;
        RECT 464.400 435.600 465.300 445.950 ;
        RECT 473.550 445.050 474.450 448.950 ;
        RECT 482.100 448.050 483.900 449.850 ;
        RECT 488.400 448.050 489.300 460.200 ;
        RECT 508.500 456.600 510.300 467.400 ;
        RECT 527.400 461.400 529.200 467.400 ;
        RECT 527.700 461.100 529.200 461.400 ;
        RECT 533.400 461.400 535.200 467.400 ;
        RECT 550.800 461.400 552.600 467.400 ;
        RECT 533.400 461.100 534.300 461.400 ;
        RECT 527.700 460.200 534.300 461.100 ;
        RECT 506.700 455.400 510.300 456.600 ;
        RECT 490.950 450.450 495.000 451.050 ;
        RECT 490.950 448.950 495.450 450.450 ;
        RECT 478.950 445.950 481.050 448.050 ;
        RECT 481.950 445.950 484.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 473.550 443.550 478.050 445.050 ;
        RECT 479.100 444.150 480.900 445.950 ;
        RECT 485.100 444.150 486.900 445.950 ;
        RECT 474.000 442.950 478.050 443.550 ;
        RECT 488.400 442.200 489.300 445.950 ;
        RECT 494.550 445.050 495.450 448.950 ;
        RECT 503.100 448.050 504.900 449.850 ;
        RECT 506.700 448.050 507.600 455.400 ;
        RECT 509.100 448.050 510.900 449.850 ;
        RECT 527.100 448.050 528.900 449.850 ;
        RECT 533.400 448.050 534.300 460.200 ;
        RECT 545.100 448.050 546.900 449.850 ;
        RECT 550.950 448.050 552.150 461.400 ;
        RECT 560.550 455.400 562.350 467.400 ;
        RECT 568.050 461.400 569.850 467.400 ;
        RECT 565.950 459.300 569.850 461.400 ;
        RECT 575.850 460.500 577.650 467.400 ;
        RECT 583.650 461.400 585.450 467.400 ;
        RECT 584.250 460.500 585.450 461.400 ;
        RECT 574.950 459.450 581.550 460.500 ;
        RECT 574.950 458.700 576.750 459.450 ;
        RECT 579.750 458.700 581.550 459.450 ;
        RECT 584.250 458.400 589.050 460.500 ;
        RECT 567.150 456.600 569.850 458.400 ;
        RECT 570.750 457.800 572.550 458.400 ;
        RECT 570.750 456.900 577.050 457.800 ;
        RECT 584.250 457.500 585.450 458.400 ;
        RECT 570.750 456.600 572.550 456.900 ;
        RECT 568.950 455.700 569.850 456.600 ;
        RECT 560.550 448.050 561.750 455.400 ;
        RECT 565.950 454.800 568.050 455.700 ;
        RECT 568.950 454.800 574.050 455.700 ;
        RECT 563.850 453.600 568.050 454.800 ;
        RECT 562.950 451.800 564.750 453.600 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 529.950 445.950 532.050 448.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 553.950 445.950 556.050 448.050 ;
        RECT 560.550 447.750 565.050 448.050 ;
        RECT 560.550 445.950 566.850 447.750 ;
        RECT 490.950 443.550 495.450 445.050 ;
        RECT 490.950 442.950 495.000 443.550 ;
        RECT 486.000 441.000 489.300 442.200 ;
        RECT 463.800 432.600 465.600 435.600 ;
        RECT 486.000 432.600 487.800 441.000 ;
        RECT 506.700 435.600 507.600 445.950 ;
        RECT 524.100 444.150 525.900 445.950 ;
        RECT 530.100 444.150 531.900 445.950 ;
        RECT 533.400 442.200 534.300 445.950 ;
        RECT 548.100 444.150 549.900 445.950 ;
        RECT 531.000 441.000 534.300 442.200 ;
        RECT 551.850 441.750 553.050 445.950 ;
        RECT 554.100 444.150 555.900 445.950 ;
        RECT 506.400 432.600 508.200 435.600 ;
        RECT 531.000 432.600 532.800 441.000 ;
        RECT 551.850 440.700 555.600 441.750 ;
        RECT 545.400 437.700 553.200 439.050 ;
        RECT 545.400 432.600 547.200 437.700 ;
        RECT 551.400 432.600 553.200 437.700 ;
        RECT 554.400 438.600 555.600 440.700 ;
        RECT 560.550 438.600 561.750 445.950 ;
        RECT 573.150 442.200 574.050 454.800 ;
        RECT 576.150 454.800 577.050 456.900 ;
        RECT 577.950 456.300 585.450 457.500 ;
        RECT 577.950 455.700 579.750 456.300 ;
        RECT 592.050 455.400 593.850 467.400 ;
        RECT 576.150 454.500 584.550 454.800 ;
        RECT 592.950 454.500 593.850 455.400 ;
        RECT 576.150 453.900 593.850 454.500 ;
        RECT 582.750 453.300 593.850 453.900 ;
        RECT 582.750 453.000 584.550 453.300 ;
        RECT 580.950 446.400 583.050 448.050 ;
        RECT 580.950 445.200 588.900 446.400 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 587.100 444.600 588.900 445.200 ;
        RECT 590.100 444.150 591.900 445.950 ;
        RECT 584.100 443.400 585.900 444.000 ;
        RECT 590.100 443.400 591.000 444.150 ;
        RECT 584.100 442.200 591.000 443.400 ;
        RECT 573.150 441.000 585.150 442.200 ;
        RECT 573.150 440.400 574.950 441.000 ;
        RECT 584.100 439.200 585.150 441.000 ;
        RECT 554.400 432.600 556.200 438.600 ;
        RECT 560.550 432.600 562.350 438.600 ;
        RECT 565.950 437.700 568.050 438.600 ;
        RECT 565.950 436.500 569.700 437.700 ;
        RECT 580.350 437.550 582.150 438.300 ;
        RECT 568.650 435.600 569.700 436.500 ;
        RECT 577.200 436.500 582.150 437.550 ;
        RECT 583.650 437.400 585.450 439.200 ;
        RECT 592.950 438.600 593.850 453.300 ;
        RECT 608.400 461.400 610.200 467.400 ;
        RECT 632.400 461.400 634.200 467.400 ;
        RECT 655.800 461.400 657.600 467.400 ;
        RECT 600.000 450.450 604.050 451.050 ;
        RECT 599.550 448.950 604.050 450.450 ;
        RECT 599.550 445.050 600.450 448.950 ;
        RECT 608.400 448.050 609.600 461.400 ;
        RECT 613.950 450.450 616.050 451.050 ;
        RECT 613.950 449.550 624.450 450.450 ;
        RECT 613.950 448.950 616.050 449.550 ;
        RECT 604.950 445.950 607.050 448.050 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 599.550 443.550 604.050 445.050 ;
        RECT 605.100 444.150 606.900 445.950 ;
        RECT 600.000 442.950 604.050 443.550 ;
        RECT 608.400 440.700 609.600 445.950 ;
        RECT 611.100 444.150 612.900 445.950 ;
        RECT 623.550 445.050 624.450 449.550 ;
        RECT 632.850 448.050 634.050 461.400 ;
        RECT 640.950 450.450 645.000 451.050 ;
        RECT 638.100 448.050 639.900 449.850 ;
        RECT 640.950 448.950 645.450 450.450 ;
        RECT 628.950 445.950 631.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 634.950 445.950 637.050 448.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 623.550 443.550 628.050 445.050 ;
        RECT 629.100 444.150 630.900 445.950 ;
        RECT 624.000 442.950 628.050 443.550 ;
        RECT 631.950 441.750 633.150 445.950 ;
        RECT 635.100 444.150 636.900 445.950 ;
        RECT 644.550 445.050 645.450 448.950 ;
        RECT 650.100 448.050 651.900 449.850 ;
        RECT 655.950 448.050 657.150 461.400 ;
        RECT 665.550 455.400 667.350 467.400 ;
        RECT 673.050 461.400 674.850 467.400 ;
        RECT 670.950 459.300 674.850 461.400 ;
        RECT 680.850 460.500 682.650 467.400 ;
        RECT 688.650 461.400 690.450 467.400 ;
        RECT 689.250 460.500 690.450 461.400 ;
        RECT 679.950 459.450 686.550 460.500 ;
        RECT 679.950 458.700 681.750 459.450 ;
        RECT 684.750 458.700 686.550 459.450 ;
        RECT 689.250 458.400 694.050 460.500 ;
        RECT 672.150 456.600 674.850 458.400 ;
        RECT 675.750 457.800 677.550 458.400 ;
        RECT 675.750 456.900 682.050 457.800 ;
        RECT 689.250 457.500 690.450 458.400 ;
        RECT 675.750 456.600 677.550 456.900 ;
        RECT 673.950 455.700 674.850 456.600 ;
        RECT 665.550 448.050 666.750 455.400 ;
        RECT 670.950 454.800 673.050 455.700 ;
        RECT 673.950 454.800 679.050 455.700 ;
        RECT 668.850 453.600 673.050 454.800 ;
        RECT 667.950 451.800 669.750 453.600 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 652.950 445.950 655.050 448.050 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 665.550 447.750 670.050 448.050 ;
        RECT 665.550 445.950 671.850 447.750 ;
        RECT 644.550 443.550 649.050 445.050 ;
        RECT 653.100 444.150 654.900 445.950 ;
        RECT 645.000 442.950 649.050 443.550 ;
        RECT 629.400 440.700 633.150 441.750 ;
        RECT 656.850 441.750 658.050 445.950 ;
        RECT 659.100 444.150 660.900 445.950 ;
        RECT 656.850 440.700 660.600 441.750 ;
        RECT 608.400 439.800 612.600 440.700 ;
        RECT 586.950 436.500 589.050 438.600 ;
        RECT 577.200 435.600 578.250 436.500 ;
        RECT 586.950 435.600 588.000 436.500 ;
        RECT 568.650 432.600 570.450 435.600 ;
        RECT 576.450 432.600 578.250 435.600 ;
        RECT 584.250 434.700 588.000 435.600 ;
        RECT 584.250 432.600 586.050 434.700 ;
        RECT 592.050 432.600 593.850 438.600 ;
        RECT 610.800 432.600 612.600 439.800 ;
        RECT 629.400 438.600 630.600 440.700 ;
        RECT 628.800 432.600 630.600 438.600 ;
        RECT 631.800 437.700 639.600 439.050 ;
        RECT 631.800 432.600 633.600 437.700 ;
        RECT 637.800 432.600 639.600 437.700 ;
        RECT 650.400 437.700 658.200 439.050 ;
        RECT 650.400 432.600 652.200 437.700 ;
        RECT 656.400 432.600 658.200 437.700 ;
        RECT 659.400 438.600 660.600 440.700 ;
        RECT 665.550 438.600 666.750 445.950 ;
        RECT 678.150 442.200 679.050 454.800 ;
        RECT 681.150 454.800 682.050 456.900 ;
        RECT 682.950 456.300 690.450 457.500 ;
        RECT 682.950 455.700 684.750 456.300 ;
        RECT 697.050 455.400 698.850 467.400 ;
        RECT 681.150 454.500 689.550 454.800 ;
        RECT 697.950 454.500 698.850 455.400 ;
        RECT 681.150 453.900 698.850 454.500 ;
        RECT 687.750 453.300 698.850 453.900 ;
        RECT 687.750 453.000 689.550 453.300 ;
        RECT 685.950 446.400 688.050 448.050 ;
        RECT 685.950 445.200 693.900 446.400 ;
        RECT 694.950 445.950 697.050 448.050 ;
        RECT 692.100 444.600 693.900 445.200 ;
        RECT 695.100 444.150 696.900 445.950 ;
        RECT 689.100 443.400 690.900 444.000 ;
        RECT 695.100 443.400 696.000 444.150 ;
        RECT 689.100 442.200 696.000 443.400 ;
        RECT 678.150 441.000 690.150 442.200 ;
        RECT 678.150 440.400 679.950 441.000 ;
        RECT 689.100 439.200 690.150 441.000 ;
        RECT 659.400 432.600 661.200 438.600 ;
        RECT 665.550 432.600 667.350 438.600 ;
        RECT 670.950 437.700 673.050 438.600 ;
        RECT 670.950 436.500 674.700 437.700 ;
        RECT 685.350 437.550 687.150 438.300 ;
        RECT 673.650 435.600 674.700 436.500 ;
        RECT 682.200 436.500 687.150 437.550 ;
        RECT 688.650 437.400 690.450 439.200 ;
        RECT 697.950 438.600 698.850 453.300 ;
        RECT 691.950 436.500 694.050 438.600 ;
        RECT 682.200 435.600 683.250 436.500 ;
        RECT 691.950 435.600 693.000 436.500 ;
        RECT 673.650 432.600 675.450 435.600 ;
        RECT 681.450 432.600 683.250 435.600 ;
        RECT 689.250 434.700 693.000 435.600 ;
        RECT 689.250 432.600 691.050 434.700 ;
        RECT 697.050 432.600 698.850 438.600 ;
        RECT 701.550 455.400 703.350 467.400 ;
        RECT 709.050 461.400 710.850 467.400 ;
        RECT 706.950 459.300 710.850 461.400 ;
        RECT 716.850 460.500 718.650 467.400 ;
        RECT 724.650 461.400 726.450 467.400 ;
        RECT 725.250 460.500 726.450 461.400 ;
        RECT 715.950 459.450 722.550 460.500 ;
        RECT 715.950 458.700 717.750 459.450 ;
        RECT 720.750 458.700 722.550 459.450 ;
        RECT 725.250 458.400 730.050 460.500 ;
        RECT 708.150 456.600 710.850 458.400 ;
        RECT 711.750 457.800 713.550 458.400 ;
        RECT 711.750 456.900 718.050 457.800 ;
        RECT 725.250 457.500 726.450 458.400 ;
        RECT 711.750 456.600 713.550 456.900 ;
        RECT 709.950 455.700 710.850 456.600 ;
        RECT 701.550 448.050 702.750 455.400 ;
        RECT 706.950 454.800 709.050 455.700 ;
        RECT 709.950 454.800 715.050 455.700 ;
        RECT 704.850 453.600 709.050 454.800 ;
        RECT 703.950 451.800 705.750 453.600 ;
        RECT 701.550 447.750 706.050 448.050 ;
        RECT 701.550 445.950 707.850 447.750 ;
        RECT 701.550 438.600 702.750 445.950 ;
        RECT 714.150 442.200 715.050 454.800 ;
        RECT 717.150 454.800 718.050 456.900 ;
        RECT 718.950 456.300 726.450 457.500 ;
        RECT 718.950 455.700 720.750 456.300 ;
        RECT 733.050 455.400 734.850 467.400 ;
        RECT 717.150 454.500 725.550 454.800 ;
        RECT 733.950 454.500 734.850 455.400 ;
        RECT 751.800 454.500 753.600 467.400 ;
        RECT 757.800 454.500 759.600 467.400 ;
        RECT 763.800 454.500 765.600 467.400 ;
        RECT 769.800 454.500 771.600 467.400 ;
        RECT 717.150 453.900 734.850 454.500 ;
        RECT 723.750 453.300 734.850 453.900 ;
        RECT 723.750 453.000 725.550 453.300 ;
        RECT 721.950 446.400 724.050 448.050 ;
        RECT 721.950 445.200 729.900 446.400 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 728.100 444.600 729.900 445.200 ;
        RECT 731.100 444.150 732.900 445.950 ;
        RECT 725.100 443.400 726.900 444.000 ;
        RECT 731.100 443.400 732.000 444.150 ;
        RECT 725.100 442.200 732.000 443.400 ;
        RECT 714.150 441.000 726.150 442.200 ;
        RECT 714.150 440.400 715.950 441.000 ;
        RECT 725.100 439.200 726.150 441.000 ;
        RECT 701.550 432.600 703.350 438.600 ;
        RECT 706.950 437.700 709.050 438.600 ;
        RECT 706.950 436.500 710.700 437.700 ;
        RECT 721.350 437.550 723.150 438.300 ;
        RECT 709.650 435.600 710.700 436.500 ;
        RECT 718.200 436.500 723.150 437.550 ;
        RECT 724.650 437.400 726.450 439.200 ;
        RECT 733.950 438.600 734.850 453.300 ;
        RECT 750.900 453.300 753.600 454.500 ;
        RECT 755.700 453.300 759.600 454.500 ;
        RECT 761.700 453.300 765.600 454.500 ;
        RECT 767.700 453.300 771.600 454.500 ;
        RECT 785.400 461.400 787.200 467.400 ;
        RECT 785.400 454.500 786.600 461.400 ;
        RECT 791.400 455.400 793.200 467.400 ;
        RECT 785.400 453.600 791.100 454.500 ;
        RECT 750.900 448.050 751.800 453.300 ;
        RECT 748.950 445.950 751.800 448.050 ;
        RECT 739.950 444.450 742.050 445.050 ;
        RECT 745.950 444.450 748.050 445.050 ;
        RECT 739.950 443.550 748.050 444.450 ;
        RECT 739.950 442.950 742.050 443.550 ;
        RECT 745.950 442.950 748.050 443.550 ;
        RECT 750.900 440.700 751.800 445.950 ;
        RECT 752.700 442.800 754.500 443.400 ;
        RECT 755.700 442.800 756.900 453.300 ;
        RECT 752.700 441.600 756.900 442.800 ;
        RECT 758.700 442.800 760.500 443.400 ;
        RECT 761.700 442.800 762.900 453.300 ;
        RECT 758.700 441.600 762.900 442.800 ;
        RECT 764.700 442.800 766.500 443.400 ;
        RECT 767.700 442.800 768.900 453.300 ;
        RECT 789.150 452.700 791.100 453.600 ;
        RECT 785.100 448.050 786.900 449.850 ;
        RECT 769.950 445.950 772.050 448.050 ;
        RECT 784.950 445.950 787.050 448.050 ;
        RECT 770.100 444.150 771.900 445.950 ;
        RECT 764.700 441.600 768.900 442.800 ;
        RECT 755.700 440.700 756.900 441.600 ;
        RECT 761.700 440.700 762.900 441.600 ;
        RECT 767.700 440.700 768.900 441.600 ;
        RECT 772.950 441.450 775.050 442.050 ;
        RECT 781.950 441.450 784.050 442.050 ;
        RECT 750.900 439.500 753.600 440.700 ;
        RECT 755.700 439.500 759.600 440.700 ;
        RECT 761.700 439.500 765.600 440.700 ;
        RECT 767.700 439.500 771.600 440.700 ;
        RECT 772.950 440.550 784.050 441.450 ;
        RECT 772.950 439.950 775.050 440.550 ;
        RECT 781.950 439.950 784.050 440.550 ;
        RECT 789.150 441.300 790.050 452.700 ;
        RECT 792.000 448.050 793.200 455.400 ;
        RECT 803.400 461.400 805.200 467.400 ;
        RECT 803.400 454.500 804.600 461.400 ;
        RECT 809.400 455.400 811.200 467.400 ;
        RECT 828.300 456.900 830.100 467.400 ;
        RECT 803.400 453.600 809.100 454.500 ;
        RECT 807.150 452.700 809.100 453.600 ;
        RECT 798.000 450.450 802.050 451.050 ;
        RECT 790.950 445.950 793.200 448.050 ;
        RECT 789.150 440.400 791.100 441.300 ;
        RECT 727.950 436.500 730.050 438.600 ;
        RECT 718.200 435.600 719.250 436.500 ;
        RECT 727.950 435.600 729.000 436.500 ;
        RECT 709.650 432.600 711.450 435.600 ;
        RECT 717.450 432.600 719.250 435.600 ;
        RECT 725.250 434.700 729.000 435.600 ;
        RECT 725.250 432.600 727.050 434.700 ;
        RECT 733.050 432.600 734.850 438.600 ;
        RECT 751.800 432.600 753.600 439.500 ;
        RECT 757.800 432.600 759.600 439.500 ;
        RECT 763.800 432.600 765.600 439.500 ;
        RECT 769.800 432.600 771.600 439.500 ;
        RECT 785.400 439.500 791.100 440.400 ;
        RECT 785.400 435.600 786.600 439.500 ;
        RECT 792.000 438.600 793.200 445.950 ;
        RECT 797.550 448.950 802.050 450.450 ;
        RECT 797.550 445.050 798.450 448.950 ;
        RECT 803.100 448.050 804.900 449.850 ;
        RECT 802.950 445.950 805.050 448.050 ;
        RECT 797.550 443.550 802.050 445.050 ;
        RECT 798.000 442.950 802.050 443.550 ;
        RECT 807.150 441.300 808.050 452.700 ;
        RECT 810.000 448.050 811.200 455.400 ;
        RECT 827.700 455.400 830.100 456.900 ;
        RECT 835.800 455.400 837.600 467.400 ;
        RECT 851.700 456.600 853.500 467.400 ;
        RECT 868.800 461.400 870.600 467.400 ;
        RECT 886.800 461.400 888.600 467.400 ;
        RECT 904.800 461.400 906.600 467.400 ;
        RECT 851.700 455.400 855.300 456.600 ;
        RECT 827.700 448.050 829.050 455.400 ;
        RECT 836.400 453.900 837.600 455.400 ;
        RECT 808.950 445.950 811.200 448.050 ;
        RECT 807.150 440.400 809.100 441.300 ;
        RECT 785.400 432.600 787.200 435.600 ;
        RECT 791.400 432.600 793.200 438.600 ;
        RECT 803.400 439.500 809.100 440.400 ;
        RECT 803.400 435.600 804.600 439.500 ;
        RECT 810.000 438.600 811.200 445.950 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 830.400 452.700 837.600 453.900 ;
        RECT 830.400 452.100 832.200 452.700 ;
        RECT 826.950 438.600 828.000 445.950 ;
        RECT 830.400 441.600 831.300 452.100 ;
        RECT 846.000 450.450 850.050 451.050 ;
        RECT 833.100 448.050 834.900 449.850 ;
        RECT 845.550 448.950 850.050 450.450 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 835.950 445.950 838.050 448.050 ;
        RECT 836.100 444.150 837.900 445.950 ;
        RECT 838.950 444.450 841.050 445.050 ;
        RECT 845.550 444.450 846.450 448.950 ;
        RECT 851.100 448.050 852.900 449.850 ;
        RECT 854.400 448.050 855.300 455.400 ;
        RECT 857.100 448.050 858.900 449.850 ;
        RECT 869.400 448.050 870.600 461.400 ;
        RECT 872.100 448.050 873.900 449.850 ;
        RECT 887.400 448.050 888.600 461.400 ;
        RECT 905.700 461.100 906.600 461.400 ;
        RECT 910.800 461.400 912.600 467.400 ;
        RECT 910.800 461.100 912.300 461.400 ;
        RECT 905.700 460.200 912.300 461.100 ;
        RECT 905.700 448.050 906.600 460.200 ;
        RECT 911.100 448.050 912.900 449.850 ;
        RECT 850.950 445.950 853.050 448.050 ;
        RECT 853.950 445.950 856.050 448.050 ;
        RECT 856.950 445.950 859.050 448.050 ;
        RECT 868.950 445.950 871.050 448.050 ;
        RECT 871.950 445.950 874.050 448.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 904.950 445.950 907.050 448.050 ;
        RECT 907.950 445.950 910.050 448.050 ;
        RECT 910.950 445.950 913.050 448.050 ;
        RECT 913.950 445.950 916.050 448.050 ;
        RECT 838.950 443.550 846.450 444.450 ;
        RECT 838.950 442.950 841.050 443.550 ;
        RECT 830.400 440.700 832.200 441.600 ;
        RECT 830.400 439.800 833.700 440.700 ;
        RECT 803.400 432.600 805.200 435.600 ;
        RECT 809.400 432.600 811.200 438.600 ;
        RECT 826.800 432.600 828.600 438.600 ;
        RECT 832.800 435.600 833.700 439.800 ;
        RECT 854.400 435.600 855.300 445.950 ;
        RECT 869.400 435.600 870.600 445.950 ;
        RECT 884.100 444.150 885.900 445.950 ;
        RECT 887.400 440.700 888.600 445.950 ;
        RECT 890.100 444.150 891.900 445.950 ;
        RECT 905.700 442.200 906.600 445.950 ;
        RECT 908.100 444.150 909.900 445.950 ;
        RECT 914.100 444.150 915.900 445.950 ;
        RECT 905.700 441.000 909.000 442.200 ;
        RECT 884.400 439.800 888.600 440.700 ;
        RECT 871.950 438.450 874.050 439.050 ;
        RECT 880.950 438.450 883.050 439.050 ;
        RECT 871.950 437.550 883.050 438.450 ;
        RECT 871.950 436.950 874.050 437.550 ;
        RECT 880.950 436.950 883.050 437.550 ;
        RECT 832.800 432.600 834.600 435.600 ;
        RECT 853.800 432.600 855.600 435.600 ;
        RECT 868.800 432.600 870.600 435.600 ;
        RECT 884.400 432.600 886.200 439.800 ;
        RECT 907.200 432.600 909.000 441.000 ;
        RECT 16.200 420.000 18.000 428.400 ;
        RECT 14.700 418.800 18.000 420.000 ;
        RECT 42.000 420.000 43.800 428.400 ;
        RECT 61.200 420.000 63.000 428.400 ;
        RECT 85.500 423.600 87.300 428.400 ;
        RECT 85.500 422.400 90.600 423.600 ;
        RECT 106.800 422.400 108.600 428.400 ;
        RECT 42.000 418.800 45.300 420.000 ;
        RECT 14.700 415.050 15.600 418.800 ;
        RECT 17.100 415.050 18.900 416.850 ;
        RECT 23.100 415.050 24.900 416.850 ;
        RECT 35.100 415.050 36.900 416.850 ;
        RECT 41.100 415.050 42.900 416.850 ;
        RECT 44.400 415.050 45.300 418.800 ;
        RECT 59.700 418.800 63.000 420.000 ;
        RECT 59.700 415.050 60.600 418.800 ;
        RECT 62.100 415.050 63.900 416.850 ;
        RECT 68.100 415.050 69.900 416.850 ;
        RECT 80.100 415.050 81.900 416.850 ;
        RECT 86.100 415.050 87.900 416.850 ;
        RECT 89.700 415.050 90.600 422.400 ;
        RECT 107.400 420.300 108.600 422.400 ;
        RECT 109.800 423.300 111.600 428.400 ;
        RECT 115.800 423.300 117.600 428.400 ;
        RECT 131.700 423.600 133.500 428.400 ;
        RECT 109.800 421.950 117.600 423.300 ;
        RECT 128.400 422.400 133.500 423.600 ;
        RECT 152.400 425.400 154.200 428.400 ;
        RECT 107.400 419.250 111.150 420.300 ;
        RECT 107.100 415.050 108.900 416.850 ;
        RECT 109.950 415.050 111.150 419.250 ;
        RECT 113.100 415.050 114.900 416.850 ;
        RECT 128.400 415.050 129.300 422.400 ;
        RECT 144.000 417.450 148.050 418.050 ;
        RECT 131.100 415.050 132.900 416.850 ;
        RECT 137.100 415.050 138.900 416.850 ;
        RECT 143.550 415.950 148.050 417.450 ;
        RECT 13.950 412.950 16.050 415.050 ;
        RECT 16.950 412.950 19.050 415.050 ;
        RECT 19.950 412.950 22.050 415.050 ;
        RECT 22.950 412.950 25.050 415.050 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 37.950 412.950 40.050 415.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 43.950 412.950 46.050 415.050 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 61.950 412.950 64.050 415.050 ;
        RECT 64.950 412.950 67.050 415.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 82.950 412.950 85.050 415.050 ;
        RECT 85.950 412.950 88.050 415.050 ;
        RECT 88.950 412.950 91.050 415.050 ;
        RECT 106.950 412.950 109.050 415.050 ;
        RECT 109.950 412.950 112.050 415.050 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 115.950 412.950 118.050 415.050 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 133.950 412.950 136.050 415.050 ;
        RECT 136.950 412.950 139.050 415.050 ;
        RECT 14.700 400.800 15.600 412.950 ;
        RECT 20.100 411.150 21.900 412.950 ;
        RECT 38.100 411.150 39.900 412.950 ;
        RECT 44.400 400.800 45.300 412.950 ;
        RECT 14.700 399.900 21.300 400.800 ;
        RECT 14.700 399.600 15.600 399.900 ;
        RECT 13.800 393.600 15.600 399.600 ;
        RECT 19.800 399.600 21.300 399.900 ;
        RECT 38.700 399.900 45.300 400.800 ;
        RECT 38.700 399.600 40.200 399.900 ;
        RECT 19.800 393.600 21.600 399.600 ;
        RECT 38.400 393.600 40.200 399.600 ;
        RECT 44.400 399.600 45.300 399.900 ;
        RECT 59.700 400.800 60.600 412.950 ;
        RECT 65.100 411.150 66.900 412.950 ;
        RECT 83.100 411.150 84.900 412.950 ;
        RECT 61.950 408.450 64.050 409.050 ;
        RECT 79.950 408.450 82.050 409.050 ;
        RECT 61.950 407.550 82.050 408.450 ;
        RECT 61.950 406.950 64.050 407.550 ;
        RECT 79.950 406.950 82.050 407.550 ;
        RECT 89.700 405.600 90.600 412.950 ;
        RECT 80.400 404.700 88.200 405.600 ;
        RECT 59.700 399.900 66.300 400.800 ;
        RECT 59.700 399.600 60.600 399.900 ;
        RECT 44.400 393.600 46.200 399.600 ;
        RECT 58.800 393.600 60.600 399.600 ;
        RECT 64.800 399.600 66.300 399.900 ;
        RECT 64.800 393.600 66.600 399.600 ;
        RECT 80.400 393.600 82.200 404.700 ;
        RECT 86.400 393.600 88.200 404.700 ;
        RECT 89.400 393.600 91.200 405.600 ;
        RECT 110.850 399.600 112.050 412.950 ;
        RECT 116.100 411.150 117.900 412.950 ;
        RECT 128.400 405.600 129.300 412.950 ;
        RECT 134.100 411.150 135.900 412.950 ;
        RECT 143.550 412.050 144.450 415.950 ;
        RECT 152.400 415.050 153.600 425.400 ;
        RECT 174.000 420.000 175.800 428.400 ;
        RECT 198.000 420.000 199.800 428.400 ;
        RECT 217.200 422.400 219.000 428.400 ;
        RECT 174.000 418.800 177.300 420.000 ;
        RECT 198.000 418.800 201.300 420.000 ;
        RECT 167.100 415.050 168.900 416.850 ;
        RECT 173.100 415.050 174.900 416.850 ;
        RECT 176.400 415.050 177.300 418.800 ;
        RECT 191.100 415.050 192.900 416.850 ;
        RECT 197.100 415.050 198.900 416.850 ;
        RECT 200.400 415.050 201.300 418.800 ;
        RECT 212.100 415.050 213.900 416.850 ;
        RECT 217.950 415.050 219.000 422.400 ;
        RECT 242.400 425.400 244.200 428.400 ;
        RECT 220.950 420.450 223.050 421.050 ;
        RECT 226.950 420.450 229.050 421.050 ;
        RECT 238.950 420.450 241.050 420.900 ;
        RECT 220.950 419.550 229.050 420.450 ;
        RECT 220.950 418.950 223.050 419.550 ;
        RECT 226.950 418.950 229.050 419.550 ;
        RECT 230.550 419.550 241.050 420.450 ;
        RECT 224.100 415.050 225.900 416.850 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 172.950 412.950 175.050 415.050 ;
        RECT 175.950 412.950 178.050 415.050 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 193.950 412.950 196.050 415.050 ;
        RECT 196.950 412.950 199.050 415.050 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 211.950 412.950 214.050 415.050 ;
        RECT 214.950 412.950 217.050 415.050 ;
        RECT 217.950 412.950 220.050 415.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 143.550 410.550 148.050 412.050 ;
        RECT 149.100 411.150 150.900 412.950 ;
        RECT 144.000 409.950 148.050 410.550 ;
        RECT 130.950 408.450 133.050 409.050 ;
        RECT 142.950 408.450 145.050 409.050 ;
        RECT 130.950 407.550 145.050 408.450 ;
        RECT 130.950 406.950 133.050 407.550 ;
        RECT 142.950 406.950 145.050 407.550 ;
        RECT 110.400 393.600 112.200 399.600 ;
        RECT 127.800 393.600 129.600 405.600 ;
        RECT 130.800 404.700 138.600 405.600 ;
        RECT 130.800 393.600 132.600 404.700 ;
        RECT 136.800 393.600 138.600 404.700 ;
        RECT 139.950 402.450 142.050 403.050 ;
        RECT 145.950 402.450 148.050 403.050 ;
        RECT 139.950 401.550 148.050 402.450 ;
        RECT 139.950 400.950 142.050 401.550 ;
        RECT 145.950 400.950 148.050 401.550 ;
        RECT 152.400 399.600 153.600 412.950 ;
        RECT 170.100 411.150 171.900 412.950 ;
        RECT 176.400 400.800 177.300 412.950 ;
        RECT 194.100 411.150 195.900 412.950 ;
        RECT 200.400 400.800 201.300 412.950 ;
        RECT 215.100 411.150 216.900 412.950 ;
        RECT 218.100 407.400 219.000 412.950 ;
        RECT 221.100 411.150 222.900 412.950 ;
        RECT 230.550 408.900 231.450 419.550 ;
        RECT 238.950 418.800 241.050 419.550 ;
        RECT 242.400 415.050 243.600 425.400 ;
        RECT 244.950 423.450 247.050 424.050 ;
        RECT 256.950 423.450 259.050 424.050 ;
        RECT 244.950 422.550 259.050 423.450 ;
        RECT 244.950 421.950 247.050 422.550 ;
        RECT 256.950 421.950 259.050 422.550 ;
        RECT 262.200 420.000 264.000 428.400 ;
        RECT 283.800 425.400 285.600 428.400 ;
        RECT 260.700 418.800 264.000 420.000 ;
        RECT 256.950 417.450 259.050 418.050 ;
        RECT 248.550 416.550 259.050 417.450 ;
        RECT 238.950 412.950 241.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 239.100 411.150 240.900 412.950 ;
        RECT 218.100 406.500 223.200 407.400 ;
        RECT 229.950 406.800 232.050 408.900 ;
        RECT 170.700 399.900 177.300 400.800 ;
        RECT 170.700 399.600 172.200 399.900 ;
        RECT 152.400 393.600 154.200 399.600 ;
        RECT 170.400 393.600 172.200 399.600 ;
        RECT 176.400 399.600 177.300 399.900 ;
        RECT 194.700 399.900 201.300 400.800 ;
        RECT 194.700 399.600 196.200 399.900 ;
        RECT 176.400 393.600 178.200 399.600 ;
        RECT 194.400 393.600 196.200 399.600 ;
        RECT 200.400 399.600 201.300 399.900 ;
        RECT 212.400 404.400 220.200 405.300 ;
        RECT 200.400 393.600 202.200 399.600 ;
        RECT 212.400 393.600 214.200 404.400 ;
        RECT 218.400 394.500 220.200 404.400 ;
        RECT 221.400 395.400 223.200 406.500 ;
        RECT 224.400 394.500 226.200 405.600 ;
        RECT 218.400 393.600 226.200 394.500 ;
        RECT 242.400 399.600 243.600 412.950 ;
        RECT 248.550 412.050 249.450 416.550 ;
        RECT 256.950 415.950 259.050 416.550 ;
        RECT 260.700 415.050 261.600 418.800 ;
        RECT 263.100 415.050 264.900 416.850 ;
        RECT 269.100 415.050 270.900 416.850 ;
        RECT 284.400 415.050 285.600 425.400 ;
        RECT 304.800 421.200 306.600 428.400 ;
        RECT 323.400 425.400 325.200 428.400 ;
        RECT 286.950 420.450 289.050 421.050 ;
        RECT 298.950 420.450 301.050 421.050 ;
        RECT 286.950 419.550 301.050 420.450 ;
        RECT 286.950 418.950 289.050 419.550 ;
        RECT 298.950 418.950 301.050 419.550 ;
        RECT 302.400 420.300 306.600 421.200 ;
        RECT 299.100 415.050 300.900 416.850 ;
        RECT 302.400 415.050 303.600 420.300 ;
        RECT 315.000 417.450 319.050 418.050 ;
        RECT 314.550 417.000 319.050 417.450 ;
        RECT 305.100 415.050 306.900 416.850 ;
        RECT 313.950 415.950 319.050 417.000 ;
        RECT 259.950 412.950 262.050 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 244.950 410.550 249.450 412.050 ;
        RECT 244.950 409.950 249.000 410.550 ;
        RECT 260.700 400.800 261.600 412.950 ;
        RECT 266.100 411.150 267.900 412.950 ;
        RECT 260.700 399.900 267.300 400.800 ;
        RECT 260.700 399.600 261.600 399.900 ;
        RECT 242.400 393.600 244.200 399.600 ;
        RECT 259.800 393.600 261.600 399.600 ;
        RECT 265.800 399.600 267.300 399.900 ;
        RECT 284.400 399.600 285.600 412.950 ;
        RECT 287.100 411.150 288.900 412.950 ;
        RECT 265.800 393.600 267.600 399.600 ;
        RECT 283.800 393.600 285.600 399.600 ;
        RECT 302.400 399.600 303.600 412.950 ;
        RECT 313.950 412.800 316.050 415.950 ;
        RECT 323.700 415.050 324.600 425.400 ;
        RECT 341.400 421.200 343.200 428.400 ;
        RECT 341.400 420.300 345.600 421.200 ;
        RECT 336.000 417.450 340.050 418.050 ;
        RECT 335.550 415.950 340.050 417.450 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 325.950 412.950 328.050 415.050 ;
        RECT 320.100 411.150 321.900 412.950 ;
        RECT 323.700 405.600 324.600 412.950 ;
        RECT 326.100 411.150 327.900 412.950 ;
        RECT 335.550 412.050 336.450 415.950 ;
        RECT 341.100 415.050 342.900 416.850 ;
        RECT 344.400 415.050 345.600 420.300 ;
        RECT 356.400 420.600 358.200 428.400 ;
        RECT 363.900 424.200 365.700 428.400 ;
        RECT 383.400 425.400 385.200 428.400 ;
        RECT 363.900 422.400 366.600 424.200 ;
        RECT 362.100 420.600 363.900 421.500 ;
        RECT 356.400 419.700 363.900 420.600 ;
        RECT 347.100 415.050 348.900 416.850 ;
        RECT 356.100 415.050 357.900 416.850 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 355.950 412.950 358.050 415.050 ;
        RECT 335.550 410.550 340.050 412.050 ;
        RECT 336.000 409.950 340.050 410.550 ;
        RECT 325.950 408.450 328.050 409.050 ;
        RECT 331.950 408.450 334.050 409.050 ;
        RECT 325.950 407.550 334.050 408.450 ;
        RECT 325.950 406.950 328.050 407.550 ;
        RECT 331.950 406.950 334.050 407.550 ;
        RECT 323.700 404.400 327.300 405.600 ;
        RECT 302.400 393.600 304.200 399.600 ;
        RECT 325.500 393.600 327.300 404.400 ;
        RECT 344.400 399.600 345.600 412.950 ;
        RECT 343.800 393.600 345.600 399.600 ;
        RECT 359.400 399.600 360.300 419.700 ;
        RECT 365.700 415.050 366.600 422.400 ;
        RECT 367.950 420.450 370.050 421.050 ;
        RECT 379.950 420.450 382.050 421.050 ;
        RECT 367.950 419.550 382.050 420.450 ;
        RECT 367.950 418.950 370.050 419.550 ;
        RECT 379.950 418.950 382.050 419.550 ;
        RECT 376.950 417.450 379.050 418.050 ;
        RECT 371.550 416.550 379.050 417.450 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 362.100 411.150 363.900 412.950 ;
        RECT 365.700 405.600 366.600 412.950 ;
        RECT 371.550 412.050 372.450 416.550 ;
        RECT 376.950 415.950 379.050 416.550 ;
        RECT 383.400 415.050 384.600 425.400 ;
        RECT 400.800 422.400 402.600 428.400 ;
        RECT 401.400 420.300 402.600 422.400 ;
        RECT 403.800 423.300 405.600 428.400 ;
        RECT 409.800 423.300 411.600 428.400 ;
        RECT 403.800 421.950 411.600 423.300 ;
        RECT 427.800 421.200 429.600 428.400 ;
        RECT 425.400 420.300 429.600 421.200 ;
        RECT 401.400 419.250 405.150 420.300 ;
        RECT 401.100 415.050 402.900 416.850 ;
        RECT 403.950 415.050 405.150 419.250 ;
        RECT 417.000 417.450 421.050 418.050 ;
        RECT 407.100 415.050 408.900 416.850 ;
        RECT 416.550 415.950 421.050 417.450 ;
        RECT 379.950 412.950 382.050 415.050 ;
        RECT 382.950 412.950 385.050 415.050 ;
        RECT 367.950 410.550 372.450 412.050 ;
        RECT 380.100 411.150 381.900 412.950 ;
        RECT 367.950 409.950 372.000 410.550 ;
        RECT 370.950 408.450 373.050 409.050 ;
        RECT 379.950 408.450 382.050 409.050 ;
        RECT 370.950 407.550 382.050 408.450 ;
        RECT 370.950 406.950 373.050 407.550 ;
        RECT 379.950 406.950 382.050 407.550 ;
        RECT 359.400 393.600 361.200 399.600 ;
        RECT 365.400 393.600 367.200 405.600 ;
        RECT 383.400 399.600 384.600 412.950 ;
        RECT 388.950 412.050 391.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 385.950 411.000 391.050 412.050 ;
        RECT 385.950 410.550 390.450 411.000 ;
        RECT 385.950 409.950 390.000 410.550 ;
        RECT 391.950 408.450 394.050 409.050 ;
        RECT 397.950 408.450 400.050 409.050 ;
        RECT 391.950 407.550 400.050 408.450 ;
        RECT 391.950 406.950 394.050 407.550 ;
        RECT 397.950 406.950 400.050 407.550 ;
        RECT 404.850 399.600 406.050 412.950 ;
        RECT 410.100 411.150 411.900 412.950 ;
        RECT 416.550 412.050 417.450 415.950 ;
        RECT 422.100 415.050 423.900 416.850 ;
        RECT 425.400 415.050 426.600 420.300 ;
        RECT 450.000 420.000 451.800 428.400 ;
        RECT 469.800 422.400 471.600 428.400 ;
        RECT 477.300 422.400 479.100 428.400 ;
        RECT 484.800 422.400 486.600 428.400 ;
        RECT 469.800 421.500 474.600 422.400 ;
        RECT 472.500 420.300 474.600 421.500 ;
        RECT 477.600 420.900 478.800 422.400 ;
        RECT 450.000 418.800 453.300 420.000 ;
        RECT 475.800 418.800 478.800 420.900 ;
        RECT 484.800 420.600 486.000 422.400 ;
        RECT 428.100 415.050 429.900 416.850 ;
        RECT 443.100 415.050 444.900 416.850 ;
        RECT 449.100 415.050 450.900 416.850 ;
        RECT 452.400 415.050 453.300 418.800 ;
        RECT 454.950 417.450 459.000 418.050 ;
        RECT 454.950 415.950 459.450 417.450 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 442.950 412.950 445.050 415.050 ;
        RECT 445.950 412.950 448.050 415.050 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 412.950 410.550 417.450 412.050 ;
        RECT 412.950 409.950 417.000 410.550 ;
        RECT 425.400 399.600 426.600 412.950 ;
        RECT 446.100 411.150 447.900 412.950 ;
        RECT 452.400 400.800 453.300 412.950 ;
        RECT 458.550 412.050 459.450 415.950 ;
        RECT 474.750 415.800 476.850 417.900 ;
        RECT 463.950 414.450 468.000 415.050 ;
        RECT 469.950 414.450 472.050 415.050 ;
        RECT 463.950 413.550 472.050 414.450 ;
        RECT 474.600 414.000 476.400 415.800 ;
        RECT 463.950 412.950 468.000 413.550 ;
        RECT 469.950 412.950 472.050 413.550 ;
        RECT 477.750 413.100 478.800 418.800 ;
        RECT 479.700 419.700 486.000 420.600 ;
        RECT 497.400 420.600 499.200 428.400 ;
        RECT 504.900 424.200 506.700 428.400 ;
        RECT 504.900 422.400 507.600 424.200 ;
        RECT 503.100 420.600 504.900 421.500 ;
        RECT 497.400 419.700 504.900 420.600 ;
        RECT 479.700 417.600 481.800 419.700 ;
        RECT 479.700 415.800 481.500 417.600 ;
        RECT 492.000 417.450 496.050 418.050 ;
        RECT 484.800 415.050 486.600 416.850 ;
        RECT 491.550 415.950 496.050 417.450 ;
        RECT 484.500 414.300 490.050 415.050 ;
        RECT 454.950 410.550 459.450 412.050 ;
        RECT 470.100 411.150 471.900 412.950 ;
        RECT 476.400 412.200 478.800 413.100 ;
        RECT 479.700 413.100 490.050 414.300 ;
        RECT 479.700 412.500 481.500 413.100 ;
        RECT 484.500 412.950 490.050 413.100 ;
        RECT 454.950 409.950 459.000 410.550 ;
        RECT 475.800 410.100 477.900 412.200 ;
        RECT 491.550 412.050 492.450 415.950 ;
        RECT 497.100 415.050 498.900 416.850 ;
        RECT 496.950 412.950 499.050 415.050 ;
        RECT 477.000 408.000 477.900 410.100 ;
        RECT 478.800 409.500 482.700 411.300 ;
        RECT 491.550 410.550 496.050 412.050 ;
        RECT 492.000 409.950 496.050 410.550 ;
        RECT 478.800 409.200 480.900 409.500 ;
        RECT 477.000 407.100 478.500 408.000 ;
        RECT 472.500 405.600 474.600 406.500 ;
        RECT 446.700 399.900 453.300 400.800 ;
        RECT 446.700 399.600 448.200 399.900 ;
        RECT 383.400 393.600 385.200 399.600 ;
        RECT 404.400 393.600 406.200 399.600 ;
        RECT 425.400 393.600 427.200 399.600 ;
        RECT 446.400 393.600 448.200 399.600 ;
        RECT 452.400 399.600 453.300 399.900 ;
        RECT 469.800 404.400 474.600 405.600 ;
        RECT 477.300 405.600 478.500 407.100 ;
        RECT 482.100 405.600 484.200 407.700 ;
        RECT 452.400 393.600 454.200 399.600 ;
        RECT 469.800 393.600 471.600 404.400 ;
        RECT 477.300 393.600 479.100 405.600 ;
        RECT 482.100 404.700 486.600 405.600 ;
        RECT 484.800 393.600 486.600 404.700 ;
        RECT 500.400 399.600 501.300 419.700 ;
        RECT 506.700 415.050 507.600 422.400 ;
        RECT 518.400 423.300 520.200 428.400 ;
        RECT 524.400 423.300 526.200 428.400 ;
        RECT 518.400 421.950 526.200 423.300 ;
        RECT 527.400 422.400 529.200 428.400 ;
        RECT 542.400 423.300 544.200 428.400 ;
        RECT 548.400 423.300 550.200 428.400 ;
        RECT 527.400 420.300 528.600 422.400 ;
        RECT 542.400 421.950 550.200 423.300 ;
        RECT 551.400 422.400 553.200 428.400 ;
        RECT 568.800 425.400 570.600 428.400 ;
        RECT 551.400 420.300 552.600 422.400 ;
        RECT 524.850 419.250 528.600 420.300 ;
        RECT 548.850 419.250 552.600 420.300 ;
        RECT 521.100 415.050 522.900 416.850 ;
        RECT 524.850 415.050 526.050 419.250 ;
        RECT 527.100 415.050 528.900 416.850 ;
        RECT 545.100 415.050 546.900 416.850 ;
        RECT 548.850 415.050 550.050 419.250 ;
        RECT 551.100 415.050 552.900 416.850 ;
        RECT 569.400 415.050 570.600 425.400 ;
        RECT 586.800 422.400 588.600 428.400 ;
        RECT 587.400 420.300 588.600 422.400 ;
        RECT 589.800 423.300 591.600 428.400 ;
        RECT 595.800 423.300 597.600 428.400 ;
        RECT 589.800 421.950 597.600 423.300 ;
        RECT 610.800 422.400 612.600 428.400 ;
        RECT 616.800 425.400 618.600 428.400 ;
        RECT 587.400 419.250 591.150 420.300 ;
        RECT 587.100 415.050 588.900 416.850 ;
        RECT 589.950 415.050 591.150 419.250 ;
        RECT 593.100 415.050 594.900 416.850 ;
        RECT 610.800 415.050 612.000 422.400 ;
        RECT 617.400 421.500 618.600 425.400 ;
        RECT 629.400 423.300 631.200 428.400 ;
        RECT 635.400 423.300 637.200 428.400 ;
        RECT 629.400 421.950 637.200 423.300 ;
        RECT 638.400 422.400 640.200 428.400 ;
        RECT 612.900 420.600 618.600 421.500 ;
        RECT 612.900 419.700 614.850 420.600 ;
        RECT 638.400 420.300 639.600 422.400 ;
        RECT 656.400 421.200 658.200 428.400 ;
        RECT 673.800 422.400 675.600 428.400 ;
        RECT 656.400 420.300 660.600 421.200 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 505.950 412.950 508.050 415.050 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 520.950 412.950 523.050 415.050 ;
        RECT 523.950 412.950 526.050 415.050 ;
        RECT 526.950 412.950 529.050 415.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 547.950 412.950 550.050 415.050 ;
        RECT 550.950 412.950 553.050 415.050 ;
        RECT 568.950 412.950 571.050 415.050 ;
        RECT 571.950 412.950 574.050 415.050 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 610.800 412.950 613.050 415.050 ;
        RECT 503.100 411.150 504.900 412.950 ;
        RECT 506.700 405.600 507.600 412.950 ;
        RECT 518.100 411.150 519.900 412.950 ;
        RECT 500.400 393.600 502.200 399.600 ;
        RECT 506.400 393.600 508.200 405.600 ;
        RECT 523.950 399.600 525.150 412.950 ;
        RECT 542.100 411.150 543.900 412.950 ;
        RECT 547.950 399.600 549.150 412.950 ;
        RECT 569.400 399.600 570.600 412.950 ;
        RECT 572.100 411.150 573.900 412.950 ;
        RECT 590.850 399.600 592.050 412.950 ;
        RECT 596.100 411.150 597.900 412.950 ;
        RECT 610.800 405.600 612.000 412.950 ;
        RECT 613.950 408.300 614.850 419.700 ;
        RECT 635.850 419.250 639.600 420.300 ;
        RECT 632.100 415.050 633.900 416.850 ;
        RECT 635.850 415.050 637.050 419.250 ;
        RECT 638.100 415.050 639.900 416.850 ;
        RECT 656.100 415.050 657.900 416.850 ;
        RECT 659.400 415.050 660.600 420.300 ;
        RECT 674.400 420.300 675.600 422.400 ;
        RECT 676.800 423.300 678.600 428.400 ;
        RECT 682.800 423.300 684.600 428.400 ;
        RECT 698.400 425.400 700.200 428.400 ;
        RECT 718.800 425.400 720.600 428.400 ;
        RECT 676.800 421.950 684.600 423.300 ;
        RECT 674.400 419.250 678.150 420.300 ;
        RECT 662.100 415.050 663.900 416.850 ;
        RECT 674.100 415.050 675.900 416.850 ;
        RECT 676.950 415.050 678.150 419.250 ;
        RECT 680.100 415.050 681.900 416.850 ;
        RECT 698.700 415.050 699.600 425.400 ;
        RECT 719.400 415.050 720.300 425.400 ;
        RECT 726.150 422.400 727.950 428.400 ;
        RECT 733.950 426.300 735.750 428.400 ;
        RECT 732.000 425.400 735.750 426.300 ;
        RECT 741.750 425.400 743.550 428.400 ;
        RECT 749.550 425.400 751.350 428.400 ;
        RECT 732.000 424.500 733.050 425.400 ;
        RECT 741.750 424.500 742.800 425.400 ;
        RECT 730.950 422.400 733.050 424.500 ;
        RECT 616.950 412.950 619.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 682.950 412.950 685.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 617.100 411.150 618.900 412.950 ;
        RECT 629.100 411.150 630.900 412.950 ;
        RECT 612.900 407.400 614.850 408.300 ;
        RECT 612.900 406.500 618.600 407.400 ;
        RECT 523.800 393.600 525.600 399.600 ;
        RECT 547.800 393.600 549.600 399.600 ;
        RECT 568.800 393.600 570.600 399.600 ;
        RECT 590.400 393.600 592.200 399.600 ;
        RECT 610.800 393.600 612.600 405.600 ;
        RECT 617.400 399.600 618.600 406.500 ;
        RECT 634.950 399.600 636.150 412.950 ;
        RECT 659.400 399.600 660.600 412.950 ;
        RECT 677.850 399.600 679.050 412.950 ;
        RECT 683.100 411.150 684.900 412.950 ;
        RECT 695.100 411.150 696.900 412.950 ;
        RECT 698.700 405.600 699.600 412.950 ;
        RECT 701.100 411.150 702.900 412.950 ;
        RECT 716.100 411.150 717.900 412.950 ;
        RECT 719.400 405.600 720.300 412.950 ;
        RECT 722.100 411.150 723.900 412.950 ;
        RECT 698.700 404.400 702.300 405.600 ;
        RECT 616.800 393.600 618.600 399.600 ;
        RECT 634.800 393.600 636.600 399.600 ;
        RECT 658.800 393.600 660.600 399.600 ;
        RECT 677.400 393.600 679.200 399.600 ;
        RECT 700.500 393.600 702.300 404.400 ;
        RECT 716.700 404.400 720.300 405.600 ;
        RECT 726.150 407.700 727.050 422.400 ;
        RECT 734.550 421.800 736.350 423.600 ;
        RECT 737.850 423.450 742.800 424.500 ;
        RECT 750.300 424.500 751.350 425.400 ;
        RECT 737.850 422.700 739.650 423.450 ;
        RECT 750.300 423.300 754.050 424.500 ;
        RECT 751.950 422.400 754.050 423.300 ;
        RECT 757.650 422.400 759.450 428.400 ;
        RECT 734.850 420.000 735.900 421.800 ;
        RECT 745.050 420.000 746.850 420.600 ;
        RECT 734.850 418.800 746.850 420.000 ;
        RECT 729.000 417.600 735.900 418.800 ;
        RECT 729.000 416.850 729.900 417.600 ;
        RECT 734.100 417.000 735.900 417.600 ;
        RECT 728.100 415.050 729.900 416.850 ;
        RECT 731.100 415.800 732.900 416.400 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 731.100 414.600 739.050 415.800 ;
        RECT 736.950 412.950 739.050 414.600 ;
        RECT 735.450 407.700 737.250 408.000 ;
        RECT 726.150 407.100 737.250 407.700 ;
        RECT 726.150 406.500 743.850 407.100 ;
        RECT 726.150 405.600 727.050 406.500 ;
        RECT 735.450 406.200 743.850 406.500 ;
        RECT 716.700 393.600 718.500 404.400 ;
        RECT 726.150 393.600 727.950 405.600 ;
        RECT 740.250 404.700 742.050 405.300 ;
        RECT 734.550 403.500 742.050 404.700 ;
        RECT 742.950 404.100 743.850 406.200 ;
        RECT 745.950 406.200 746.850 418.800 ;
        RECT 758.250 415.050 759.450 422.400 ;
        RECT 770.400 423.300 772.200 428.400 ;
        RECT 776.400 423.300 778.200 428.400 ;
        RECT 770.400 421.950 778.200 423.300 ;
        RECT 779.400 422.400 781.200 428.400 ;
        RECT 779.400 420.300 780.600 422.400 ;
        RECT 796.800 421.200 798.600 428.400 ;
        RECT 814.800 427.500 822.600 428.400 ;
        RECT 814.800 422.400 816.600 427.500 ;
        RECT 817.800 422.400 819.600 426.600 ;
        RECT 820.800 423.000 822.600 427.500 ;
        RECT 826.800 423.000 828.600 428.400 ;
        RECT 829.950 424.950 832.050 427.050 ;
        RECT 838.800 425.400 840.600 428.400 ;
        RECT 776.850 419.250 780.600 420.300 ;
        RECT 794.400 420.300 798.600 421.200 ;
        RECT 802.950 420.450 805.050 421.050 ;
        RECT 818.400 420.900 819.300 422.400 ;
        RECT 820.800 422.100 828.600 423.000 ;
        RECT 830.550 421.050 831.450 424.950 ;
        RECT 832.950 421.950 835.050 424.050 ;
        RECT 814.950 420.450 817.050 420.900 ;
        RECT 765.000 417.450 769.050 418.050 ;
        RECT 764.550 415.950 769.050 417.450 ;
        RECT 764.550 415.050 765.450 415.950 ;
        RECT 773.100 415.050 774.900 416.850 ;
        RECT 776.850 415.050 778.050 419.250 ;
        RECT 781.950 417.450 786.000 418.050 ;
        RECT 779.100 415.050 780.900 416.850 ;
        RECT 781.950 415.950 786.450 417.450 ;
        RECT 753.150 413.250 759.450 415.050 ;
        RECT 762.000 414.900 765.450 415.050 ;
        RECT 754.950 412.950 759.450 413.250 ;
        RECT 755.250 407.400 757.050 409.200 ;
        RECT 751.950 406.200 756.150 407.400 ;
        RECT 745.950 405.300 751.050 406.200 ;
        RECT 751.950 405.300 754.050 406.200 ;
        RECT 758.250 405.600 759.450 412.950 ;
        RECT 760.950 413.550 765.450 414.900 ;
        RECT 760.950 412.950 765.000 413.550 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 778.950 412.950 781.050 415.050 ;
        RECT 760.950 412.800 763.050 412.950 ;
        RECT 763.950 411.450 768.000 412.050 ;
        RECT 763.950 411.000 768.450 411.450 ;
        RECT 770.100 411.150 771.900 412.950 ;
        RECT 763.950 409.950 769.050 411.000 ;
        RECT 766.950 406.950 769.050 409.950 ;
        RECT 750.150 404.400 751.050 405.300 ;
        RECT 747.450 404.100 749.250 404.400 ;
        RECT 734.550 402.600 735.750 403.500 ;
        RECT 742.950 403.200 749.250 404.100 ;
        RECT 747.450 402.600 749.250 403.200 ;
        RECT 750.150 402.600 752.850 404.400 ;
        RECT 730.950 400.500 735.750 402.600 ;
        RECT 738.450 401.550 740.250 402.300 ;
        RECT 743.250 401.550 745.050 402.300 ;
        RECT 738.450 400.500 745.050 401.550 ;
        RECT 734.550 399.600 735.750 400.500 ;
        RECT 734.550 393.600 736.350 399.600 ;
        RECT 742.350 393.600 744.150 400.500 ;
        RECT 750.150 399.600 754.050 401.700 ;
        RECT 750.150 393.600 751.950 399.600 ;
        RECT 757.650 393.600 759.450 405.600 ;
        RECT 775.950 399.600 777.150 412.950 ;
        RECT 785.550 412.050 786.450 415.950 ;
        RECT 791.100 415.050 792.900 416.850 ;
        RECT 794.400 415.050 795.600 420.300 ;
        RECT 802.950 419.550 817.050 420.450 ;
        RECT 818.400 419.700 823.050 420.900 ;
        RECT 802.950 418.950 805.050 419.550 ;
        RECT 814.950 418.800 817.050 419.550 ;
        RECT 799.950 417.450 804.000 418.050 ;
        RECT 811.950 417.450 814.050 418.050 ;
        RECT 797.100 415.050 798.900 416.850 ;
        RECT 799.950 415.950 804.450 417.450 ;
        RECT 806.550 417.000 814.050 417.450 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 796.950 412.950 799.050 415.050 ;
        RECT 785.550 410.550 790.050 412.050 ;
        RECT 786.000 409.950 790.050 410.550 ;
        RECT 794.400 399.600 795.600 412.950 ;
        RECT 803.550 412.050 804.450 415.950 ;
        RECT 805.950 416.550 814.050 417.000 ;
        RECT 805.950 412.950 808.050 416.550 ;
        RECT 811.950 415.950 814.050 416.550 ;
        RECT 818.100 415.050 819.900 416.850 ;
        RECT 821.700 415.050 823.050 419.700 ;
        RECT 826.950 419.550 831.450 421.050 ;
        RECT 826.950 418.950 831.000 419.550 ;
        RECT 824.100 415.050 825.900 416.850 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 817.950 412.950 820.050 415.050 ;
        RECT 820.950 412.950 823.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 799.950 410.550 804.450 412.050 ;
        RECT 815.100 411.150 816.900 412.950 ;
        RECT 799.950 409.950 804.000 410.550 ;
        RECT 796.950 408.450 799.050 408.750 ;
        RECT 805.950 408.450 808.050 409.050 ;
        RECT 796.950 407.550 808.050 408.450 ;
        RECT 796.950 406.650 799.050 407.550 ;
        RECT 805.950 406.950 808.050 407.550 ;
        RECT 821.700 405.600 822.900 412.950 ;
        RECT 827.100 411.150 828.900 412.950 ;
        RECT 833.550 412.050 834.450 421.950 ;
        RECT 839.400 415.050 840.600 425.400 ;
        RECT 850.950 424.050 853.050 427.050 ;
        RECT 847.950 423.000 853.050 424.050 ;
        RECT 847.950 422.550 852.450 423.000 ;
        RECT 847.950 421.950 852.000 422.550 ;
        RECT 859.200 422.400 861.000 428.400 ;
        RECT 881.400 425.400 883.200 428.400 ;
        RECT 902.400 425.400 904.200 428.400 ;
        RECT 854.100 415.050 855.900 416.850 ;
        RECT 859.950 415.050 861.000 422.400 ;
        RECT 862.950 420.450 865.050 421.050 ;
        RECT 871.950 420.450 874.050 421.050 ;
        RECT 862.950 419.550 874.050 420.450 ;
        RECT 862.950 418.950 865.050 419.550 ;
        RECT 871.950 418.950 874.050 419.550 ;
        RECT 868.950 417.450 873.000 418.050 ;
        RECT 866.100 415.050 867.900 416.850 ;
        RECT 868.950 415.950 873.450 417.450 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 841.950 412.950 844.050 415.050 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 865.950 412.950 868.050 415.050 ;
        RECT 829.950 410.550 834.450 412.050 ;
        RECT 829.950 409.950 834.000 410.550 ;
        RECT 775.800 393.600 777.600 399.600 ;
        RECT 794.400 393.600 796.200 399.600 ;
        RECT 820.800 393.600 824.100 405.600 ;
        RECT 839.400 399.600 840.600 412.950 ;
        RECT 842.100 411.150 843.900 412.950 ;
        RECT 857.100 411.150 858.900 412.950 ;
        RECT 860.100 407.400 861.000 412.950 ;
        RECT 863.100 411.150 864.900 412.950 ;
        RECT 872.550 412.050 873.450 415.950 ;
        RECT 881.700 415.050 882.600 425.400 ;
        RECT 883.950 420.450 886.050 421.200 ;
        RECT 883.950 419.550 891.450 420.450 ;
        RECT 883.950 419.100 886.050 419.550 ;
        RECT 877.950 412.950 880.050 415.050 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 883.950 412.950 886.050 415.050 ;
        RECT 868.950 410.550 873.450 412.050 ;
        RECT 878.100 411.150 879.900 412.950 ;
        RECT 868.950 409.950 873.000 410.550 ;
        RECT 860.100 406.500 865.200 407.400 ;
        RECT 838.800 393.600 840.600 399.600 ;
        RECT 854.400 404.400 862.200 405.300 ;
        RECT 854.400 393.600 856.200 404.400 ;
        RECT 860.400 394.500 862.200 404.400 ;
        RECT 863.400 395.400 865.200 406.500 ;
        RECT 881.700 405.600 882.600 412.950 ;
        RECT 884.100 411.150 885.900 412.950 ;
        RECT 890.550 412.050 891.450 419.550 ;
        RECT 902.400 415.050 903.600 425.400 ;
        RECT 898.950 412.950 901.050 415.050 ;
        RECT 901.950 412.950 904.050 415.050 ;
        RECT 886.950 410.550 891.450 412.050 ;
        RECT 899.100 411.150 900.900 412.950 ;
        RECT 886.950 409.950 891.000 410.550 ;
        RECT 866.400 394.500 868.200 405.600 ;
        RECT 881.700 404.400 885.300 405.600 ;
        RECT 860.400 393.600 868.200 394.500 ;
        RECT 883.500 393.600 885.300 404.400 ;
        RECT 902.400 399.600 903.600 412.950 ;
        RECT 902.400 393.600 904.200 399.600 ;
        RECT 10.800 377.400 12.600 389.400 ;
        RECT 16.800 383.400 18.600 389.400 ;
        RECT 11.400 370.050 12.300 377.400 ;
        RECT 14.100 370.050 15.900 371.850 ;
        RECT 10.950 367.950 13.050 370.050 ;
        RECT 13.950 367.950 16.050 370.050 ;
        RECT 11.400 360.600 12.300 367.950 ;
        RECT 17.700 363.300 18.600 383.400 ;
        RECT 35.400 383.400 37.200 389.400 ;
        RECT 22.950 372.450 27.000 373.050 ;
        RECT 22.950 370.950 27.450 372.450 ;
        RECT 19.950 367.950 22.050 370.050 ;
        RECT 20.100 366.150 21.900 367.950 ;
        RECT 26.550 367.050 27.450 370.950 ;
        RECT 35.400 370.050 36.600 383.400 ;
        RECT 53.400 378.300 55.200 389.400 ;
        RECT 59.400 378.300 61.200 389.400 ;
        RECT 53.400 377.400 61.200 378.300 ;
        RECT 62.400 377.400 64.200 389.400 ;
        RECT 76.800 383.400 78.600 389.400 ;
        RECT 97.800 383.400 99.600 389.400 ;
        RECT 56.100 370.050 57.900 371.850 ;
        RECT 62.700 370.050 63.600 377.400 ;
        RECT 77.400 370.050 78.600 383.400 ;
        RECT 80.100 370.050 81.900 371.850 ;
        RECT 92.100 370.050 93.900 371.850 ;
        RECT 97.950 370.050 99.150 383.400 ;
        RECT 119.700 378.600 121.500 389.400 ;
        RECT 142.800 383.400 144.600 389.400 ;
        RECT 160.800 383.400 162.600 389.400 ;
        RECT 119.700 377.400 123.300 378.600 ;
        RECT 119.100 370.050 120.900 371.850 ;
        RECT 122.400 370.050 123.300 377.400 ;
        RECT 125.100 370.050 126.900 371.850 ;
        RECT 143.400 370.050 144.600 383.400 ;
        RECT 153.000 372.450 157.050 373.050 ;
        RECT 152.550 370.950 157.050 372.450 ;
        RECT 31.950 367.950 34.050 370.050 ;
        RECT 34.950 367.950 37.050 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 76.950 367.950 79.050 370.050 ;
        RECT 79.950 367.950 82.050 370.050 ;
        RECT 91.950 367.950 94.050 370.050 ;
        RECT 94.950 367.950 97.050 370.050 ;
        RECT 97.950 367.950 100.050 370.050 ;
        RECT 100.950 367.950 103.050 370.050 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 124.950 367.950 127.050 370.050 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 26.550 365.550 31.050 367.050 ;
        RECT 32.100 366.150 33.900 367.950 ;
        RECT 27.000 364.950 31.050 365.550 ;
        RECT 14.100 362.400 21.600 363.300 ;
        RECT 14.100 361.500 15.900 362.400 ;
        RECT 11.400 358.800 14.100 360.600 ;
        RECT 12.300 354.600 14.100 358.800 ;
        RECT 19.800 354.600 21.600 362.400 ;
        RECT 35.400 362.700 36.600 367.950 ;
        RECT 38.100 366.150 39.900 367.950 ;
        RECT 53.100 366.150 54.900 367.950 ;
        RECT 59.100 366.150 60.900 367.950 ;
        RECT 35.400 361.800 39.600 362.700 ;
        RECT 37.800 354.600 39.600 361.800 ;
        RECT 62.700 360.600 63.600 367.950 ;
        RECT 58.500 359.400 63.600 360.600 ;
        RECT 58.500 354.600 60.300 359.400 ;
        RECT 77.400 357.600 78.600 367.950 ;
        RECT 95.100 366.150 96.900 367.950 ;
        RECT 98.850 363.750 100.050 367.950 ;
        RECT 101.100 366.150 102.900 367.950 ;
        RECT 98.850 362.700 102.600 363.750 ;
        RECT 76.800 354.600 78.600 357.600 ;
        RECT 92.400 359.700 100.200 361.050 ;
        RECT 92.400 354.600 94.200 359.700 ;
        RECT 98.400 354.600 100.200 359.700 ;
        RECT 101.400 360.600 102.600 362.700 ;
        RECT 101.400 354.600 103.200 360.600 ;
        RECT 122.400 357.600 123.300 367.950 ;
        RECT 140.100 366.150 141.900 367.950 ;
        RECT 143.400 362.700 144.600 367.950 ;
        RECT 146.100 366.150 147.900 367.950 ;
        RECT 140.400 361.800 144.600 362.700 ;
        RECT 145.950 363.450 148.050 364.050 ;
        RECT 152.550 363.450 153.450 370.950 ;
        RECT 161.400 370.050 162.600 383.400 ;
        RECT 179.400 383.400 181.200 389.400 ;
        RECT 199.800 383.400 201.600 389.400 ;
        RECT 220.800 383.400 222.600 389.400 ;
        RECT 163.950 378.450 166.050 379.050 ;
        RECT 175.950 378.450 178.050 379.050 ;
        RECT 163.950 377.550 178.050 378.450 ;
        RECT 163.950 376.950 166.050 377.550 ;
        RECT 175.950 376.950 178.050 377.550 ;
        RECT 176.100 370.050 177.900 371.850 ;
        RECT 179.400 370.050 180.600 383.400 ;
        RECT 181.950 372.450 186.000 373.050 ;
        RECT 181.950 372.000 186.450 372.450 ;
        RECT 181.950 370.950 187.050 372.000 ;
        RECT 187.950 370.950 190.050 373.050 ;
        RECT 157.950 367.950 160.050 370.050 ;
        RECT 160.950 367.950 163.050 370.050 ;
        RECT 163.950 367.950 166.050 370.050 ;
        RECT 175.950 367.950 178.050 370.050 ;
        RECT 178.950 367.950 181.050 370.050 ;
        RECT 158.100 366.150 159.900 367.950 ;
        RECT 145.950 362.550 153.450 363.450 ;
        RECT 161.400 362.700 162.600 367.950 ;
        RECT 164.100 366.150 165.900 367.950 ;
        RECT 145.950 361.950 148.050 362.550 ;
        RECT 158.400 361.800 162.600 362.700 ;
        RECT 121.800 354.600 123.600 357.600 ;
        RECT 140.400 354.600 142.200 361.800 ;
        RECT 158.400 354.600 160.200 361.800 ;
        RECT 179.400 357.600 180.600 367.950 ;
        RECT 184.950 367.800 187.050 370.950 ;
        RECT 188.550 367.050 189.450 370.950 ;
        RECT 194.100 370.050 195.900 371.850 ;
        RECT 199.950 370.050 201.150 383.400 ;
        RECT 221.700 383.100 222.600 383.400 ;
        RECT 226.800 383.400 228.600 389.400 ;
        RECT 245.400 383.400 247.200 389.400 ;
        RECT 269.400 383.400 271.200 389.400 ;
        RECT 290.400 383.400 292.200 389.400 ;
        RECT 226.800 383.100 228.300 383.400 ;
        RECT 221.700 382.200 228.300 383.100 ;
        RECT 202.950 375.450 205.050 376.050 ;
        RECT 214.950 375.450 217.050 376.050 ;
        RECT 202.950 374.550 217.050 375.450 ;
        RECT 202.950 373.950 205.050 374.550 ;
        RECT 214.950 373.950 217.050 374.550 ;
        RECT 221.700 370.050 222.600 382.200 ;
        RECT 227.100 370.050 228.900 371.850 ;
        RECT 245.850 370.050 247.050 383.400 ;
        RECT 251.100 370.050 252.900 371.850 ;
        RECT 269.850 370.050 271.050 383.400 ;
        RECT 275.100 370.050 276.900 371.850 ;
        RECT 290.400 370.050 291.600 383.400 ;
        RECT 292.950 381.450 295.050 382.050 ;
        RECT 304.950 381.450 307.050 382.050 ;
        RECT 292.950 380.550 307.050 381.450 ;
        RECT 292.950 379.950 295.050 380.550 ;
        RECT 304.950 379.950 307.050 380.550 ;
        RECT 310.800 377.400 312.600 389.400 ;
        RECT 316.800 383.400 318.600 389.400 ;
        RECT 292.950 375.450 295.050 376.050 ;
        RECT 307.950 375.450 310.050 376.050 ;
        RECT 292.950 374.550 310.050 375.450 ;
        RECT 292.950 373.950 295.050 374.550 ;
        RECT 307.950 373.950 310.050 374.550 ;
        RECT 311.400 370.050 312.300 377.400 ;
        RECT 314.100 370.050 315.900 371.850 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 199.950 367.950 202.050 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 220.950 367.950 223.050 370.050 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 226.950 367.950 229.050 370.050 ;
        RECT 229.950 367.950 232.050 370.050 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 244.950 367.950 247.050 370.050 ;
        RECT 247.950 367.950 250.050 370.050 ;
        RECT 250.950 367.950 253.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 274.950 367.950 277.050 370.050 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 289.950 367.950 292.050 370.050 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 188.550 365.550 193.050 367.050 ;
        RECT 197.100 366.150 198.900 367.950 ;
        RECT 189.000 364.950 193.050 365.550 ;
        RECT 200.850 363.750 202.050 367.950 ;
        RECT 203.100 366.150 204.900 367.950 ;
        RECT 221.700 364.200 222.600 367.950 ;
        RECT 224.100 366.150 225.900 367.950 ;
        RECT 230.100 366.150 231.900 367.950 ;
        RECT 242.100 366.150 243.900 367.950 ;
        RECT 200.850 362.700 204.600 363.750 ;
        RECT 221.700 363.000 225.000 364.200 ;
        RECT 244.950 363.750 246.150 367.950 ;
        RECT 248.100 366.150 249.900 367.950 ;
        RECT 266.100 366.150 267.900 367.950 ;
        RECT 268.950 363.750 270.150 367.950 ;
        RECT 272.100 366.150 273.900 367.950 ;
        RECT 287.100 366.150 288.900 367.950 ;
        RECT 194.400 359.700 202.200 361.050 ;
        RECT 179.400 354.600 181.200 357.600 ;
        RECT 194.400 354.600 196.200 359.700 ;
        RECT 200.400 354.600 202.200 359.700 ;
        RECT 203.400 360.600 204.600 362.700 ;
        RECT 203.400 354.600 205.200 360.600 ;
        RECT 223.200 354.600 225.000 363.000 ;
        RECT 242.400 362.700 246.150 363.750 ;
        RECT 266.400 362.700 270.150 363.750 ;
        RECT 290.400 362.700 291.600 367.950 ;
        RECT 293.100 366.150 294.900 367.950 ;
        RECT 242.400 360.600 243.600 362.700 ;
        RECT 241.800 354.600 243.600 360.600 ;
        RECT 244.800 359.700 252.600 361.050 ;
        RECT 266.400 360.600 267.600 362.700 ;
        RECT 290.400 361.800 294.600 362.700 ;
        RECT 244.800 354.600 246.600 359.700 ;
        RECT 250.800 354.600 252.600 359.700 ;
        RECT 265.800 354.600 267.600 360.600 ;
        RECT 268.800 359.700 276.600 361.050 ;
        RECT 268.800 354.600 270.600 359.700 ;
        RECT 274.800 354.600 276.600 359.700 ;
        RECT 292.800 354.600 294.600 361.800 ;
        RECT 311.400 360.600 312.300 367.950 ;
        RECT 317.700 363.300 318.600 383.400 ;
        RECT 334.800 377.400 336.600 389.400 ;
        RECT 340.800 383.400 342.600 389.400 ;
        RECT 334.800 370.050 336.000 377.400 ;
        RECT 341.400 376.500 342.600 383.400 ;
        RECT 336.900 375.600 342.600 376.500 ;
        RECT 352.800 377.400 354.600 389.400 ;
        RECT 358.800 383.400 360.600 389.400 ;
        RECT 336.900 374.700 338.850 375.600 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 334.800 367.950 337.050 370.050 ;
        RECT 320.100 366.150 321.900 367.950 ;
        RECT 314.100 362.400 321.600 363.300 ;
        RECT 314.100 361.500 315.900 362.400 ;
        RECT 311.400 358.800 314.100 360.600 ;
        RECT 312.300 354.600 314.100 358.800 ;
        RECT 319.800 354.600 321.600 362.400 ;
        RECT 334.800 360.600 336.000 367.950 ;
        RECT 337.950 363.300 338.850 374.700 ;
        RECT 341.100 370.050 342.900 371.850 ;
        RECT 352.800 370.050 354.000 377.400 ;
        RECT 359.400 376.500 360.600 383.400 ;
        RECT 373.800 377.400 375.600 389.400 ;
        RECT 376.800 378.300 378.600 389.400 ;
        RECT 382.800 378.300 384.600 389.400 ;
        RECT 398.400 383.400 400.200 389.400 ;
        RECT 376.800 377.400 384.600 378.300 ;
        RECT 354.900 375.600 360.600 376.500 ;
        RECT 354.900 374.700 356.850 375.600 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 352.800 367.950 355.050 370.050 ;
        RECT 336.900 362.400 338.850 363.300 ;
        RECT 336.900 361.500 342.600 362.400 ;
        RECT 334.800 354.600 336.600 360.600 ;
        RECT 341.400 357.600 342.600 361.500 ;
        RECT 340.800 354.600 342.600 357.600 ;
        RECT 352.800 360.600 354.000 367.950 ;
        RECT 355.950 363.300 356.850 374.700 ;
        RECT 361.950 372.450 364.050 373.050 ;
        RECT 359.100 370.050 360.900 371.850 ;
        RECT 361.950 371.550 369.450 372.450 ;
        RECT 361.950 370.950 364.050 371.550 ;
        RECT 358.950 367.950 361.050 370.050 ;
        RECT 368.550 367.050 369.450 371.550 ;
        RECT 374.400 370.050 375.300 377.400 ;
        RECT 380.100 370.050 381.900 371.850 ;
        RECT 398.850 370.050 400.050 383.400 ;
        RECT 416.400 379.500 418.200 389.400 ;
        RECT 422.400 388.500 430.200 389.400 ;
        RECT 422.400 379.500 424.200 388.500 ;
        RECT 416.400 378.600 424.200 379.500 ;
        RECT 425.400 379.800 427.200 387.600 ;
        RECT 428.400 380.700 430.200 388.500 ;
        RECT 432.000 388.500 439.800 389.400 ;
        RECT 432.000 379.800 433.800 388.500 ;
        RECT 425.400 378.900 433.800 379.800 ;
        RECT 435.000 379.800 436.800 387.600 ;
        RECT 435.000 377.400 436.200 379.800 ;
        RECT 438.000 379.200 439.800 388.500 ;
        RECT 452.400 378.300 454.200 389.400 ;
        RECT 458.400 378.300 460.200 389.400 ;
        RECT 452.400 377.400 460.200 378.300 ;
        RECT 461.400 377.400 463.200 389.400 ;
        RECT 476.400 383.400 478.200 389.400 ;
        RECT 496.800 383.400 498.600 389.400 ;
        RECT 512.400 383.400 514.200 389.400 ;
        RECT 432.750 376.200 436.200 377.400 ;
        RECT 403.950 375.450 406.050 376.050 ;
        RECT 427.950 375.450 430.050 376.050 ;
        RECT 403.950 374.550 430.050 375.450 ;
        RECT 403.950 373.950 406.050 374.550 ;
        RECT 427.950 373.950 430.050 374.550 ;
        RECT 414.000 372.450 418.050 373.050 ;
        RECT 404.100 370.050 405.900 371.850 ;
        RECT 413.550 370.950 418.050 372.450 ;
        RECT 373.950 367.950 376.050 370.050 ;
        RECT 376.950 367.950 379.050 370.050 ;
        RECT 379.950 367.950 382.050 370.050 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 394.950 367.950 397.050 370.050 ;
        RECT 397.950 367.950 400.050 370.050 ;
        RECT 400.950 367.950 403.050 370.050 ;
        RECT 403.950 367.950 406.050 370.050 ;
        RECT 368.550 365.550 373.050 367.050 ;
        RECT 369.000 364.950 373.050 365.550 ;
        RECT 354.900 362.400 356.850 363.300 ;
        RECT 354.900 361.500 360.600 362.400 ;
        RECT 352.800 354.600 354.600 360.600 ;
        RECT 359.400 357.600 360.600 361.500 ;
        RECT 374.400 360.600 375.300 367.950 ;
        RECT 377.100 366.150 378.900 367.950 ;
        RECT 383.100 366.150 384.900 367.950 ;
        RECT 395.100 366.150 396.900 367.950 ;
        RECT 397.950 363.750 399.150 367.950 ;
        RECT 401.100 366.150 402.900 367.950 ;
        RECT 406.950 366.450 409.050 367.050 ;
        RECT 413.550 366.450 414.450 370.950 ;
        RECT 419.100 369.900 420.900 371.700 ;
        RECT 428.100 369.900 429.900 371.700 ;
        RECT 432.750 369.900 433.950 376.200 ;
        RECT 436.950 372.450 441.000 373.050 ;
        RECT 436.950 370.950 441.450 372.450 ;
        RECT 418.950 367.800 421.050 369.900 ;
        RECT 424.950 367.800 427.050 369.900 ;
        RECT 427.950 367.800 430.050 369.900 ;
        RECT 432.750 367.800 436.050 369.900 ;
        RECT 406.950 365.550 414.450 366.450 ;
        RECT 425.100 366.000 426.900 367.800 ;
        RECT 406.950 364.950 409.050 365.550 ;
        RECT 395.400 362.700 399.150 363.750 ;
        RECT 406.950 363.450 409.050 363.900 ;
        RECT 421.950 363.450 424.050 364.050 ;
        RECT 395.400 360.600 396.600 362.700 ;
        RECT 406.950 362.550 424.050 363.450 ;
        RECT 406.950 361.800 409.050 362.550 ;
        RECT 421.950 361.950 424.050 362.550 ;
        RECT 374.400 359.400 379.500 360.600 ;
        RECT 358.800 354.600 360.600 357.600 ;
        RECT 377.700 354.600 379.500 359.400 ;
        RECT 394.800 354.600 396.600 360.600 ;
        RECT 397.800 359.700 405.600 361.050 ;
        RECT 397.800 354.600 399.600 359.700 ;
        RECT 403.800 354.600 405.600 359.700 ;
        RECT 432.750 359.400 433.950 367.800 ;
        RECT 440.550 367.050 441.450 370.950 ;
        RECT 455.100 370.050 456.900 371.850 ;
        RECT 461.700 370.050 462.600 377.400 ;
        RECT 463.950 372.450 468.000 373.050 ;
        RECT 463.950 370.950 468.450 372.450 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 460.950 367.950 463.050 370.050 ;
        RECT 436.950 365.550 441.450 367.050 ;
        RECT 452.100 366.150 453.900 367.950 ;
        RECT 458.100 366.150 459.900 367.950 ;
        RECT 436.950 364.950 441.000 365.550 ;
        RECT 461.700 360.600 462.600 367.950 ;
        RECT 467.550 367.050 468.450 370.950 ;
        RECT 473.100 370.050 474.900 371.850 ;
        RECT 476.400 370.050 477.600 383.400 ;
        RECT 491.100 370.050 492.900 371.850 ;
        RECT 496.950 370.050 498.150 383.400 ;
        RECT 512.400 376.500 513.600 383.400 ;
        RECT 518.400 377.400 520.200 389.400 ;
        RECT 538.800 383.400 540.600 389.400 ;
        RECT 563.400 383.400 565.200 389.400 ;
        RECT 583.800 383.400 585.600 389.400 ;
        RECT 512.400 375.600 518.100 376.500 ;
        RECT 516.150 374.700 518.100 375.600 ;
        RECT 502.950 372.450 507.000 373.050 ;
        RECT 502.950 370.950 507.450 372.450 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 490.950 367.950 493.050 370.050 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 467.550 365.550 472.050 367.050 ;
        RECT 468.000 364.950 472.050 365.550 ;
        RECT 423.150 358.500 433.950 359.400 ;
        RECT 457.500 359.400 462.600 360.600 ;
        RECT 423.150 357.600 424.200 358.500 ;
        RECT 429.150 357.600 430.200 358.500 ;
        RECT 422.400 354.600 424.200 357.600 ;
        RECT 428.400 354.600 430.200 357.600 ;
        RECT 457.500 354.600 459.300 359.400 ;
        RECT 476.400 357.600 477.600 367.950 ;
        RECT 494.100 366.150 495.900 367.950 ;
        RECT 497.850 363.750 499.050 367.950 ;
        RECT 500.100 366.150 501.900 367.950 ;
        RECT 506.550 367.050 507.450 370.950 ;
        RECT 512.100 370.050 513.900 371.850 ;
        RECT 511.950 367.950 514.050 370.050 ;
        RECT 506.550 365.550 511.050 367.050 ;
        RECT 507.000 364.950 511.050 365.550 ;
        RECT 497.850 362.700 501.600 363.750 ;
        RECT 491.400 359.700 499.200 361.050 ;
        RECT 476.400 354.600 478.200 357.600 ;
        RECT 491.400 354.600 493.200 359.700 ;
        RECT 497.400 354.600 499.200 359.700 ;
        RECT 500.400 360.600 501.600 362.700 ;
        RECT 516.150 363.300 517.050 374.700 ;
        RECT 519.000 370.050 520.200 377.400 ;
        RECT 533.100 370.050 534.900 371.850 ;
        RECT 538.950 370.050 540.150 383.400 ;
        RECT 547.950 375.450 550.050 376.050 ;
        RECT 559.950 375.450 562.050 376.200 ;
        RECT 547.950 374.550 562.050 375.450 ;
        RECT 547.950 373.950 550.050 374.550 ;
        RECT 559.950 374.100 562.050 374.550 ;
        RECT 563.850 370.050 565.050 383.400 ;
        RECT 569.100 370.050 570.900 371.850 ;
        RECT 584.400 370.050 585.600 383.400 ;
        RECT 599.400 378.300 601.200 389.400 ;
        RECT 605.400 378.300 607.200 389.400 ;
        RECT 599.400 377.400 607.200 378.300 ;
        RECT 608.400 377.400 610.200 389.400 ;
        RECT 628.800 383.400 630.600 389.400 ;
        RECT 587.100 370.050 588.900 371.850 ;
        RECT 602.100 370.050 603.900 371.850 ;
        RECT 608.700 370.050 609.600 377.400 ;
        RECT 623.100 370.050 624.900 371.850 ;
        RECT 628.950 370.050 630.150 383.400 ;
        RECT 650.700 378.600 652.500 389.400 ;
        RECT 671.400 383.400 673.200 389.400 ;
        RECT 692.400 383.400 694.200 389.400 ;
        RECT 650.700 377.400 654.300 378.600 ;
        RECT 650.100 370.050 651.900 371.850 ;
        RECT 653.400 370.050 654.300 377.400 ;
        RECT 655.950 375.450 658.050 376.050 ;
        RECT 655.950 374.550 663.450 375.450 ;
        RECT 655.950 373.950 658.050 374.550 ;
        RECT 656.100 370.050 657.900 371.850 ;
        RECT 517.950 367.950 520.200 370.050 ;
        RECT 532.950 367.950 535.050 370.050 ;
        RECT 535.950 367.950 538.050 370.050 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 559.950 367.950 562.050 370.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 565.950 367.950 568.050 370.050 ;
        RECT 568.950 367.950 571.050 370.050 ;
        RECT 583.950 367.950 586.050 370.050 ;
        RECT 586.950 367.950 589.050 370.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 516.150 362.400 518.100 363.300 ;
        RECT 512.400 361.500 518.100 362.400 ;
        RECT 500.400 354.600 502.200 360.600 ;
        RECT 512.400 357.600 513.600 361.500 ;
        RECT 519.000 360.600 520.200 367.950 ;
        RECT 536.100 366.150 537.900 367.950 ;
        RECT 539.850 363.750 541.050 367.950 ;
        RECT 542.100 366.150 543.900 367.950 ;
        RECT 560.100 366.150 561.900 367.950 ;
        RECT 562.950 363.750 564.150 367.950 ;
        RECT 566.100 366.150 567.900 367.950 ;
        RECT 539.850 362.700 543.600 363.750 ;
        RECT 512.400 354.600 514.200 357.600 ;
        RECT 518.400 354.600 520.200 360.600 ;
        RECT 533.400 359.700 541.200 361.050 ;
        RECT 533.400 354.600 535.200 359.700 ;
        RECT 539.400 354.600 541.200 359.700 ;
        RECT 542.400 360.600 543.600 362.700 ;
        RECT 560.400 362.700 564.150 363.750 ;
        RECT 560.400 360.600 561.600 362.700 ;
        RECT 542.400 354.600 544.200 360.600 ;
        RECT 559.800 354.600 561.600 360.600 ;
        RECT 562.800 359.700 570.600 361.050 ;
        RECT 562.800 354.600 564.600 359.700 ;
        RECT 568.800 354.600 570.600 359.700 ;
        RECT 584.400 357.600 585.600 367.950 ;
        RECT 599.100 366.150 600.900 367.950 ;
        RECT 605.100 366.150 606.900 367.950 ;
        RECT 608.700 360.600 609.600 367.950 ;
        RECT 626.100 366.150 627.900 367.950 ;
        RECT 629.850 363.750 631.050 367.950 ;
        RECT 632.100 366.150 633.900 367.950 ;
        RECT 629.850 362.700 633.600 363.750 ;
        RECT 583.800 354.600 585.600 357.600 ;
        RECT 604.500 359.400 609.600 360.600 ;
        RECT 623.400 359.700 631.200 361.050 ;
        RECT 604.500 354.600 606.300 359.400 ;
        RECT 623.400 354.600 625.200 359.700 ;
        RECT 629.400 354.600 631.200 359.700 ;
        RECT 632.400 360.600 633.600 362.700 ;
        RECT 632.400 354.600 634.200 360.600 ;
        RECT 653.400 357.600 654.300 367.950 ;
        RECT 662.550 367.050 663.450 374.550 ;
        RECT 671.400 370.050 672.600 383.400 ;
        RECT 692.850 370.050 694.050 383.400 ;
        RECT 713.700 378.600 715.500 389.400 ;
        RECT 733.800 383.400 735.600 389.400 ;
        RECT 751.800 383.400 753.600 389.400 ;
        RECT 713.700 377.400 717.300 378.600 ;
        RECT 700.950 372.450 705.000 373.050 ;
        RECT 698.100 370.050 699.900 371.850 ;
        RECT 700.950 370.950 705.450 372.450 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 670.950 367.950 673.050 370.050 ;
        RECT 673.950 367.950 676.050 370.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 691.950 367.950 694.050 370.050 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 697.950 367.950 700.050 370.050 ;
        RECT 658.950 365.550 663.450 367.050 ;
        RECT 668.100 366.150 669.900 367.950 ;
        RECT 658.950 364.950 663.000 365.550 ;
        RECT 671.400 362.700 672.600 367.950 ;
        RECT 674.100 366.150 675.900 367.950 ;
        RECT 689.100 366.150 690.900 367.950 ;
        RECT 691.950 363.750 693.150 367.950 ;
        RECT 695.100 366.150 696.900 367.950 ;
        RECT 704.550 366.450 705.450 370.950 ;
        RECT 713.100 370.050 714.900 371.850 ;
        RECT 716.400 370.050 717.300 377.400 ;
        RECT 721.950 372.450 726.000 373.050 ;
        RECT 719.100 370.050 720.900 371.850 ;
        RECT 721.950 370.950 726.450 372.450 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 715.950 367.950 718.050 370.050 ;
        RECT 718.950 367.950 721.050 370.050 ;
        RECT 709.950 366.450 712.050 367.050 ;
        RECT 704.550 365.550 712.050 366.450 ;
        RECT 709.950 364.950 712.050 365.550 ;
        RECT 689.400 362.700 693.150 363.750 ;
        RECT 671.400 361.800 675.600 362.700 ;
        RECT 652.800 354.600 654.600 357.600 ;
        RECT 673.800 354.600 675.600 361.800 ;
        RECT 689.400 360.600 690.600 362.700 ;
        RECT 688.800 354.600 690.600 360.600 ;
        RECT 691.800 359.700 699.600 361.050 ;
        RECT 691.800 354.600 693.600 359.700 ;
        RECT 697.800 354.600 699.600 359.700 ;
        RECT 716.400 357.600 717.300 367.950 ;
        RECT 725.550 367.050 726.450 370.950 ;
        RECT 734.400 370.050 735.600 383.400 ;
        RECT 752.700 383.100 753.600 383.400 ;
        RECT 757.800 383.400 759.600 389.400 ;
        RECT 776.400 383.400 778.200 389.400 ;
        RECT 797.400 383.400 799.200 389.400 ;
        RECT 757.800 383.100 759.300 383.400 ;
        RECT 752.700 382.200 759.300 383.100 ;
        RECT 752.700 370.050 753.600 382.200 ;
        RECT 763.950 372.450 768.000 373.050 ;
        RECT 758.100 370.050 759.900 371.850 ;
        RECT 763.950 370.950 768.450 372.450 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 721.950 365.550 726.450 367.050 ;
        RECT 731.100 366.150 732.900 367.950 ;
        RECT 721.950 364.950 726.000 365.550 ;
        RECT 734.400 362.700 735.600 367.950 ;
        RECT 737.100 366.150 738.900 367.950 ;
        RECT 752.700 364.200 753.600 367.950 ;
        RECT 755.100 366.150 756.900 367.950 ;
        RECT 761.100 366.150 762.900 367.950 ;
        RECT 767.550 367.050 768.450 370.950 ;
        RECT 773.100 370.050 774.900 371.850 ;
        RECT 776.400 370.050 777.600 383.400 ;
        RECT 797.850 370.050 799.050 383.400 ;
        RECT 815.400 377.400 817.200 389.400 ;
        RECT 822.900 378.900 824.700 389.400 ;
        RECT 842.400 383.400 844.200 389.400 ;
        RECT 863.400 383.400 865.200 389.400 ;
        RECT 822.900 377.400 825.300 378.900 ;
        RECT 815.400 375.900 816.600 377.400 ;
        RECT 815.400 374.700 822.600 375.900 ;
        RECT 820.800 374.100 822.600 374.700 ;
        RECT 803.100 370.050 804.900 371.850 ;
        RECT 818.100 370.050 819.900 371.850 ;
        RECT 772.950 367.950 775.050 370.050 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 793.950 367.950 796.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 799.950 367.950 802.050 370.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 814.950 367.950 817.050 370.050 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 767.550 365.550 772.050 367.050 ;
        RECT 768.000 364.950 772.050 365.550 ;
        RECT 752.700 363.000 756.000 364.200 ;
        RECT 731.400 361.800 735.600 362.700 ;
        RECT 715.800 354.600 717.600 357.600 ;
        RECT 731.400 354.600 733.200 361.800 ;
        RECT 754.200 354.600 756.000 363.000 ;
        RECT 776.400 357.600 777.600 367.950 ;
        RECT 794.100 366.150 795.900 367.950 ;
        RECT 796.950 363.750 798.150 367.950 ;
        RECT 800.100 366.150 801.900 367.950 ;
        RECT 815.100 366.150 816.900 367.950 ;
        RECT 794.400 362.700 798.150 363.750 ;
        RECT 821.700 363.600 822.600 374.100 ;
        RECT 823.950 370.050 825.300 377.400 ;
        RECT 842.850 370.050 844.050 383.400 ;
        RECT 848.100 370.050 849.900 371.850 ;
        RECT 863.850 370.050 865.050 383.400 ;
        RECT 884.700 378.600 886.500 389.400 ;
        RECT 905.400 383.400 907.200 389.400 ;
        RECT 884.700 377.400 888.300 378.600 ;
        RECT 880.950 372.450 883.050 373.050 ;
        RECT 869.100 370.050 870.900 371.850 ;
        RECT 875.550 371.550 883.050 372.450 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 859.950 367.950 862.050 370.050 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 865.950 367.950 868.050 370.050 ;
        RECT 868.950 367.950 871.050 370.050 ;
        RECT 820.800 362.700 822.600 363.600 ;
        RECT 794.400 360.600 795.600 362.700 ;
        RECT 819.300 361.800 822.600 362.700 ;
        RECT 776.400 354.600 778.200 357.600 ;
        RECT 793.800 354.600 795.600 360.600 ;
        RECT 796.800 359.700 804.600 361.050 ;
        RECT 796.800 354.600 798.600 359.700 ;
        RECT 802.800 354.600 804.600 359.700 ;
        RECT 819.300 357.600 820.200 361.800 ;
        RECT 825.000 360.600 826.050 367.950 ;
        RECT 839.100 366.150 840.900 367.950 ;
        RECT 841.950 363.750 843.150 367.950 ;
        RECT 845.100 366.150 846.900 367.950 ;
        RECT 860.100 366.150 861.900 367.950 ;
        RECT 862.950 363.750 864.150 367.950 ;
        RECT 866.100 366.150 867.900 367.950 ;
        RECT 875.550 367.050 876.450 371.550 ;
        RECT 880.950 370.950 883.050 371.550 ;
        RECT 884.100 370.050 885.900 371.850 ;
        RECT 887.400 370.050 888.300 377.400 ;
        RECT 901.950 375.450 904.050 376.050 ;
        RECT 896.550 374.550 904.050 375.450 ;
        RECT 890.100 370.050 891.900 371.850 ;
        RECT 883.950 367.950 886.050 370.050 ;
        RECT 886.950 367.950 889.050 370.050 ;
        RECT 889.950 367.950 892.050 370.050 ;
        RECT 871.950 365.550 876.450 367.050 ;
        RECT 871.950 364.950 876.000 365.550 ;
        RECT 839.400 362.700 843.150 363.750 ;
        RECT 860.400 362.700 864.150 363.750 ;
        RECT 839.400 360.600 840.600 362.700 ;
        RECT 818.400 354.600 820.200 357.600 ;
        RECT 824.400 354.600 826.200 360.600 ;
        RECT 838.800 354.600 840.600 360.600 ;
        RECT 841.800 359.700 849.600 361.050 ;
        RECT 860.400 360.600 861.600 362.700 ;
        RECT 841.800 354.600 843.600 359.700 ;
        RECT 847.800 354.600 849.600 359.700 ;
        RECT 859.800 354.600 861.600 360.600 ;
        RECT 862.800 359.700 870.600 361.050 ;
        RECT 862.800 354.600 864.600 359.700 ;
        RECT 868.800 354.600 870.600 359.700 ;
        RECT 887.400 357.600 888.300 367.950 ;
        RECT 896.550 367.050 897.450 374.550 ;
        RECT 901.950 373.950 904.050 374.550 ;
        RECT 905.400 370.050 906.600 383.400 ;
        RECT 901.950 367.950 904.050 370.050 ;
        RECT 904.950 367.950 907.050 370.050 ;
        RECT 907.950 367.950 910.050 370.050 ;
        RECT 892.950 365.550 897.450 367.050 ;
        RECT 902.100 366.150 903.900 367.950 ;
        RECT 892.950 364.950 897.000 365.550 ;
        RECT 905.400 362.700 906.600 367.950 ;
        RECT 908.100 366.150 909.900 367.950 ;
        RECT 905.400 361.800 909.600 362.700 ;
        RECT 886.800 354.600 888.600 357.600 ;
        RECT 907.800 354.600 909.600 361.800 ;
        RECT 13.800 344.400 15.600 350.400 ;
        RECT 14.400 342.300 15.600 344.400 ;
        RECT 16.800 345.300 18.600 350.400 ;
        RECT 22.800 345.300 24.600 350.400 ;
        RECT 16.800 343.950 24.600 345.300 ;
        RECT 14.400 341.250 18.150 342.300 ;
        RECT 40.200 342.000 42.000 350.400 ;
        RECT 61.800 344.400 63.600 350.400 ;
        RECT 9.000 339.450 13.050 340.050 ;
        RECT 8.550 337.950 13.050 339.450 ;
        RECT 8.550 333.450 9.450 337.950 ;
        RECT 14.100 337.050 15.900 338.850 ;
        RECT 16.950 337.050 18.150 341.250 ;
        RECT 38.700 340.800 42.000 342.000 ;
        RECT 62.400 342.300 63.600 344.400 ;
        RECT 64.800 345.300 66.600 350.400 ;
        RECT 70.800 345.300 72.600 350.400 ;
        RECT 64.800 343.950 72.600 345.300 ;
        RECT 62.400 341.250 66.150 342.300 ;
        RECT 20.100 337.050 21.900 338.850 ;
        RECT 38.700 337.050 39.600 340.800 ;
        RECT 41.100 337.050 42.900 338.850 ;
        RECT 47.100 337.050 48.900 338.850 ;
        RECT 62.100 337.050 63.900 338.850 ;
        RECT 64.950 337.050 66.150 341.250 ;
        RECT 90.000 342.000 91.800 350.400 ;
        RECT 107.400 345.300 109.200 350.400 ;
        RECT 113.400 345.300 115.200 350.400 ;
        RECT 107.400 343.950 115.200 345.300 ;
        RECT 116.400 344.400 118.200 350.400 ;
        RECT 133.800 347.400 135.600 350.400 ;
        RECT 116.400 342.300 117.600 344.400 ;
        RECT 90.000 340.800 93.300 342.000 ;
        RECT 73.950 339.450 78.000 340.050 ;
        RECT 68.100 337.050 69.900 338.850 ;
        RECT 73.950 337.950 78.450 339.450 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 16.950 334.950 19.050 337.050 ;
        RECT 19.950 334.950 22.050 337.050 ;
        RECT 22.950 334.950 25.050 337.050 ;
        RECT 30.000 336.450 34.050 337.050 ;
        RECT 29.550 334.950 34.050 336.450 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 46.950 334.950 49.050 337.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 64.950 334.950 67.050 337.050 ;
        RECT 67.950 334.950 70.050 337.050 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 8.550 332.550 12.450 333.450 ;
        RECT 11.550 331.050 12.450 332.550 ;
        RECT 11.550 330.750 15.000 331.050 ;
        RECT 11.550 329.550 16.050 330.750 ;
        RECT 12.000 328.950 16.050 329.550 ;
        RECT 13.950 328.650 16.050 328.950 ;
        RECT 17.850 321.600 19.050 334.950 ;
        RECT 23.100 333.150 24.900 334.950 ;
        RECT 29.550 334.050 30.450 334.950 ;
        RECT 25.950 332.550 30.450 334.050 ;
        RECT 25.950 331.950 30.000 332.550 ;
        RECT 38.700 322.800 39.600 334.950 ;
        RECT 44.100 333.150 45.900 334.950 ;
        RECT 38.700 321.900 45.300 322.800 ;
        RECT 38.700 321.600 39.600 321.900 ;
        RECT 17.400 315.600 19.200 321.600 ;
        RECT 37.800 315.600 39.600 321.600 ;
        RECT 43.800 321.600 45.300 321.900 ;
        RECT 65.850 321.600 67.050 334.950 ;
        RECT 71.100 333.150 72.900 334.950 ;
        RECT 77.550 334.050 78.450 337.950 ;
        RECT 83.100 337.050 84.900 338.850 ;
        RECT 89.100 337.050 90.900 338.850 ;
        RECT 92.400 337.050 93.300 340.800 ;
        RECT 113.850 341.250 117.600 342.300 ;
        RECT 110.100 337.050 111.900 338.850 ;
        RECT 113.850 337.050 115.050 341.250 ;
        RECT 116.100 337.050 117.900 338.850 ;
        RECT 134.400 337.050 135.600 347.400 ;
        RECT 154.200 342.000 156.000 350.400 ;
        RECT 178.200 344.400 180.000 350.400 ;
        RECT 202.200 344.400 204.000 350.400 ;
        RECT 152.700 340.800 156.000 342.000 ;
        RECT 152.700 337.050 153.600 340.800 ;
        RECT 168.000 339.450 172.050 340.050 ;
        RECT 155.100 337.050 156.900 338.850 ;
        RECT 161.100 337.050 162.900 338.850 ;
        RECT 167.550 337.950 172.050 339.450 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 88.950 334.950 91.050 337.050 ;
        RECT 91.950 334.950 94.050 337.050 ;
        RECT 106.950 334.950 109.050 337.050 ;
        RECT 109.950 334.950 112.050 337.050 ;
        RECT 112.950 334.950 115.050 337.050 ;
        RECT 115.950 334.950 118.050 337.050 ;
        RECT 133.950 334.950 136.050 337.050 ;
        RECT 136.950 334.950 139.050 337.050 ;
        RECT 151.950 334.950 154.050 337.050 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 77.550 332.550 82.050 334.050 ;
        RECT 86.100 333.150 87.900 334.950 ;
        RECT 78.000 331.950 82.050 332.550 ;
        RECT 92.400 322.800 93.300 334.950 ;
        RECT 107.100 333.150 108.900 334.950 ;
        RECT 86.700 321.900 93.300 322.800 ;
        RECT 86.700 321.600 88.200 321.900 ;
        RECT 43.800 315.600 45.600 321.600 ;
        RECT 65.400 315.600 67.200 321.600 ;
        RECT 86.400 315.600 88.200 321.600 ;
        RECT 92.400 321.600 93.300 321.900 ;
        RECT 112.950 321.600 114.150 334.950 ;
        RECT 124.950 333.450 127.050 334.050 ;
        RECT 130.950 333.450 133.050 334.050 ;
        RECT 124.950 332.550 133.050 333.450 ;
        RECT 124.950 331.950 127.050 332.550 ;
        RECT 130.950 331.950 133.050 332.550 ;
        RECT 134.400 321.600 135.600 334.950 ;
        RECT 137.100 333.150 138.900 334.950 ;
        RECT 152.700 322.800 153.600 334.950 ;
        RECT 158.100 333.150 159.900 334.950 ;
        RECT 167.550 333.450 168.450 337.950 ;
        RECT 173.100 337.050 174.900 338.850 ;
        RECT 178.950 337.050 180.000 344.400 ;
        RECT 185.100 337.050 186.900 338.850 ;
        RECT 197.100 337.050 198.900 338.850 ;
        RECT 202.950 337.050 204.000 344.400 ;
        RECT 226.800 343.200 228.600 350.400 ;
        RECT 247.800 347.400 249.600 350.400 ;
        RECT 224.400 342.300 228.600 343.200 ;
        RECT 209.100 337.050 210.900 338.850 ;
        RECT 221.100 337.050 222.900 338.850 ;
        RECT 224.400 337.050 225.600 342.300 ;
        RECT 227.100 337.050 228.900 338.850 ;
        RECT 248.400 337.050 249.300 347.400 ;
        RECT 250.950 345.450 253.050 346.050 ;
        RECT 259.950 345.450 262.050 346.050 ;
        RECT 250.950 344.550 262.050 345.450 ;
        RECT 250.950 343.950 253.050 344.550 ;
        RECT 259.950 343.950 262.050 344.550 ;
        RECT 270.000 344.400 271.800 350.400 ;
        RECT 288.300 346.200 290.100 350.400 ;
        RECT 287.400 344.400 290.100 346.200 ;
        RECT 253.950 339.450 258.000 340.050 ;
        RECT 253.950 337.950 258.450 339.450 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 164.550 332.550 168.450 333.450 ;
        RECT 176.100 333.150 177.900 334.950 ;
        RECT 154.950 330.450 157.050 331.050 ;
        RECT 164.550 330.450 165.450 332.550 ;
        RECT 154.950 329.550 165.450 330.450 ;
        RECT 154.950 328.950 157.050 329.550 ;
        RECT 179.100 329.400 180.000 334.950 ;
        RECT 182.100 333.150 183.900 334.950 ;
        RECT 200.100 333.150 201.900 334.950 ;
        RECT 203.100 329.400 204.000 334.950 ;
        RECT 206.100 333.150 207.900 334.950 ;
        RECT 179.100 328.500 184.200 329.400 ;
        RECT 203.100 328.500 208.200 329.400 ;
        RECT 173.400 326.400 181.200 327.300 ;
        RECT 152.700 321.900 159.300 322.800 ;
        RECT 152.700 321.600 153.600 321.900 ;
        RECT 92.400 315.600 94.200 321.600 ;
        RECT 112.800 315.600 114.600 321.600 ;
        RECT 133.800 315.600 135.600 321.600 ;
        RECT 151.800 315.600 153.600 321.600 ;
        RECT 157.800 321.600 159.300 321.900 ;
        RECT 157.800 315.600 159.600 321.600 ;
        RECT 173.400 315.600 175.200 326.400 ;
        RECT 179.400 316.500 181.200 326.400 ;
        RECT 182.400 317.400 184.200 328.500 ;
        RECT 185.400 316.500 187.200 327.600 ;
        RECT 179.400 315.600 187.200 316.500 ;
        RECT 197.400 326.400 205.200 327.300 ;
        RECT 197.400 315.600 199.200 326.400 ;
        RECT 203.400 316.500 205.200 326.400 ;
        RECT 206.400 317.400 208.200 328.500 ;
        RECT 209.400 316.500 211.200 327.600 ;
        RECT 203.400 315.600 211.200 316.500 ;
        RECT 224.400 321.600 225.600 334.950 ;
        RECT 232.950 333.450 235.050 334.050 ;
        RECT 241.950 333.450 244.050 334.050 ;
        RECT 232.950 332.550 244.050 333.450 ;
        RECT 245.100 333.150 246.900 334.950 ;
        RECT 232.950 331.950 235.050 332.550 ;
        RECT 241.950 331.950 244.050 332.550 ;
        RECT 248.400 327.600 249.300 334.950 ;
        RECT 251.100 333.150 252.900 334.950 ;
        RECT 257.550 334.050 258.450 337.950 ;
        RECT 263.100 337.050 264.900 338.850 ;
        RECT 270.000 337.050 271.050 344.400 ;
        RECT 275.100 337.050 276.900 338.850 ;
        RECT 280.950 337.950 283.050 340.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 265.950 334.950 268.050 337.050 ;
        RECT 268.950 334.950 271.050 337.050 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 257.550 332.550 262.050 334.050 ;
        RECT 266.100 333.150 267.900 334.950 ;
        RECT 258.000 331.950 262.050 332.550 ;
        RECT 270.000 329.400 270.900 334.950 ;
        RECT 272.100 333.150 273.900 334.950 ;
        RECT 281.550 333.450 282.450 337.950 ;
        RECT 287.400 337.050 288.300 344.400 ;
        RECT 290.100 342.600 291.900 343.500 ;
        RECT 295.800 342.600 297.600 350.400 ;
        RECT 290.100 341.700 297.600 342.600 ;
        RECT 311.400 343.200 313.200 350.400 ;
        RECT 334.800 347.400 336.600 350.400 ;
        RECT 311.400 342.300 315.600 343.200 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 289.950 334.950 292.050 337.050 ;
        RECT 278.550 332.550 282.450 333.450 ;
        RECT 265.800 328.500 270.900 329.400 ;
        RECT 271.950 330.450 274.050 331.050 ;
        RECT 278.550 330.450 279.450 332.550 ;
        RECT 283.950 330.450 286.050 331.050 ;
        RECT 271.950 329.550 286.050 330.450 ;
        RECT 271.950 328.950 274.050 329.550 ;
        RECT 283.950 328.950 286.050 329.550 ;
        RECT 245.700 326.400 249.300 327.600 ;
        RECT 224.400 315.600 226.200 321.600 ;
        RECT 245.700 315.600 247.500 326.400 ;
        RECT 262.800 316.500 264.600 327.600 ;
        RECT 265.800 317.400 267.600 328.500 ;
        RECT 287.400 327.600 288.300 334.950 ;
        RECT 290.100 333.150 291.900 334.950 ;
        RECT 268.800 326.400 276.600 327.300 ;
        RECT 268.800 316.500 270.600 326.400 ;
        RECT 262.800 315.600 270.600 316.500 ;
        RECT 274.800 315.600 276.600 326.400 ;
        RECT 286.800 315.600 288.600 327.600 ;
        RECT 293.700 321.600 294.600 341.700 ;
        RECT 306.000 339.450 310.050 340.050 ;
        RECT 296.100 337.050 297.900 338.850 ;
        RECT 305.550 337.950 310.050 339.450 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 305.550 334.050 306.450 337.950 ;
        RECT 311.100 337.050 312.900 338.850 ;
        RECT 314.400 337.050 315.600 342.300 ;
        RECT 325.950 340.950 328.050 343.050 ;
        RECT 317.100 337.050 318.900 338.850 ;
        RECT 310.950 334.950 313.050 337.050 ;
        RECT 313.950 334.950 316.050 337.050 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 305.550 332.550 310.050 334.050 ;
        RECT 306.000 331.950 310.050 332.550 ;
        RECT 295.950 324.450 298.050 325.050 ;
        RECT 310.950 324.450 313.050 325.050 ;
        RECT 295.950 323.550 313.050 324.450 ;
        RECT 295.950 322.950 298.050 323.550 ;
        RECT 310.950 322.950 313.050 323.550 ;
        RECT 314.400 321.600 315.600 334.950 ;
        RECT 326.550 334.050 327.450 340.950 ;
        RECT 335.400 337.050 336.300 347.400 ;
        RECT 353.400 344.400 355.200 350.400 ;
        RECT 372.300 346.200 374.100 350.400 ;
        RECT 371.400 344.400 374.100 346.200 ;
        RECT 350.100 337.050 351.900 338.850 ;
        RECT 353.400 337.050 354.600 344.400 ;
        RECT 358.950 342.450 361.050 343.050 ;
        RECT 367.950 342.450 370.050 343.050 ;
        RECT 358.950 341.550 370.050 342.450 ;
        RECT 358.950 340.950 361.050 341.550 ;
        RECT 367.950 340.950 370.050 341.550 ;
        RECT 355.950 339.450 360.000 340.050 ;
        RECT 355.950 337.950 360.450 339.450 ;
        RECT 331.950 334.950 334.050 337.050 ;
        RECT 334.950 334.950 337.050 337.050 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 326.550 332.550 331.050 334.050 ;
        RECT 332.100 333.150 333.900 334.950 ;
        RECT 327.000 331.950 331.050 332.550 ;
        RECT 335.400 327.600 336.300 334.950 ;
        RECT 338.100 333.150 339.900 334.950 ;
        RECT 292.800 315.600 294.600 321.600 ;
        RECT 313.800 315.600 315.600 321.600 ;
        RECT 332.700 326.400 336.300 327.600 ;
        RECT 353.400 327.600 354.600 334.950 ;
        RECT 359.550 333.450 360.450 337.950 ;
        RECT 371.400 337.050 372.300 344.400 ;
        RECT 374.100 342.600 375.900 343.500 ;
        RECT 379.800 342.600 381.600 350.400 ;
        RECT 374.100 341.700 381.600 342.600 ;
        RECT 394.800 344.400 396.600 350.400 ;
        RECT 400.800 347.400 402.600 350.400 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 364.950 333.450 367.050 333.900 ;
        RECT 359.550 332.550 367.050 333.450 ;
        RECT 364.950 331.800 367.050 332.550 ;
        RECT 371.400 327.600 372.300 334.950 ;
        RECT 374.100 333.150 375.900 334.950 ;
        RECT 332.700 315.600 334.500 326.400 ;
        RECT 353.400 315.600 355.200 327.600 ;
        RECT 370.800 315.600 372.600 327.600 ;
        RECT 377.700 321.600 378.600 341.700 ;
        RECT 380.100 337.050 381.900 338.850 ;
        RECT 394.800 337.050 396.000 344.400 ;
        RECT 401.400 343.500 402.600 347.400 ;
        RECT 396.900 342.600 402.600 343.500 ;
        RECT 415.800 344.400 417.600 350.400 ;
        RECT 421.800 347.400 423.600 350.400 ;
        RECT 396.900 341.700 398.850 342.600 ;
        RECT 379.950 334.950 382.050 337.050 ;
        RECT 394.800 334.950 397.050 337.050 ;
        RECT 376.800 315.600 378.600 321.600 ;
        RECT 394.800 327.600 396.000 334.950 ;
        RECT 397.950 330.300 398.850 341.700 ;
        RECT 403.950 339.450 408.000 340.050 ;
        RECT 403.950 337.950 408.450 339.450 ;
        RECT 400.950 334.950 403.050 337.050 ;
        RECT 401.100 333.150 402.900 334.950 ;
        RECT 407.550 333.900 408.450 337.950 ;
        RECT 415.800 337.050 417.000 344.400 ;
        RECT 422.400 343.500 423.600 347.400 ;
        RECT 417.900 342.600 423.600 343.500 ;
        RECT 437.400 347.400 439.200 350.400 ;
        RECT 457.800 347.400 459.600 350.400 ;
        RECT 417.900 341.700 419.850 342.600 ;
        RECT 415.800 334.950 418.050 337.050 ;
        RECT 406.950 331.800 409.050 333.900 ;
        RECT 396.900 329.400 398.850 330.300 ;
        RECT 396.900 328.500 402.600 329.400 ;
        RECT 394.800 315.600 396.600 327.600 ;
        RECT 401.400 321.600 402.600 328.500 ;
        RECT 400.800 315.600 402.600 321.600 ;
        RECT 415.800 327.600 417.000 334.950 ;
        RECT 418.950 330.300 419.850 341.700 ;
        RECT 437.400 337.050 438.600 347.400 ;
        RECT 458.400 337.050 459.300 347.400 ;
        RECT 470.400 345.300 472.200 350.400 ;
        RECT 476.400 345.300 478.200 350.400 ;
        RECT 470.400 343.950 478.200 345.300 ;
        RECT 479.400 344.400 481.200 350.400 ;
        RECT 496.800 344.400 498.600 350.400 ;
        RECT 502.800 347.400 504.600 350.400 ;
        RECT 479.400 342.300 480.600 344.400 ;
        RECT 476.850 341.250 480.600 342.300 ;
        RECT 473.100 337.050 474.900 338.850 ;
        RECT 476.850 337.050 478.050 341.250 ;
        RECT 479.100 337.050 480.900 338.850 ;
        RECT 496.800 337.050 498.000 344.400 ;
        RECT 503.400 343.500 504.600 347.400 ;
        RECT 498.900 342.600 504.600 343.500 ;
        RECT 517.800 344.400 519.600 350.400 ;
        RECT 523.800 347.400 525.600 350.400 ;
        RECT 538.800 347.400 540.600 350.400 ;
        RECT 498.900 341.700 500.850 342.600 ;
        RECT 421.950 334.950 424.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 436.950 334.950 439.050 337.050 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 460.950 334.950 463.050 337.050 ;
        RECT 469.950 334.950 472.050 337.050 ;
        RECT 472.950 334.950 475.050 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 478.950 334.950 481.050 337.050 ;
        RECT 496.800 334.950 499.050 337.050 ;
        RECT 422.100 333.150 423.900 334.950 ;
        RECT 434.100 333.150 435.900 334.950 ;
        RECT 417.900 329.400 419.850 330.300 ;
        RECT 417.900 328.500 423.600 329.400 ;
        RECT 415.800 315.600 417.600 327.600 ;
        RECT 422.400 321.600 423.600 328.500 ;
        RECT 421.800 315.600 423.600 321.600 ;
        RECT 437.400 321.600 438.600 334.950 ;
        RECT 455.100 333.150 456.900 334.950 ;
        RECT 458.400 327.600 459.300 334.950 ;
        RECT 461.100 333.150 462.900 334.950 ;
        RECT 470.100 333.150 471.900 334.950 ;
        RECT 455.700 326.400 459.300 327.600 ;
        RECT 437.400 315.600 439.200 321.600 ;
        RECT 455.700 315.600 457.500 326.400 ;
        RECT 475.950 321.600 477.150 334.950 ;
        RECT 496.800 327.600 498.000 334.950 ;
        RECT 499.950 330.300 500.850 341.700 ;
        RECT 517.800 337.050 519.000 344.400 ;
        RECT 524.400 343.500 525.600 347.400 ;
        RECT 519.900 342.600 525.600 343.500 ;
        RECT 519.900 341.700 521.850 342.600 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 517.800 334.950 520.050 337.050 ;
        RECT 503.100 333.150 504.900 334.950 ;
        RECT 498.900 329.400 500.850 330.300 ;
        RECT 498.900 328.500 504.600 329.400 ;
        RECT 475.800 315.600 477.600 321.600 ;
        RECT 496.800 315.600 498.600 327.600 ;
        RECT 503.400 321.600 504.600 328.500 ;
        RECT 502.800 315.600 504.600 321.600 ;
        RECT 517.800 327.600 519.000 334.950 ;
        RECT 520.950 330.300 521.850 341.700 ;
        RECT 539.400 337.050 540.600 347.400 ;
        RECT 545.550 344.400 547.350 350.400 ;
        RECT 553.650 347.400 555.450 350.400 ;
        RECT 561.450 347.400 563.250 350.400 ;
        RECT 569.250 348.300 571.050 350.400 ;
        RECT 569.250 347.400 573.000 348.300 ;
        RECT 553.650 346.500 554.700 347.400 ;
        RECT 550.950 345.300 554.700 346.500 ;
        RECT 562.200 346.500 563.250 347.400 ;
        RECT 571.950 346.500 573.000 347.400 ;
        RECT 562.200 345.450 567.150 346.500 ;
        RECT 550.950 344.400 553.050 345.300 ;
        RECT 565.350 344.700 567.150 345.450 ;
        RECT 545.550 337.050 546.750 344.400 ;
        RECT 568.650 343.800 570.450 345.600 ;
        RECT 571.950 344.400 574.050 346.500 ;
        RECT 577.050 344.400 578.850 350.400 ;
        RECT 592.200 344.400 594.000 350.400 ;
        RECT 613.800 344.400 615.600 350.400 ;
        RECT 558.150 342.000 559.950 342.600 ;
        RECT 569.100 342.000 570.150 343.800 ;
        RECT 558.150 340.800 570.150 342.000 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 545.550 335.250 551.850 337.050 ;
        RECT 545.550 334.950 550.050 335.250 ;
        RECT 524.100 333.150 525.900 334.950 ;
        RECT 519.900 329.400 521.850 330.300 ;
        RECT 519.900 328.500 525.600 329.400 ;
        RECT 517.800 315.600 519.600 327.600 ;
        RECT 524.400 321.600 525.600 328.500 ;
        RECT 539.400 321.600 540.600 334.950 ;
        RECT 542.100 333.150 543.900 334.950 ;
        RECT 523.800 315.600 525.600 321.600 ;
        RECT 538.800 315.600 540.600 321.600 ;
        RECT 545.550 327.600 546.750 334.950 ;
        RECT 547.950 329.400 549.750 331.200 ;
        RECT 548.850 328.200 553.050 329.400 ;
        RECT 558.150 328.200 559.050 340.800 ;
        RECT 569.100 339.600 576.000 340.800 ;
        RECT 569.100 339.000 570.900 339.600 ;
        RECT 575.100 338.850 576.000 339.600 ;
        RECT 572.100 337.800 573.900 338.400 ;
        RECT 565.950 336.600 573.900 337.800 ;
        RECT 575.100 337.050 576.900 338.850 ;
        RECT 565.950 334.950 568.050 336.600 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 567.750 329.700 569.550 330.000 ;
        RECT 577.950 329.700 578.850 344.400 ;
        RECT 580.950 337.950 583.050 340.050 ;
        RECT 581.550 333.450 582.450 337.950 ;
        RECT 587.100 337.050 588.900 338.850 ;
        RECT 592.950 337.050 594.000 344.400 ;
        RECT 614.400 342.300 615.600 344.400 ;
        RECT 616.800 345.300 618.600 350.400 ;
        RECT 622.800 345.300 624.600 350.400 ;
        RECT 640.800 347.400 642.600 350.400 ;
        RECT 616.800 343.950 624.600 345.300 ;
        RECT 614.400 341.250 618.150 342.300 ;
        RECT 601.950 339.450 606.000 340.050 ;
        RECT 609.000 339.450 613.050 340.050 ;
        RECT 599.100 337.050 600.900 338.850 ;
        RECT 601.950 337.950 606.450 339.450 ;
        RECT 586.950 334.950 589.050 337.050 ;
        RECT 589.950 334.950 592.050 337.050 ;
        RECT 592.950 334.950 595.050 337.050 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 581.550 332.550 585.450 333.450 ;
        RECT 590.100 333.150 591.900 334.950 ;
        RECT 567.750 329.100 578.850 329.700 ;
        RECT 584.550 330.450 585.450 332.550 ;
        RECT 589.950 330.450 592.050 331.050 ;
        RECT 584.550 329.550 592.050 330.450 ;
        RECT 545.550 315.600 547.350 327.600 ;
        RECT 550.950 327.300 553.050 328.200 ;
        RECT 553.950 327.300 559.050 328.200 ;
        RECT 561.150 328.500 578.850 329.100 ;
        RECT 589.950 328.950 592.050 329.550 ;
        RECT 593.100 329.400 594.000 334.950 ;
        RECT 596.100 333.150 597.900 334.950 ;
        RECT 605.550 334.050 606.450 337.950 ;
        RECT 601.950 332.550 606.450 334.050 ;
        RECT 608.550 337.950 613.050 339.450 ;
        RECT 608.550 334.050 609.450 337.950 ;
        RECT 614.100 337.050 615.900 338.850 ;
        RECT 616.950 337.050 618.150 341.250 ;
        RECT 620.100 337.050 621.900 338.850 ;
        RECT 641.400 337.050 642.300 347.400 ;
        RECT 663.000 344.400 664.800 350.400 ;
        RECT 671.550 344.400 673.350 350.400 ;
        RECT 679.650 347.400 681.450 350.400 ;
        RECT 687.450 347.400 689.250 350.400 ;
        RECT 695.250 348.300 697.050 350.400 ;
        RECT 695.250 347.400 699.000 348.300 ;
        RECT 679.650 346.500 680.700 347.400 ;
        RECT 676.950 345.300 680.700 346.500 ;
        RECT 688.200 346.500 689.250 347.400 ;
        RECT 697.950 346.500 699.000 347.400 ;
        RECT 688.200 345.450 693.150 346.500 ;
        RECT 676.950 344.400 679.050 345.300 ;
        RECT 691.350 344.700 693.150 345.450 ;
        RECT 656.100 337.050 657.900 338.850 ;
        RECT 663.000 337.050 664.050 344.400 ;
        RECT 668.100 337.050 669.900 338.850 ;
        RECT 671.550 337.050 672.750 344.400 ;
        RECT 694.650 343.800 696.450 345.600 ;
        RECT 697.950 344.400 700.050 346.500 ;
        RECT 703.050 344.400 704.850 350.400 ;
        RECT 719.400 347.400 721.200 350.400 ;
        RECT 740.400 347.400 742.200 350.400 ;
        RECT 755.400 347.400 757.200 350.400 ;
        RECT 760.950 348.450 763.050 349.050 ;
        RECT 766.950 348.450 769.050 349.050 ;
        RECT 760.950 347.550 769.050 348.450 ;
        RECT 684.150 342.000 685.950 342.600 ;
        RECT 695.100 342.000 696.150 343.800 ;
        RECT 684.150 340.800 696.150 342.000 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 616.950 334.950 619.050 337.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 637.950 334.950 640.050 337.050 ;
        RECT 640.950 334.950 643.050 337.050 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 655.950 334.950 658.050 337.050 ;
        RECT 658.950 334.950 661.050 337.050 ;
        RECT 661.950 334.950 664.050 337.050 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 671.550 335.250 677.850 337.050 ;
        RECT 671.550 334.950 676.050 335.250 ;
        RECT 608.550 332.550 613.050 334.050 ;
        RECT 601.950 331.950 606.000 332.550 ;
        RECT 609.000 331.950 613.050 332.550 ;
        RECT 593.100 328.500 598.200 329.400 ;
        RECT 561.150 328.200 569.550 328.500 ;
        RECT 553.950 326.400 554.850 327.300 ;
        RECT 552.150 324.600 554.850 326.400 ;
        RECT 555.750 326.100 557.550 326.400 ;
        RECT 561.150 326.100 562.050 328.200 ;
        RECT 577.950 327.600 578.850 328.500 ;
        RECT 555.750 325.200 562.050 326.100 ;
        RECT 562.950 326.700 564.750 327.300 ;
        RECT 562.950 325.500 570.450 326.700 ;
        RECT 555.750 324.600 557.550 325.200 ;
        RECT 569.250 324.600 570.450 325.500 ;
        RECT 550.950 321.600 554.850 323.700 ;
        RECT 559.950 323.550 561.750 324.300 ;
        RECT 564.750 323.550 566.550 324.300 ;
        RECT 559.950 322.500 566.550 323.550 ;
        RECT 569.250 322.500 574.050 324.600 ;
        RECT 553.050 315.600 554.850 321.600 ;
        RECT 560.850 315.600 562.650 322.500 ;
        RECT 569.250 321.600 570.450 322.500 ;
        RECT 568.650 315.600 570.450 321.600 ;
        RECT 577.050 315.600 578.850 327.600 ;
        RECT 587.400 326.400 595.200 327.300 ;
        RECT 587.400 315.600 589.200 326.400 ;
        RECT 593.400 316.500 595.200 326.400 ;
        RECT 596.400 317.400 598.200 328.500 ;
        RECT 599.400 316.500 601.200 327.600 ;
        RECT 617.850 321.600 619.050 334.950 ;
        RECT 623.100 333.150 624.900 334.950 ;
        RECT 638.100 333.150 639.900 334.950 ;
        RECT 641.400 327.600 642.300 334.950 ;
        RECT 644.100 333.150 645.900 334.950 ;
        RECT 659.100 333.150 660.900 334.950 ;
        RECT 663.000 329.400 663.900 334.950 ;
        RECT 665.100 333.150 666.900 334.950 ;
        RECT 658.800 328.500 663.900 329.400 ;
        RECT 638.700 326.400 642.300 327.600 ;
        RECT 593.400 315.600 601.200 316.500 ;
        RECT 617.400 315.600 619.200 321.600 ;
        RECT 638.700 315.600 640.500 326.400 ;
        RECT 655.800 316.500 657.600 327.600 ;
        RECT 658.800 317.400 660.600 328.500 ;
        RECT 671.550 327.600 672.750 334.950 ;
        RECT 673.950 329.400 675.750 331.200 ;
        RECT 674.850 328.200 679.050 329.400 ;
        RECT 684.150 328.200 685.050 340.800 ;
        RECT 695.100 339.600 702.000 340.800 ;
        RECT 695.100 339.000 696.900 339.600 ;
        RECT 701.100 338.850 702.000 339.600 ;
        RECT 698.100 337.800 699.900 338.400 ;
        RECT 691.950 336.600 699.900 337.800 ;
        RECT 701.100 337.050 702.900 338.850 ;
        RECT 691.950 334.950 694.050 336.600 ;
        RECT 700.950 334.950 703.050 337.050 ;
        RECT 693.750 329.700 695.550 330.000 ;
        RECT 703.950 329.700 704.850 344.400 ;
        RECT 719.700 337.050 720.600 347.400 ;
        RECT 727.950 339.450 730.050 340.050 ;
        RECT 733.950 339.450 736.050 340.050 ;
        RECT 727.950 338.550 736.050 339.450 ;
        RECT 727.950 337.950 730.050 338.550 ;
        RECT 733.950 337.950 736.050 338.550 ;
        RECT 740.400 337.050 741.600 347.400 ;
        RECT 755.400 337.050 756.600 347.400 ;
        RECT 760.950 346.950 763.050 347.550 ;
        RECT 766.950 346.950 769.050 347.550 ;
        RECT 775.800 347.400 777.600 350.400 ;
        RECT 757.950 339.450 760.050 340.050 ;
        RECT 757.950 338.550 768.450 339.450 ;
        RECT 757.950 337.950 760.050 338.550 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 754.950 334.950 757.050 337.050 ;
        RECT 716.100 333.150 717.900 334.950 ;
        RECT 693.750 329.100 704.850 329.700 ;
        RECT 661.800 326.400 669.600 327.300 ;
        RECT 661.800 316.500 663.600 326.400 ;
        RECT 655.800 315.600 663.600 316.500 ;
        RECT 667.800 315.600 669.600 326.400 ;
        RECT 671.550 315.600 673.350 327.600 ;
        RECT 676.950 327.300 679.050 328.200 ;
        RECT 679.950 327.300 685.050 328.200 ;
        RECT 687.150 328.500 704.850 329.100 ;
        RECT 687.150 328.200 695.550 328.500 ;
        RECT 679.950 326.400 680.850 327.300 ;
        RECT 678.150 324.600 680.850 326.400 ;
        RECT 681.750 326.100 683.550 326.400 ;
        RECT 687.150 326.100 688.050 328.200 ;
        RECT 703.950 327.600 704.850 328.500 ;
        RECT 681.750 325.200 688.050 326.100 ;
        RECT 688.950 326.700 690.750 327.300 ;
        RECT 688.950 325.500 696.450 326.700 ;
        RECT 681.750 324.600 683.550 325.200 ;
        RECT 695.250 324.600 696.450 325.500 ;
        RECT 676.950 321.600 680.850 323.700 ;
        RECT 685.950 323.550 687.750 324.300 ;
        RECT 690.750 323.550 692.550 324.300 ;
        RECT 685.950 322.500 692.550 323.550 ;
        RECT 695.250 322.500 700.050 324.600 ;
        RECT 679.050 315.600 680.850 321.600 ;
        RECT 686.850 315.600 688.650 322.500 ;
        RECT 695.250 321.600 696.450 322.500 ;
        RECT 694.650 315.600 696.450 321.600 ;
        RECT 703.050 315.600 704.850 327.600 ;
        RECT 719.700 327.600 720.600 334.950 ;
        RECT 722.100 333.150 723.900 334.950 ;
        RECT 737.100 333.150 738.900 334.950 ;
        RECT 719.700 326.400 723.300 327.600 ;
        RECT 721.500 315.600 723.300 326.400 ;
        RECT 740.400 321.600 741.600 334.950 ;
        RECT 752.100 333.150 753.900 334.950 ;
        RECT 755.400 321.600 756.600 334.950 ;
        RECT 767.550 334.050 768.450 338.550 ;
        RECT 776.400 337.050 777.300 347.400 ;
        RECT 796.800 343.200 798.600 350.400 ;
        RECT 794.400 342.300 798.600 343.200 ;
        RECT 791.100 337.050 792.900 338.850 ;
        RECT 794.400 337.050 795.600 342.300 ;
        RECT 819.000 342.000 820.800 350.400 ;
        RECT 833.400 345.300 835.200 350.400 ;
        RECT 839.400 345.300 841.200 350.400 ;
        RECT 833.400 343.950 841.200 345.300 ;
        RECT 842.400 344.400 844.200 350.400 ;
        RECT 859.800 347.400 861.600 350.400 ;
        RECT 842.400 342.300 843.600 344.400 ;
        RECT 819.000 340.800 822.300 342.000 ;
        RECT 797.100 337.050 798.900 338.850 ;
        RECT 812.100 337.050 813.900 338.850 ;
        RECT 818.100 337.050 819.900 338.850 ;
        RECT 821.400 337.050 822.300 340.800 ;
        RECT 839.850 341.250 843.600 342.300 ;
        RECT 836.100 337.050 837.900 338.850 ;
        RECT 839.850 337.050 841.050 341.250 ;
        RECT 842.100 337.050 843.900 338.850 ;
        RECT 860.400 337.050 861.600 347.400 ;
        RECT 878.400 347.400 880.200 350.400 ;
        RECT 878.400 337.050 879.600 347.400 ;
        RECT 890.400 342.600 892.200 350.400 ;
        RECT 897.900 346.200 899.700 350.400 ;
        RECT 897.900 344.400 900.600 346.200 ;
        RECT 896.100 342.600 897.900 343.500 ;
        RECT 890.400 341.700 897.900 342.600 ;
        RECT 890.100 337.050 891.900 338.850 ;
        RECT 772.950 334.950 775.050 337.050 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 814.950 334.950 817.050 337.050 ;
        RECT 817.950 334.950 820.050 337.050 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 859.950 334.950 862.050 337.050 ;
        RECT 862.950 334.950 865.050 337.050 ;
        RECT 874.950 334.950 877.050 337.050 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 889.950 334.950 892.050 337.050 ;
        RECT 767.550 332.550 772.050 334.050 ;
        RECT 773.100 333.150 774.900 334.950 ;
        RECT 768.000 331.950 772.050 332.550 ;
        RECT 776.400 327.600 777.300 334.950 ;
        RECT 779.100 333.150 780.900 334.950 ;
        RECT 773.700 326.400 777.300 327.600 ;
        RECT 740.400 315.600 742.200 321.600 ;
        RECT 755.400 315.600 757.200 321.600 ;
        RECT 773.700 315.600 775.500 326.400 ;
        RECT 794.400 321.600 795.600 334.950 ;
        RECT 815.100 333.150 816.900 334.950 ;
        RECT 799.950 327.450 802.050 328.050 ;
        RECT 811.950 327.450 814.050 328.050 ;
        RECT 799.950 326.550 814.050 327.450 ;
        RECT 799.950 325.950 802.050 326.550 ;
        RECT 811.950 325.950 814.050 326.550 ;
        RECT 821.400 322.800 822.300 334.950 ;
        RECT 833.100 333.150 834.900 334.950 ;
        RECT 815.700 321.900 822.300 322.800 ;
        RECT 815.700 321.600 817.200 321.900 ;
        RECT 794.400 315.600 796.200 321.600 ;
        RECT 815.400 315.600 817.200 321.600 ;
        RECT 821.400 321.600 822.300 321.900 ;
        RECT 838.950 321.600 840.150 334.950 ;
        RECT 860.400 321.600 861.600 334.950 ;
        RECT 863.100 333.150 864.900 334.950 ;
        RECT 875.100 333.150 876.900 334.950 ;
        RECT 821.400 315.600 823.200 321.600 ;
        RECT 838.800 315.600 840.600 321.600 ;
        RECT 859.800 315.600 861.600 321.600 ;
        RECT 878.400 321.600 879.600 334.950 ;
        RECT 893.400 321.600 894.300 341.700 ;
        RECT 899.700 337.050 900.600 344.400 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 896.100 333.150 897.900 334.950 ;
        RECT 899.700 327.600 900.600 334.950 ;
        RECT 878.400 315.600 880.200 321.600 ;
        RECT 893.400 315.600 895.200 321.600 ;
        RECT 899.400 315.600 901.200 327.600 ;
        RECT 13.800 305.400 15.600 311.400 ;
        RECT 14.700 305.100 15.600 305.400 ;
        RECT 19.800 305.400 21.600 311.400 ;
        RECT 19.800 305.100 21.300 305.400 ;
        RECT 14.700 304.200 21.300 305.100 ;
        RECT 14.700 292.050 15.600 304.200 ;
        RECT 34.800 299.400 36.600 311.400 ;
        RECT 37.800 300.300 39.600 311.400 ;
        RECT 43.800 300.300 45.600 311.400 ;
        RECT 37.800 299.400 45.600 300.300 ;
        RECT 55.800 299.400 57.600 311.400 ;
        RECT 58.800 300.300 60.600 311.400 ;
        RECT 64.800 300.300 66.600 311.400 ;
        RECT 77.400 305.400 79.200 311.400 ;
        RECT 77.700 305.100 79.200 305.400 ;
        RECT 83.400 305.400 85.200 311.400 ;
        RECT 101.400 305.400 103.200 311.400 ;
        RECT 83.400 305.100 84.300 305.400 ;
        RECT 77.700 304.200 84.300 305.100 ;
        RECT 101.700 305.100 103.200 305.400 ;
        RECT 107.400 305.400 109.200 311.400 ;
        RECT 125.400 305.400 127.200 311.400 ;
        RECT 107.400 305.100 108.300 305.400 ;
        RECT 101.700 304.200 108.300 305.100 ;
        RECT 58.800 299.400 66.600 300.300 ;
        RECT 20.100 292.050 21.900 293.850 ;
        RECT 35.400 292.050 36.300 299.400 ;
        RECT 41.100 292.050 42.900 293.850 ;
        RECT 56.400 292.050 57.300 299.400 ;
        RECT 62.100 292.050 63.900 293.850 ;
        RECT 77.100 292.050 78.900 293.850 ;
        RECT 83.400 292.050 84.300 304.200 ;
        RECT 94.950 297.450 97.050 298.050 ;
        RECT 100.950 297.450 103.050 298.050 ;
        RECT 94.950 296.550 103.050 297.450 ;
        RECT 94.950 295.950 97.050 296.550 ;
        RECT 100.950 295.950 103.050 296.550 ;
        RECT 101.100 292.050 102.900 293.850 ;
        RECT 107.400 292.050 108.300 304.200 ;
        RECT 125.850 292.050 127.050 305.400 ;
        RECT 145.800 299.400 147.600 311.400 ;
        RECT 148.800 300.300 150.600 311.400 ;
        RECT 154.800 300.300 156.600 311.400 ;
        RECT 170.400 305.400 172.200 311.400 ;
        RECT 194.400 305.400 196.200 311.400 ;
        RECT 214.800 305.400 216.600 311.400 ;
        RECT 148.800 299.400 156.600 300.300 ;
        RECT 130.950 297.450 135.000 298.050 ;
        RECT 130.950 295.950 135.450 297.450 ;
        RECT 134.550 294.450 135.450 295.950 ;
        RECT 131.100 292.050 132.900 293.850 ;
        RECT 134.550 293.550 138.450 294.450 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 22.950 289.950 25.050 292.050 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 43.950 289.950 46.050 292.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 61.950 289.950 64.050 292.050 ;
        RECT 64.950 289.950 67.050 292.050 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 100.950 289.950 103.050 292.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 14.700 286.200 15.600 289.950 ;
        RECT 17.100 288.150 18.900 289.950 ;
        RECT 23.100 288.150 24.900 289.950 ;
        RECT 14.700 285.000 18.000 286.200 ;
        RECT 16.200 276.600 18.000 285.000 ;
        RECT 35.400 282.600 36.300 289.950 ;
        RECT 38.100 288.150 39.900 289.950 ;
        RECT 44.100 288.150 45.900 289.950 ;
        RECT 56.400 282.600 57.300 289.950 ;
        RECT 59.100 288.150 60.900 289.950 ;
        RECT 65.100 288.150 66.900 289.950 ;
        RECT 74.100 288.150 75.900 289.950 ;
        RECT 80.100 288.150 81.900 289.950 ;
        RECT 83.400 286.200 84.300 289.950 ;
        RECT 98.100 288.150 99.900 289.950 ;
        RECT 104.100 288.150 105.900 289.950 ;
        RECT 107.400 286.200 108.300 289.950 ;
        RECT 122.100 288.150 123.900 289.950 ;
        RECT 81.000 285.000 84.300 286.200 ;
        RECT 105.000 285.000 108.300 286.200 ;
        RECT 124.950 285.750 126.150 289.950 ;
        RECT 128.100 288.150 129.900 289.950 ;
        RECT 137.550 289.050 138.450 293.550 ;
        RECT 146.400 292.050 147.300 299.400 ;
        RECT 154.950 297.450 157.050 298.050 ;
        RECT 160.950 297.450 163.050 298.050 ;
        RECT 154.950 296.550 163.050 297.450 ;
        RECT 154.950 295.950 157.050 296.550 ;
        RECT 160.950 295.950 163.050 296.550 ;
        RECT 152.100 292.050 153.900 293.850 ;
        RECT 170.850 292.050 172.050 305.400 ;
        RECT 176.100 292.050 177.900 293.850 ;
        RECT 194.850 292.050 196.050 305.400 ;
        RECT 200.100 292.050 201.900 293.850 ;
        RECT 215.400 292.050 216.600 305.400 ;
        RECT 233.400 305.400 235.200 311.400 ;
        RECT 251.400 305.400 253.200 311.400 ;
        RECT 271.800 305.400 273.600 311.400 ;
        RECT 293.400 305.400 295.200 311.400 ;
        RECT 233.400 292.050 234.600 305.400 ;
        RECT 235.950 303.450 238.050 304.050 ;
        RECT 247.950 303.450 250.050 304.050 ;
        RECT 235.950 302.550 250.050 303.450 ;
        RECT 235.950 301.950 238.050 302.550 ;
        RECT 247.950 301.950 250.050 302.550 ;
        RECT 251.400 292.050 252.600 305.400 ;
        RECT 261.000 294.450 265.050 295.050 ;
        RECT 260.550 292.950 265.050 294.450 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 166.950 289.950 169.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 199.950 289.950 202.050 292.050 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 250.950 289.950 253.050 292.050 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 133.950 287.550 138.450 289.050 ;
        RECT 133.950 286.950 138.000 287.550 ;
        RECT 35.400 281.400 40.500 282.600 ;
        RECT 56.400 281.400 61.500 282.600 ;
        RECT 38.700 276.600 40.500 281.400 ;
        RECT 59.700 276.600 61.500 281.400 ;
        RECT 81.000 276.600 82.800 285.000 ;
        RECT 105.000 276.600 106.800 285.000 ;
        RECT 122.400 284.700 126.150 285.750 ;
        RECT 122.400 282.600 123.600 284.700 ;
        RECT 121.800 276.600 123.600 282.600 ;
        RECT 124.800 281.700 132.600 283.050 ;
        RECT 124.800 276.600 126.600 281.700 ;
        RECT 130.800 276.600 132.600 281.700 ;
        RECT 146.400 282.600 147.300 289.950 ;
        RECT 149.100 288.150 150.900 289.950 ;
        RECT 155.100 288.150 156.900 289.950 ;
        RECT 167.100 288.150 168.900 289.950 ;
        RECT 169.950 285.750 171.150 289.950 ;
        RECT 173.100 288.150 174.900 289.950 ;
        RECT 191.100 288.150 192.900 289.950 ;
        RECT 193.950 285.750 195.150 289.950 ;
        RECT 197.100 288.150 198.900 289.950 ;
        RECT 212.100 288.150 213.900 289.950 ;
        RECT 167.400 284.700 171.150 285.750 ;
        RECT 191.400 284.700 195.150 285.750 ;
        RECT 215.400 284.700 216.600 289.950 ;
        RECT 218.100 288.150 219.900 289.950 ;
        RECT 230.100 288.150 231.900 289.950 ;
        RECT 167.400 282.600 168.600 284.700 ;
        RECT 146.400 281.400 151.500 282.600 ;
        RECT 149.700 276.600 151.500 281.400 ;
        RECT 166.800 276.600 168.600 282.600 ;
        RECT 169.800 281.700 177.600 283.050 ;
        RECT 191.400 282.600 192.600 284.700 ;
        RECT 212.400 283.800 216.600 284.700 ;
        RECT 233.400 284.700 234.600 289.950 ;
        RECT 236.100 288.150 237.900 289.950 ;
        RECT 248.100 288.150 249.900 289.950 ;
        RECT 251.400 284.700 252.600 289.950 ;
        RECT 254.100 288.150 255.900 289.950 ;
        RECT 260.550 289.050 261.450 292.950 ;
        RECT 266.100 292.050 267.900 293.850 ;
        RECT 271.950 292.050 273.150 305.400 ;
        RECT 274.950 297.450 277.050 298.050 ;
        RECT 289.950 297.450 292.050 298.050 ;
        RECT 274.950 296.550 292.050 297.450 ;
        RECT 274.950 295.950 277.050 296.550 ;
        RECT 289.950 295.950 292.050 296.550 ;
        RECT 293.400 292.050 294.600 305.400 ;
        RECT 313.800 299.400 315.600 311.400 ;
        RECT 319.800 305.400 321.600 311.400 ;
        RECT 298.950 294.450 303.000 295.050 ;
        RECT 298.950 292.950 303.450 294.450 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 268.950 289.950 271.050 292.050 ;
        RECT 271.950 289.950 274.050 292.050 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 256.950 287.550 261.450 289.050 ;
        RECT 269.100 288.150 270.900 289.950 ;
        RECT 256.950 286.950 261.000 287.550 ;
        RECT 272.850 285.750 274.050 289.950 ;
        RECT 275.100 288.150 276.900 289.950 ;
        RECT 290.100 288.150 291.900 289.950 ;
        RECT 272.850 284.700 276.600 285.750 ;
        RECT 233.400 283.800 237.600 284.700 ;
        RECT 251.400 283.800 255.600 284.700 ;
        RECT 169.800 276.600 171.600 281.700 ;
        RECT 175.800 276.600 177.600 281.700 ;
        RECT 190.800 276.600 192.600 282.600 ;
        RECT 193.800 281.700 201.600 283.050 ;
        RECT 193.800 276.600 195.600 281.700 ;
        RECT 199.800 276.600 201.600 281.700 ;
        RECT 212.400 276.600 214.200 283.800 ;
        RECT 235.800 276.600 237.600 283.800 ;
        RECT 253.800 276.600 255.600 283.800 ;
        RECT 266.400 281.700 274.200 283.050 ;
        RECT 266.400 276.600 268.200 281.700 ;
        RECT 272.400 276.600 274.200 281.700 ;
        RECT 275.400 282.600 276.600 284.700 ;
        RECT 293.400 284.700 294.600 289.950 ;
        RECT 296.100 288.150 297.900 289.950 ;
        RECT 302.550 289.050 303.450 292.950 ;
        RECT 314.400 292.050 315.300 299.400 ;
        RECT 317.100 292.050 318.900 293.850 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 298.950 287.550 303.450 289.050 ;
        RECT 298.950 286.950 303.000 287.550 ;
        RECT 293.400 283.800 297.600 284.700 ;
        RECT 275.400 276.600 277.200 282.600 ;
        RECT 295.800 276.600 297.600 283.800 ;
        RECT 314.400 282.600 315.300 289.950 ;
        RECT 320.700 285.300 321.600 305.400 ;
        RECT 338.400 305.400 340.200 311.400 ;
        RECT 358.800 305.400 360.600 311.400 ;
        RECT 338.400 292.050 339.600 305.400 ;
        RECT 359.700 305.100 360.600 305.400 ;
        RECT 364.800 305.400 366.600 311.400 ;
        RECT 383.400 305.400 385.200 311.400 ;
        RECT 403.800 305.400 405.600 311.400 ;
        RECT 425.400 305.400 427.200 311.400 ;
        RECT 442.800 305.400 444.600 311.400 ;
        RECT 463.800 305.400 465.600 311.400 ;
        RECT 485.400 305.400 487.200 311.400 ;
        RECT 508.800 305.400 510.600 311.400 ;
        RECT 364.800 305.100 366.300 305.400 ;
        RECT 359.700 304.200 366.300 305.100 ;
        RECT 340.950 297.450 343.050 298.050 ;
        RECT 349.950 297.450 352.050 298.050 ;
        RECT 340.950 296.550 352.050 297.450 ;
        RECT 340.950 295.950 343.050 296.550 ;
        RECT 349.950 295.950 352.050 296.550 ;
        RECT 359.700 292.050 360.600 304.200 ;
        RECT 370.950 300.450 373.050 301.050 ;
        RECT 376.950 300.450 379.050 301.050 ;
        RECT 370.950 299.550 379.050 300.450 ;
        RECT 370.950 298.950 373.050 299.550 ;
        RECT 376.950 298.950 379.050 299.550 ;
        RECT 364.950 297.450 367.050 298.050 ;
        RECT 376.950 297.450 379.050 297.900 ;
        RECT 364.950 296.550 379.050 297.450 ;
        RECT 364.950 295.950 367.050 296.550 ;
        RECT 376.950 295.800 379.050 296.550 ;
        RECT 365.100 292.050 366.900 293.850 ;
        RECT 383.400 292.050 384.600 305.400 ;
        RECT 404.400 292.050 405.600 305.400 ;
        RECT 409.950 294.450 414.000 295.050 ;
        RECT 417.000 294.450 421.050 295.050 ;
        RECT 409.950 292.950 414.450 294.450 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 361.950 289.950 364.050 292.050 ;
        RECT 364.950 289.950 367.050 292.050 ;
        RECT 367.950 289.950 370.050 292.050 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 385.950 289.950 388.050 292.050 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 406.950 289.950 409.050 292.050 ;
        RECT 323.100 288.150 324.900 289.950 ;
        RECT 335.100 288.150 336.900 289.950 ;
        RECT 317.100 284.400 324.600 285.300 ;
        RECT 317.100 283.500 318.900 284.400 ;
        RECT 314.400 280.800 317.100 282.600 ;
        RECT 315.300 276.600 317.100 280.800 ;
        RECT 322.800 276.600 324.600 284.400 ;
        RECT 338.400 284.700 339.600 289.950 ;
        RECT 341.100 288.150 342.900 289.950 ;
        RECT 359.700 286.200 360.600 289.950 ;
        RECT 362.100 288.150 363.900 289.950 ;
        RECT 368.100 288.150 369.900 289.950 ;
        RECT 380.100 288.150 381.900 289.950 ;
        RECT 359.700 285.000 363.000 286.200 ;
        RECT 338.400 283.800 342.600 284.700 ;
        RECT 340.800 276.600 342.600 283.800 ;
        RECT 361.200 276.600 363.000 285.000 ;
        RECT 383.400 284.700 384.600 289.950 ;
        RECT 386.100 288.150 387.900 289.950 ;
        RECT 401.100 288.150 402.900 289.950 ;
        RECT 404.400 284.700 405.600 289.950 ;
        RECT 407.100 288.150 408.900 289.950 ;
        RECT 383.400 283.800 387.600 284.700 ;
        RECT 385.800 276.600 387.600 283.800 ;
        RECT 401.400 283.800 405.600 284.700 ;
        RECT 413.550 286.050 414.450 292.950 ;
        RECT 416.550 292.950 421.050 294.450 ;
        RECT 416.550 289.050 417.450 292.950 ;
        RECT 425.850 292.050 427.050 305.400 ;
        RECT 431.100 292.050 432.900 293.850 ;
        RECT 443.400 292.050 444.600 305.400 ;
        RECT 446.100 292.050 447.900 293.850 ;
        RECT 458.100 292.050 459.900 293.850 ;
        RECT 463.950 292.050 465.150 305.400 ;
        RECT 485.400 292.050 486.600 305.400 ;
        RECT 509.400 292.050 510.600 305.400 ;
        RECT 526.800 310.500 534.600 311.400 ;
        RECT 511.950 300.450 514.050 301.050 ;
        RECT 517.950 300.450 520.050 301.050 ;
        RECT 511.950 299.550 520.050 300.450 ;
        RECT 511.950 298.950 514.050 299.550 ;
        RECT 517.950 298.950 520.050 299.550 ;
        RECT 526.800 299.400 528.600 310.500 ;
        RECT 529.800 298.500 531.600 309.600 ;
        RECT 532.800 300.600 534.600 310.500 ;
        RECT 538.800 300.600 540.600 311.400 ;
        RECT 553.800 305.400 555.600 311.400 ;
        RECT 572.400 305.400 574.200 311.400 ;
        RECT 595.800 305.400 597.600 311.400 ;
        RECT 532.800 299.700 540.600 300.600 ;
        RECT 529.800 297.600 534.900 298.500 ;
        RECT 530.100 292.050 531.900 293.850 ;
        RECT 534.000 292.050 534.900 297.600 ;
        RECT 536.100 292.050 537.900 293.850 ;
        RECT 554.400 292.050 555.600 305.400 ;
        RECT 557.100 292.050 558.900 293.850 ;
        RECT 572.850 292.050 574.050 305.400 ;
        RECT 578.100 292.050 579.900 293.850 ;
        RECT 596.400 292.050 597.600 305.400 ;
        RECT 613.800 299.400 615.600 311.400 ;
        RECT 616.800 300.300 618.600 311.400 ;
        RECT 622.800 300.300 624.600 311.400 ;
        RECT 638.400 305.400 640.200 311.400 ;
        RECT 661.800 305.400 663.600 311.400 ;
        RECT 683.400 305.400 685.200 311.400 ;
        RECT 703.800 305.400 705.600 311.400 ;
        RECT 616.800 299.400 624.600 300.300 ;
        RECT 614.400 292.050 615.300 299.400 ;
        RECT 620.100 292.050 621.900 293.850 ;
        RECT 638.850 292.050 640.050 305.400 ;
        RECT 646.950 294.450 651.000 295.050 ;
        RECT 644.100 292.050 645.900 293.850 ;
        RECT 646.950 292.950 651.450 294.450 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 427.950 289.950 430.050 292.050 ;
        RECT 430.950 289.950 433.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 457.950 289.950 460.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 508.950 289.950 511.050 292.050 ;
        RECT 511.950 289.950 514.050 292.050 ;
        RECT 526.950 289.950 529.050 292.050 ;
        RECT 529.950 289.950 532.050 292.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 535.950 289.950 538.050 292.050 ;
        RECT 538.950 289.950 541.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 556.950 289.950 559.050 292.050 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 577.950 289.950 580.050 292.050 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 598.950 289.950 601.050 292.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 616.950 289.950 619.050 292.050 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 622.950 289.950 625.050 292.050 ;
        RECT 634.950 289.950 637.050 292.050 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 416.550 287.550 421.050 289.050 ;
        RECT 422.100 288.150 423.900 289.950 ;
        RECT 417.000 286.950 421.050 287.550 ;
        RECT 413.550 284.550 418.050 286.050 ;
        RECT 424.950 285.750 426.150 289.950 ;
        RECT 428.100 288.150 429.900 289.950 ;
        RECT 414.000 283.950 418.050 284.550 ;
        RECT 422.400 284.700 426.150 285.750 ;
        RECT 401.400 276.600 403.200 283.800 ;
        RECT 422.400 282.600 423.600 284.700 ;
        RECT 421.800 276.600 423.600 282.600 ;
        RECT 424.800 281.700 432.600 283.050 ;
        RECT 424.800 276.600 426.600 281.700 ;
        RECT 430.800 276.600 432.600 281.700 ;
        RECT 443.400 279.600 444.600 289.950 ;
        RECT 461.100 288.150 462.900 289.950 ;
        RECT 454.950 285.450 457.050 286.050 ;
        RECT 446.550 285.000 457.050 285.450 ;
        RECT 445.950 284.550 457.050 285.000 ;
        RECT 464.850 285.750 466.050 289.950 ;
        RECT 467.100 288.150 468.900 289.950 ;
        RECT 482.100 288.150 483.900 289.950 ;
        RECT 464.850 284.700 468.600 285.750 ;
        RECT 445.950 280.950 448.050 284.550 ;
        RECT 454.950 283.950 457.050 284.550 ;
        RECT 458.400 281.700 466.200 283.050 ;
        RECT 442.800 276.600 444.600 279.600 ;
        RECT 458.400 276.600 460.200 281.700 ;
        RECT 464.400 276.600 466.200 281.700 ;
        RECT 467.400 282.600 468.600 284.700 ;
        RECT 485.400 284.700 486.600 289.950 ;
        RECT 488.100 288.150 489.900 289.950 ;
        RECT 506.100 288.150 507.900 289.950 ;
        RECT 509.400 284.700 510.600 289.950 ;
        RECT 512.100 288.150 513.900 289.950 ;
        RECT 527.100 288.150 528.900 289.950 ;
        RECT 485.400 283.800 489.600 284.700 ;
        RECT 467.400 276.600 469.200 282.600 ;
        RECT 487.800 276.600 489.600 283.800 ;
        RECT 506.400 283.800 510.600 284.700 ;
        RECT 506.400 276.600 508.200 283.800 ;
        RECT 534.000 282.600 535.050 289.950 ;
        RECT 539.100 288.150 540.900 289.950 ;
        RECT 534.000 276.600 535.800 282.600 ;
        RECT 554.400 279.600 555.600 289.950 ;
        RECT 569.100 288.150 570.900 289.950 ;
        RECT 571.950 285.750 573.150 289.950 ;
        RECT 575.100 288.150 576.900 289.950 ;
        RECT 593.100 288.150 594.900 289.950 ;
        RECT 569.400 284.700 573.150 285.750 ;
        RECT 596.400 284.700 597.600 289.950 ;
        RECT 599.100 288.150 600.900 289.950 ;
        RECT 569.400 282.600 570.600 284.700 ;
        RECT 593.400 283.800 597.600 284.700 ;
        RECT 553.800 276.600 555.600 279.600 ;
        RECT 568.800 276.600 570.600 282.600 ;
        RECT 571.800 281.700 579.600 283.050 ;
        RECT 571.800 276.600 573.600 281.700 ;
        RECT 577.800 276.600 579.600 281.700 ;
        RECT 593.400 276.600 595.200 283.800 ;
        RECT 614.400 282.600 615.300 289.950 ;
        RECT 617.100 288.150 618.900 289.950 ;
        RECT 623.100 288.150 624.900 289.950 ;
        RECT 635.100 288.150 636.900 289.950 ;
        RECT 637.950 285.750 639.150 289.950 ;
        RECT 641.100 288.150 642.900 289.950 ;
        RECT 650.550 288.900 651.450 292.950 ;
        RECT 656.100 292.050 657.900 293.850 ;
        RECT 661.950 292.050 663.150 305.400 ;
        RECT 670.950 303.450 673.050 304.050 ;
        RECT 679.950 303.450 682.050 304.050 ;
        RECT 670.950 302.550 682.050 303.450 ;
        RECT 670.950 301.950 673.050 302.550 ;
        RECT 679.950 301.950 682.050 302.550 ;
        RECT 683.400 292.050 684.600 305.400 ;
        RECT 685.950 297.450 688.050 298.050 ;
        RECT 685.950 296.550 693.450 297.450 ;
        RECT 685.950 295.950 688.050 296.550 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 649.950 286.800 652.050 288.900 ;
        RECT 659.100 288.150 660.900 289.950 ;
        RECT 635.400 284.700 639.150 285.750 ;
        RECT 662.850 285.750 664.050 289.950 ;
        RECT 665.100 288.150 666.900 289.950 ;
        RECT 680.100 288.150 681.900 289.950 ;
        RECT 662.850 284.700 666.600 285.750 ;
        RECT 635.400 282.600 636.600 284.700 ;
        RECT 614.400 281.400 619.500 282.600 ;
        RECT 617.700 276.600 619.500 281.400 ;
        RECT 634.800 276.600 636.600 282.600 ;
        RECT 637.800 281.700 645.600 283.050 ;
        RECT 637.800 276.600 639.600 281.700 ;
        RECT 643.800 276.600 645.600 281.700 ;
        RECT 656.400 281.700 664.200 283.050 ;
        RECT 656.400 276.600 658.200 281.700 ;
        RECT 662.400 276.600 664.200 281.700 ;
        RECT 665.400 282.600 666.600 284.700 ;
        RECT 673.950 285.450 676.050 286.050 ;
        RECT 679.950 285.450 682.050 286.050 ;
        RECT 673.950 284.550 682.050 285.450 ;
        RECT 673.950 283.950 676.050 284.550 ;
        RECT 679.950 283.950 682.050 284.550 ;
        RECT 683.400 284.700 684.600 289.950 ;
        RECT 686.100 288.150 687.900 289.950 ;
        RECT 692.550 289.050 693.450 296.550 ;
        RECT 704.400 292.050 705.600 305.400 ;
        RECT 722.400 305.400 724.200 311.400 ;
        RECT 707.100 292.050 708.900 293.850 ;
        RECT 722.400 292.050 723.600 305.400 ;
        RECT 743.400 299.400 745.200 311.400 ;
        RECT 763.800 305.400 765.600 311.400 ;
        RECT 743.700 292.050 744.750 299.400 ;
        RECT 764.400 292.050 765.600 305.400 ;
        RECT 779.400 305.400 781.200 311.400 ;
        RECT 767.100 292.050 768.900 293.850 ;
        RECT 776.100 292.050 777.900 293.850 ;
        RECT 779.400 292.050 780.600 305.400 ;
        RECT 794.400 300.300 796.200 311.400 ;
        RECT 800.400 300.300 802.200 311.400 ;
        RECT 794.400 299.400 802.200 300.300 ;
        RECT 803.400 299.400 805.200 311.400 ;
        RECT 818.400 300.600 820.200 311.400 ;
        RECT 824.400 310.500 832.200 311.400 ;
        RECT 824.400 300.600 826.200 310.500 ;
        RECT 818.400 299.700 826.200 300.600 ;
        RECT 796.950 297.450 799.050 298.050 ;
        RECT 791.550 296.550 799.050 297.450 ;
        RECT 791.550 294.450 792.450 296.550 ;
        RECT 796.950 295.950 799.050 296.550 ;
        RECT 788.550 293.550 792.450 294.450 ;
        RECT 703.950 289.950 706.050 292.050 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 743.700 289.950 748.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 775.950 289.950 778.050 292.050 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 688.950 287.550 693.450 289.050 ;
        RECT 688.950 286.950 693.000 287.550 ;
        RECT 683.400 283.800 687.600 284.700 ;
        RECT 665.400 276.600 667.200 282.600 ;
        RECT 685.800 276.600 687.600 283.800 ;
        RECT 704.400 279.600 705.600 289.950 ;
        RECT 719.100 288.150 720.900 289.950 ;
        RECT 722.400 284.700 723.600 289.950 ;
        RECT 725.100 288.150 726.900 289.950 ;
        RECT 740.100 288.150 741.900 289.950 ;
        RECT 722.400 283.800 726.600 284.700 ;
        RECT 703.800 276.600 705.600 279.600 ;
        RECT 724.800 276.600 726.600 283.800 ;
        RECT 743.700 282.600 744.750 289.950 ;
        RECT 743.400 276.600 745.200 282.600 ;
        RECT 764.400 279.600 765.600 289.950 ;
        RECT 763.800 276.600 765.600 279.600 ;
        RECT 779.400 279.600 780.600 289.950 ;
        RECT 788.550 285.450 789.450 293.550 ;
        RECT 797.100 292.050 798.900 293.850 ;
        RECT 803.700 292.050 804.600 299.400 ;
        RECT 827.400 298.500 829.200 309.600 ;
        RECT 830.400 299.400 832.200 310.500 ;
        RECT 850.800 305.400 852.600 311.400 ;
        RECT 872.400 305.400 874.200 311.400 ;
        RECT 895.800 305.400 897.600 311.400 ;
        RECT 824.100 297.600 829.200 298.500 ;
        RECT 805.950 294.450 810.000 295.050 ;
        RECT 805.950 292.950 810.450 294.450 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 796.950 289.950 799.050 292.050 ;
        RECT 799.950 289.950 802.050 292.050 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 794.100 288.150 795.900 289.950 ;
        RECT 800.100 288.150 801.900 289.950 ;
        RECT 796.950 285.450 799.050 286.050 ;
        RECT 788.550 284.550 799.050 285.450 ;
        RECT 796.950 283.950 799.050 284.550 ;
        RECT 803.700 282.600 804.600 289.950 ;
        RECT 809.550 289.050 810.450 292.950 ;
        RECT 821.100 292.050 822.900 293.850 ;
        RECT 824.100 292.050 825.000 297.600 ;
        RECT 832.950 297.450 835.050 298.050 ;
        RECT 844.950 297.450 847.050 298.050 ;
        RECT 832.950 296.550 847.050 297.450 ;
        RECT 832.950 295.950 835.050 296.550 ;
        RECT 844.950 295.950 847.050 296.550 ;
        RECT 840.000 294.450 844.050 295.050 ;
        RECT 827.100 292.050 828.900 293.850 ;
        RECT 839.550 292.950 844.050 294.450 ;
        RECT 817.950 289.950 820.050 292.050 ;
        RECT 820.950 289.950 823.050 292.050 ;
        RECT 823.950 289.950 826.050 292.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 805.950 287.550 810.450 289.050 ;
        RECT 818.100 288.150 819.900 289.950 ;
        RECT 805.950 286.950 810.000 287.550 ;
        RECT 823.950 282.600 825.000 289.950 ;
        RECT 830.100 288.150 831.900 289.950 ;
        RECT 839.550 288.450 840.450 292.950 ;
        RECT 845.100 292.050 846.900 293.850 ;
        RECT 850.950 292.050 852.150 305.400 ;
        RECT 853.950 300.450 856.050 301.050 ;
        RECT 865.950 300.450 868.050 300.900 ;
        RECT 853.950 299.550 868.050 300.450 ;
        RECT 853.950 298.950 856.050 299.550 ;
        RECT 865.950 298.800 868.050 299.550 ;
        RECT 853.950 297.450 856.050 297.900 ;
        RECT 862.950 297.450 865.050 298.050 ;
        RECT 853.950 296.550 865.050 297.450 ;
        RECT 853.950 295.800 856.050 296.550 ;
        RECT 862.950 295.950 865.050 296.550 ;
        RECT 872.400 292.050 873.600 305.400 ;
        RECT 877.950 294.450 880.050 295.050 ;
        RECT 877.950 293.550 885.450 294.450 ;
        RECT 877.950 292.950 880.050 293.550 ;
        RECT 844.950 289.950 847.050 292.050 ;
        RECT 847.950 289.950 850.050 292.050 ;
        RECT 850.950 289.950 853.050 292.050 ;
        RECT 853.950 289.950 856.050 292.050 ;
        RECT 868.950 289.950 871.050 292.050 ;
        RECT 871.950 289.950 874.050 292.050 ;
        RECT 874.950 289.950 877.050 292.050 ;
        RECT 839.550 288.000 843.450 288.450 ;
        RECT 848.100 288.150 849.900 289.950 ;
        RECT 839.550 287.550 844.050 288.000 ;
        RECT 841.950 283.950 844.050 287.550 ;
        RECT 851.850 285.750 853.050 289.950 ;
        RECT 854.100 288.150 855.900 289.950 ;
        RECT 869.100 288.150 870.900 289.950 ;
        RECT 851.850 284.700 855.600 285.750 ;
        RECT 799.500 281.400 804.600 282.600 ;
        RECT 779.400 276.600 781.200 279.600 ;
        RECT 799.500 276.600 801.300 281.400 ;
        RECT 823.200 276.600 825.000 282.600 ;
        RECT 845.400 281.700 853.200 283.050 ;
        RECT 845.400 276.600 847.200 281.700 ;
        RECT 851.400 276.600 853.200 281.700 ;
        RECT 854.400 282.600 855.600 284.700 ;
        RECT 856.950 285.450 859.050 286.050 ;
        RECT 865.950 285.450 868.050 286.050 ;
        RECT 856.950 284.550 868.050 285.450 ;
        RECT 856.950 283.950 859.050 284.550 ;
        RECT 865.950 283.950 868.050 284.550 ;
        RECT 872.400 284.700 873.600 289.950 ;
        RECT 875.100 288.150 876.900 289.950 ;
        RECT 884.550 289.050 885.450 293.550 ;
        RECT 890.100 292.050 891.900 293.850 ;
        RECT 895.950 292.050 897.150 305.400 ;
        RECT 889.950 289.950 892.050 292.050 ;
        RECT 892.950 289.950 895.050 292.050 ;
        RECT 895.950 289.950 898.050 292.050 ;
        RECT 898.950 289.950 901.050 292.050 ;
        RECT 884.550 287.550 889.050 289.050 ;
        RECT 893.100 288.150 894.900 289.950 ;
        RECT 885.000 286.950 889.050 287.550 ;
        RECT 896.850 285.750 898.050 289.950 ;
        RECT 899.100 288.150 900.900 289.950 ;
        RECT 896.850 284.700 900.600 285.750 ;
        RECT 872.400 283.800 876.600 284.700 ;
        RECT 854.400 276.600 856.200 282.600 ;
        RECT 874.800 276.600 876.600 283.800 ;
        RECT 890.400 281.700 898.200 283.050 ;
        RECT 890.400 276.600 892.200 281.700 ;
        RECT 896.400 276.600 898.200 281.700 ;
        RECT 899.400 282.600 900.600 284.700 ;
        RECT 899.400 276.600 901.200 282.600 ;
        RECT 13.800 266.400 15.600 272.400 ;
        RECT 14.400 264.300 15.600 266.400 ;
        RECT 16.800 267.300 18.600 272.400 ;
        RECT 22.800 267.300 24.600 272.400 ;
        RECT 16.800 265.950 24.600 267.300 ;
        RECT 34.800 266.400 36.600 272.400 ;
        RECT 35.400 264.300 36.600 266.400 ;
        RECT 37.800 267.300 39.600 272.400 ;
        RECT 43.800 267.300 45.600 272.400 ;
        RECT 37.800 265.950 45.600 267.300 ;
        RECT 14.400 263.250 18.150 264.300 ;
        RECT 35.400 263.250 39.150 264.300 ;
        RECT 61.200 264.000 63.000 272.400 ;
        RECT 82.800 269.400 84.600 272.400 ;
        RECT 14.100 259.050 15.900 260.850 ;
        RECT 16.950 259.050 18.150 263.250 ;
        RECT 25.950 261.450 30.000 262.050 ;
        RECT 20.100 259.050 21.900 260.850 ;
        RECT 25.950 259.950 30.450 261.450 ;
        RECT 13.950 256.950 16.050 259.050 ;
        RECT 16.950 256.950 19.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 22.950 256.950 25.050 259.050 ;
        RECT 17.850 243.600 19.050 256.950 ;
        RECT 23.100 255.150 24.900 256.950 ;
        RECT 29.550 256.050 30.450 259.950 ;
        RECT 35.100 259.050 36.900 260.850 ;
        RECT 37.950 259.050 39.150 263.250 ;
        RECT 59.700 262.800 63.000 264.000 ;
        RECT 49.950 261.450 52.050 262.050 ;
        RECT 55.950 261.450 58.050 262.050 ;
        RECT 41.100 259.050 42.900 260.850 ;
        RECT 49.950 260.550 58.050 261.450 ;
        RECT 49.950 259.950 52.050 260.550 ;
        RECT 55.950 259.950 58.050 260.550 ;
        RECT 59.700 259.050 60.600 262.800 ;
        RECT 62.100 259.050 63.900 260.850 ;
        RECT 68.100 259.050 69.900 260.850 ;
        RECT 83.400 259.050 84.600 269.400 ;
        RECT 105.000 266.400 106.800 272.400 ;
        RECT 98.100 259.050 99.900 260.850 ;
        RECT 105.000 259.050 106.050 266.400 ;
        RECT 124.800 265.200 126.600 272.400 ;
        RECT 122.400 264.300 126.600 265.200 ;
        RECT 110.100 259.050 111.900 260.850 ;
        RECT 119.100 259.050 120.900 260.850 ;
        RECT 122.400 259.050 123.600 264.300 ;
        RECT 145.200 264.000 147.000 272.400 ;
        RECT 143.700 262.800 147.000 264.000 ;
        RECT 164.400 269.400 166.200 272.400 ;
        RECT 125.100 259.050 126.900 260.850 ;
        RECT 143.700 259.050 144.600 262.800 ;
        RECT 146.100 259.050 147.900 260.850 ;
        RECT 152.100 259.050 153.900 260.850 ;
        RECT 164.400 259.050 165.600 269.400 ;
        RECT 184.200 264.000 186.000 272.400 ;
        RECT 205.800 269.400 207.600 272.400 ;
        RECT 182.700 262.800 186.000 264.000 ;
        RECT 182.700 259.050 183.600 262.800 ;
        RECT 185.100 259.050 186.900 260.850 ;
        RECT 191.100 259.050 192.900 260.850 ;
        RECT 206.400 259.050 207.600 269.400 ;
        RECT 226.200 264.000 228.000 272.400 ;
        RECT 241.950 265.950 244.050 268.050 ;
        RECT 224.700 262.800 228.000 264.000 ;
        RECT 224.700 259.050 225.600 262.800 ;
        RECT 227.100 259.050 228.900 260.850 ;
        RECT 233.100 259.050 234.900 260.850 ;
        RECT 34.950 256.950 37.050 259.050 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 67.950 256.950 70.050 259.050 ;
        RECT 82.950 256.950 85.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 142.950 256.950 145.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 160.950 256.950 163.050 259.050 ;
        RECT 163.950 256.950 166.050 259.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 29.550 254.550 34.050 256.050 ;
        RECT 30.000 253.950 34.050 254.550 ;
        RECT 38.850 243.600 40.050 256.950 ;
        RECT 44.100 255.150 45.900 256.950 ;
        RECT 59.700 244.800 60.600 256.950 ;
        RECT 65.100 255.150 66.900 256.950 ;
        RECT 59.700 243.900 66.300 244.800 ;
        RECT 59.700 243.600 60.600 243.900 ;
        RECT 17.400 237.600 19.200 243.600 ;
        RECT 38.400 237.600 40.200 243.600 ;
        RECT 58.800 237.600 60.600 243.600 ;
        RECT 64.800 243.600 66.300 243.900 ;
        RECT 83.400 243.600 84.600 256.950 ;
        RECT 86.100 255.150 87.900 256.950 ;
        RECT 101.100 255.150 102.900 256.950 ;
        RECT 105.000 251.400 105.900 256.950 ;
        RECT 107.100 255.150 108.900 256.950 ;
        RECT 100.800 250.500 105.900 251.400 ;
        RECT 64.800 237.600 66.600 243.600 ;
        RECT 82.800 237.600 84.600 243.600 ;
        RECT 97.800 238.500 99.600 249.600 ;
        RECT 100.800 239.400 102.600 250.500 ;
        RECT 103.800 248.400 111.600 249.300 ;
        RECT 103.800 238.500 105.600 248.400 ;
        RECT 97.800 237.600 105.600 238.500 ;
        RECT 109.800 237.600 111.600 248.400 ;
        RECT 122.400 243.600 123.600 256.950 ;
        RECT 143.700 244.800 144.600 256.950 ;
        RECT 149.100 255.150 150.900 256.950 ;
        RECT 161.100 255.150 162.900 256.950 ;
        RECT 143.700 243.900 150.300 244.800 ;
        RECT 143.700 243.600 144.600 243.900 ;
        RECT 122.400 237.600 124.200 243.600 ;
        RECT 142.800 237.600 144.600 243.600 ;
        RECT 148.800 243.600 150.300 243.900 ;
        RECT 164.400 243.600 165.600 256.950 ;
        RECT 182.700 244.800 183.600 256.950 ;
        RECT 188.100 255.150 189.900 256.950 ;
        RECT 182.700 243.900 189.300 244.800 ;
        RECT 182.700 243.600 183.600 243.900 ;
        RECT 148.800 237.600 150.600 243.600 ;
        RECT 164.400 237.600 166.200 243.600 ;
        RECT 181.800 237.600 183.600 243.600 ;
        RECT 187.800 243.600 189.300 243.900 ;
        RECT 206.400 243.600 207.600 256.950 ;
        RECT 209.100 255.150 210.900 256.950 ;
        RECT 224.700 244.800 225.600 256.950 ;
        RECT 230.100 255.150 231.900 256.950 ;
        RECT 242.550 256.050 243.450 265.950 ;
        RECT 250.200 264.000 252.000 272.400 ;
        RECT 248.700 262.800 252.000 264.000 ;
        RECT 279.000 266.400 280.800 272.400 ;
        RECT 298.800 266.400 300.600 272.400 ;
        RECT 248.700 259.050 249.600 262.800 ;
        RECT 251.100 259.050 252.900 260.850 ;
        RECT 257.100 259.050 258.900 260.850 ;
        RECT 262.950 259.950 265.050 262.050 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 242.550 254.550 247.050 256.050 ;
        RECT 243.000 253.950 247.050 254.550 ;
        RECT 248.700 244.800 249.600 256.950 ;
        RECT 254.100 255.150 255.900 256.950 ;
        RECT 263.550 256.050 264.450 259.950 ;
        RECT 272.100 259.050 273.900 260.850 ;
        RECT 279.000 259.050 280.050 266.400 ;
        RECT 299.400 264.300 300.600 266.400 ;
        RECT 301.800 267.300 303.600 272.400 ;
        RECT 307.800 267.300 309.600 272.400 ;
        RECT 301.800 265.950 309.600 267.300 ;
        RECT 320.400 267.300 322.200 272.400 ;
        RECT 326.400 267.300 328.200 272.400 ;
        RECT 320.400 265.950 328.200 267.300 ;
        RECT 329.400 266.400 331.200 272.400 ;
        RECT 329.400 264.300 330.600 266.400 ;
        RECT 346.800 265.200 348.600 272.400 ;
        RECT 364.800 269.400 366.600 272.400 ;
        RECT 299.400 263.250 303.150 264.300 ;
        RECT 295.950 261.450 298.050 262.050 ;
        RECT 284.100 259.050 285.900 260.850 ;
        RECT 290.550 260.550 298.050 261.450 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 283.950 256.950 286.050 259.050 ;
        RECT 259.950 254.550 264.450 256.050 ;
        RECT 275.100 255.150 276.900 256.950 ;
        RECT 259.950 253.950 264.000 254.550 ;
        RECT 279.000 251.400 279.900 256.950 ;
        RECT 281.100 255.150 282.900 256.950 ;
        RECT 290.550 255.450 291.450 260.550 ;
        RECT 295.950 259.950 298.050 260.550 ;
        RECT 299.100 259.050 300.900 260.850 ;
        RECT 301.950 259.050 303.150 263.250 ;
        RECT 326.850 263.250 330.600 264.300 ;
        RECT 344.400 264.300 348.600 265.200 ;
        RECT 315.000 261.450 319.050 262.050 ;
        RECT 305.100 259.050 306.900 260.850 ;
        RECT 314.550 259.950 319.050 261.450 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 304.950 256.950 307.050 259.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 287.550 254.550 291.450 255.450 ;
        RECT 274.800 250.500 279.900 251.400 ;
        RECT 280.950 252.450 283.050 253.050 ;
        RECT 287.550 252.450 288.450 254.550 ;
        RECT 280.950 251.550 288.450 252.450 ;
        RECT 280.950 250.950 283.050 251.550 ;
        RECT 250.950 249.450 253.050 250.050 ;
        RECT 265.950 249.450 268.050 250.050 ;
        RECT 250.950 248.550 268.050 249.450 ;
        RECT 250.950 247.950 253.050 248.550 ;
        RECT 265.950 247.950 268.050 248.550 ;
        RECT 224.700 243.900 231.300 244.800 ;
        RECT 224.700 243.600 225.600 243.900 ;
        RECT 187.800 237.600 189.600 243.600 ;
        RECT 205.800 237.600 207.600 243.600 ;
        RECT 223.800 237.600 225.600 243.600 ;
        RECT 229.800 243.600 231.300 243.900 ;
        RECT 248.700 243.900 255.300 244.800 ;
        RECT 248.700 243.600 249.600 243.900 ;
        RECT 229.800 237.600 231.600 243.600 ;
        RECT 247.800 237.600 249.600 243.600 ;
        RECT 253.800 243.600 255.300 243.900 ;
        RECT 253.800 237.600 255.600 243.600 ;
        RECT 271.800 238.500 273.600 249.600 ;
        RECT 274.800 239.400 276.600 250.500 ;
        RECT 277.800 248.400 285.600 249.300 ;
        RECT 277.800 238.500 279.600 248.400 ;
        RECT 271.800 237.600 279.600 238.500 ;
        RECT 283.800 237.600 285.600 248.400 ;
        RECT 302.850 243.600 304.050 256.950 ;
        RECT 308.100 255.150 309.900 256.950 ;
        RECT 314.550 256.050 315.450 259.950 ;
        RECT 323.100 259.050 324.900 260.850 ;
        RECT 326.850 259.050 328.050 263.250 ;
        RECT 336.000 261.450 340.050 262.050 ;
        RECT 329.100 259.050 330.900 260.850 ;
        RECT 335.550 259.950 340.050 261.450 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 322.950 256.950 325.050 259.050 ;
        RECT 325.950 256.950 328.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 310.950 254.550 315.450 256.050 ;
        RECT 320.100 255.150 321.900 256.950 ;
        RECT 310.950 253.950 315.000 254.550 ;
        RECT 307.950 252.450 310.050 253.050 ;
        RECT 319.950 252.450 322.050 253.050 ;
        RECT 307.950 251.550 322.050 252.450 ;
        RECT 307.950 250.950 310.050 251.550 ;
        RECT 319.950 250.950 322.050 251.550 ;
        RECT 325.950 243.600 327.150 256.950 ;
        RECT 335.550 256.050 336.450 259.950 ;
        RECT 341.100 259.050 342.900 260.850 ;
        RECT 344.400 259.050 345.600 264.300 ;
        RECT 347.100 259.050 348.900 260.850 ;
        RECT 365.400 259.050 366.300 269.400 ;
        RECT 385.800 265.200 387.600 272.400 ;
        RECT 402.300 268.200 404.100 272.400 ;
        RECT 383.400 264.300 387.600 265.200 ;
        RECT 401.400 266.400 404.100 268.200 ;
        RECT 380.100 259.050 381.900 260.850 ;
        RECT 383.400 259.050 384.600 264.300 ;
        RECT 386.100 259.050 387.900 260.850 ;
        RECT 401.400 259.050 402.300 266.400 ;
        RECT 404.100 264.600 405.900 265.500 ;
        RECT 409.800 264.600 411.600 272.400 ;
        RECT 404.100 263.700 411.600 264.600 ;
        RECT 422.400 264.600 424.200 272.400 ;
        RECT 429.900 268.200 431.700 272.400 ;
        RECT 445.800 269.400 447.600 272.400 ;
        RECT 464.400 269.400 466.200 272.400 ;
        RECT 429.900 266.400 432.600 268.200 ;
        RECT 428.100 264.600 429.900 265.500 ;
        RECT 422.400 263.700 429.900 264.600 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 367.950 256.950 370.050 259.050 ;
        RECT 379.950 256.950 382.050 259.050 ;
        RECT 382.950 256.950 385.050 259.050 ;
        RECT 385.950 256.950 388.050 259.050 ;
        RECT 400.950 256.950 403.050 259.050 ;
        RECT 403.950 256.950 406.050 259.050 ;
        RECT 335.550 254.550 340.050 256.050 ;
        RECT 336.000 253.950 340.050 254.550 ;
        RECT 344.400 243.600 345.600 256.950 ;
        RECT 362.100 255.150 363.900 256.950 ;
        RECT 365.400 249.600 366.300 256.950 ;
        RECT 368.100 255.150 369.900 256.950 ;
        RECT 362.700 248.400 366.300 249.600 ;
        RECT 302.400 237.600 304.200 243.600 ;
        RECT 325.800 237.600 327.600 243.600 ;
        RECT 344.400 237.600 346.200 243.600 ;
        RECT 362.700 237.600 364.500 248.400 ;
        RECT 383.400 243.600 384.600 256.950 ;
        RECT 401.400 249.600 402.300 256.950 ;
        RECT 404.100 255.150 405.900 256.950 ;
        RECT 383.400 237.600 385.200 243.600 ;
        RECT 400.800 237.600 402.600 249.600 ;
        RECT 407.700 243.600 408.600 263.700 ;
        RECT 410.100 259.050 411.900 260.850 ;
        RECT 422.100 259.050 423.900 260.850 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 421.950 256.950 424.050 259.050 ;
        RECT 409.950 252.450 412.050 252.750 ;
        RECT 415.950 252.450 418.050 253.050 ;
        RECT 409.950 251.550 418.050 252.450 ;
        RECT 409.950 250.650 412.050 251.550 ;
        RECT 415.950 250.950 418.050 251.550 ;
        RECT 406.800 237.600 408.600 243.600 ;
        RECT 425.400 243.600 426.300 263.700 ;
        RECT 431.700 259.050 432.600 266.400 ;
        RECT 446.400 259.050 447.600 269.400 ;
        RECT 464.700 259.050 465.600 269.400 ;
        RECT 486.300 268.200 488.100 272.400 ;
        RECT 485.400 266.400 488.100 268.200 ;
        RECT 485.400 259.050 486.300 266.400 ;
        RECT 488.100 264.600 489.900 265.500 ;
        RECT 493.800 264.600 495.600 272.400 ;
        RECT 509.400 269.400 511.200 272.400 ;
        RECT 488.100 263.700 495.600 264.600 ;
        RECT 510.300 265.200 511.200 269.400 ;
        RECT 515.400 266.400 517.200 272.400 ;
        RECT 510.300 264.300 513.600 265.200 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 430.950 256.950 433.050 259.050 ;
        RECT 445.950 256.950 448.050 259.050 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 463.950 256.950 466.050 259.050 ;
        RECT 466.950 256.950 469.050 259.050 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 428.100 255.150 429.900 256.950 ;
        RECT 431.700 249.600 432.600 256.950 ;
        RECT 425.400 237.600 427.200 243.600 ;
        RECT 431.400 237.600 433.200 249.600 ;
        RECT 446.400 243.600 447.600 256.950 ;
        RECT 449.100 255.150 450.900 256.950 ;
        RECT 461.100 255.150 462.900 256.950 ;
        RECT 464.700 249.600 465.600 256.950 ;
        RECT 467.100 255.150 468.900 256.950 ;
        RECT 485.400 249.600 486.300 256.950 ;
        RECT 488.100 255.150 489.900 256.950 ;
        RECT 464.700 248.400 468.300 249.600 ;
        RECT 445.800 237.600 447.600 243.600 ;
        RECT 466.500 237.600 468.300 248.400 ;
        RECT 484.800 237.600 486.600 249.600 ;
        RECT 491.700 243.600 492.600 263.700 ;
        RECT 511.800 263.400 513.600 264.300 ;
        RECT 494.100 259.050 495.900 260.850 ;
        RECT 506.100 259.050 507.900 260.850 ;
        RECT 493.950 256.950 496.050 259.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 509.100 255.150 510.900 256.950 ;
        RECT 512.700 252.900 513.600 263.400 ;
        RECT 516.000 259.050 517.050 266.400 ;
        RECT 532.800 265.200 534.600 272.400 ;
        RECT 551.400 269.400 553.200 272.400 ;
        RECT 523.950 261.450 526.050 265.050 ;
        RECT 511.800 252.300 513.600 252.900 ;
        RECT 490.800 237.600 492.600 243.600 ;
        RECT 506.400 251.100 513.600 252.300 ;
        RECT 514.950 256.950 517.050 259.050 ;
        RECT 521.550 261.000 526.050 261.450 ;
        RECT 530.400 264.300 534.600 265.200 ;
        RECT 552.300 265.200 553.200 269.400 ;
        RECT 557.400 266.400 559.200 272.400 ;
        RECT 535.950 264.450 538.050 265.050 ;
        RECT 547.950 264.450 550.050 265.050 ;
        RECT 521.550 260.550 525.450 261.000 ;
        RECT 506.400 249.600 507.600 251.100 ;
        RECT 514.950 249.600 516.300 256.950 ;
        RECT 521.550 256.050 522.450 260.550 ;
        RECT 527.100 259.050 528.900 260.850 ;
        RECT 530.400 259.050 531.600 264.300 ;
        RECT 535.950 263.550 550.050 264.450 ;
        RECT 552.300 264.300 555.600 265.200 ;
        RECT 535.950 262.950 538.050 263.550 ;
        RECT 547.950 262.950 550.050 263.550 ;
        RECT 553.800 263.400 555.600 264.300 ;
        RECT 533.100 259.050 534.900 260.850 ;
        RECT 548.100 259.050 549.900 260.850 ;
        RECT 526.950 256.950 529.050 259.050 ;
        RECT 529.950 256.950 532.050 259.050 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 547.950 256.950 550.050 259.050 ;
        RECT 550.950 256.950 553.050 259.050 ;
        RECT 521.550 254.550 526.050 256.050 ;
        RECT 522.000 253.950 526.050 254.550 ;
        RECT 506.400 237.600 508.200 249.600 ;
        RECT 513.900 248.100 516.300 249.600 ;
        RECT 513.900 237.600 515.700 248.100 ;
        RECT 530.400 243.600 531.600 256.950 ;
        RECT 551.100 255.150 552.900 256.950 ;
        RECT 554.700 252.900 555.600 263.400 ;
        RECT 558.000 259.050 559.050 266.400 ;
        RECT 577.800 265.200 579.600 272.400 ;
        RECT 575.400 264.300 579.600 265.200 ;
        RECT 593.400 269.400 595.200 272.400 ;
        RECT 567.000 261.450 571.050 262.050 ;
        RECT 553.800 252.300 555.600 252.900 ;
        RECT 548.400 251.100 555.600 252.300 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 566.550 259.950 571.050 261.450 ;
        RECT 548.400 249.600 549.600 251.100 ;
        RECT 556.950 249.600 558.300 256.950 ;
        RECT 566.550 256.050 567.450 259.950 ;
        RECT 572.100 259.050 573.900 260.850 ;
        RECT 575.400 259.050 576.600 264.300 ;
        RECT 578.100 259.050 579.900 260.850 ;
        RECT 593.400 259.050 594.600 269.400 ;
        RECT 605.400 267.300 607.200 272.400 ;
        RECT 611.400 267.300 613.200 272.400 ;
        RECT 605.400 265.950 613.200 267.300 ;
        RECT 614.400 266.400 616.200 272.400 ;
        RECT 629.400 269.400 631.200 272.400 ;
        RECT 614.400 264.300 615.600 266.400 ;
        RECT 630.300 265.200 631.200 269.400 ;
        RECT 635.400 266.400 637.200 272.400 ;
        RECT 630.300 264.300 633.600 265.200 ;
        RECT 611.850 263.250 615.600 264.300 ;
        RECT 631.800 263.400 633.600 264.300 ;
        RECT 608.100 259.050 609.900 260.850 ;
        RECT 611.850 259.050 613.050 263.250 ;
        RECT 621.000 261.450 625.050 262.050 ;
        RECT 614.100 259.050 615.900 260.850 ;
        RECT 620.550 259.950 625.050 261.450 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 589.950 256.950 592.050 259.050 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 566.550 254.550 571.050 256.050 ;
        RECT 567.000 253.950 571.050 254.550 ;
        RECT 530.400 237.600 532.200 243.600 ;
        RECT 548.400 237.600 550.200 249.600 ;
        RECT 555.900 248.100 558.300 249.600 ;
        RECT 555.900 237.600 557.700 248.100 ;
        RECT 575.400 243.600 576.600 256.950 ;
        RECT 590.100 255.150 591.900 256.950 ;
        RECT 593.400 243.600 594.600 256.950 ;
        RECT 605.100 255.150 606.900 256.950 ;
        RECT 610.950 243.600 612.150 256.950 ;
        RECT 620.550 256.050 621.450 259.950 ;
        RECT 626.100 259.050 627.900 260.850 ;
        RECT 625.950 256.950 628.050 259.050 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 620.550 254.550 625.050 256.050 ;
        RECT 629.100 255.150 630.900 256.950 ;
        RECT 621.000 253.950 625.050 254.550 ;
        RECT 632.700 252.900 633.600 263.400 ;
        RECT 636.000 259.050 637.050 266.400 ;
        RECT 655.800 265.200 657.600 272.400 ;
        RECT 673.800 269.400 675.600 272.400 ;
        RECT 653.400 264.300 657.600 265.200 ;
        RECT 650.100 259.050 651.900 260.850 ;
        RECT 653.400 259.050 654.600 264.300 ;
        RECT 656.100 259.050 657.900 260.850 ;
        RECT 674.400 259.050 675.300 269.400 ;
        RECT 689.400 264.600 691.200 272.400 ;
        RECT 696.900 268.200 698.700 272.400 ;
        RECT 696.900 266.400 699.600 268.200 ;
        RECT 695.100 264.600 696.900 265.500 ;
        RECT 689.400 263.700 696.900 264.600 ;
        RECT 679.950 261.450 684.000 262.050 ;
        RECT 679.950 259.950 684.450 261.450 ;
        RECT 631.800 252.300 633.600 252.900 ;
        RECT 626.400 251.100 633.600 252.300 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 626.400 249.600 627.600 251.100 ;
        RECT 634.950 249.600 636.300 256.950 ;
        RECT 575.400 237.600 577.200 243.600 ;
        RECT 593.400 237.600 595.200 243.600 ;
        RECT 610.800 237.600 612.600 243.600 ;
        RECT 626.400 237.600 628.200 249.600 ;
        RECT 633.900 248.100 636.300 249.600 ;
        RECT 633.900 237.600 635.700 248.100 ;
        RECT 653.400 243.600 654.600 256.950 ;
        RECT 671.100 255.150 672.900 256.950 ;
        RECT 664.950 252.450 667.050 253.050 ;
        RECT 670.950 252.450 673.050 253.050 ;
        RECT 664.950 251.550 673.050 252.450 ;
        RECT 664.950 250.950 667.050 251.550 ;
        RECT 670.950 250.950 673.050 251.550 ;
        RECT 674.400 249.600 675.300 256.950 ;
        RECT 677.100 255.150 678.900 256.950 ;
        RECT 683.550 252.450 684.450 259.950 ;
        RECT 689.100 259.050 690.900 260.850 ;
        RECT 688.950 256.950 691.050 259.050 ;
        RECT 688.950 252.450 691.050 252.750 ;
        RECT 683.550 251.550 691.050 252.450 ;
        RECT 688.950 250.650 691.050 251.550 ;
        RECT 671.700 248.400 675.300 249.600 ;
        RECT 653.400 237.600 655.200 243.600 ;
        RECT 671.700 237.600 673.500 248.400 ;
        RECT 692.400 243.600 693.300 263.700 ;
        RECT 698.700 259.050 699.600 266.400 ;
        RECT 710.400 267.300 712.200 272.400 ;
        RECT 716.400 267.300 718.200 272.400 ;
        RECT 710.400 265.950 718.200 267.300 ;
        RECT 719.400 266.400 721.200 272.400 ;
        RECT 725.550 266.400 727.350 272.400 ;
        RECT 733.650 269.400 735.450 272.400 ;
        RECT 741.450 269.400 743.250 272.400 ;
        RECT 749.250 270.300 751.050 272.400 ;
        RECT 749.250 269.400 753.000 270.300 ;
        RECT 733.650 268.500 734.700 269.400 ;
        RECT 730.950 267.300 734.700 268.500 ;
        RECT 742.200 268.500 743.250 269.400 ;
        RECT 751.950 268.500 753.000 269.400 ;
        RECT 742.200 267.450 747.150 268.500 ;
        RECT 730.950 266.400 733.050 267.300 ;
        RECT 745.350 266.700 747.150 267.450 ;
        RECT 719.400 264.300 720.600 266.400 ;
        RECT 716.850 263.250 720.600 264.300 ;
        RECT 713.100 259.050 714.900 260.850 ;
        RECT 716.850 259.050 718.050 263.250 ;
        RECT 719.100 259.050 720.900 260.850 ;
        RECT 725.550 259.050 726.750 266.400 ;
        RECT 748.650 265.800 750.450 267.600 ;
        RECT 751.950 266.400 754.050 268.500 ;
        RECT 757.050 266.400 758.850 272.400 ;
        RECT 738.150 264.000 739.950 264.600 ;
        RECT 749.100 264.000 750.150 265.800 ;
        RECT 738.150 262.800 750.150 264.000 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 709.950 256.950 712.050 259.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 725.550 257.250 731.850 259.050 ;
        RECT 725.550 256.950 730.050 257.250 ;
        RECT 695.100 255.150 696.900 256.950 ;
        RECT 698.700 249.600 699.600 256.950 ;
        RECT 710.100 255.150 711.900 256.950 ;
        RECT 692.400 237.600 694.200 243.600 ;
        RECT 698.400 237.600 700.200 249.600 ;
        RECT 715.950 243.600 717.150 256.950 ;
        RECT 725.550 249.600 726.750 256.950 ;
        RECT 727.950 251.400 729.750 253.200 ;
        RECT 728.850 250.200 733.050 251.400 ;
        RECT 738.150 250.200 739.050 262.800 ;
        RECT 749.100 261.600 756.000 262.800 ;
        RECT 749.100 261.000 750.900 261.600 ;
        RECT 755.100 260.850 756.000 261.600 ;
        RECT 752.100 259.800 753.900 260.400 ;
        RECT 745.950 258.600 753.900 259.800 ;
        RECT 755.100 259.050 756.900 260.850 ;
        RECT 745.950 256.950 748.050 258.600 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 747.750 251.700 749.550 252.000 ;
        RECT 757.950 251.700 758.850 266.400 ;
        RECT 773.400 265.200 775.200 272.400 ;
        RECT 793.800 269.400 795.600 272.400 ;
        RECT 812.400 269.400 814.200 272.400 ;
        RECT 829.800 269.400 831.600 272.400 ;
        RECT 841.200 269.400 843.000 272.400 ;
        RECT 773.400 264.300 777.600 265.200 ;
        RECT 773.100 259.050 774.900 260.850 ;
        RECT 776.400 259.050 777.600 264.300 ;
        RECT 784.950 264.450 787.050 264.900 ;
        RECT 790.950 264.450 793.050 265.050 ;
        RECT 784.950 263.550 793.050 264.450 ;
        RECT 784.950 262.800 787.050 263.550 ;
        RECT 790.950 262.950 793.050 263.550 ;
        RECT 779.100 259.050 780.900 260.850 ;
        RECT 794.400 259.050 795.300 269.400 ;
        RECT 802.950 267.450 805.050 268.050 ;
        RECT 808.950 267.450 811.050 268.050 ;
        RECT 802.950 266.550 811.050 267.450 ;
        RECT 802.950 265.950 805.050 266.550 ;
        RECT 808.950 265.950 811.050 266.550 ;
        RECT 812.400 259.050 813.600 269.400 ;
        RECT 823.950 261.450 826.050 262.050 ;
        RECT 818.550 260.550 826.050 261.450 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 796.950 256.950 799.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 747.750 251.100 758.850 251.700 ;
        RECT 715.800 237.600 717.600 243.600 ;
        RECT 725.550 237.600 727.350 249.600 ;
        RECT 730.950 249.300 733.050 250.200 ;
        RECT 733.950 249.300 739.050 250.200 ;
        RECT 741.150 250.500 758.850 251.100 ;
        RECT 741.150 250.200 749.550 250.500 ;
        RECT 733.950 248.400 734.850 249.300 ;
        RECT 732.150 246.600 734.850 248.400 ;
        RECT 735.750 248.100 737.550 248.400 ;
        RECT 741.150 248.100 742.050 250.200 ;
        RECT 757.950 249.600 758.850 250.500 ;
        RECT 735.750 247.200 742.050 248.100 ;
        RECT 742.950 248.700 744.750 249.300 ;
        RECT 742.950 247.500 750.450 248.700 ;
        RECT 735.750 246.600 737.550 247.200 ;
        RECT 749.250 246.600 750.450 247.500 ;
        RECT 730.950 243.600 734.850 245.700 ;
        RECT 739.950 245.550 741.750 246.300 ;
        RECT 744.750 245.550 746.550 246.300 ;
        RECT 739.950 244.500 746.550 245.550 ;
        RECT 749.250 244.500 754.050 246.600 ;
        RECT 733.050 237.600 734.850 243.600 ;
        RECT 740.850 237.600 742.650 244.500 ;
        RECT 749.250 243.600 750.450 244.500 ;
        RECT 748.650 237.600 750.450 243.600 ;
        RECT 757.050 237.600 758.850 249.600 ;
        RECT 776.400 243.600 777.600 256.950 ;
        RECT 791.100 255.150 792.900 256.950 ;
        RECT 794.400 249.600 795.300 256.950 ;
        RECT 797.100 255.150 798.900 256.950 ;
        RECT 809.100 255.150 810.900 256.950 ;
        RECT 775.800 237.600 777.600 243.600 ;
        RECT 791.700 248.400 795.300 249.600 ;
        RECT 791.700 237.600 793.500 248.400 ;
        RECT 812.400 243.600 813.600 256.950 ;
        RECT 818.550 256.050 819.450 260.550 ;
        RECT 823.950 259.950 826.050 260.550 ;
        RECT 830.400 259.050 831.300 269.400 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 814.950 254.550 819.450 256.050 ;
        RECT 827.100 255.150 828.900 256.950 ;
        RECT 814.950 253.950 819.000 254.550 ;
        RECT 830.400 249.600 831.300 256.950 ;
        RECT 833.100 255.150 834.900 256.950 ;
        RECT 841.500 256.050 843.000 269.400 ;
        RECT 838.950 253.950 843.000 256.050 ;
        RECT 827.700 248.400 831.300 249.600 ;
        RECT 812.400 237.600 814.200 243.600 ;
        RECT 827.700 237.600 829.500 248.400 ;
        RECT 841.500 243.600 843.000 253.950 ;
        RECT 845.100 266.400 846.900 272.400 ;
        RECT 855.600 267.600 857.400 272.400 ;
        RECT 860.400 269.400 862.200 272.400 ;
        RECT 863.400 269.400 865.200 272.400 ;
        RECT 866.400 269.400 868.200 272.400 ;
        RECT 870.000 269.400 871.800 272.400 ;
        RECT 876.000 269.400 877.800 272.400 ;
        RECT 883.500 269.400 885.300 272.400 ;
        RECT 886.500 269.400 888.300 272.400 ;
        RECT 889.500 269.400 891.300 272.400 ;
        RECT 860.400 268.500 862.050 269.400 ;
        RECT 863.400 268.500 865.050 269.400 ;
        RECT 866.400 268.500 868.050 269.400 ;
        RECT 870.000 268.500 871.050 269.400 ;
        RECT 876.000 268.500 877.050 269.400 ;
        RECT 853.200 266.400 857.400 267.600 ;
        RECT 859.950 266.400 862.050 268.500 ;
        RECT 862.950 266.400 865.050 268.500 ;
        RECT 865.950 266.400 868.050 268.500 ;
        RECT 868.950 266.400 871.050 268.500 ;
        RECT 874.950 266.400 877.050 268.500 ;
        RECT 883.950 268.500 885.300 269.400 ;
        RECT 886.950 268.500 888.300 269.400 ;
        RECT 889.950 268.500 891.300 269.400 ;
        RECT 878.700 266.400 880.500 268.200 ;
        RECT 883.950 266.400 886.050 268.500 ;
        RECT 886.950 266.400 889.050 268.500 ;
        RECT 889.950 266.400 892.050 268.500 ;
        RECT 845.100 249.600 846.000 266.400 ;
        RECT 853.200 262.800 854.700 266.400 ;
        RECT 879.600 265.200 880.500 266.400 ;
        RECT 859.500 262.800 866.100 264.600 ;
        RECT 846.900 261.300 854.700 262.800 ;
        RECT 872.100 261.900 873.900 264.300 ;
        RECT 879.600 264.000 889.500 265.200 ;
        RECT 881.400 262.050 883.200 262.650 ;
        RECT 884.400 262.200 886.200 264.000 ;
        RECT 846.900 261.000 848.700 261.300 ;
        RECT 851.700 261.000 853.500 261.300 ;
        RECT 855.600 260.400 873.900 261.900 ;
        RECT 877.950 260.850 883.200 262.050 ;
        RECT 855.600 260.100 857.100 260.400 ;
        RECT 850.200 258.900 857.100 260.100 ;
        RECT 877.950 259.950 880.050 260.850 ;
        RECT 888.450 258.900 889.500 264.000 ;
        RECT 891.000 262.800 892.050 266.400 ;
        RECT 893.700 266.400 895.500 272.400 ;
        RECT 904.500 266.400 906.300 272.400 ;
        RECT 893.700 265.500 895.200 266.400 ;
        RECT 893.700 264.300 902.100 265.500 ;
        RECT 900.300 263.700 902.100 264.300 ;
        RECT 905.100 262.800 906.300 266.400 ;
        RECT 891.000 261.600 906.300 262.800 ;
        RECT 850.200 256.050 851.400 258.900 ;
        RECT 858.300 257.700 887.550 258.900 ;
        RECT 858.300 256.200 859.200 257.700 ;
        RECT 847.950 253.950 851.400 256.050 ;
        RECT 854.100 254.400 859.200 256.200 ;
        RECT 862.500 255.900 877.050 256.800 ;
        RECT 883.800 255.900 885.600 256.500 ;
        RECT 862.500 254.700 863.400 255.900 ;
        RECT 874.950 254.700 885.600 255.900 ;
        RECT 886.500 256.200 887.550 257.700 ;
        RECT 888.450 257.100 890.250 258.900 ;
        RECT 892.050 257.550 903.900 258.750 ;
        RECT 892.050 256.200 893.250 257.550 ;
        RECT 886.500 255.150 893.250 256.200 ;
        RECT 902.100 256.050 903.900 257.550 ;
        RECT 895.950 255.750 898.050 256.050 ;
        RECT 862.500 252.900 864.300 254.700 ;
        RECT 868.950 252.900 872.850 254.700 ;
        RECT 868.950 252.600 871.050 252.900 ;
        RECT 874.950 252.600 877.050 254.700 ;
        RECT 894.150 253.950 898.050 255.750 ;
        RECT 901.950 253.950 904.050 256.050 ;
        RECT 894.150 253.200 895.950 253.950 ;
        RECT 882.600 252.300 895.950 253.200 ;
        RECT 846.900 251.700 848.700 252.300 ;
        RECT 882.600 251.700 883.800 252.300 ;
        RECT 894.150 252.150 895.950 252.300 ;
        RECT 846.900 250.500 883.800 251.700 ;
        RECT 886.950 250.500 889.050 250.800 ;
        RECT 845.100 248.700 862.050 249.600 ;
        RECT 841.200 237.600 843.000 243.600 ;
        RECT 847.800 243.600 849.000 248.700 ;
        RECT 859.950 247.500 862.050 248.700 ;
        RECT 865.950 248.400 883.800 249.600 ;
        RECT 886.950 249.300 898.500 250.500 ;
        RECT 886.950 248.700 889.050 249.300 ;
        RECT 896.700 248.700 898.500 249.300 ;
        RECT 865.950 247.500 868.050 248.400 ;
        RECT 882.600 247.800 883.800 248.400 ;
        RECT 900.000 247.800 901.800 248.100 ;
        RECT 849.900 245.700 851.700 246.300 ;
        RECT 856.500 245.700 858.300 246.300 ;
        RECT 869.100 245.700 871.800 247.500 ;
        RECT 849.900 244.500 855.600 245.700 ;
        RECT 856.500 244.500 864.150 245.700 ;
        RECT 847.800 237.600 849.600 243.600 ;
        RECT 853.800 237.600 855.600 244.500 ;
        RECT 863.100 242.700 864.150 244.500 ;
        RECT 868.950 243.600 871.800 245.700 ;
        RECT 874.950 245.100 877.800 247.200 ;
        RECT 882.600 246.600 901.800 247.800 ;
        RECT 859.950 240.600 862.050 242.700 ;
        RECT 863.100 240.600 865.200 242.700 ;
        RECT 866.100 240.600 868.200 242.700 ;
        RECT 860.400 237.600 862.200 240.600 ;
        RECT 863.400 237.600 865.200 240.600 ;
        RECT 866.400 237.600 868.200 240.600 ;
        RECT 870.000 237.600 871.800 243.600 ;
        RECT 876.000 237.600 877.800 245.100 ;
        RECT 883.650 243.300 886.050 245.400 ;
        RECT 886.950 243.300 889.050 245.400 ;
        RECT 889.950 243.300 892.050 245.400 ;
        RECT 883.650 240.600 884.850 243.300 ;
        RECT 886.950 240.600 888.000 243.300 ;
        RECT 889.950 240.600 891.000 243.300 ;
        RECT 882.900 237.600 884.850 240.600 ;
        RECT 885.900 237.600 888.000 240.600 ;
        RECT 888.900 237.600 891.000 240.600 ;
        RECT 895.500 237.600 897.300 246.600 ;
        RECT 900.000 246.300 901.800 246.600 ;
        RECT 905.100 245.400 906.300 261.600 ;
        RECT 902.250 244.500 906.300 245.400 ;
        RECT 902.250 243.600 903.300 244.500 ;
        RECT 901.500 237.600 903.300 243.600 ;
        RECT 13.800 227.400 15.600 233.400 ;
        RECT 14.700 227.100 15.600 227.400 ;
        RECT 19.800 227.400 21.600 233.400 ;
        RECT 19.800 227.100 21.300 227.400 ;
        RECT 14.700 226.200 21.300 227.100 ;
        RECT 14.700 214.050 15.600 226.200 ;
        RECT 32.400 222.300 34.200 233.400 ;
        RECT 38.400 222.300 40.200 233.400 ;
        RECT 32.400 221.400 40.200 222.300 ;
        RECT 41.400 221.400 43.200 233.400 ;
        RECT 61.800 227.400 63.600 233.400 ;
        RECT 20.100 214.050 21.900 215.850 ;
        RECT 35.100 214.050 36.900 215.850 ;
        RECT 41.700 214.050 42.600 221.400 ;
        RECT 62.400 214.050 63.600 227.400 ;
        RECT 80.400 227.400 82.200 233.400 ;
        RECT 101.400 227.400 103.200 233.400 ;
        RECT 80.400 214.050 81.600 227.400 ;
        RECT 101.850 214.050 103.050 227.400 ;
        RECT 124.500 222.600 126.300 233.400 ;
        RECT 145.800 227.400 147.600 233.400 ;
        RECT 122.700 221.400 126.300 222.600 ;
        RECT 107.100 214.050 108.900 215.850 ;
        RECT 119.100 214.050 120.900 215.850 ;
        RECT 122.700 214.050 123.600 221.400 ;
        RECT 125.100 214.050 126.900 215.850 ;
        RECT 140.100 214.050 141.900 215.850 ;
        RECT 145.950 214.050 147.150 227.400 ;
        RECT 166.800 221.400 168.600 233.400 ;
        RECT 169.800 222.300 171.600 233.400 ;
        RECT 175.800 222.300 177.600 233.400 ;
        RECT 188.400 227.400 190.200 233.400 ;
        RECT 188.700 227.100 190.200 227.400 ;
        RECT 194.400 227.400 196.200 233.400 ;
        RECT 214.800 227.400 216.600 233.400 ;
        RECT 236.400 227.400 238.200 233.400 ;
        RECT 256.800 227.400 258.600 233.400 ;
        RECT 277.800 227.400 279.600 233.400 ;
        RECT 298.800 227.400 300.600 233.400 ;
        RECT 194.400 227.100 195.300 227.400 ;
        RECT 188.700 226.200 195.300 227.100 ;
        RECT 169.800 221.400 177.600 222.300 ;
        RECT 167.400 214.050 168.300 221.400 ;
        RECT 169.950 219.450 172.050 220.050 ;
        RECT 184.950 219.450 187.050 220.050 ;
        RECT 169.950 218.550 187.050 219.450 ;
        RECT 169.950 217.950 172.050 218.550 ;
        RECT 184.950 217.950 187.050 218.550 ;
        RECT 173.100 214.050 174.900 215.850 ;
        RECT 188.100 214.050 189.900 215.850 ;
        RECT 194.400 214.050 195.300 226.200 ;
        RECT 215.400 214.050 216.600 227.400 ;
        RECT 236.850 214.050 238.050 227.400 ;
        RECT 241.950 219.450 244.050 220.050 ;
        RECT 247.950 219.450 250.050 220.050 ;
        RECT 241.950 218.550 250.050 219.450 ;
        RECT 241.950 217.950 244.050 218.550 ;
        RECT 247.950 217.950 250.050 218.550 ;
        RECT 242.100 214.050 243.900 215.850 ;
        RECT 257.400 214.050 258.600 227.400 ;
        RECT 259.950 219.450 262.050 220.050 ;
        RECT 271.950 219.450 274.050 220.050 ;
        RECT 259.950 218.550 274.050 219.450 ;
        RECT 259.950 217.950 262.050 218.550 ;
        RECT 271.950 217.950 274.050 218.550 ;
        RECT 260.100 214.050 261.900 215.850 ;
        RECT 272.100 214.050 273.900 215.850 ;
        RECT 277.950 214.050 279.150 227.400 ;
        RECT 299.700 227.100 300.600 227.400 ;
        RECT 304.800 227.400 306.600 233.400 ;
        RECT 322.800 227.400 324.600 233.400 ;
        RECT 341.400 227.400 343.200 233.400 ;
        RECT 359.400 227.400 361.200 233.400 ;
        RECT 304.800 227.100 306.300 227.400 ;
        RECT 299.700 226.200 306.300 227.100 ;
        RECT 280.950 222.450 283.050 223.050 ;
        RECT 295.950 222.450 298.050 223.050 ;
        RECT 280.950 221.550 298.050 222.450 ;
        RECT 280.950 220.950 283.050 221.550 ;
        RECT 295.950 220.950 298.050 221.550 ;
        RECT 294.000 216.450 298.050 217.050 ;
        RECT 293.550 214.950 298.050 216.450 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 19.950 211.950 22.050 214.050 ;
        RECT 22.950 211.950 25.050 214.050 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 79.950 211.950 82.050 214.050 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 121.950 211.950 124.050 214.050 ;
        RECT 124.950 211.950 127.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 142.950 211.950 145.050 214.050 ;
        RECT 145.950 211.950 148.050 214.050 ;
        RECT 148.950 211.950 151.050 214.050 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 184.950 211.950 187.050 214.050 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 214.950 211.950 217.050 214.050 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 232.950 211.950 235.050 214.050 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 256.950 211.950 259.050 214.050 ;
        RECT 259.950 211.950 262.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 280.950 211.950 283.050 214.050 ;
        RECT 14.700 208.200 15.600 211.950 ;
        RECT 17.100 210.150 18.900 211.950 ;
        RECT 23.100 210.150 24.900 211.950 ;
        RECT 32.100 210.150 33.900 211.950 ;
        RECT 38.100 210.150 39.900 211.950 ;
        RECT 14.700 207.000 18.000 208.200 ;
        RECT 16.200 198.600 18.000 207.000 ;
        RECT 41.700 204.600 42.600 211.950 ;
        RECT 59.100 210.150 60.900 211.950 ;
        RECT 62.400 206.700 63.600 211.950 ;
        RECT 65.100 210.150 66.900 211.950 ;
        RECT 77.100 210.150 78.900 211.950 ;
        RECT 37.500 203.400 42.600 204.600 ;
        RECT 59.400 205.800 63.600 206.700 ;
        RECT 80.400 206.700 81.600 211.950 ;
        RECT 83.100 210.150 84.900 211.950 ;
        RECT 85.950 210.450 88.050 211.050 ;
        RECT 91.950 210.450 94.050 211.050 ;
        RECT 85.950 209.550 94.050 210.450 ;
        RECT 98.100 210.150 99.900 211.950 ;
        RECT 85.950 208.950 88.050 209.550 ;
        RECT 91.950 208.950 94.050 209.550 ;
        RECT 100.950 207.750 102.150 211.950 ;
        RECT 104.100 210.150 105.900 211.950 ;
        RECT 98.400 206.700 102.150 207.750 ;
        RECT 80.400 205.800 84.600 206.700 ;
        RECT 37.500 198.600 39.300 203.400 ;
        RECT 59.400 198.600 61.200 205.800 ;
        RECT 82.800 198.600 84.600 205.800 ;
        RECT 98.400 204.600 99.600 206.700 ;
        RECT 97.800 198.600 99.600 204.600 ;
        RECT 100.800 203.700 108.600 205.050 ;
        RECT 100.800 198.600 102.600 203.700 ;
        RECT 106.800 198.600 108.600 203.700 ;
        RECT 122.700 201.600 123.600 211.950 ;
        RECT 143.100 210.150 144.900 211.950 ;
        RECT 146.850 207.750 148.050 211.950 ;
        RECT 149.100 210.150 150.900 211.950 ;
        RECT 146.850 206.700 150.600 207.750 ;
        RECT 140.400 203.700 148.200 205.050 ;
        RECT 122.400 198.600 124.200 201.600 ;
        RECT 140.400 198.600 142.200 203.700 ;
        RECT 146.400 198.600 148.200 203.700 ;
        RECT 149.400 204.600 150.600 206.700 ;
        RECT 167.400 204.600 168.300 211.950 ;
        RECT 170.100 210.150 171.900 211.950 ;
        RECT 176.100 210.150 177.900 211.950 ;
        RECT 185.100 210.150 186.900 211.950 ;
        RECT 191.100 210.150 192.900 211.950 ;
        RECT 194.400 208.200 195.300 211.950 ;
        RECT 212.100 210.150 213.900 211.950 ;
        RECT 192.000 207.000 195.300 208.200 ;
        RECT 149.400 198.600 151.200 204.600 ;
        RECT 167.400 203.400 172.500 204.600 ;
        RECT 170.700 198.600 172.500 203.400 ;
        RECT 192.000 198.600 193.800 207.000 ;
        RECT 215.400 206.700 216.600 211.950 ;
        RECT 218.100 210.150 219.900 211.950 ;
        RECT 233.100 210.150 234.900 211.950 ;
        RECT 212.400 205.800 216.600 206.700 ;
        RECT 220.950 207.450 223.050 208.050 ;
        RECT 229.950 207.450 232.050 208.050 ;
        RECT 235.950 207.750 237.150 211.950 ;
        RECT 239.100 210.150 240.900 211.950 ;
        RECT 220.950 206.550 232.050 207.450 ;
        RECT 220.950 205.950 223.050 206.550 ;
        RECT 229.950 205.950 232.050 206.550 ;
        RECT 233.400 206.700 237.150 207.750 ;
        RECT 212.400 198.600 214.200 205.800 ;
        RECT 233.400 204.600 234.600 206.700 ;
        RECT 232.800 198.600 234.600 204.600 ;
        RECT 235.800 203.700 243.600 205.050 ;
        RECT 235.800 198.600 237.600 203.700 ;
        RECT 241.800 198.600 243.600 203.700 ;
        RECT 257.400 201.600 258.600 211.950 ;
        RECT 275.100 210.150 276.900 211.950 ;
        RECT 278.850 207.750 280.050 211.950 ;
        RECT 281.100 210.150 282.900 211.950 ;
        RECT 293.550 211.050 294.450 214.950 ;
        RECT 299.700 214.050 300.600 226.200 ;
        RECT 305.100 214.050 306.900 215.850 ;
        RECT 317.100 214.050 318.900 215.850 ;
        RECT 322.950 214.050 324.150 227.400 ;
        RECT 328.950 216.450 333.000 217.050 ;
        RECT 328.950 214.950 333.450 216.450 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 307.950 211.950 310.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 293.550 209.550 298.050 211.050 ;
        RECT 294.000 208.950 298.050 209.550 ;
        RECT 299.700 208.200 300.600 211.950 ;
        RECT 302.100 210.150 303.900 211.950 ;
        RECT 308.100 210.150 309.900 211.950 ;
        RECT 320.100 210.150 321.900 211.950 ;
        RECT 278.850 206.700 282.600 207.750 ;
        RECT 299.700 207.000 303.000 208.200 ;
        RECT 256.800 198.600 258.600 201.600 ;
        RECT 272.400 203.700 280.200 205.050 ;
        RECT 272.400 198.600 274.200 203.700 ;
        RECT 278.400 198.600 280.200 203.700 ;
        RECT 281.400 204.600 282.600 206.700 ;
        RECT 281.400 198.600 283.200 204.600 ;
        RECT 301.200 198.600 303.000 207.000 ;
        RECT 323.850 207.750 325.050 211.950 ;
        RECT 326.100 210.150 327.900 211.950 ;
        RECT 332.550 211.050 333.450 214.950 ;
        RECT 338.100 214.050 339.900 215.850 ;
        RECT 341.400 214.050 342.600 227.400 ;
        RECT 359.400 214.050 360.600 227.400 ;
        RECT 376.800 221.400 378.600 233.400 ;
        RECT 382.800 227.400 384.600 233.400 ;
        RECT 377.400 214.050 378.300 221.400 ;
        RECT 380.100 214.050 381.900 215.850 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 379.950 211.950 382.050 214.050 ;
        RECT 328.950 209.550 333.450 211.050 ;
        RECT 328.950 208.950 333.000 209.550 ;
        RECT 323.850 206.700 327.600 207.750 ;
        RECT 317.400 203.700 325.200 205.050 ;
        RECT 317.400 198.600 319.200 203.700 ;
        RECT 323.400 198.600 325.200 203.700 ;
        RECT 326.400 204.600 327.600 206.700 ;
        RECT 326.400 198.600 328.200 204.600 ;
        RECT 341.400 201.600 342.600 211.950 ;
        RECT 356.100 210.150 357.900 211.950 ;
        RECT 359.400 206.700 360.600 211.950 ;
        RECT 362.100 210.150 363.900 211.950 ;
        RECT 359.400 205.800 363.600 206.700 ;
        RECT 341.400 198.600 343.200 201.600 ;
        RECT 361.800 198.600 363.600 205.800 ;
        RECT 377.400 204.600 378.300 211.950 ;
        RECT 383.700 207.300 384.600 227.400 ;
        RECT 398.400 227.400 400.200 233.400 ;
        RECT 422.400 227.400 424.200 233.400 ;
        RECT 443.400 227.400 445.200 233.400 ;
        RECT 463.800 227.400 465.600 233.400 ;
        RECT 482.400 227.400 484.200 233.400 ;
        RECT 398.400 214.050 399.600 227.400 ;
        RECT 422.850 214.050 424.050 227.400 ;
        RECT 435.000 216.450 439.050 217.050 ;
        RECT 428.100 214.050 429.900 215.850 ;
        RECT 434.550 214.950 439.050 216.450 ;
        RECT 385.950 211.950 388.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 400.950 211.950 403.050 214.050 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 424.950 211.950 427.050 214.050 ;
        RECT 427.950 211.950 430.050 214.050 ;
        RECT 386.100 210.150 387.900 211.950 ;
        RECT 395.100 210.150 396.900 211.950 ;
        RECT 380.100 206.400 387.600 207.300 ;
        RECT 380.100 205.500 381.900 206.400 ;
        RECT 377.400 202.800 380.100 204.600 ;
        RECT 378.300 198.600 380.100 202.800 ;
        RECT 385.800 198.600 387.600 206.400 ;
        RECT 398.400 206.700 399.600 211.950 ;
        RECT 401.100 210.150 402.900 211.950 ;
        RECT 419.100 210.150 420.900 211.950 ;
        RECT 421.950 207.750 423.150 211.950 ;
        RECT 425.100 210.150 426.900 211.950 ;
        RECT 434.550 211.050 435.450 214.950 ;
        RECT 443.850 214.050 445.050 227.400 ;
        RECT 449.100 214.050 450.900 215.850 ;
        RECT 458.100 214.050 459.900 215.850 ;
        RECT 463.950 214.050 465.150 227.400 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 448.950 211.950 451.050 214.050 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 434.550 209.550 439.050 211.050 ;
        RECT 440.100 210.150 441.900 211.950 ;
        RECT 435.000 208.950 439.050 209.550 ;
        RECT 442.950 207.750 444.150 211.950 ;
        RECT 446.100 210.150 447.900 211.950 ;
        RECT 461.100 210.150 462.900 211.950 ;
        RECT 419.400 206.700 423.150 207.750 ;
        RECT 440.400 206.700 444.150 207.750 ;
        RECT 464.850 207.750 466.050 211.950 ;
        RECT 467.100 210.150 468.900 211.950 ;
        RECT 479.100 210.150 480.900 211.950 ;
        RECT 464.850 206.700 468.600 207.750 ;
        RECT 482.400 207.300 483.300 227.400 ;
        RECT 488.400 221.400 490.200 233.400 ;
        RECT 508.500 222.600 510.300 233.400 ;
        RECT 514.950 231.450 517.050 232.050 ;
        RECT 523.950 231.450 526.050 232.050 ;
        RECT 514.950 230.550 526.050 231.450 ;
        RECT 514.950 229.950 517.050 230.550 ;
        RECT 523.950 229.950 526.050 230.550 ;
        RECT 530.400 227.400 532.200 233.400 ;
        RECT 551.400 227.400 553.200 233.400 ;
        RECT 572.400 227.400 574.200 233.400 ;
        RECT 592.800 227.400 594.600 233.400 ;
        RECT 506.700 221.400 510.300 222.600 ;
        RECT 485.100 214.050 486.900 215.850 ;
        RECT 488.700 214.050 489.600 221.400 ;
        RECT 490.950 216.450 495.000 217.050 ;
        RECT 490.950 214.950 495.450 216.450 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 398.400 205.800 402.600 206.700 ;
        RECT 400.800 198.600 402.600 205.800 ;
        RECT 419.400 204.600 420.600 206.700 ;
        RECT 418.800 198.600 420.600 204.600 ;
        RECT 421.800 203.700 429.600 205.050 ;
        RECT 440.400 204.600 441.600 206.700 ;
        RECT 421.800 198.600 423.600 203.700 ;
        RECT 427.800 198.600 429.600 203.700 ;
        RECT 439.800 198.600 441.600 204.600 ;
        RECT 442.800 203.700 450.600 205.050 ;
        RECT 442.800 198.600 444.600 203.700 ;
        RECT 448.800 198.600 450.600 203.700 ;
        RECT 458.400 203.700 466.200 205.050 ;
        RECT 458.400 198.600 460.200 203.700 ;
        RECT 464.400 198.600 466.200 203.700 ;
        RECT 467.400 204.600 468.600 206.700 ;
        RECT 479.400 206.400 486.900 207.300 ;
        RECT 467.400 198.600 469.200 204.600 ;
        RECT 479.400 198.600 481.200 206.400 ;
        RECT 485.100 205.500 486.900 206.400 ;
        RECT 488.700 204.600 489.600 211.950 ;
        RECT 494.550 210.450 495.450 214.950 ;
        RECT 503.100 214.050 504.900 215.850 ;
        RECT 506.700 214.050 507.600 221.400 ;
        RECT 511.950 216.450 516.000 217.050 ;
        RECT 509.100 214.050 510.900 215.850 ;
        RECT 511.950 214.950 516.450 216.450 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 505.950 211.950 508.050 214.050 ;
        RECT 508.950 211.950 511.050 214.050 ;
        RECT 491.550 210.000 495.450 210.450 ;
        RECT 490.950 209.550 495.450 210.000 ;
        RECT 490.950 205.950 493.050 209.550 ;
        RECT 486.900 202.800 489.600 204.600 ;
        RECT 486.900 198.600 488.700 202.800 ;
        RECT 506.700 201.600 507.600 211.950 ;
        RECT 515.550 211.050 516.450 214.950 ;
        RECT 530.850 214.050 532.050 227.400 ;
        RECT 536.100 214.050 537.900 215.850 ;
        RECT 551.400 214.050 552.600 227.400 ;
        RECT 569.100 214.050 570.900 215.850 ;
        RECT 572.400 214.050 573.600 227.400 ;
        RECT 587.100 214.050 588.900 215.850 ;
        RECT 592.950 214.050 594.150 227.400 ;
        RECT 611.400 221.400 613.200 233.400 ;
        RECT 618.900 222.900 620.700 233.400 ;
        RECT 634.800 227.400 636.600 233.400 ;
        RECT 635.700 227.100 636.600 227.400 ;
        RECT 640.800 227.400 642.600 233.400 ;
        RECT 640.800 227.100 642.300 227.400 ;
        RECT 635.700 226.200 642.300 227.100 ;
        RECT 618.900 221.400 621.300 222.900 ;
        RECT 611.400 219.900 612.600 221.400 ;
        RECT 611.400 218.700 618.600 219.900 ;
        RECT 616.800 218.100 618.600 218.700 ;
        RECT 614.100 214.050 615.900 215.850 ;
        RECT 526.950 211.950 529.050 214.050 ;
        RECT 529.950 211.950 532.050 214.050 ;
        RECT 532.950 211.950 535.050 214.050 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 547.950 211.950 550.050 214.050 ;
        RECT 550.950 211.950 553.050 214.050 ;
        RECT 553.950 211.950 556.050 214.050 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 571.950 211.950 574.050 214.050 ;
        RECT 586.950 211.950 589.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 595.950 211.950 598.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 511.950 209.550 516.450 211.050 ;
        RECT 527.100 210.150 528.900 211.950 ;
        RECT 511.950 208.950 516.000 209.550 ;
        RECT 514.950 207.450 517.050 207.900 ;
        RECT 523.950 207.450 526.050 208.050 ;
        RECT 529.950 207.750 531.150 211.950 ;
        RECT 533.100 210.150 534.900 211.950 ;
        RECT 548.100 210.150 549.900 211.950 ;
        RECT 514.950 206.550 526.050 207.450 ;
        RECT 514.950 205.800 517.050 206.550 ;
        RECT 523.950 205.950 526.050 206.550 ;
        RECT 527.400 206.700 531.150 207.750 ;
        RECT 551.400 206.700 552.600 211.950 ;
        RECT 554.100 210.150 555.900 211.950 ;
        RECT 527.400 204.600 528.600 206.700 ;
        RECT 551.400 205.800 555.600 206.700 ;
        RECT 506.400 198.600 508.200 201.600 ;
        RECT 526.800 198.600 528.600 204.600 ;
        RECT 529.800 203.700 537.600 205.050 ;
        RECT 529.800 198.600 531.600 203.700 ;
        RECT 535.800 198.600 537.600 203.700 ;
        RECT 553.800 198.600 555.600 205.800 ;
        RECT 572.400 201.600 573.600 211.950 ;
        RECT 590.100 210.150 591.900 211.950 ;
        RECT 593.850 207.750 595.050 211.950 ;
        RECT 596.100 210.150 597.900 211.950 ;
        RECT 611.100 210.150 612.900 211.950 ;
        RECT 593.850 206.700 597.600 207.750 ;
        RECT 617.700 207.600 618.600 218.100 ;
        RECT 619.950 214.050 621.300 221.400 ;
        RECT 635.700 214.050 636.600 226.200 ;
        RECT 656.400 222.300 658.200 233.400 ;
        RECT 662.400 222.300 664.200 233.400 ;
        RECT 656.400 221.400 664.200 222.300 ;
        RECT 665.400 221.400 667.200 233.400 ;
        RECT 682.800 227.400 684.600 233.400 ;
        RECT 706.800 227.400 708.600 233.400 ;
        RECT 731.400 227.400 733.200 233.400 ;
        RECT 637.950 219.450 640.050 220.050 ;
        RECT 655.950 219.450 658.050 220.050 ;
        RECT 637.950 218.550 658.050 219.450 ;
        RECT 637.950 217.950 640.050 218.550 ;
        RECT 655.950 217.950 658.050 218.550 ;
        RECT 641.100 214.050 642.900 215.850 ;
        RECT 659.100 214.050 660.900 215.850 ;
        RECT 665.700 214.050 666.600 221.400 ;
        RECT 677.100 214.050 678.900 215.850 ;
        RECT 682.950 214.050 684.150 227.400 ;
        RECT 697.950 216.450 700.050 217.050 ;
        RECT 692.550 215.550 700.050 216.450 ;
        RECT 619.950 211.950 622.050 214.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 640.950 211.950 643.050 214.050 ;
        RECT 643.950 211.950 646.050 214.050 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 676.950 211.950 679.050 214.050 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 616.800 206.700 618.600 207.600 ;
        RECT 587.400 203.700 595.200 205.050 ;
        RECT 572.400 198.600 574.200 201.600 ;
        RECT 587.400 198.600 589.200 203.700 ;
        RECT 593.400 198.600 595.200 203.700 ;
        RECT 596.400 204.600 597.600 206.700 ;
        RECT 615.300 205.800 618.600 206.700 ;
        RECT 596.400 198.600 598.200 204.600 ;
        RECT 615.300 201.600 616.200 205.800 ;
        RECT 621.000 204.600 622.050 211.950 ;
        RECT 635.700 208.200 636.600 211.950 ;
        RECT 638.100 210.150 639.900 211.950 ;
        RECT 644.100 210.150 645.900 211.950 ;
        RECT 656.100 210.150 657.900 211.950 ;
        RECT 662.100 210.150 663.900 211.950 ;
        RECT 635.700 207.000 639.000 208.200 ;
        RECT 614.400 198.600 616.200 201.600 ;
        RECT 620.400 198.600 622.200 204.600 ;
        RECT 637.200 198.600 639.000 207.000 ;
        RECT 665.700 204.600 666.600 211.950 ;
        RECT 680.100 210.150 681.900 211.950 ;
        RECT 683.850 207.750 685.050 211.950 ;
        RECT 686.100 210.150 687.900 211.950 ;
        RECT 692.550 211.050 693.450 215.550 ;
        RECT 697.950 214.950 700.050 215.550 ;
        RECT 701.100 214.050 702.900 215.850 ;
        RECT 706.950 214.050 708.150 227.400 ;
        RECT 709.950 219.450 712.050 220.050 ;
        RECT 718.950 219.450 721.050 220.050 ;
        RECT 709.950 218.550 721.050 219.450 ;
        RECT 709.950 217.950 712.050 218.550 ;
        RECT 718.950 217.950 721.050 218.550 ;
        RECT 731.850 214.050 733.050 227.400 ;
        RECT 752.700 222.600 754.500 233.400 ;
        RECT 772.800 227.400 774.600 233.400 ;
        RECT 790.800 227.400 792.600 233.400 ;
        RECT 809.400 227.400 811.200 233.400 ;
        RECT 823.200 227.400 825.000 233.400 ;
        RECT 752.700 221.400 756.300 222.600 ;
        RECT 737.100 214.050 738.900 215.850 ;
        RECT 752.100 214.050 753.900 215.850 ;
        RECT 755.400 214.050 756.300 221.400 ;
        RECT 758.100 214.050 759.900 215.850 ;
        RECT 773.400 214.050 774.600 227.400 ;
        RECT 778.950 216.450 781.050 217.050 ;
        RECT 778.950 215.550 786.450 216.450 ;
        RECT 778.950 214.950 781.050 215.550 ;
        RECT 700.950 211.950 703.050 214.050 ;
        RECT 703.950 211.950 706.050 214.050 ;
        RECT 706.950 211.950 709.050 214.050 ;
        RECT 709.950 211.950 712.050 214.050 ;
        RECT 727.950 211.950 730.050 214.050 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 751.950 211.950 754.050 214.050 ;
        RECT 754.950 211.950 757.050 214.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 769.950 211.950 772.050 214.050 ;
        RECT 772.950 211.950 775.050 214.050 ;
        RECT 775.950 211.950 778.050 214.050 ;
        RECT 688.950 209.550 693.450 211.050 ;
        RECT 704.100 210.150 705.900 211.950 ;
        RECT 688.950 208.950 693.000 209.550 ;
        RECT 707.850 207.750 709.050 211.950 ;
        RECT 710.100 210.150 711.900 211.950 ;
        RECT 728.100 210.150 729.900 211.950 ;
        RECT 730.950 207.750 732.150 211.950 ;
        RECT 734.100 210.150 735.900 211.950 ;
        RECT 683.850 206.700 687.600 207.750 ;
        RECT 707.850 206.700 711.600 207.750 ;
        RECT 661.500 203.400 666.600 204.600 ;
        RECT 677.400 203.700 685.200 205.050 ;
        RECT 661.500 198.600 663.300 203.400 ;
        RECT 677.400 198.600 679.200 203.700 ;
        RECT 683.400 198.600 685.200 203.700 ;
        RECT 686.400 204.600 687.600 206.700 ;
        RECT 686.400 198.600 688.200 204.600 ;
        RECT 701.400 203.700 709.200 205.050 ;
        RECT 701.400 198.600 703.200 203.700 ;
        RECT 707.400 198.600 709.200 203.700 ;
        RECT 710.400 204.600 711.600 206.700 ;
        RECT 728.400 206.700 732.150 207.750 ;
        RECT 728.400 204.600 729.600 206.700 ;
        RECT 710.400 198.600 712.200 204.600 ;
        RECT 727.800 198.600 729.600 204.600 ;
        RECT 730.800 203.700 738.600 205.050 ;
        RECT 730.800 198.600 732.600 203.700 ;
        RECT 736.800 198.600 738.600 203.700 ;
        RECT 755.400 201.600 756.300 211.950 ;
        RECT 770.100 210.150 771.900 211.950 ;
        RECT 773.400 206.700 774.600 211.950 ;
        RECT 776.100 210.150 777.900 211.950 ;
        RECT 785.550 211.050 786.450 215.550 ;
        RECT 791.400 214.050 792.600 227.400 ;
        RECT 796.950 216.450 801.000 217.050 ;
        RECT 794.100 214.050 795.900 215.850 ;
        RECT 796.950 214.950 801.450 216.450 ;
        RECT 790.950 211.950 793.050 214.050 ;
        RECT 793.950 211.950 796.050 214.050 ;
        RECT 785.550 209.550 790.050 211.050 ;
        RECT 786.000 208.950 790.050 209.550 ;
        RECT 770.400 205.800 774.600 206.700 ;
        RECT 754.800 198.600 756.600 201.600 ;
        RECT 770.400 198.600 772.200 205.800 ;
        RECT 791.400 201.600 792.600 211.950 ;
        RECT 800.550 211.050 801.450 214.950 ;
        RECT 809.850 214.050 811.050 227.400 ;
        RECT 823.500 217.050 825.000 227.400 ;
        RECT 829.800 227.400 831.600 233.400 ;
        RECT 829.800 222.300 831.000 227.400 ;
        RECT 835.800 226.500 837.600 233.400 ;
        RECT 842.400 230.400 844.200 233.400 ;
        RECT 845.400 230.400 847.200 233.400 ;
        RECT 848.400 230.400 850.200 233.400 ;
        RECT 841.950 228.300 844.050 230.400 ;
        RECT 845.100 228.300 847.200 230.400 ;
        RECT 848.100 228.300 850.200 230.400 ;
        RECT 845.100 226.500 846.150 228.300 ;
        RECT 852.000 227.400 853.800 233.400 ;
        RECT 831.900 225.300 837.600 226.500 ;
        RECT 838.500 225.300 846.150 226.500 ;
        RECT 850.950 225.300 853.800 227.400 ;
        RECT 858.000 225.900 859.800 233.400 ;
        RECT 864.900 230.400 866.850 233.400 ;
        RECT 867.900 230.400 870.000 233.400 ;
        RECT 870.900 230.400 873.000 233.400 ;
        RECT 831.900 224.700 833.700 225.300 ;
        RECT 838.500 224.700 840.300 225.300 ;
        RECT 851.100 223.500 853.800 225.300 ;
        RECT 856.950 223.800 859.800 225.900 ;
        RECT 865.650 227.700 866.850 230.400 ;
        RECT 868.950 227.700 870.000 230.400 ;
        RECT 871.950 227.700 873.000 230.400 ;
        RECT 865.650 225.600 868.050 227.700 ;
        RECT 868.950 225.600 871.050 227.700 ;
        RECT 871.950 225.600 874.050 227.700 ;
        RECT 877.500 224.400 879.300 233.400 ;
        RECT 883.500 227.400 885.300 233.400 ;
        RECT 901.800 227.400 903.600 233.400 ;
        RECT 884.250 226.500 885.300 227.400 ;
        RECT 884.250 225.600 888.300 226.500 ;
        RECT 882.000 224.400 883.800 224.700 ;
        RECT 841.950 222.300 844.050 223.500 ;
        RECT 815.100 214.050 816.900 215.850 ;
        RECT 820.950 214.950 825.000 217.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 811.950 211.950 814.050 214.050 ;
        RECT 814.950 211.950 817.050 214.050 ;
        RECT 800.550 209.550 805.050 211.050 ;
        RECT 806.100 210.150 807.900 211.950 ;
        RECT 801.000 208.950 805.050 209.550 ;
        RECT 808.950 207.750 810.150 211.950 ;
        RECT 812.100 210.150 813.900 211.950 ;
        RECT 806.400 206.700 810.150 207.750 ;
        RECT 806.400 204.600 807.600 206.700 ;
        RECT 790.800 198.600 792.600 201.600 ;
        RECT 805.800 198.600 807.600 204.600 ;
        RECT 808.800 203.700 816.600 205.050 ;
        RECT 808.800 198.600 810.600 203.700 ;
        RECT 814.800 198.600 816.600 203.700 ;
        RECT 823.500 201.600 825.000 214.950 ;
        RECT 823.200 198.600 825.000 201.600 ;
        RECT 827.100 221.400 844.050 222.300 ;
        RECT 847.950 222.600 850.050 223.500 ;
        RECT 864.600 223.200 883.800 224.400 ;
        RECT 864.600 222.600 865.800 223.200 ;
        RECT 882.000 222.900 883.800 223.200 ;
        RECT 847.950 221.400 865.800 222.600 ;
        RECT 868.950 221.700 871.050 222.300 ;
        RECT 878.700 221.700 880.500 222.300 ;
        RECT 827.100 204.600 828.000 221.400 ;
        RECT 868.950 220.500 880.500 221.700 ;
        RECT 828.900 219.300 865.800 220.500 ;
        RECT 868.950 220.200 871.050 220.500 ;
        RECT 828.900 218.700 830.700 219.300 ;
        RECT 864.600 218.700 865.800 219.300 ;
        RECT 876.150 218.700 877.950 218.850 ;
        RECT 850.950 218.100 853.050 218.400 ;
        RECT 829.950 214.950 833.400 217.050 ;
        RECT 832.200 212.100 833.400 214.950 ;
        RECT 836.100 214.800 841.200 216.600 ;
        RECT 840.300 213.300 841.200 214.800 ;
        RECT 844.500 216.300 846.300 218.100 ;
        RECT 850.950 216.300 854.850 218.100 ;
        RECT 856.950 216.300 859.050 218.400 ;
        RECT 864.600 217.800 877.950 218.700 ;
        RECT 876.150 217.050 877.950 217.800 ;
        RECT 844.500 215.100 845.400 216.300 ;
        RECT 856.950 215.100 867.600 216.300 ;
        RECT 844.500 214.200 859.050 215.100 ;
        RECT 865.800 214.500 867.600 215.100 ;
        RECT 868.500 214.800 875.250 215.850 ;
        RECT 876.150 215.250 880.050 217.050 ;
        RECT 877.950 214.950 880.050 215.250 ;
        RECT 883.950 214.950 886.050 217.050 ;
        RECT 868.500 213.300 869.550 214.800 ;
        RECT 840.300 212.100 869.550 213.300 ;
        RECT 870.450 212.100 872.250 213.900 ;
        RECT 874.050 213.450 875.250 214.800 ;
        RECT 884.100 213.450 885.900 214.950 ;
        RECT 874.050 212.250 885.900 213.450 ;
        RECT 832.200 210.900 839.100 212.100 ;
        RECT 837.600 210.600 839.100 210.900 ;
        RECT 828.900 209.700 830.700 210.000 ;
        RECT 833.700 209.700 835.500 210.000 ;
        RECT 828.900 208.200 836.700 209.700 ;
        RECT 837.600 209.100 855.900 210.600 ;
        RECT 835.200 204.600 836.700 208.200 ;
        RECT 841.500 206.400 848.100 208.200 ;
        RECT 854.100 206.700 855.900 209.100 ;
        RECT 859.950 210.150 862.050 211.050 ;
        RECT 859.950 208.950 865.200 210.150 ;
        RECT 863.400 208.350 865.200 208.950 ;
        RECT 866.400 207.000 868.200 208.800 ;
        RECT 870.450 207.000 871.500 212.100 ;
        RECT 887.100 209.400 888.300 225.600 ;
        RECT 902.400 214.050 903.600 227.400 ;
        RECT 904.950 219.450 907.050 220.050 ;
        RECT 910.950 219.450 913.050 220.050 ;
        RECT 904.950 218.550 913.050 219.450 ;
        RECT 904.950 217.950 907.050 218.550 ;
        RECT 910.950 217.950 913.050 218.550 ;
        RECT 905.100 214.050 906.900 215.850 ;
        RECT 901.950 211.950 904.050 214.050 ;
        RECT 904.950 211.950 907.050 214.050 ;
        RECT 861.600 205.800 871.500 207.000 ;
        RECT 873.000 208.200 888.300 209.400 ;
        RECT 861.600 204.600 862.500 205.800 ;
        RECT 873.000 204.600 874.050 208.200 ;
        RECT 882.300 206.700 884.100 207.300 ;
        RECT 827.100 198.600 828.900 204.600 ;
        RECT 835.200 203.400 839.400 204.600 ;
        RECT 837.600 198.600 839.400 203.400 ;
        RECT 841.950 202.500 844.050 204.600 ;
        RECT 844.950 202.500 847.050 204.600 ;
        RECT 847.950 202.500 850.050 204.600 ;
        RECT 850.950 202.500 853.050 204.600 ;
        RECT 856.950 202.500 859.050 204.600 ;
        RECT 860.700 202.800 862.500 204.600 ;
        RECT 842.400 201.600 844.050 202.500 ;
        RECT 845.400 201.600 847.050 202.500 ;
        RECT 848.400 201.600 850.050 202.500 ;
        RECT 852.000 201.600 853.050 202.500 ;
        RECT 858.000 201.600 859.050 202.500 ;
        RECT 865.950 202.500 868.050 204.600 ;
        RECT 868.950 202.500 871.050 204.600 ;
        RECT 871.950 202.500 874.050 204.600 ;
        RECT 875.700 205.500 884.100 206.700 ;
        RECT 875.700 204.600 877.200 205.500 ;
        RECT 887.100 204.600 888.300 208.200 ;
        RECT 865.950 201.600 867.300 202.500 ;
        RECT 868.950 201.600 870.300 202.500 ;
        RECT 871.950 201.600 873.300 202.500 ;
        RECT 842.400 198.600 844.200 201.600 ;
        RECT 845.400 198.600 847.200 201.600 ;
        RECT 848.400 198.600 850.200 201.600 ;
        RECT 852.000 198.600 853.800 201.600 ;
        RECT 858.000 198.600 859.800 201.600 ;
        RECT 865.500 198.600 867.300 201.600 ;
        RECT 868.500 198.600 870.300 201.600 ;
        RECT 871.500 198.600 873.300 201.600 ;
        RECT 875.700 198.600 877.500 204.600 ;
        RECT 886.500 198.600 888.300 204.600 ;
        RECT 889.950 204.450 892.050 205.050 ;
        RECT 898.950 204.450 901.050 205.050 ;
        RECT 889.950 203.550 901.050 204.450 ;
        RECT 889.950 202.950 892.050 203.550 ;
        RECT 898.950 202.950 901.050 203.550 ;
        RECT 902.400 201.600 903.600 211.950 ;
        RECT 907.950 210.450 910.050 211.050 ;
        RECT 916.950 210.450 919.050 211.050 ;
        RECT 907.950 209.550 919.050 210.450 ;
        RECT 907.950 208.950 910.050 209.550 ;
        RECT 916.950 208.950 919.050 209.550 ;
        RECT 901.800 198.600 903.600 201.600 ;
        RECT 13.800 188.400 15.600 194.400 ;
        RECT 14.400 186.300 15.600 188.400 ;
        RECT 16.800 189.300 18.600 194.400 ;
        RECT 22.800 189.300 24.600 194.400 ;
        RECT 16.800 187.950 24.600 189.300 ;
        RECT 35.400 187.200 37.200 194.400 ;
        RECT 35.400 186.300 39.600 187.200 ;
        RECT 14.400 185.250 18.150 186.300 ;
        RECT 14.100 181.050 15.900 182.850 ;
        RECT 16.950 181.050 18.150 185.250 ;
        RECT 20.100 181.050 21.900 182.850 ;
        RECT 35.100 181.050 36.900 182.850 ;
        RECT 38.400 181.050 39.600 186.300 ;
        RECT 58.200 186.000 60.000 194.400 ;
        RECT 56.700 184.800 60.000 186.000 ;
        RECT 77.400 191.400 79.200 194.400 ;
        RECT 41.100 181.050 42.900 182.850 ;
        RECT 56.700 181.050 57.600 184.800 ;
        RECT 59.100 181.050 60.900 182.850 ;
        RECT 65.100 181.050 66.900 182.850 ;
        RECT 77.400 181.050 78.600 191.400 ;
        RECT 99.000 186.000 100.800 194.400 ;
        RECT 118.200 186.000 120.000 194.400 ;
        RECT 137.400 189.300 139.200 194.400 ;
        RECT 143.400 189.300 145.200 194.400 ;
        RECT 137.400 187.950 145.200 189.300 ;
        RECT 146.400 188.400 148.200 194.400 ;
        RECT 167.700 189.600 169.500 194.400 ;
        RECT 164.400 188.400 169.500 189.600 ;
        RECT 146.400 186.300 147.600 188.400 ;
        RECT 99.000 184.800 102.300 186.000 ;
        RECT 92.100 181.050 93.900 182.850 ;
        RECT 98.100 181.050 99.900 182.850 ;
        RECT 101.400 181.050 102.300 184.800 ;
        RECT 116.700 184.800 120.000 186.000 ;
        RECT 143.850 185.250 147.600 186.300 ;
        RECT 116.700 181.050 117.600 184.800 ;
        RECT 119.100 181.050 120.900 182.850 ;
        RECT 125.100 181.050 126.900 182.850 ;
        RECT 140.100 181.050 141.900 182.850 ;
        RECT 143.850 181.050 145.050 185.250 ;
        RECT 146.100 181.050 147.900 182.850 ;
        RECT 164.400 181.050 165.300 188.400 ;
        RECT 192.000 186.000 193.800 194.400 ;
        RECT 212.400 187.200 214.200 194.400 ;
        RECT 212.400 186.300 216.600 187.200 ;
        RECT 192.000 184.800 195.300 186.000 ;
        RECT 167.100 181.050 168.900 182.850 ;
        RECT 173.100 181.050 174.900 182.850 ;
        RECT 185.100 181.050 186.900 182.850 ;
        RECT 191.100 181.050 192.900 182.850 ;
        RECT 194.400 181.050 195.300 184.800 ;
        RECT 212.100 181.050 213.900 182.850 ;
        RECT 215.400 181.050 216.600 186.300 ;
        RECT 227.400 186.600 229.200 194.400 ;
        RECT 234.900 190.200 236.700 194.400 ;
        RECT 234.900 188.400 237.600 190.200 ;
        RECT 257.700 189.600 259.500 194.400 ;
        RECT 274.800 191.400 276.600 194.400 ;
        RECT 295.800 191.400 297.600 194.400 ;
        RECT 233.100 186.600 234.900 187.500 ;
        RECT 227.400 185.700 234.900 186.600 ;
        RECT 218.100 181.050 219.900 182.850 ;
        RECT 227.100 181.050 228.900 182.850 ;
        RECT 4.950 180.450 9.000 181.050 ;
        RECT 4.950 178.950 9.450 180.450 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 22.950 178.950 25.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 73.950 178.950 76.050 181.050 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 145.950 178.950 148.050 181.050 ;
        RECT 163.950 178.950 166.050 181.050 ;
        RECT 166.950 178.950 169.050 181.050 ;
        RECT 169.950 178.950 172.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 8.550 178.050 9.450 178.950 ;
        RECT 8.550 176.550 13.050 178.050 ;
        RECT 9.000 175.950 13.050 176.550 ;
        RECT 17.850 165.600 19.050 178.950 ;
        RECT 23.100 177.150 24.900 178.950 ;
        RECT 38.400 165.600 39.600 178.950 ;
        RECT 56.700 166.800 57.600 178.950 ;
        RECT 62.100 177.150 63.900 178.950 ;
        RECT 74.100 177.150 75.900 178.950 ;
        RECT 56.700 165.900 63.300 166.800 ;
        RECT 56.700 165.600 57.600 165.900 ;
        RECT 17.400 159.600 19.200 165.600 ;
        RECT 37.800 159.600 39.600 165.600 ;
        RECT 55.800 159.600 57.600 165.600 ;
        RECT 61.800 165.600 63.300 165.900 ;
        RECT 77.400 165.600 78.600 178.950 ;
        RECT 95.100 177.150 96.900 178.950 ;
        RECT 85.950 174.450 88.050 175.050 ;
        RECT 91.950 174.450 94.050 174.750 ;
        RECT 85.950 173.550 94.050 174.450 ;
        RECT 85.950 172.950 88.050 173.550 ;
        RECT 91.950 172.650 94.050 173.550 ;
        RECT 101.400 166.800 102.300 178.950 ;
        RECT 95.700 165.900 102.300 166.800 ;
        RECT 95.700 165.600 97.200 165.900 ;
        RECT 61.800 159.600 63.600 165.600 ;
        RECT 77.400 159.600 79.200 165.600 ;
        RECT 95.400 159.600 97.200 165.600 ;
        RECT 101.400 165.600 102.300 165.900 ;
        RECT 116.700 166.800 117.600 178.950 ;
        RECT 122.100 177.150 123.900 178.950 ;
        RECT 137.100 177.150 138.900 178.950 ;
        RECT 116.700 165.900 123.300 166.800 ;
        RECT 116.700 165.600 117.600 165.900 ;
        RECT 101.400 159.600 103.200 165.600 ;
        RECT 115.800 159.600 117.600 165.600 ;
        RECT 121.800 165.600 123.300 165.900 ;
        RECT 142.950 165.600 144.150 178.950 ;
        RECT 164.400 171.600 165.300 178.950 ;
        RECT 170.100 177.150 171.900 178.950 ;
        RECT 188.100 177.150 189.900 178.950 ;
        RECT 178.950 174.450 181.050 175.050 ;
        RECT 184.950 174.450 187.050 175.050 ;
        RECT 178.950 173.550 187.050 174.450 ;
        RECT 178.950 172.950 181.050 173.550 ;
        RECT 184.950 172.950 187.050 173.550 ;
        RECT 121.800 159.600 123.600 165.600 ;
        RECT 142.800 159.600 144.600 165.600 ;
        RECT 163.800 159.600 165.600 171.600 ;
        RECT 166.800 170.700 174.600 171.600 ;
        RECT 166.800 159.600 168.600 170.700 ;
        RECT 172.800 159.600 174.600 170.700 ;
        RECT 194.400 166.800 195.300 178.950 ;
        RECT 188.700 165.900 195.300 166.800 ;
        RECT 188.700 165.600 190.200 165.900 ;
        RECT 188.400 159.600 190.200 165.600 ;
        RECT 194.400 165.600 195.300 165.900 ;
        RECT 215.400 165.600 216.600 178.950 ;
        RECT 194.400 159.600 196.200 165.600 ;
        RECT 214.800 159.600 216.600 165.600 ;
        RECT 230.400 165.600 231.300 185.700 ;
        RECT 236.700 181.050 237.600 188.400 ;
        RECT 254.400 188.400 259.500 189.600 ;
        RECT 254.400 181.050 255.300 188.400 ;
        RECT 257.100 181.050 258.900 182.850 ;
        RECT 263.100 181.050 264.900 182.850 ;
        RECT 275.400 181.050 276.600 191.400 ;
        RECT 296.400 181.050 297.300 191.400 ;
        RECT 308.400 189.300 310.200 194.400 ;
        RECT 314.400 189.300 316.200 194.400 ;
        RECT 308.400 187.950 316.200 189.300 ;
        RECT 317.400 188.400 319.200 194.400 ;
        RECT 329.400 189.300 331.200 194.400 ;
        RECT 335.400 189.300 337.200 194.400 ;
        RECT 317.400 186.300 318.600 188.400 ;
        RECT 329.400 187.950 337.200 189.300 ;
        RECT 338.400 188.400 340.200 194.400 ;
        RECT 338.400 186.300 339.600 188.400 ;
        RECT 314.850 185.250 318.600 186.300 ;
        RECT 335.850 185.250 339.600 186.300 ;
        RECT 358.200 186.000 360.000 194.400 ;
        RECT 377.400 189.300 379.200 194.400 ;
        RECT 383.400 189.300 385.200 194.400 ;
        RECT 377.400 187.950 385.200 189.300 ;
        RECT 386.400 188.400 388.200 194.400 ;
        RECT 404.400 191.400 406.200 194.400 ;
        RECT 386.400 186.300 387.600 188.400 ;
        RECT 311.100 181.050 312.900 182.850 ;
        RECT 314.850 181.050 316.050 185.250 ;
        RECT 317.100 181.050 318.900 182.850 ;
        RECT 332.100 181.050 333.900 182.850 ;
        RECT 335.850 181.050 337.050 185.250 ;
        RECT 356.700 184.800 360.000 186.000 ;
        RECT 383.850 185.250 387.600 186.300 ;
        RECT 340.950 183.450 345.000 184.050 ;
        RECT 338.100 181.050 339.900 182.850 ;
        RECT 340.950 181.950 345.450 183.450 ;
        RECT 232.950 178.950 235.050 181.050 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 253.950 178.950 256.050 181.050 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 259.950 178.950 262.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 277.950 178.950 280.050 181.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 334.950 178.950 337.050 181.050 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 233.100 177.150 234.900 178.950 ;
        RECT 236.700 171.600 237.600 178.950 ;
        RECT 254.400 171.600 255.300 178.950 ;
        RECT 260.100 177.150 261.900 178.950 ;
        RECT 230.400 159.600 232.200 165.600 ;
        RECT 236.400 159.600 238.200 171.600 ;
        RECT 253.800 159.600 255.600 171.600 ;
        RECT 256.800 170.700 264.600 171.600 ;
        RECT 256.800 159.600 258.600 170.700 ;
        RECT 262.800 159.600 264.600 170.700 ;
        RECT 275.400 165.600 276.600 178.950 ;
        RECT 278.100 177.150 279.900 178.950 ;
        RECT 293.100 177.150 294.900 178.950 ;
        RECT 296.400 171.600 297.300 178.950 ;
        RECT 299.100 177.150 300.900 178.950 ;
        RECT 308.100 177.150 309.900 178.950 ;
        RECT 274.800 159.600 276.600 165.600 ;
        RECT 293.700 170.400 297.300 171.600 ;
        RECT 293.700 159.600 295.500 170.400 ;
        RECT 313.950 165.600 315.150 178.950 ;
        RECT 329.100 177.150 330.900 178.950 ;
        RECT 334.950 165.600 336.150 178.950 ;
        RECT 344.550 177.450 345.450 181.950 ;
        RECT 356.700 181.050 357.600 184.800 ;
        RECT 359.100 181.050 360.900 182.850 ;
        RECT 365.100 181.050 366.900 182.850 ;
        RECT 380.100 181.050 381.900 182.850 ;
        RECT 383.850 181.050 385.050 185.250 ;
        RECT 386.100 181.050 387.900 182.850 ;
        RECT 404.700 181.050 405.600 191.400 ;
        RECT 425.700 189.600 427.500 194.400 ;
        RECT 422.400 188.400 427.500 189.600 ;
        RECT 446.400 191.400 448.200 194.400 ;
        RECT 422.400 181.050 423.300 188.400 ;
        RECT 425.100 181.050 426.900 182.850 ;
        RECT 431.100 181.050 432.900 182.850 ;
        RECT 446.400 181.050 447.600 191.400 ;
        RECT 465.000 186.000 466.800 194.400 ;
        RECT 489.000 186.000 490.800 194.400 ;
        RECT 512.700 189.600 514.500 194.400 ;
        RECT 509.400 188.400 514.500 189.600 ;
        RECT 530.400 189.300 532.200 194.400 ;
        RECT 536.400 189.300 538.200 194.400 ;
        RECT 465.000 184.800 468.300 186.000 ;
        RECT 489.000 184.800 492.300 186.000 ;
        RECT 453.000 183.450 457.050 184.050 ;
        RECT 452.550 181.950 457.050 183.450 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 358.950 178.950 361.050 181.050 ;
        RECT 361.950 178.950 364.050 181.050 ;
        RECT 364.950 178.950 367.050 181.050 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 382.950 178.950 385.050 181.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 421.950 178.950 424.050 181.050 ;
        RECT 424.950 178.950 427.050 181.050 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 442.950 178.950 445.050 181.050 ;
        RECT 445.950 178.950 448.050 181.050 ;
        RECT 352.950 177.450 355.050 178.050 ;
        RECT 344.550 176.550 355.050 177.450 ;
        RECT 352.950 175.950 355.050 176.550 ;
        RECT 356.700 166.800 357.600 178.950 ;
        RECT 362.100 177.150 363.900 178.950 ;
        RECT 377.100 177.150 378.900 178.950 ;
        RECT 356.700 165.900 363.300 166.800 ;
        RECT 356.700 165.600 357.600 165.900 ;
        RECT 313.800 159.600 315.600 165.600 ;
        RECT 334.800 159.600 336.600 165.600 ;
        RECT 355.800 159.600 357.600 165.600 ;
        RECT 361.800 165.600 363.300 165.900 ;
        RECT 382.950 165.600 384.150 178.950 ;
        RECT 401.100 177.150 402.900 178.950 ;
        RECT 404.700 171.600 405.600 178.950 ;
        RECT 407.100 177.150 408.900 178.950 ;
        RECT 422.400 171.600 423.300 178.950 ;
        RECT 428.100 177.150 429.900 178.950 ;
        RECT 443.100 177.150 444.900 178.950 ;
        RECT 404.700 170.400 408.300 171.600 ;
        RECT 361.800 159.600 363.600 165.600 ;
        RECT 382.800 159.600 384.600 165.600 ;
        RECT 406.500 159.600 408.300 170.400 ;
        RECT 421.800 159.600 423.600 171.600 ;
        RECT 424.800 170.700 432.600 171.600 ;
        RECT 424.800 159.600 426.600 170.700 ;
        RECT 430.800 159.600 432.600 170.700 ;
        RECT 446.400 165.600 447.600 178.950 ;
        RECT 452.550 178.050 453.450 181.950 ;
        RECT 458.100 181.050 459.900 182.850 ;
        RECT 464.100 181.050 465.900 182.850 ;
        RECT 467.400 181.050 468.300 184.800 ;
        RECT 482.100 181.050 483.900 182.850 ;
        RECT 488.100 181.050 489.900 182.850 ;
        RECT 491.400 181.050 492.300 184.800 ;
        RECT 509.400 181.050 510.300 188.400 ;
        RECT 530.400 187.950 538.200 189.300 ;
        RECT 539.400 188.400 541.200 194.400 ;
        RECT 554.400 191.400 556.200 194.400 ;
        RECT 539.400 186.300 540.600 188.400 ;
        RECT 536.850 185.250 540.600 186.300 ;
        RECT 512.100 181.050 513.900 182.850 ;
        RECT 518.100 181.050 519.900 182.850 ;
        RECT 533.100 181.050 534.900 182.850 ;
        RECT 536.850 181.050 538.050 185.250 ;
        RECT 541.950 183.450 546.000 184.050 ;
        RECT 539.100 181.050 540.900 182.850 ;
        RECT 541.950 181.950 546.450 183.450 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 460.950 178.950 463.050 181.050 ;
        RECT 463.950 178.950 466.050 181.050 ;
        RECT 466.950 178.950 469.050 181.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 484.950 178.950 487.050 181.050 ;
        RECT 487.950 178.950 490.050 181.050 ;
        RECT 490.950 178.950 493.050 181.050 ;
        RECT 508.950 178.950 511.050 181.050 ;
        RECT 511.950 178.950 514.050 181.050 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 517.950 178.950 520.050 181.050 ;
        RECT 529.950 178.950 532.050 181.050 ;
        RECT 532.950 178.950 535.050 181.050 ;
        RECT 535.950 178.950 538.050 181.050 ;
        RECT 538.950 178.950 541.050 181.050 ;
        RECT 452.550 176.550 457.050 178.050 ;
        RECT 461.100 177.150 462.900 178.950 ;
        RECT 453.000 175.950 457.050 176.550 ;
        RECT 467.400 166.800 468.300 178.950 ;
        RECT 485.100 177.150 486.900 178.950 ;
        RECT 491.400 166.800 492.300 178.950 ;
        RECT 509.400 171.600 510.300 178.950 ;
        RECT 515.100 177.150 516.900 178.950 ;
        RECT 530.100 177.150 531.900 178.950 ;
        RECT 461.700 165.900 468.300 166.800 ;
        RECT 461.700 165.600 463.200 165.900 ;
        RECT 446.400 159.600 448.200 165.600 ;
        RECT 461.400 159.600 463.200 165.600 ;
        RECT 467.400 165.600 468.300 165.900 ;
        RECT 485.700 165.900 492.300 166.800 ;
        RECT 485.700 165.600 487.200 165.900 ;
        RECT 467.400 159.600 469.200 165.600 ;
        RECT 485.400 159.600 487.200 165.600 ;
        RECT 491.400 165.600 492.300 165.900 ;
        RECT 491.400 159.600 493.200 165.600 ;
        RECT 508.800 159.600 510.600 171.600 ;
        RECT 511.800 170.700 519.600 171.600 ;
        RECT 511.800 159.600 513.600 170.700 ;
        RECT 517.800 159.600 519.600 170.700 ;
        RECT 535.950 165.600 537.150 178.950 ;
        RECT 545.550 178.050 546.450 181.950 ;
        RECT 554.400 181.050 555.600 191.400 ;
        RECT 576.000 186.000 577.800 194.400 ;
        RECT 595.500 189.600 597.300 194.400 ;
        RECT 595.500 188.400 600.600 189.600 ;
        RECT 576.000 184.800 579.300 186.000 ;
        RECT 556.950 183.450 561.000 184.050 ;
        RECT 564.000 183.450 568.050 184.050 ;
        RECT 556.950 181.950 561.450 183.450 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 545.550 176.550 550.050 178.050 ;
        RECT 551.100 177.150 552.900 178.950 ;
        RECT 546.000 175.950 550.050 176.550 ;
        RECT 554.400 165.600 555.600 178.950 ;
        RECT 560.550 174.450 561.450 181.950 ;
        RECT 563.550 181.950 568.050 183.450 ;
        RECT 563.550 178.050 564.450 181.950 ;
        RECT 569.100 181.050 570.900 182.850 ;
        RECT 575.100 181.050 576.900 182.850 ;
        RECT 578.400 181.050 579.300 184.800 ;
        RECT 590.100 181.050 591.900 182.850 ;
        RECT 596.100 181.050 597.900 182.850 ;
        RECT 599.700 181.050 600.600 188.400 ;
        RECT 621.000 186.000 622.800 194.400 ;
        RECT 638.400 187.200 640.200 194.400 ;
        RECT 659.400 187.200 661.200 194.400 ;
        RECT 680.400 191.400 682.200 194.400 ;
        RECT 638.400 186.300 642.600 187.200 ;
        RECT 659.400 186.300 663.600 187.200 ;
        RECT 621.000 184.800 624.300 186.000 ;
        RECT 614.100 181.050 615.900 182.850 ;
        RECT 620.100 181.050 621.900 182.850 ;
        RECT 623.400 181.050 624.300 184.800 ;
        RECT 638.100 181.050 639.900 182.850 ;
        RECT 641.400 181.050 642.600 186.300 ;
        RECT 644.100 181.050 645.900 182.850 ;
        RECT 659.100 181.050 660.900 182.850 ;
        RECT 662.400 181.050 663.600 186.300 ;
        RECT 664.950 186.450 667.050 187.050 ;
        RECT 670.950 186.450 673.050 187.050 ;
        RECT 664.950 185.550 673.050 186.450 ;
        RECT 664.950 184.950 667.050 185.550 ;
        RECT 670.950 184.950 673.050 185.550 ;
        RECT 665.100 181.050 666.900 182.850 ;
        RECT 680.400 181.050 681.600 191.400 ;
        RECT 694.800 188.400 696.600 194.400 ;
        RECT 700.800 191.400 702.600 194.400 ;
        RECT 694.800 181.050 696.000 188.400 ;
        RECT 701.400 187.500 702.600 191.400 ;
        RECT 696.900 186.600 702.600 187.500 ;
        RECT 704.550 188.400 706.350 194.400 ;
        RECT 712.650 191.400 714.450 194.400 ;
        RECT 720.450 191.400 722.250 194.400 ;
        RECT 728.250 192.300 730.050 194.400 ;
        RECT 728.250 191.400 732.000 192.300 ;
        RECT 712.650 190.500 713.700 191.400 ;
        RECT 709.950 189.300 713.700 190.500 ;
        RECT 721.200 190.500 722.250 191.400 ;
        RECT 730.950 190.500 732.000 191.400 ;
        RECT 721.200 189.450 726.150 190.500 ;
        RECT 709.950 188.400 712.050 189.300 ;
        RECT 724.350 188.700 726.150 189.450 ;
        RECT 696.900 185.700 698.850 186.600 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 571.950 178.950 574.050 181.050 ;
        RECT 574.950 178.950 577.050 181.050 ;
        RECT 577.950 178.950 580.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 598.950 178.950 601.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 619.950 178.950 622.050 181.050 ;
        RECT 622.950 178.950 625.050 181.050 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 664.950 178.950 667.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 694.800 178.950 697.050 181.050 ;
        RECT 563.550 176.550 568.050 178.050 ;
        RECT 572.100 177.150 573.900 178.950 ;
        RECT 564.000 175.950 568.050 176.550 ;
        RECT 568.950 174.450 571.050 175.050 ;
        RECT 560.550 173.550 571.050 174.450 ;
        RECT 568.950 172.950 571.050 173.550 ;
        RECT 578.400 166.800 579.300 178.950 ;
        RECT 593.100 177.150 594.900 178.950 ;
        RECT 583.950 174.450 586.050 175.050 ;
        RECT 592.950 174.450 595.050 175.050 ;
        RECT 583.950 173.550 595.050 174.450 ;
        RECT 583.950 172.950 586.050 173.550 ;
        RECT 592.950 172.950 595.050 173.550 ;
        RECT 599.700 171.600 600.600 178.950 ;
        RECT 617.100 177.150 618.900 178.950 ;
        RECT 572.700 165.900 579.300 166.800 ;
        RECT 572.700 165.600 574.200 165.900 ;
        RECT 535.800 159.600 537.600 165.600 ;
        RECT 554.400 159.600 556.200 165.600 ;
        RECT 572.400 159.600 574.200 165.600 ;
        RECT 578.400 165.600 579.300 165.900 ;
        RECT 590.400 170.700 598.200 171.600 ;
        RECT 578.400 159.600 580.200 165.600 ;
        RECT 590.400 159.600 592.200 170.700 ;
        RECT 596.400 159.600 598.200 170.700 ;
        RECT 599.400 159.600 601.200 171.600 ;
        RECT 623.400 166.800 624.300 178.950 ;
        RECT 617.700 165.900 624.300 166.800 ;
        RECT 617.700 165.600 619.200 165.900 ;
        RECT 617.400 159.600 619.200 165.600 ;
        RECT 623.400 165.600 624.300 165.900 ;
        RECT 641.400 165.600 642.600 178.950 ;
        RECT 662.400 165.600 663.600 178.950 ;
        RECT 677.100 177.150 678.900 178.950 ;
        RECT 623.400 159.600 625.200 165.600 ;
        RECT 640.800 159.600 642.600 165.600 ;
        RECT 661.800 159.600 663.600 165.600 ;
        RECT 680.400 165.600 681.600 178.950 ;
        RECT 694.800 171.600 696.000 178.950 ;
        RECT 697.950 174.300 698.850 185.700 ;
        RECT 704.550 181.050 705.750 188.400 ;
        RECT 727.650 187.800 729.450 189.600 ;
        RECT 730.950 188.400 733.050 190.500 ;
        RECT 736.050 188.400 737.850 194.400 ;
        RECT 717.150 186.000 718.950 186.600 ;
        RECT 728.100 186.000 729.150 187.800 ;
        RECT 717.150 184.800 729.150 186.000 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 704.550 179.250 710.850 181.050 ;
        RECT 704.550 178.950 709.050 179.250 ;
        RECT 701.100 177.150 702.900 178.950 ;
        RECT 696.900 173.400 698.850 174.300 ;
        RECT 696.900 172.500 702.600 173.400 ;
        RECT 680.400 159.600 682.200 165.600 ;
        RECT 694.800 159.600 696.600 171.600 ;
        RECT 701.400 165.600 702.600 172.500 ;
        RECT 700.800 159.600 702.600 165.600 ;
        RECT 704.550 171.600 705.750 178.950 ;
        RECT 706.950 173.400 708.750 175.200 ;
        RECT 707.850 172.200 712.050 173.400 ;
        RECT 717.150 172.200 718.050 184.800 ;
        RECT 728.100 183.600 735.000 184.800 ;
        RECT 728.100 183.000 729.900 183.600 ;
        RECT 734.100 182.850 735.000 183.600 ;
        RECT 731.100 181.800 732.900 182.400 ;
        RECT 724.950 180.600 732.900 181.800 ;
        RECT 734.100 181.050 735.900 182.850 ;
        RECT 724.950 178.950 727.050 180.600 ;
        RECT 733.950 178.950 736.050 181.050 ;
        RECT 726.750 173.700 728.550 174.000 ;
        RECT 736.950 173.700 737.850 188.400 ;
        RECT 754.800 187.500 756.600 194.400 ;
        RECT 760.800 187.500 762.600 194.400 ;
        RECT 766.800 187.500 768.600 194.400 ;
        RECT 772.800 187.500 774.600 194.400 ;
        RECT 793.500 189.600 795.300 194.400 ;
        RECT 815.400 191.400 817.200 194.400 ;
        RECT 793.500 188.400 798.600 189.600 ;
        RECT 753.900 186.300 756.600 187.500 ;
        RECT 758.700 186.300 762.600 187.500 ;
        RECT 764.700 186.300 768.600 187.500 ;
        RECT 770.700 186.300 774.600 187.500 ;
        RECT 753.900 181.050 754.800 186.300 ;
        RECT 758.700 185.400 759.900 186.300 ;
        RECT 764.700 185.400 765.900 186.300 ;
        RECT 770.700 185.400 771.900 186.300 ;
        RECT 755.700 184.200 759.900 185.400 ;
        RECT 755.700 183.600 757.500 184.200 ;
        RECT 751.950 178.950 754.800 181.050 ;
        RECT 726.750 173.100 737.850 173.700 ;
        RECT 704.550 159.600 706.350 171.600 ;
        RECT 709.950 171.300 712.050 172.200 ;
        RECT 712.950 171.300 718.050 172.200 ;
        RECT 720.150 172.500 737.850 173.100 ;
        RECT 753.900 173.700 754.800 178.950 ;
        RECT 758.700 173.700 759.900 184.200 ;
        RECT 761.700 184.200 765.900 185.400 ;
        RECT 761.700 183.600 763.500 184.200 ;
        RECT 764.700 173.700 765.900 184.200 ;
        RECT 767.700 184.200 771.900 185.400 ;
        RECT 767.700 183.600 769.500 184.200 ;
        RECT 770.700 173.700 771.900 184.200 ;
        RECT 773.100 181.050 774.900 182.850 ;
        RECT 788.100 181.050 789.900 182.850 ;
        RECT 794.100 181.050 795.900 182.850 ;
        RECT 797.700 181.050 798.600 188.400 ;
        RECT 815.400 181.050 816.600 191.400 ;
        RECT 833.400 188.400 835.200 194.400 ;
        RECT 844.200 191.400 846.000 194.400 ;
        RECT 826.950 183.450 829.050 187.050 ;
        RECT 824.550 183.000 829.050 183.450 ;
        RECT 824.550 182.550 828.450 183.000 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 793.950 178.950 796.050 181.050 ;
        RECT 796.950 178.950 799.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 814.950 178.950 817.050 181.050 ;
        RECT 791.100 177.150 792.900 178.950 ;
        RECT 781.950 174.450 784.050 175.050 ;
        RECT 793.950 174.450 796.050 175.050 ;
        RECT 753.900 172.500 756.600 173.700 ;
        RECT 758.700 172.500 762.600 173.700 ;
        RECT 764.700 172.500 768.600 173.700 ;
        RECT 770.700 172.500 774.600 173.700 ;
        RECT 781.950 173.550 796.050 174.450 ;
        RECT 781.950 172.950 784.050 173.550 ;
        RECT 793.950 172.950 796.050 173.550 ;
        RECT 720.150 172.200 728.550 172.500 ;
        RECT 712.950 170.400 713.850 171.300 ;
        RECT 711.150 168.600 713.850 170.400 ;
        RECT 714.750 170.100 716.550 170.400 ;
        RECT 720.150 170.100 721.050 172.200 ;
        RECT 736.950 171.600 737.850 172.500 ;
        RECT 714.750 169.200 721.050 170.100 ;
        RECT 721.950 170.700 723.750 171.300 ;
        RECT 721.950 169.500 729.450 170.700 ;
        RECT 714.750 168.600 716.550 169.200 ;
        RECT 728.250 168.600 729.450 169.500 ;
        RECT 709.950 165.600 713.850 167.700 ;
        RECT 718.950 167.550 720.750 168.300 ;
        RECT 723.750 167.550 725.550 168.300 ;
        RECT 718.950 166.500 725.550 167.550 ;
        RECT 728.250 166.500 733.050 168.600 ;
        RECT 712.050 159.600 713.850 165.600 ;
        RECT 719.850 159.600 721.650 166.500 ;
        RECT 728.250 165.600 729.450 166.500 ;
        RECT 727.650 159.600 729.450 165.600 ;
        RECT 736.050 159.600 737.850 171.600 ;
        RECT 754.800 159.600 756.600 172.500 ;
        RECT 760.800 159.600 762.600 172.500 ;
        RECT 766.800 159.600 768.600 172.500 ;
        RECT 772.800 159.600 774.600 172.500 ;
        RECT 797.700 171.600 798.600 178.950 ;
        RECT 812.100 177.150 813.900 178.950 ;
        RECT 788.400 170.700 796.200 171.600 ;
        RECT 788.400 159.600 790.200 170.700 ;
        RECT 794.400 159.600 796.200 170.700 ;
        RECT 797.400 159.600 799.200 171.600 ;
        RECT 815.400 165.600 816.600 178.950 ;
        RECT 817.950 177.450 820.050 178.050 ;
        RECT 824.550 177.450 825.450 182.550 ;
        RECT 830.100 181.050 831.900 182.850 ;
        RECT 833.400 181.050 834.600 188.400 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 817.950 176.550 825.450 177.450 ;
        RECT 817.950 175.950 820.050 176.550 ;
        RECT 833.400 171.600 834.600 178.950 ;
        RECT 844.500 178.050 846.000 191.400 ;
        RECT 841.950 175.950 846.000 178.050 ;
        RECT 815.400 159.600 817.200 165.600 ;
        RECT 833.400 159.600 835.200 171.600 ;
        RECT 844.500 165.600 846.000 175.950 ;
        RECT 848.100 188.400 849.900 194.400 ;
        RECT 858.600 189.600 860.400 194.400 ;
        RECT 863.400 191.400 865.200 194.400 ;
        RECT 866.400 191.400 868.200 194.400 ;
        RECT 869.400 191.400 871.200 194.400 ;
        RECT 873.000 191.400 874.800 194.400 ;
        RECT 879.000 191.400 880.800 194.400 ;
        RECT 886.500 191.400 888.300 194.400 ;
        RECT 889.500 191.400 891.300 194.400 ;
        RECT 892.500 191.400 894.300 194.400 ;
        RECT 863.400 190.500 865.050 191.400 ;
        RECT 866.400 190.500 868.050 191.400 ;
        RECT 869.400 190.500 871.050 191.400 ;
        RECT 873.000 190.500 874.050 191.400 ;
        RECT 879.000 190.500 880.050 191.400 ;
        RECT 856.200 188.400 860.400 189.600 ;
        RECT 862.950 188.400 865.050 190.500 ;
        RECT 865.950 188.400 868.050 190.500 ;
        RECT 868.950 188.400 871.050 190.500 ;
        RECT 871.950 188.400 874.050 190.500 ;
        RECT 877.950 188.400 880.050 190.500 ;
        RECT 886.950 190.500 888.300 191.400 ;
        RECT 889.950 190.500 891.300 191.400 ;
        RECT 892.950 190.500 894.300 191.400 ;
        RECT 881.700 188.400 883.500 190.200 ;
        RECT 886.950 188.400 889.050 190.500 ;
        RECT 889.950 188.400 892.050 190.500 ;
        RECT 892.950 188.400 895.050 190.500 ;
        RECT 848.100 171.600 849.000 188.400 ;
        RECT 856.200 184.800 857.700 188.400 ;
        RECT 882.600 187.200 883.500 188.400 ;
        RECT 862.500 184.800 869.100 186.600 ;
        RECT 849.900 183.300 857.700 184.800 ;
        RECT 875.100 183.900 876.900 186.300 ;
        RECT 882.600 186.000 892.500 187.200 ;
        RECT 884.400 184.050 886.200 184.650 ;
        RECT 887.400 184.200 889.200 186.000 ;
        RECT 849.900 183.000 851.700 183.300 ;
        RECT 854.700 183.000 856.500 183.300 ;
        RECT 858.600 182.400 876.900 183.900 ;
        RECT 880.950 182.850 886.200 184.050 ;
        RECT 858.600 182.100 860.100 182.400 ;
        RECT 853.200 180.900 860.100 182.100 ;
        RECT 880.950 181.950 883.050 182.850 ;
        RECT 891.450 180.900 892.500 186.000 ;
        RECT 894.000 184.800 895.050 188.400 ;
        RECT 896.700 188.400 898.500 194.400 ;
        RECT 907.500 188.400 909.300 194.400 ;
        RECT 896.700 187.500 898.200 188.400 ;
        RECT 896.700 186.300 905.100 187.500 ;
        RECT 903.300 185.700 905.100 186.300 ;
        RECT 908.100 184.800 909.300 188.400 ;
        RECT 894.000 183.600 909.300 184.800 ;
        RECT 853.200 178.050 854.400 180.900 ;
        RECT 861.300 179.700 890.550 180.900 ;
        RECT 861.300 178.200 862.200 179.700 ;
        RECT 850.950 175.950 854.400 178.050 ;
        RECT 857.100 176.400 862.200 178.200 ;
        RECT 865.500 177.900 880.050 178.800 ;
        RECT 886.800 177.900 888.600 178.500 ;
        RECT 865.500 176.700 866.400 177.900 ;
        RECT 877.950 176.700 888.600 177.900 ;
        RECT 889.500 178.200 890.550 179.700 ;
        RECT 891.450 179.100 893.250 180.900 ;
        RECT 895.050 179.550 906.900 180.750 ;
        RECT 895.050 178.200 896.250 179.550 ;
        RECT 889.500 177.150 896.250 178.200 ;
        RECT 905.100 178.050 906.900 179.550 ;
        RECT 898.950 177.750 901.050 178.050 ;
        RECT 865.500 174.900 867.300 176.700 ;
        RECT 871.950 174.900 875.850 176.700 ;
        RECT 871.950 174.600 874.050 174.900 ;
        RECT 877.950 174.600 880.050 176.700 ;
        RECT 897.150 175.950 901.050 177.750 ;
        RECT 904.950 175.950 907.050 178.050 ;
        RECT 897.150 175.200 898.950 175.950 ;
        RECT 885.600 174.300 898.950 175.200 ;
        RECT 849.900 173.700 851.700 174.300 ;
        RECT 885.600 173.700 886.800 174.300 ;
        RECT 897.150 174.150 898.950 174.300 ;
        RECT 849.900 172.500 886.800 173.700 ;
        RECT 889.950 172.500 892.050 172.800 ;
        RECT 848.100 170.700 865.050 171.600 ;
        RECT 844.200 159.600 846.000 165.600 ;
        RECT 850.800 165.600 852.000 170.700 ;
        RECT 862.950 169.500 865.050 170.700 ;
        RECT 868.950 170.400 886.800 171.600 ;
        RECT 889.950 171.300 901.500 172.500 ;
        RECT 889.950 170.700 892.050 171.300 ;
        RECT 899.700 170.700 901.500 171.300 ;
        RECT 868.950 169.500 871.050 170.400 ;
        RECT 885.600 169.800 886.800 170.400 ;
        RECT 903.000 169.800 904.800 170.100 ;
        RECT 852.900 167.700 854.700 168.300 ;
        RECT 859.500 167.700 861.300 168.300 ;
        RECT 872.100 167.700 874.800 169.500 ;
        RECT 852.900 166.500 858.600 167.700 ;
        RECT 859.500 166.500 867.150 167.700 ;
        RECT 850.800 159.600 852.600 165.600 ;
        RECT 856.800 159.600 858.600 166.500 ;
        RECT 866.100 164.700 867.150 166.500 ;
        RECT 871.950 165.600 874.800 167.700 ;
        RECT 877.950 167.100 880.800 169.200 ;
        RECT 885.600 168.600 904.800 169.800 ;
        RECT 862.950 162.600 865.050 164.700 ;
        RECT 866.100 162.600 868.200 164.700 ;
        RECT 869.100 162.600 871.200 164.700 ;
        RECT 863.400 159.600 865.200 162.600 ;
        RECT 866.400 159.600 868.200 162.600 ;
        RECT 869.400 159.600 871.200 162.600 ;
        RECT 873.000 159.600 874.800 165.600 ;
        RECT 879.000 159.600 880.800 167.100 ;
        RECT 886.650 165.300 889.050 167.400 ;
        RECT 889.950 165.300 892.050 167.400 ;
        RECT 892.950 165.300 895.050 167.400 ;
        RECT 886.650 162.600 887.850 165.300 ;
        RECT 889.950 162.600 891.000 165.300 ;
        RECT 892.950 162.600 894.000 165.300 ;
        RECT 885.900 159.600 887.850 162.600 ;
        RECT 888.900 159.600 891.000 162.600 ;
        RECT 891.900 159.600 894.000 162.600 ;
        RECT 898.500 159.600 900.300 168.600 ;
        RECT 903.000 168.300 904.800 168.600 ;
        RECT 908.100 167.400 909.300 183.600 ;
        RECT 910.950 178.950 913.050 181.050 ;
        RECT 911.550 172.050 912.450 178.950 ;
        RECT 910.950 169.950 913.050 172.050 ;
        RECT 905.250 166.500 909.300 167.400 ;
        RECT 905.250 165.600 906.300 166.500 ;
        RECT 904.500 159.600 906.300 165.600 ;
        RECT 13.800 143.400 15.600 155.400 ;
        RECT 16.800 144.300 18.600 155.400 ;
        RECT 22.800 144.300 24.600 155.400 ;
        RECT 35.400 149.400 37.200 155.400 ;
        RECT 35.700 149.100 37.200 149.400 ;
        RECT 41.400 149.400 43.200 155.400 ;
        RECT 41.400 149.100 42.300 149.400 ;
        RECT 35.700 148.200 42.300 149.100 ;
        RECT 16.800 143.400 24.600 144.300 ;
        RECT 14.400 136.050 15.300 143.400 ;
        RECT 16.950 141.450 19.050 142.050 ;
        RECT 37.950 141.450 40.050 142.050 ;
        RECT 16.950 140.550 40.050 141.450 ;
        RECT 16.950 139.950 19.050 140.550 ;
        RECT 37.950 139.950 40.050 140.550 ;
        RECT 20.100 136.050 21.900 137.850 ;
        RECT 35.100 136.050 36.900 137.850 ;
        RECT 41.400 136.050 42.300 148.200 ;
        RECT 56.400 144.300 58.200 155.400 ;
        RECT 62.400 144.300 64.200 155.400 ;
        RECT 56.400 143.400 64.200 144.300 ;
        RECT 65.400 143.400 67.200 155.400 ;
        RECT 80.400 149.400 82.200 155.400 ;
        RECT 80.700 149.100 82.200 149.400 ;
        RECT 86.400 149.400 88.200 155.400 ;
        RECT 106.800 149.400 108.600 155.400 ;
        RECT 86.400 149.100 87.300 149.400 ;
        RECT 80.700 148.200 87.300 149.100 ;
        RECT 59.100 136.050 60.900 137.850 ;
        RECT 65.700 136.050 66.600 143.400 ;
        RECT 80.100 136.050 81.900 137.850 ;
        RECT 86.400 136.050 87.300 148.200 ;
        RECT 107.400 136.050 108.600 149.400 ;
        RECT 124.800 143.400 126.600 155.400 ;
        RECT 127.800 144.300 129.600 155.400 ;
        RECT 133.800 144.300 135.600 155.400 ;
        RECT 148.800 149.400 150.600 155.400 ;
        RECT 127.800 143.400 135.600 144.300 ;
        RECT 149.700 149.100 150.600 149.400 ;
        RECT 154.800 149.400 156.600 155.400 ;
        RECT 175.800 149.400 177.600 155.400 ;
        RECT 197.400 149.400 199.200 155.400 ;
        RECT 154.800 149.100 156.300 149.400 ;
        RECT 149.700 148.200 156.300 149.100 ;
        RECT 125.400 136.050 126.300 143.400 ;
        RECT 131.100 136.050 132.900 137.850 ;
        RECT 149.700 136.050 150.600 148.200 ;
        RECT 151.950 141.450 154.050 142.050 ;
        RECT 160.950 141.450 163.050 142.050 ;
        RECT 151.950 140.550 163.050 141.450 ;
        RECT 151.950 139.950 154.050 140.550 ;
        RECT 160.950 139.950 163.050 140.550 ;
        RECT 155.100 136.050 156.900 137.850 ;
        RECT 170.100 136.050 171.900 137.850 ;
        RECT 175.950 136.050 177.150 149.400 ;
        RECT 197.700 149.100 199.200 149.400 ;
        RECT 203.400 149.400 205.200 155.400 ;
        RECT 220.800 149.400 222.600 155.400 ;
        RECT 203.400 149.100 204.300 149.400 ;
        RECT 197.700 148.200 204.300 149.100 ;
        RECT 178.950 141.450 181.050 142.050 ;
        RECT 196.950 141.450 199.050 142.050 ;
        RECT 178.950 140.550 199.050 141.450 ;
        RECT 178.950 139.950 181.050 140.550 ;
        RECT 196.950 139.950 199.050 140.550 ;
        RECT 197.100 136.050 198.900 137.850 ;
        RECT 203.400 136.050 204.300 148.200 ;
        RECT 221.700 149.100 222.600 149.400 ;
        RECT 226.800 149.400 228.600 155.400 ;
        RECT 244.800 149.400 246.600 155.400 ;
        RECT 265.800 149.400 267.600 155.400 ;
        RECT 287.400 149.400 289.200 155.400 ;
        RECT 226.800 149.100 228.300 149.400 ;
        RECT 221.700 148.200 228.300 149.100 ;
        RECT 221.700 136.050 222.600 148.200 ;
        RECT 223.950 141.450 226.050 142.050 ;
        RECT 232.950 141.450 235.050 142.050 ;
        RECT 223.950 140.550 235.050 141.450 ;
        RECT 223.950 139.950 226.050 140.550 ;
        RECT 232.950 139.950 235.050 140.550 ;
        RECT 235.950 138.450 238.050 138.900 ;
        RECT 241.950 138.450 244.050 139.050 ;
        RECT 227.100 136.050 228.900 137.850 ;
        RECT 235.950 137.550 244.050 138.450 ;
        RECT 235.950 136.800 238.050 137.550 ;
        RECT 241.950 136.950 244.050 137.550 ;
        RECT 245.400 136.050 246.600 149.400 ;
        RECT 248.100 136.050 249.900 137.850 ;
        RECT 260.100 136.050 261.900 137.850 ;
        RECT 265.950 136.050 267.150 149.400 ;
        RECT 287.700 149.100 289.200 149.400 ;
        RECT 293.400 149.400 295.200 155.400 ;
        RECT 313.800 149.400 315.600 155.400 ;
        RECT 337.800 149.400 339.600 155.400 ;
        RECT 293.400 149.100 294.300 149.400 ;
        RECT 287.700 148.200 294.300 149.100 ;
        RECT 287.100 136.050 288.900 137.850 ;
        RECT 293.400 136.050 294.300 148.200 ;
        RECT 295.950 138.450 298.050 139.050 ;
        RECT 301.950 138.450 304.050 139.050 ;
        RECT 295.950 137.550 304.050 138.450 ;
        RECT 295.950 136.950 298.050 137.550 ;
        RECT 301.950 136.950 304.050 137.550 ;
        RECT 308.100 136.050 309.900 137.850 ;
        RECT 313.950 136.050 315.150 149.400 ;
        RECT 316.950 144.450 319.050 145.050 ;
        RECT 325.950 144.450 328.050 148.050 ;
        RECT 316.950 144.000 328.050 144.450 ;
        RECT 316.950 143.550 327.450 144.000 ;
        RECT 316.950 142.950 319.050 143.550 ;
        RECT 338.400 136.050 339.600 149.400 ;
        RECT 353.400 149.400 355.200 155.400 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 31.950 133.950 34.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 55.950 133.950 58.050 136.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 157.950 133.950 160.050 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 292.950 133.950 295.050 136.050 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 310.950 133.950 313.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 14.400 126.600 15.300 133.950 ;
        RECT 17.100 132.150 18.900 133.950 ;
        RECT 23.100 132.150 24.900 133.950 ;
        RECT 32.100 132.150 33.900 133.950 ;
        RECT 38.100 132.150 39.900 133.950 ;
        RECT 41.400 130.200 42.300 133.950 ;
        RECT 56.100 132.150 57.900 133.950 ;
        RECT 62.100 132.150 63.900 133.950 ;
        RECT 39.000 129.000 42.300 130.200 ;
        RECT 14.400 125.400 19.500 126.600 ;
        RECT 17.700 120.600 19.500 125.400 ;
        RECT 39.000 120.600 40.800 129.000 ;
        RECT 65.700 126.600 66.600 133.950 ;
        RECT 77.100 132.150 78.900 133.950 ;
        RECT 83.100 132.150 84.900 133.950 ;
        RECT 86.400 130.200 87.300 133.950 ;
        RECT 104.100 132.150 105.900 133.950 ;
        RECT 61.500 125.400 66.600 126.600 ;
        RECT 84.000 129.000 87.300 130.200 ;
        RECT 61.500 120.600 63.300 125.400 ;
        RECT 84.000 120.600 85.800 129.000 ;
        RECT 107.400 128.700 108.600 133.950 ;
        RECT 110.100 132.150 111.900 133.950 ;
        RECT 104.400 127.800 108.600 128.700 ;
        RECT 104.400 120.600 106.200 127.800 ;
        RECT 125.400 126.600 126.300 133.950 ;
        RECT 128.100 132.150 129.900 133.950 ;
        RECT 134.100 132.150 135.900 133.950 ;
        RECT 149.700 130.200 150.600 133.950 ;
        RECT 152.100 132.150 153.900 133.950 ;
        RECT 158.100 132.150 159.900 133.950 ;
        RECT 173.100 132.150 174.900 133.950 ;
        RECT 149.700 129.000 153.000 130.200 ;
        RECT 125.400 125.400 130.500 126.600 ;
        RECT 128.700 120.600 130.500 125.400 ;
        RECT 151.200 120.600 153.000 129.000 ;
        RECT 176.850 129.750 178.050 133.950 ;
        RECT 179.100 132.150 180.900 133.950 ;
        RECT 194.100 132.150 195.900 133.950 ;
        RECT 200.100 132.150 201.900 133.950 ;
        RECT 203.400 130.200 204.300 133.950 ;
        RECT 176.850 128.700 180.600 129.750 ;
        RECT 170.400 125.700 178.200 127.050 ;
        RECT 170.400 120.600 172.200 125.700 ;
        RECT 176.400 120.600 178.200 125.700 ;
        RECT 179.400 126.600 180.600 128.700 ;
        RECT 201.000 129.000 204.300 130.200 ;
        RECT 221.700 130.200 222.600 133.950 ;
        RECT 224.100 132.150 225.900 133.950 ;
        RECT 230.100 132.150 231.900 133.950 ;
        RECT 221.700 129.000 225.000 130.200 ;
        RECT 179.400 120.600 181.200 126.600 ;
        RECT 201.000 120.600 202.800 129.000 ;
        RECT 223.200 120.600 225.000 129.000 ;
        RECT 245.400 123.600 246.600 133.950 ;
        RECT 263.100 132.150 264.900 133.950 ;
        RECT 266.850 129.750 268.050 133.950 ;
        RECT 269.100 132.150 270.900 133.950 ;
        RECT 284.100 132.150 285.900 133.950 ;
        RECT 290.100 132.150 291.900 133.950 ;
        RECT 293.400 130.200 294.300 133.950 ;
        RECT 311.100 132.150 312.900 133.950 ;
        RECT 266.850 128.700 270.600 129.750 ;
        RECT 244.800 120.600 246.600 123.600 ;
        RECT 260.400 125.700 268.200 127.050 ;
        RECT 260.400 120.600 262.200 125.700 ;
        RECT 266.400 120.600 268.200 125.700 ;
        RECT 269.400 126.600 270.600 128.700 ;
        RECT 291.000 129.000 294.300 130.200 ;
        RECT 314.850 129.750 316.050 133.950 ;
        RECT 317.100 132.150 318.900 133.950 ;
        RECT 335.100 132.150 336.900 133.950 ;
        RECT 269.400 120.600 271.200 126.600 ;
        RECT 291.000 120.600 292.800 129.000 ;
        RECT 314.850 128.700 318.600 129.750 ;
        RECT 338.400 128.700 339.600 133.950 ;
        RECT 341.100 132.150 342.900 133.950 ;
        RECT 350.100 132.150 351.900 133.950 ;
        RECT 353.400 129.300 354.300 149.400 ;
        RECT 359.400 143.400 361.200 155.400 ;
        RECT 373.800 143.400 375.600 155.400 ;
        RECT 376.800 144.300 378.600 155.400 ;
        RECT 382.800 144.300 384.600 155.400 ;
        RECT 398.400 149.400 400.200 155.400 ;
        RECT 398.700 149.100 400.200 149.400 ;
        RECT 404.400 149.400 406.200 155.400 ;
        RECT 422.400 149.400 424.200 155.400 ;
        RECT 445.800 149.400 447.600 155.400 ;
        RECT 467.400 149.400 469.200 155.400 ;
        RECT 472.950 153.450 475.050 153.900 ;
        RECT 478.950 153.450 481.050 154.050 ;
        RECT 472.950 152.550 481.050 153.450 ;
        RECT 472.950 151.800 475.050 152.550 ;
        RECT 478.950 151.950 481.050 152.550 ;
        RECT 404.400 149.100 405.300 149.400 ;
        RECT 398.700 148.200 405.300 149.100 ;
        RECT 376.800 143.400 384.600 144.300 ;
        RECT 356.100 136.050 357.900 137.850 ;
        RECT 359.700 136.050 360.600 143.400 ;
        RECT 374.400 136.050 375.300 143.400 ;
        RECT 379.950 141.450 382.050 142.050 ;
        RECT 394.950 141.450 397.050 142.050 ;
        RECT 379.950 140.550 397.050 141.450 ;
        RECT 379.950 139.950 382.050 140.550 ;
        RECT 394.950 139.950 397.050 140.550 ;
        RECT 380.100 136.050 381.900 137.850 ;
        RECT 398.100 136.050 399.900 137.850 ;
        RECT 404.400 136.050 405.300 148.200 ;
        RECT 422.400 136.050 423.600 149.400 ;
        RECT 440.100 136.050 441.900 137.850 ;
        RECT 445.950 136.050 447.150 149.400 ;
        RECT 464.100 136.050 465.900 137.850 ;
        RECT 467.400 136.050 468.600 149.400 ;
        RECT 484.800 143.400 486.600 155.400 ;
        RECT 487.800 144.300 489.600 155.400 ;
        RECT 493.800 144.300 495.600 155.400 ;
        RECT 506.400 149.400 508.200 155.400 ;
        RECT 506.700 149.100 508.200 149.400 ;
        RECT 512.400 149.400 514.200 155.400 ;
        RECT 529.800 149.400 531.600 155.400 ;
        RECT 512.400 149.100 513.300 149.400 ;
        RECT 506.700 148.200 513.300 149.100 ;
        RECT 487.800 143.400 495.600 144.300 ;
        RECT 485.400 136.050 486.300 143.400 ;
        RECT 491.100 136.050 492.900 137.850 ;
        RECT 506.100 136.050 507.900 137.850 ;
        RECT 512.400 136.050 513.300 148.200 ;
        RECT 530.700 149.100 531.600 149.400 ;
        RECT 535.800 149.400 537.600 155.400 ;
        RECT 535.800 149.100 537.300 149.400 ;
        RECT 530.700 148.200 537.300 149.100 ;
        RECT 530.700 136.050 531.600 148.200 ;
        RECT 551.400 144.300 553.200 155.400 ;
        RECT 557.400 144.300 559.200 155.400 ;
        RECT 551.400 143.400 559.200 144.300 ;
        RECT 560.400 143.400 562.200 155.400 ;
        RECT 578.400 149.400 580.200 155.400 ;
        RECT 578.700 149.100 580.200 149.400 ;
        RECT 584.400 149.400 586.200 155.400 ;
        RECT 598.800 149.400 600.600 155.400 ;
        RECT 619.800 149.400 621.600 155.400 ;
        RECT 640.800 149.400 642.600 155.400 ;
        RECT 662.400 149.400 664.200 155.400 ;
        RECT 680.400 149.400 682.200 155.400 ;
        RECT 584.400 149.100 585.300 149.400 ;
        RECT 578.700 148.200 585.300 149.100 ;
        RECT 536.100 136.050 537.900 137.850 ;
        RECT 554.100 136.050 555.900 137.850 ;
        RECT 560.700 136.050 561.600 143.400 ;
        RECT 578.100 136.050 579.900 137.850 ;
        RECT 584.400 136.050 585.300 148.200 ;
        RECT 599.400 136.050 600.600 149.400 ;
        RECT 604.950 138.450 609.000 139.050 ;
        RECT 602.100 136.050 603.900 137.850 ;
        RECT 604.950 136.950 609.450 138.450 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 382.950 133.950 385.050 136.050 ;
        RECT 394.950 133.950 397.050 136.050 ;
        RECT 397.950 133.950 400.050 136.050 ;
        RECT 400.950 133.950 403.050 136.050 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 424.950 133.950 427.050 136.050 ;
        RECT 439.950 133.950 442.050 136.050 ;
        RECT 442.950 133.950 445.050 136.050 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 508.950 133.950 511.050 136.050 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 535.950 133.950 538.050 136.050 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 550.950 133.950 553.050 136.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 556.950 133.950 559.050 136.050 ;
        RECT 559.950 133.950 562.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 577.950 133.950 580.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 308.400 125.700 316.200 127.050 ;
        RECT 308.400 120.600 310.200 125.700 ;
        RECT 314.400 120.600 316.200 125.700 ;
        RECT 317.400 126.600 318.600 128.700 ;
        RECT 335.400 127.800 339.600 128.700 ;
        RECT 350.400 128.400 357.900 129.300 ;
        RECT 317.400 120.600 319.200 126.600 ;
        RECT 335.400 120.600 337.200 127.800 ;
        RECT 350.400 120.600 352.200 128.400 ;
        RECT 356.100 127.500 357.900 128.400 ;
        RECT 359.700 126.600 360.600 133.950 ;
        RECT 357.900 124.800 360.600 126.600 ;
        RECT 374.400 126.600 375.300 133.950 ;
        RECT 377.100 132.150 378.900 133.950 ;
        RECT 383.100 132.150 384.900 133.950 ;
        RECT 395.100 132.150 396.900 133.950 ;
        RECT 401.100 132.150 402.900 133.950 ;
        RECT 404.400 130.200 405.300 133.950 ;
        RECT 419.100 132.150 420.900 133.950 ;
        RECT 402.000 129.000 405.300 130.200 ;
        RECT 374.400 125.400 379.500 126.600 ;
        RECT 357.900 120.600 359.700 124.800 ;
        RECT 377.700 120.600 379.500 125.400 ;
        RECT 402.000 120.600 403.800 129.000 ;
        RECT 422.400 128.700 423.600 133.950 ;
        RECT 425.100 132.150 426.900 133.950 ;
        RECT 443.100 132.150 444.900 133.950 ;
        RECT 446.850 129.750 448.050 133.950 ;
        RECT 449.100 132.150 450.900 133.950 ;
        RECT 446.850 128.700 450.600 129.750 ;
        RECT 422.400 127.800 426.600 128.700 ;
        RECT 424.800 120.600 426.600 127.800 ;
        RECT 440.400 125.700 448.200 127.050 ;
        RECT 440.400 120.600 442.200 125.700 ;
        RECT 446.400 120.600 448.200 125.700 ;
        RECT 449.400 126.600 450.600 128.700 ;
        RECT 449.400 120.600 451.200 126.600 ;
        RECT 467.400 123.600 468.600 133.950 ;
        RECT 485.400 126.600 486.300 133.950 ;
        RECT 488.100 132.150 489.900 133.950 ;
        RECT 494.100 132.150 495.900 133.950 ;
        RECT 503.100 132.150 504.900 133.950 ;
        RECT 509.100 132.150 510.900 133.950 ;
        RECT 512.400 130.200 513.300 133.950 ;
        RECT 490.950 129.450 493.050 130.050 ;
        RECT 499.950 129.450 502.050 130.050 ;
        RECT 490.950 128.550 502.050 129.450 ;
        RECT 490.950 127.950 493.050 128.550 ;
        RECT 499.950 127.950 502.050 128.550 ;
        RECT 510.000 129.000 513.300 130.200 ;
        RECT 530.700 130.200 531.600 133.950 ;
        RECT 533.100 132.150 534.900 133.950 ;
        RECT 539.100 132.150 540.900 133.950 ;
        RECT 551.100 132.150 552.900 133.950 ;
        RECT 557.100 132.150 558.900 133.950 ;
        RECT 530.700 129.000 534.000 130.200 ;
        RECT 485.400 125.400 490.500 126.600 ;
        RECT 467.400 120.600 469.200 123.600 ;
        RECT 488.700 120.600 490.500 125.400 ;
        RECT 510.000 120.600 511.800 129.000 ;
        RECT 532.200 120.600 534.000 129.000 ;
        RECT 560.700 126.600 561.600 133.950 ;
        RECT 575.100 132.150 576.900 133.950 ;
        RECT 581.100 132.150 582.900 133.950 ;
        RECT 584.400 130.200 585.300 133.950 ;
        RECT 556.500 125.400 561.600 126.600 ;
        RECT 582.000 129.000 585.300 130.200 ;
        RECT 556.500 120.600 558.300 125.400 ;
        RECT 582.000 120.600 583.800 129.000 ;
        RECT 599.400 123.600 600.600 133.950 ;
        RECT 608.550 132.450 609.450 136.950 ;
        RECT 614.100 136.050 615.900 137.850 ;
        RECT 619.950 136.050 621.150 149.400 ;
        RECT 622.950 141.450 625.050 142.050 ;
        RECT 631.950 141.450 634.050 142.050 ;
        RECT 622.950 140.550 634.050 141.450 ;
        RECT 622.950 139.950 625.050 140.550 ;
        RECT 631.950 139.950 634.050 140.550 ;
        RECT 635.100 136.050 636.900 137.850 ;
        RECT 640.950 136.050 642.150 149.400 ;
        RECT 643.950 141.450 646.050 142.200 ;
        RECT 658.950 141.450 661.050 142.050 ;
        RECT 643.950 140.550 661.050 141.450 ;
        RECT 643.950 140.100 646.050 140.550 ;
        RECT 658.950 139.950 661.050 140.550 ;
        RECT 659.100 136.050 660.900 137.850 ;
        RECT 662.400 136.050 663.600 149.400 ;
        RECT 680.700 149.100 682.200 149.400 ;
        RECT 686.400 149.400 688.200 155.400 ;
        RECT 704.400 149.400 706.200 155.400 ;
        RECT 727.800 149.400 729.600 155.400 ;
        RECT 746.400 149.400 748.200 155.400 ;
        RECT 770.400 149.400 772.200 155.400 ;
        RECT 686.400 149.100 687.300 149.400 ;
        RECT 680.700 148.200 687.300 149.100 ;
        RECT 680.100 136.050 681.900 137.850 ;
        RECT 686.400 136.050 687.300 148.200 ;
        RECT 704.400 136.050 705.600 149.400 ;
        RECT 722.100 136.050 723.900 137.850 ;
        RECT 727.950 136.050 729.150 149.400 ;
        RECT 746.400 136.050 747.600 149.400 ;
        RECT 757.950 144.450 760.050 145.050 ;
        RECT 763.950 144.450 766.050 145.050 ;
        RECT 757.950 143.550 766.050 144.450 ;
        RECT 757.950 142.950 760.050 143.550 ;
        RECT 763.950 142.950 766.050 143.550 ;
        RECT 762.000 138.450 766.050 139.050 ;
        RECT 761.550 136.950 766.050 138.450 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 634.950 133.950 637.050 136.050 ;
        RECT 637.950 133.950 640.050 136.050 ;
        RECT 640.950 133.950 643.050 136.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 658.950 133.950 661.050 136.050 ;
        RECT 661.950 133.950 664.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 679.950 133.950 682.050 136.050 ;
        RECT 682.950 133.950 685.050 136.050 ;
        RECT 685.950 133.950 688.050 136.050 ;
        RECT 700.950 133.950 703.050 136.050 ;
        RECT 703.950 133.950 706.050 136.050 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 724.950 133.950 727.050 136.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 742.950 133.950 745.050 136.050 ;
        RECT 745.950 133.950 748.050 136.050 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 608.550 132.000 612.450 132.450 ;
        RECT 617.100 132.150 618.900 133.950 ;
        RECT 608.550 131.550 613.050 132.000 ;
        RECT 610.950 127.950 613.050 131.550 ;
        RECT 620.850 129.750 622.050 133.950 ;
        RECT 623.100 132.150 624.900 133.950 ;
        RECT 638.100 132.150 639.900 133.950 ;
        RECT 641.850 129.750 643.050 133.950 ;
        RECT 644.100 132.150 645.900 133.950 ;
        RECT 620.850 128.700 624.600 129.750 ;
        RECT 641.850 128.700 645.600 129.750 ;
        RECT 598.800 120.600 600.600 123.600 ;
        RECT 614.400 125.700 622.200 127.050 ;
        RECT 614.400 120.600 616.200 125.700 ;
        RECT 620.400 120.600 622.200 125.700 ;
        RECT 623.400 126.600 624.600 128.700 ;
        RECT 623.400 120.600 625.200 126.600 ;
        RECT 635.400 125.700 643.200 127.050 ;
        RECT 635.400 120.600 637.200 125.700 ;
        RECT 641.400 120.600 643.200 125.700 ;
        RECT 644.400 126.600 645.600 128.700 ;
        RECT 644.400 120.600 646.200 126.600 ;
        RECT 662.400 123.600 663.600 133.950 ;
        RECT 677.100 132.150 678.900 133.950 ;
        RECT 683.100 132.150 684.900 133.950 ;
        RECT 686.400 130.200 687.300 133.950 ;
        RECT 701.100 132.150 702.900 133.950 ;
        RECT 684.000 129.000 687.300 130.200 ;
        RECT 662.400 120.600 664.200 123.600 ;
        RECT 684.000 120.600 685.800 129.000 ;
        RECT 704.400 128.700 705.600 133.950 ;
        RECT 707.100 132.150 708.900 133.950 ;
        RECT 725.100 132.150 726.900 133.950 ;
        RECT 728.850 129.750 730.050 133.950 ;
        RECT 731.100 132.150 732.900 133.950 ;
        RECT 743.100 132.150 744.900 133.950 ;
        RECT 728.850 128.700 732.600 129.750 ;
        RECT 704.400 127.800 708.600 128.700 ;
        RECT 706.800 120.600 708.600 127.800 ;
        RECT 722.400 125.700 730.200 127.050 ;
        RECT 722.400 120.600 724.200 125.700 ;
        RECT 728.400 120.600 730.200 125.700 ;
        RECT 731.400 126.600 732.600 128.700 ;
        RECT 746.400 128.700 747.600 133.950 ;
        RECT 749.100 132.150 750.900 133.950 ;
        RECT 761.550 133.050 762.450 136.950 ;
        RECT 770.850 136.050 772.050 149.400 ;
        RECT 788.400 144.300 790.200 155.400 ;
        RECT 794.400 144.300 796.200 155.400 ;
        RECT 788.400 143.400 796.200 144.300 ;
        RECT 797.400 143.400 799.200 155.400 ;
        RECT 812.400 149.400 814.200 155.400 ;
        RECT 836.400 149.400 838.200 155.400 ;
        RECT 783.000 138.450 787.050 139.050 ;
        RECT 776.100 136.050 777.900 137.850 ;
        RECT 782.550 136.950 787.050 138.450 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 761.550 131.550 766.050 133.050 ;
        RECT 767.100 132.150 768.900 133.950 ;
        RECT 762.000 130.950 766.050 131.550 ;
        RECT 769.950 129.750 771.150 133.950 ;
        RECT 773.100 132.150 774.900 133.950 ;
        RECT 782.550 133.050 783.450 136.950 ;
        RECT 791.100 136.050 792.900 137.850 ;
        RECT 797.700 136.050 798.600 143.400 ;
        RECT 812.400 136.050 813.600 149.400 ;
        RECT 817.950 138.450 822.000 139.050 ;
        RECT 817.950 136.950 822.450 138.450 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 778.950 131.550 783.450 133.050 ;
        RECT 788.100 132.150 789.900 133.950 ;
        RECT 794.100 132.150 795.900 133.950 ;
        RECT 778.950 130.950 783.000 131.550 ;
        RECT 767.400 128.700 771.150 129.750 ;
        RECT 746.400 127.800 750.600 128.700 ;
        RECT 731.400 120.600 733.200 126.600 ;
        RECT 748.800 120.600 750.600 127.800 ;
        RECT 767.400 126.600 768.600 128.700 ;
        RECT 766.800 120.600 768.600 126.600 ;
        RECT 769.800 125.700 777.600 127.050 ;
        RECT 797.700 126.600 798.600 133.950 ;
        RECT 809.100 132.150 810.900 133.950 ;
        RECT 812.400 128.700 813.600 133.950 ;
        RECT 815.100 132.150 816.900 133.950 ;
        RECT 821.550 133.050 822.450 136.950 ;
        RECT 836.850 136.050 838.050 149.400 ;
        RECT 857.400 143.400 859.200 155.400 ;
        RECT 847.950 141.450 850.050 142.050 ;
        RECT 853.950 141.450 856.050 142.200 ;
        RECT 847.950 140.550 856.050 141.450 ;
        RECT 847.950 139.950 850.050 140.550 ;
        RECT 853.950 140.100 856.050 140.550 ;
        RECT 842.100 136.050 843.900 137.850 ;
        RECT 857.700 136.050 858.750 143.400 ;
        RECT 880.800 142.500 882.600 155.400 ;
        RECT 886.800 142.500 888.600 155.400 ;
        RECT 892.800 142.500 894.600 155.400 ;
        RECT 898.800 142.500 900.600 155.400 ;
        RECT 879.900 141.300 882.600 142.500 ;
        RECT 884.700 141.300 888.600 142.500 ;
        RECT 890.700 141.300 894.600 142.500 ;
        RECT 896.700 141.300 900.600 142.500 ;
        RECT 879.900 136.050 880.800 141.300 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 853.950 133.950 856.050 136.050 ;
        RECT 857.700 133.950 862.050 136.050 ;
        RECT 877.950 133.950 880.800 136.050 ;
        RECT 817.950 131.550 822.450 133.050 ;
        RECT 833.100 132.150 834.900 133.950 ;
        RECT 817.950 130.950 822.000 131.550 ;
        RECT 835.950 129.750 837.150 133.950 ;
        RECT 839.100 132.150 840.900 133.950 ;
        RECT 854.100 132.150 855.900 133.950 ;
        RECT 833.400 128.700 837.150 129.750 ;
        RECT 812.400 127.800 816.600 128.700 ;
        RECT 769.800 120.600 771.600 125.700 ;
        RECT 775.800 120.600 777.600 125.700 ;
        RECT 793.500 125.400 798.600 126.600 ;
        RECT 793.500 120.600 795.300 125.400 ;
        RECT 814.800 120.600 816.600 127.800 ;
        RECT 833.400 126.600 834.600 128.700 ;
        RECT 832.800 120.600 834.600 126.600 ;
        RECT 835.800 125.700 843.600 127.050 ;
        RECT 857.700 126.600 858.750 133.950 ;
        RECT 879.900 128.700 880.800 133.950 ;
        RECT 881.700 130.800 883.500 131.400 ;
        RECT 884.700 130.800 885.900 141.300 ;
        RECT 881.700 129.600 885.900 130.800 ;
        RECT 887.700 130.800 889.500 131.400 ;
        RECT 890.700 130.800 891.900 141.300 ;
        RECT 887.700 129.600 891.900 130.800 ;
        RECT 893.700 130.800 895.500 131.400 ;
        RECT 896.700 130.800 897.900 141.300 ;
        RECT 898.950 133.950 901.050 136.050 ;
        RECT 899.100 132.150 900.900 133.950 ;
        RECT 893.700 129.600 897.900 130.800 ;
        RECT 884.700 128.700 885.900 129.600 ;
        RECT 890.700 128.700 891.900 129.600 ;
        RECT 896.700 128.700 897.900 129.600 ;
        RECT 879.900 127.500 882.600 128.700 ;
        RECT 884.700 127.500 888.600 128.700 ;
        RECT 890.700 127.500 894.600 128.700 ;
        RECT 896.700 127.500 900.600 128.700 ;
        RECT 835.800 120.600 837.600 125.700 ;
        RECT 841.800 120.600 843.600 125.700 ;
        RECT 857.400 120.600 859.200 126.600 ;
        RECT 880.800 120.600 882.600 127.500 ;
        RECT 886.800 120.600 888.600 127.500 ;
        RECT 892.800 120.600 894.600 127.500 ;
        RECT 898.800 120.600 900.600 127.500 ;
        RECT 13.800 110.400 15.600 116.400 ;
        RECT 14.400 108.300 15.600 110.400 ;
        RECT 16.800 111.300 18.600 116.400 ;
        RECT 22.800 111.300 24.600 116.400 ;
        RECT 16.800 109.950 24.600 111.300 ;
        RECT 14.400 107.250 18.150 108.300 ;
        RECT 40.200 108.000 42.000 116.400 ;
        RECT 59.400 111.300 61.200 116.400 ;
        RECT 65.400 111.300 67.200 116.400 ;
        RECT 59.400 109.950 67.200 111.300 ;
        RECT 68.400 110.400 70.200 116.400 ;
        RECT 68.400 108.300 69.600 110.400 ;
        RECT 14.100 103.050 15.900 104.850 ;
        RECT 16.950 103.050 18.150 107.250 ;
        RECT 38.700 106.800 42.000 108.000 ;
        RECT 65.850 107.250 69.600 108.300 ;
        RECT 90.000 108.000 91.800 116.400 ;
        RECT 109.800 110.400 111.600 116.400 ;
        RECT 110.400 108.300 111.600 110.400 ;
        RECT 112.800 111.300 114.600 116.400 ;
        RECT 118.800 111.300 120.600 116.400 ;
        RECT 137.700 111.600 139.500 116.400 ;
        RECT 112.800 109.950 120.600 111.300 ;
        RECT 134.400 110.400 139.500 111.600 ;
        RECT 20.100 103.050 21.900 104.850 ;
        RECT 38.700 103.050 39.600 106.800 ;
        RECT 41.100 103.050 42.900 104.850 ;
        RECT 47.100 103.050 48.900 104.850 ;
        RECT 62.100 103.050 63.900 104.850 ;
        RECT 65.850 103.050 67.050 107.250 ;
        RECT 90.000 106.800 93.300 108.000 ;
        RECT 110.400 107.250 114.150 108.300 ;
        RECT 68.100 103.050 69.900 104.850 ;
        RECT 83.100 103.050 84.900 104.850 ;
        RECT 89.100 103.050 90.900 104.850 ;
        RECT 92.400 103.050 93.300 106.800 ;
        RECT 110.100 103.050 111.900 104.850 ;
        RECT 112.950 103.050 114.150 107.250 ;
        RECT 116.100 103.050 117.900 104.850 ;
        RECT 134.400 103.050 135.300 110.400 ;
        RECT 162.000 108.000 163.800 116.400 ;
        RECT 181.200 108.000 183.000 116.400 ;
        RECT 205.500 111.600 207.300 116.400 ;
        RECT 230.700 111.600 232.500 116.400 ;
        RECT 205.500 110.400 210.600 111.600 ;
        RECT 162.000 106.800 165.300 108.000 ;
        RECT 137.100 103.050 138.900 104.850 ;
        RECT 143.100 103.050 144.900 104.850 ;
        RECT 155.100 103.050 156.900 104.850 ;
        RECT 161.100 103.050 162.900 104.850 ;
        RECT 164.400 103.050 165.300 106.800 ;
        RECT 179.700 106.800 183.000 108.000 ;
        RECT 179.700 103.050 180.600 106.800 ;
        RECT 190.950 105.450 195.000 106.050 ;
        RECT 182.100 103.050 183.900 104.850 ;
        RECT 188.100 103.050 189.900 104.850 ;
        RECT 190.950 103.950 195.450 105.450 ;
        RECT 13.950 100.950 16.050 103.050 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 22.950 100.950 25.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 136.950 100.950 139.050 103.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 154.950 100.950 157.050 103.050 ;
        RECT 157.950 100.950 160.050 103.050 ;
        RECT 160.950 100.950 163.050 103.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 17.850 87.600 19.050 100.950 ;
        RECT 23.100 99.150 24.900 100.950 ;
        RECT 38.700 88.800 39.600 100.950 ;
        RECT 44.100 99.150 45.900 100.950 ;
        RECT 59.100 99.150 60.900 100.950 ;
        RECT 38.700 87.900 45.300 88.800 ;
        RECT 38.700 87.600 39.600 87.900 ;
        RECT 17.400 81.600 19.200 87.600 ;
        RECT 37.800 81.600 39.600 87.600 ;
        RECT 43.800 87.600 45.300 87.900 ;
        RECT 64.950 87.600 66.150 100.950 ;
        RECT 86.100 99.150 87.900 100.950 ;
        RECT 92.400 88.800 93.300 100.950 ;
        RECT 86.700 87.900 93.300 88.800 ;
        RECT 86.700 87.600 88.200 87.900 ;
        RECT 43.800 81.600 45.600 87.600 ;
        RECT 64.800 81.600 66.600 87.600 ;
        RECT 86.400 81.600 88.200 87.600 ;
        RECT 92.400 87.600 93.300 87.900 ;
        RECT 113.850 87.600 115.050 100.950 ;
        RECT 119.100 99.150 120.900 100.950 ;
        RECT 134.400 93.600 135.300 100.950 ;
        RECT 140.100 99.150 141.900 100.950 ;
        RECT 158.100 99.150 159.900 100.950 ;
        RECT 92.400 81.600 94.200 87.600 ;
        RECT 113.400 81.600 115.200 87.600 ;
        RECT 133.800 81.600 135.600 93.600 ;
        RECT 136.800 92.700 144.600 93.600 ;
        RECT 136.800 81.600 138.600 92.700 ;
        RECT 142.800 81.600 144.600 92.700 ;
        RECT 164.400 88.800 165.300 100.950 ;
        RECT 158.700 87.900 165.300 88.800 ;
        RECT 158.700 87.600 160.200 87.900 ;
        RECT 158.400 81.600 160.200 87.600 ;
        RECT 164.400 87.600 165.300 87.900 ;
        RECT 179.700 88.800 180.600 100.950 ;
        RECT 185.100 99.150 186.900 100.950 ;
        RECT 194.550 100.050 195.450 103.950 ;
        RECT 200.100 103.050 201.900 104.850 ;
        RECT 206.100 103.050 207.900 104.850 ;
        RECT 209.700 103.050 210.600 110.400 ;
        RECT 227.400 110.400 232.500 111.600 ;
        RECT 227.400 103.050 228.300 110.400 ;
        RECT 252.000 108.000 253.800 116.400 ;
        RECT 272.700 111.600 274.500 116.400 ;
        RECT 269.400 110.400 274.500 111.600 ;
        RECT 289.800 110.400 291.600 116.400 ;
        RECT 252.000 106.800 255.300 108.000 ;
        RECT 230.100 103.050 231.900 104.850 ;
        RECT 236.100 103.050 237.900 104.850 ;
        RECT 245.100 103.050 246.900 104.850 ;
        RECT 251.100 103.050 252.900 104.850 ;
        RECT 254.400 103.050 255.300 106.800 ;
        RECT 256.950 105.450 261.000 106.050 ;
        RECT 256.950 103.950 261.450 105.450 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 226.950 100.950 229.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 194.550 98.550 199.050 100.050 ;
        RECT 203.100 99.150 204.900 100.950 ;
        RECT 195.000 97.950 199.050 98.550 ;
        RECT 209.700 93.600 210.600 100.950 ;
        RECT 227.400 93.600 228.300 100.950 ;
        RECT 233.100 99.150 234.900 100.950 ;
        RECT 248.100 99.150 249.900 100.950 ;
        RECT 229.950 96.450 232.050 97.050 ;
        RECT 250.950 96.450 253.050 97.050 ;
        RECT 229.950 95.550 253.050 96.450 ;
        RECT 229.950 94.950 232.050 95.550 ;
        RECT 250.950 94.950 253.050 95.550 ;
        RECT 200.400 92.700 208.200 93.600 ;
        RECT 179.700 87.900 186.300 88.800 ;
        RECT 179.700 87.600 180.600 87.900 ;
        RECT 164.400 81.600 166.200 87.600 ;
        RECT 178.800 81.600 180.600 87.600 ;
        RECT 184.800 87.600 186.300 87.900 ;
        RECT 184.800 81.600 186.600 87.600 ;
        RECT 200.400 81.600 202.200 92.700 ;
        RECT 206.400 81.600 208.200 92.700 ;
        RECT 209.400 81.600 211.200 93.600 ;
        RECT 226.800 81.600 228.600 93.600 ;
        RECT 229.800 92.700 237.600 93.600 ;
        RECT 229.800 81.600 231.600 92.700 ;
        RECT 235.800 81.600 237.600 92.700 ;
        RECT 254.400 88.800 255.300 100.950 ;
        RECT 260.550 99.450 261.450 103.950 ;
        RECT 269.400 103.050 270.300 110.400 ;
        RECT 277.950 108.450 280.050 109.050 ;
        RECT 283.950 108.450 286.050 109.050 ;
        RECT 277.950 107.550 286.050 108.450 ;
        RECT 277.950 106.950 280.050 107.550 ;
        RECT 283.950 106.950 286.050 107.550 ;
        RECT 290.400 108.300 291.600 110.400 ;
        RECT 292.800 111.300 294.600 116.400 ;
        RECT 298.800 111.300 300.600 116.400 ;
        RECT 292.800 109.950 300.600 111.300 ;
        RECT 313.800 110.400 315.600 116.400 ;
        RECT 314.400 108.300 315.600 110.400 ;
        RECT 316.800 111.300 318.600 116.400 ;
        RECT 322.800 111.300 324.600 116.400 ;
        RECT 316.800 109.950 324.600 111.300 ;
        RECT 290.400 107.250 294.150 108.300 ;
        RECT 314.400 107.250 318.150 108.300 ;
        RECT 340.200 108.000 342.000 116.400 ;
        RECT 359.400 111.300 361.200 116.400 ;
        RECT 365.400 111.300 367.200 116.400 ;
        RECT 359.400 109.950 367.200 111.300 ;
        RECT 368.400 110.400 370.200 116.400 ;
        RECT 368.400 108.300 369.600 110.400 ;
        RECT 272.100 103.050 273.900 104.850 ;
        RECT 278.100 103.050 279.900 104.850 ;
        RECT 290.100 103.050 291.900 104.850 ;
        RECT 292.950 103.050 294.150 107.250 ;
        RECT 310.950 105.450 313.050 106.050 ;
        RECT 296.100 103.050 297.900 104.850 ;
        RECT 305.550 104.550 313.050 105.450 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 274.950 100.950 277.050 103.050 ;
        RECT 277.950 100.950 280.050 103.050 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 295.950 100.950 298.050 103.050 ;
        RECT 298.950 100.950 301.050 103.050 ;
        RECT 260.550 99.000 267.450 99.450 ;
        RECT 260.550 98.550 268.050 99.000 ;
        RECT 265.950 94.950 268.050 98.550 ;
        RECT 269.400 93.600 270.300 100.950 ;
        RECT 275.100 99.150 276.900 100.950 ;
        RECT 248.700 87.900 255.300 88.800 ;
        RECT 248.700 87.600 250.200 87.900 ;
        RECT 248.400 81.600 250.200 87.600 ;
        RECT 254.400 87.600 255.300 87.900 ;
        RECT 254.400 81.600 256.200 87.600 ;
        RECT 268.800 81.600 270.600 93.600 ;
        RECT 271.800 92.700 279.600 93.600 ;
        RECT 271.800 81.600 273.600 92.700 ;
        RECT 277.800 81.600 279.600 92.700 ;
        RECT 293.850 87.600 295.050 100.950 ;
        RECT 299.100 99.150 300.900 100.950 ;
        RECT 305.550 100.050 306.450 104.550 ;
        RECT 310.950 103.950 313.050 104.550 ;
        RECT 314.100 103.050 315.900 104.850 ;
        RECT 316.950 103.050 318.150 107.250 ;
        RECT 338.700 106.800 342.000 108.000 ;
        RECT 365.850 107.250 369.600 108.300 ;
        RECT 387.000 108.000 388.800 116.400 ;
        RECT 411.000 108.000 412.800 116.400 ;
        RECT 428.400 108.600 430.200 116.400 ;
        RECT 435.900 112.200 437.700 116.400 ;
        RECT 435.900 110.400 438.600 112.200 ;
        RECT 434.100 108.600 435.900 109.500 ;
        RECT 333.000 105.450 337.050 106.050 ;
        RECT 320.100 103.050 321.900 104.850 ;
        RECT 332.550 103.950 337.050 105.450 ;
        RECT 313.950 100.950 316.050 103.050 ;
        RECT 316.950 100.950 319.050 103.050 ;
        RECT 319.950 100.950 322.050 103.050 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 332.550 102.450 333.450 103.950 ;
        RECT 338.700 103.050 339.600 106.800 ;
        RECT 341.100 103.050 342.900 104.850 ;
        RECT 347.100 103.050 348.900 104.850 ;
        RECT 362.100 103.050 363.900 104.850 ;
        RECT 365.850 103.050 367.050 107.250 ;
        RECT 387.000 106.800 390.300 108.000 ;
        RECT 411.000 106.800 414.300 108.000 ;
        RECT 428.400 107.700 435.900 108.600 ;
        RECT 368.100 103.050 369.900 104.850 ;
        RECT 380.100 103.050 381.900 104.850 ;
        RECT 386.100 103.050 387.900 104.850 ;
        RECT 389.400 103.050 390.300 106.800 ;
        RECT 404.100 103.050 405.900 104.850 ;
        RECT 410.100 103.050 411.900 104.850 ;
        RECT 413.400 103.050 414.300 106.800 ;
        RECT 428.100 103.050 429.900 104.850 ;
        RECT 329.550 101.550 333.450 102.450 ;
        RECT 301.950 98.550 306.450 100.050 ;
        RECT 301.950 97.950 306.000 98.550 ;
        RECT 317.850 87.600 319.050 100.950 ;
        RECT 323.100 99.150 324.900 100.950 ;
        RECT 329.550 100.050 330.450 101.550 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 340.950 100.950 343.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 358.950 100.950 361.050 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 403.950 100.950 406.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 325.950 98.550 330.450 100.050 ;
        RECT 325.950 97.950 330.000 98.550 ;
        RECT 338.700 88.800 339.600 100.950 ;
        RECT 344.100 99.150 345.900 100.950 ;
        RECT 359.100 99.150 360.900 100.950 ;
        RECT 338.700 87.900 345.300 88.800 ;
        RECT 338.700 87.600 339.600 87.900 ;
        RECT 293.400 81.600 295.200 87.600 ;
        RECT 317.400 81.600 319.200 87.600 ;
        RECT 337.800 81.600 339.600 87.600 ;
        RECT 343.800 87.600 345.300 87.900 ;
        RECT 364.950 87.600 366.150 100.950 ;
        RECT 383.100 99.150 384.900 100.950 ;
        RECT 389.400 88.800 390.300 100.950 ;
        RECT 407.100 99.150 408.900 100.950 ;
        RECT 413.400 88.800 414.300 100.950 ;
        RECT 383.700 87.900 390.300 88.800 ;
        RECT 383.700 87.600 385.200 87.900 ;
        RECT 343.800 81.600 345.600 87.600 ;
        RECT 364.800 81.600 366.600 87.600 ;
        RECT 383.400 81.600 385.200 87.600 ;
        RECT 389.400 87.600 390.300 87.900 ;
        RECT 407.700 87.900 414.300 88.800 ;
        RECT 407.700 87.600 409.200 87.900 ;
        RECT 389.400 81.600 391.200 87.600 ;
        RECT 407.400 81.600 409.200 87.600 ;
        RECT 413.400 87.600 414.300 87.900 ;
        RECT 431.400 87.600 432.300 107.700 ;
        RECT 437.700 103.050 438.600 110.400 ;
        RECT 462.000 110.400 463.800 116.400 ;
        RECT 485.700 111.600 487.500 116.400 ;
        RECT 482.400 110.400 487.500 111.600 ;
        RECT 445.950 108.450 448.050 109.050 ;
        RECT 457.950 108.450 460.050 109.050 ;
        RECT 445.950 107.550 460.050 108.450 ;
        RECT 445.950 106.950 448.050 107.550 ;
        RECT 457.950 106.950 460.050 107.550 ;
        RECT 442.950 105.450 445.050 106.050 ;
        RECT 451.950 105.450 454.050 106.050 ;
        RECT 442.950 104.550 454.050 105.450 ;
        RECT 442.950 103.950 445.050 104.550 ;
        RECT 451.950 103.950 454.050 104.550 ;
        RECT 455.100 103.050 456.900 104.850 ;
        RECT 462.000 103.050 463.050 110.400 ;
        RECT 467.100 103.050 468.900 104.850 ;
        RECT 475.950 103.950 478.050 106.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 463.950 100.950 466.050 103.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 434.100 99.150 435.900 100.950 ;
        RECT 437.700 93.600 438.600 100.950 ;
        RECT 458.100 99.150 459.900 100.950 ;
        RECT 462.000 95.400 462.900 100.950 ;
        RECT 464.100 99.150 465.900 100.950 ;
        RECT 472.950 100.050 475.050 103.050 ;
        RECT 476.550 100.050 477.450 103.950 ;
        RECT 482.400 103.050 483.300 110.400 ;
        RECT 507.000 108.000 508.800 116.400 ;
        RECT 523.800 110.400 525.600 116.400 ;
        RECT 524.400 108.300 525.600 110.400 ;
        RECT 526.800 111.300 528.600 116.400 ;
        RECT 532.800 111.300 534.600 116.400 ;
        RECT 526.800 109.950 534.600 111.300 ;
        RECT 545.400 111.300 547.200 116.400 ;
        RECT 551.400 111.300 553.200 116.400 ;
        RECT 545.400 109.950 553.200 111.300 ;
        RECT 554.400 110.400 556.200 116.400 ;
        RECT 554.400 108.300 555.600 110.400 ;
        RECT 507.000 106.800 510.300 108.000 ;
        RECT 524.400 107.250 528.150 108.300 ;
        RECT 485.100 103.050 486.900 104.850 ;
        RECT 491.100 103.050 492.900 104.850 ;
        RECT 500.100 103.050 501.900 104.850 ;
        RECT 506.100 103.050 507.900 104.850 ;
        RECT 509.400 103.050 510.300 106.800 ;
        RECT 524.100 103.050 525.900 104.850 ;
        RECT 526.950 103.050 528.150 107.250 ;
        RECT 551.850 107.250 555.600 108.300 ;
        RECT 574.200 108.000 576.000 116.400 ;
        RECT 598.500 111.600 600.300 116.400 ;
        RECT 628.800 113.400 630.600 116.400 ;
        RECT 634.800 113.400 636.600 116.400 ;
        RECT 628.800 112.500 629.850 113.400 ;
        RECT 634.800 112.500 635.850 113.400 ;
        RECT 625.050 111.600 635.850 112.500 ;
        RECT 598.500 110.400 603.600 111.600 ;
        RECT 530.100 103.050 531.900 104.850 ;
        RECT 548.100 103.050 549.900 104.850 ;
        RECT 551.850 103.050 553.050 107.250 ;
        RECT 572.700 106.800 576.000 108.000 ;
        RECT 586.950 108.450 589.050 109.050 ;
        RECT 595.950 108.450 598.050 109.050 ;
        RECT 586.950 107.550 598.050 108.450 ;
        RECT 586.950 106.950 589.050 107.550 ;
        RECT 595.950 106.950 598.050 107.550 ;
        RECT 554.100 103.050 555.900 104.850 ;
        RECT 572.700 103.050 573.600 106.800 ;
        RECT 575.100 103.050 576.900 104.850 ;
        RECT 581.100 103.050 582.900 104.850 ;
        RECT 593.100 103.050 594.900 104.850 ;
        RECT 599.100 103.050 600.900 104.850 ;
        RECT 602.700 103.050 603.600 110.400 ;
        RECT 625.050 103.200 626.250 111.600 ;
        RECT 653.400 111.300 655.200 116.400 ;
        RECT 659.400 111.300 661.200 116.400 ;
        RECT 653.400 109.950 661.200 111.300 ;
        RECT 662.400 110.400 664.200 116.400 ;
        RECT 677.400 113.400 679.200 116.400 ;
        RECT 637.950 108.450 640.050 109.050 ;
        RECT 649.950 108.450 652.050 109.050 ;
        RECT 637.950 107.550 652.050 108.450 ;
        RECT 662.400 108.300 663.600 110.400 ;
        RECT 637.950 106.950 640.050 107.550 ;
        RECT 649.950 106.950 652.050 107.550 ;
        RECT 659.850 107.250 663.600 108.300 ;
        RECT 632.100 103.200 633.900 105.000 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 499.950 100.950 502.050 103.050 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 523.950 100.950 526.050 103.050 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 544.950 100.950 547.050 103.050 ;
        RECT 547.950 100.950 550.050 103.050 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 565.950 100.950 568.050 103.050 ;
        RECT 571.950 100.950 574.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 598.950 100.950 601.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 622.950 101.100 626.250 103.200 ;
        RECT 628.950 101.100 631.050 103.200 ;
        RECT 631.950 101.100 634.050 103.200 ;
        RECT 637.950 101.100 640.050 103.200 ;
        RECT 656.100 103.050 657.900 104.850 ;
        RECT 659.850 103.050 661.050 107.250 ;
        RECT 662.100 103.050 663.900 104.850 ;
        RECT 677.400 103.050 678.600 113.400 ;
        RECT 697.800 109.200 699.600 116.400 ;
        RECT 719.700 111.600 721.500 116.400 ;
        RECT 695.400 108.300 699.600 109.200 ;
        RECT 716.400 110.400 721.500 111.600 ;
        RECT 742.200 110.400 744.000 116.400 ;
        RECT 767.700 111.600 769.500 116.400 ;
        RECT 692.100 103.050 693.900 104.850 ;
        RECT 695.400 103.050 696.600 108.300 ;
        RECT 698.100 103.050 699.900 104.850 ;
        RECT 716.400 103.050 717.300 110.400 ;
        RECT 735.000 108.450 739.050 109.050 ;
        RECT 734.550 106.950 739.050 108.450 ;
        RECT 734.550 105.450 735.450 106.950 ;
        RECT 719.100 103.050 720.900 104.850 ;
        RECT 725.100 103.050 726.900 104.850 ;
        RECT 731.550 104.550 735.450 105.450 ;
        RECT 469.950 99.000 475.050 100.050 ;
        RECT 469.950 98.550 474.450 99.000 ;
        RECT 469.950 97.950 474.000 98.550 ;
        RECT 475.950 97.950 478.050 100.050 ;
        RECT 457.800 94.500 462.900 95.400 ;
        RECT 413.400 81.600 415.200 87.600 ;
        RECT 431.400 81.600 433.200 87.600 ;
        RECT 437.400 81.600 439.200 93.600 ;
        RECT 454.800 82.500 456.600 93.600 ;
        RECT 457.800 83.400 459.600 94.500 ;
        RECT 482.400 93.600 483.300 100.950 ;
        RECT 488.100 99.150 489.900 100.950 ;
        RECT 503.100 99.150 504.900 100.950 ;
        RECT 460.800 92.400 468.600 93.300 ;
        RECT 460.800 82.500 462.600 92.400 ;
        RECT 454.800 81.600 462.600 82.500 ;
        RECT 466.800 81.600 468.600 92.400 ;
        RECT 481.800 81.600 483.600 93.600 ;
        RECT 484.800 92.700 492.600 93.600 ;
        RECT 484.800 81.600 486.600 92.700 ;
        RECT 490.800 81.600 492.600 92.700 ;
        RECT 509.400 88.800 510.300 100.950 ;
        RECT 503.700 87.900 510.300 88.800 ;
        RECT 503.700 87.600 505.200 87.900 ;
        RECT 503.400 81.600 505.200 87.600 ;
        RECT 509.400 87.600 510.300 87.900 ;
        RECT 527.850 87.600 529.050 100.950 ;
        RECT 533.100 99.150 534.900 100.950 ;
        RECT 545.100 99.150 546.900 100.950 ;
        RECT 550.950 87.600 552.150 100.950 ;
        RECT 556.950 99.450 559.050 100.050 ;
        RECT 562.950 99.450 565.050 100.050 ;
        RECT 556.950 98.550 565.050 99.450 ;
        RECT 556.950 97.950 559.050 98.550 ;
        RECT 562.950 97.950 565.050 98.550 ;
        RECT 566.550 97.050 567.450 100.950 ;
        RECT 565.950 94.950 568.050 97.050 ;
        RECT 572.700 88.800 573.600 100.950 ;
        RECT 578.100 99.150 579.900 100.950 ;
        RECT 596.100 99.150 597.900 100.950 ;
        RECT 574.950 96.450 577.050 97.050 ;
        RECT 592.950 96.450 595.050 97.050 ;
        RECT 574.950 95.550 595.050 96.450 ;
        RECT 574.950 94.950 577.050 95.550 ;
        RECT 592.950 94.950 595.050 95.550 ;
        RECT 602.700 93.600 603.600 100.950 ;
        RECT 625.050 94.800 626.250 101.100 ;
        RECT 629.100 99.300 630.900 101.100 ;
        RECT 638.100 99.300 639.900 101.100 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 718.950 100.950 721.050 103.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 724.950 100.950 727.050 103.050 ;
        RECT 653.100 99.150 654.900 100.950 ;
        RECT 622.800 93.600 626.250 94.800 ;
        RECT 593.400 92.700 601.200 93.600 ;
        RECT 572.700 87.900 579.300 88.800 ;
        RECT 572.700 87.600 573.600 87.900 ;
        RECT 509.400 81.600 511.200 87.600 ;
        RECT 527.400 81.600 529.200 87.600 ;
        RECT 550.800 81.600 552.600 87.600 ;
        RECT 571.800 81.600 573.600 87.600 ;
        RECT 577.800 87.600 579.300 87.900 ;
        RECT 577.800 81.600 579.600 87.600 ;
        RECT 593.400 81.600 595.200 92.700 ;
        RECT 599.400 81.600 601.200 92.700 ;
        RECT 602.400 81.600 604.200 93.600 ;
        RECT 619.200 82.500 621.000 91.800 ;
        RECT 622.800 91.200 624.000 93.600 ;
        RECT 622.200 83.400 624.000 91.200 ;
        RECT 625.200 91.200 633.600 92.100 ;
        RECT 625.200 82.500 627.000 91.200 ;
        RECT 619.200 81.600 627.000 82.500 ;
        RECT 628.800 82.500 630.600 90.300 ;
        RECT 631.800 83.400 633.600 91.200 ;
        RECT 634.800 91.500 642.600 92.400 ;
        RECT 634.800 82.500 636.600 91.500 ;
        RECT 628.800 81.600 636.600 82.500 ;
        RECT 640.800 81.600 642.600 91.500 ;
        RECT 658.950 87.600 660.150 100.950 ;
        RECT 674.100 99.150 675.900 100.950 ;
        RECT 677.400 87.600 678.600 100.950 ;
        RECT 695.400 87.600 696.600 100.950 ;
        RECT 716.400 93.600 717.300 100.950 ;
        RECT 722.100 99.150 723.900 100.950 ;
        RECT 731.550 100.050 732.450 104.550 ;
        RECT 737.100 103.050 738.900 104.850 ;
        RECT 742.950 103.050 744.000 110.400 ;
        RECT 764.400 110.400 769.500 111.600 ;
        RECT 787.500 111.600 789.300 116.400 ;
        RECT 787.500 110.400 792.600 111.600 ;
        RECT 749.100 103.050 750.900 104.850 ;
        RECT 764.400 103.050 765.300 110.400 ;
        RECT 767.100 103.050 768.900 104.850 ;
        RECT 773.100 103.050 774.900 104.850 ;
        RECT 782.100 103.050 783.900 104.850 ;
        RECT 788.100 103.050 789.900 104.850 ;
        RECT 791.700 103.050 792.600 110.400 ;
        RECT 813.000 110.400 814.800 116.400 ;
        RECT 835.500 111.600 837.300 116.400 ;
        RECT 835.500 110.400 840.600 111.600 ;
        RECT 806.100 103.050 807.900 104.850 ;
        RECT 813.000 103.050 814.050 110.400 ;
        RECT 818.100 103.050 819.900 104.850 ;
        RECT 830.100 103.050 831.900 104.850 ;
        RECT 836.100 103.050 837.900 104.850 ;
        RECT 839.700 103.050 840.600 110.400 ;
        RECT 861.000 110.400 862.800 116.400 ;
        RECT 881.400 113.400 883.200 116.400 ;
        RECT 899.400 113.400 901.200 116.400 ;
        RECT 854.100 103.050 855.900 104.850 ;
        RECT 861.000 103.050 862.050 110.400 ;
        RECT 873.000 105.450 877.050 106.050 ;
        RECT 866.100 103.050 867.900 104.850 ;
        RECT 872.550 103.950 877.050 105.450 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 742.950 100.950 745.050 103.050 ;
        RECT 745.950 100.950 748.050 103.050 ;
        RECT 748.950 100.950 751.050 103.050 ;
        RECT 763.950 100.950 766.050 103.050 ;
        RECT 766.950 100.950 769.050 103.050 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 808.950 100.950 811.050 103.050 ;
        RECT 811.950 100.950 814.050 103.050 ;
        RECT 814.950 100.950 817.050 103.050 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 856.950 100.950 859.050 103.050 ;
        RECT 859.950 100.950 862.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 865.950 100.950 868.050 103.050 ;
        RECT 727.950 98.550 732.450 100.050 ;
        RECT 740.100 99.150 741.900 100.950 ;
        RECT 727.950 97.950 732.000 98.550 ;
        RECT 743.100 95.400 744.000 100.950 ;
        RECT 746.100 99.150 747.900 100.950 ;
        RECT 743.100 94.500 748.200 95.400 ;
        RECT 658.800 81.600 660.600 87.600 ;
        RECT 677.400 81.600 679.200 87.600 ;
        RECT 695.400 81.600 697.200 87.600 ;
        RECT 715.800 81.600 717.600 93.600 ;
        RECT 718.800 92.700 726.600 93.600 ;
        RECT 718.800 81.600 720.600 92.700 ;
        RECT 724.800 81.600 726.600 92.700 ;
        RECT 737.400 92.400 745.200 93.300 ;
        RECT 737.400 81.600 739.200 92.400 ;
        RECT 743.400 82.500 745.200 92.400 ;
        RECT 746.400 83.400 748.200 94.500 ;
        RECT 764.400 93.600 765.300 100.950 ;
        RECT 770.100 99.150 771.900 100.950 ;
        RECT 785.100 99.150 786.900 100.950 ;
        RECT 791.700 93.600 792.600 100.950 ;
        RECT 809.100 99.150 810.900 100.950 ;
        RECT 813.000 95.400 813.900 100.950 ;
        RECT 815.100 99.150 816.900 100.950 ;
        RECT 833.100 99.150 834.900 100.950 ;
        RECT 808.800 94.500 813.900 95.400 ;
        RECT 749.400 82.500 751.200 93.600 ;
        RECT 743.400 81.600 751.200 82.500 ;
        RECT 763.800 81.600 765.600 93.600 ;
        RECT 766.800 92.700 774.600 93.600 ;
        RECT 766.800 81.600 768.600 92.700 ;
        RECT 772.800 81.600 774.600 92.700 ;
        RECT 782.400 92.700 790.200 93.600 ;
        RECT 782.400 81.600 784.200 92.700 ;
        RECT 788.400 81.600 790.200 92.700 ;
        RECT 791.400 81.600 793.200 93.600 ;
        RECT 805.800 82.500 807.600 93.600 ;
        RECT 808.800 83.400 810.600 94.500 ;
        RECT 839.700 93.600 840.600 100.950 ;
        RECT 857.100 99.150 858.900 100.950 ;
        RECT 861.000 95.400 861.900 100.950 ;
        RECT 863.100 99.150 864.900 100.950 ;
        RECT 872.550 100.050 873.450 103.950 ;
        RECT 881.400 103.050 882.600 113.400 ;
        RECT 899.400 103.050 900.600 113.400 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 880.950 100.950 883.050 103.050 ;
        RECT 895.950 100.950 898.050 103.050 ;
        RECT 898.950 100.950 901.050 103.050 ;
        RECT 868.950 98.550 873.450 100.050 ;
        RECT 878.100 99.150 879.900 100.950 ;
        RECT 868.950 97.950 873.000 98.550 ;
        RECT 856.800 94.500 861.900 95.400 ;
        RECT 811.800 92.400 819.600 93.300 ;
        RECT 811.800 82.500 813.600 92.400 ;
        RECT 805.800 81.600 813.600 82.500 ;
        RECT 817.800 81.600 819.600 92.400 ;
        RECT 830.400 92.700 838.200 93.600 ;
        RECT 830.400 81.600 832.200 92.700 ;
        RECT 836.400 81.600 838.200 92.700 ;
        RECT 839.400 81.600 841.200 93.600 ;
        RECT 853.800 82.500 855.600 93.600 ;
        RECT 856.800 83.400 858.600 94.500 ;
        RECT 859.800 92.400 867.600 93.300 ;
        RECT 859.800 82.500 861.600 92.400 ;
        RECT 853.800 81.600 861.600 82.500 ;
        RECT 865.800 81.600 867.600 92.400 ;
        RECT 881.400 87.600 882.600 100.950 ;
        RECT 896.100 99.150 897.900 100.950 ;
        RECT 899.400 87.600 900.600 100.950 ;
        RECT 881.400 81.600 883.200 87.600 ;
        RECT 899.400 81.600 901.200 87.600 ;
        RECT 13.800 71.400 15.600 77.400 ;
        RECT 14.700 71.100 15.600 71.400 ;
        RECT 19.800 71.400 21.600 77.400 ;
        RECT 19.800 71.100 21.300 71.400 ;
        RECT 14.700 70.200 21.300 71.100 ;
        RECT 14.700 58.050 15.600 70.200 ;
        RECT 32.400 66.300 34.200 77.400 ;
        RECT 38.400 66.300 40.200 77.400 ;
        RECT 32.400 65.400 40.200 66.300 ;
        RECT 41.400 65.400 43.200 77.400 ;
        RECT 58.800 65.400 60.600 77.400 ;
        RECT 61.800 66.300 63.600 77.400 ;
        RECT 67.800 66.300 69.600 77.400 ;
        RECT 80.400 71.400 82.200 77.400 ;
        RECT 80.700 71.100 82.200 71.400 ;
        RECT 86.400 71.400 88.200 77.400 ;
        RECT 107.400 71.400 109.200 77.400 ;
        RECT 86.400 71.100 87.300 71.400 ;
        RECT 80.700 70.200 87.300 71.100 ;
        RECT 61.800 65.400 69.600 66.300 ;
        RECT 20.100 58.050 21.900 59.850 ;
        RECT 35.100 58.050 36.900 59.850 ;
        RECT 41.700 58.050 42.600 65.400 ;
        RECT 59.400 58.050 60.300 65.400 ;
        RECT 67.950 63.450 70.050 64.050 ;
        RECT 73.950 63.450 76.050 64.050 ;
        RECT 67.950 62.550 76.050 63.450 ;
        RECT 67.950 61.950 70.050 62.550 ;
        RECT 73.950 61.950 76.050 62.550 ;
        RECT 65.100 58.050 66.900 59.850 ;
        RECT 80.100 58.050 81.900 59.850 ;
        RECT 86.400 58.050 87.300 70.200 ;
        RECT 107.850 58.050 109.050 71.400 ;
        RECT 124.800 65.400 126.600 77.400 ;
        RECT 127.800 66.300 129.600 77.400 ;
        RECT 133.800 66.300 135.600 77.400 ;
        RECT 152.400 71.400 154.200 77.400 ;
        RECT 173.400 71.400 175.200 77.400 ;
        RECT 193.800 71.400 195.600 77.400 ;
        RECT 127.800 65.400 135.600 66.300 ;
        RECT 113.100 58.050 114.900 59.850 ;
        RECT 125.400 58.050 126.300 65.400 ;
        RECT 131.100 58.050 132.900 59.850 ;
        RECT 152.850 58.050 154.050 71.400 ;
        RECT 158.100 58.050 159.900 59.850 ;
        RECT 173.850 58.050 175.050 71.400 ;
        RECT 179.100 58.050 180.900 59.850 ;
        RECT 188.100 58.050 189.900 59.850 ;
        RECT 193.950 58.050 195.150 71.400 ;
        RECT 212.400 66.300 214.200 77.400 ;
        RECT 219.900 66.300 221.700 77.400 ;
        RECT 227.400 66.600 229.200 77.400 ;
        RECT 212.400 65.100 217.200 66.300 ;
        RECT 219.900 65.400 223.200 66.300 ;
        RECT 215.100 64.200 217.200 65.100 ;
        RECT 215.100 63.300 220.500 64.200 ;
        RECT 218.700 61.200 220.500 63.300 ;
        RECT 222.000 60.900 223.200 65.400 ;
        RECT 224.100 65.400 229.200 66.600 ;
        RECT 245.400 71.400 247.200 77.400 ;
        RECT 265.800 76.500 273.600 77.400 ;
        RECT 224.100 64.500 226.200 65.400 ;
        RECT 221.400 60.300 223.500 60.900 ;
        RECT 238.950 60.450 241.050 61.050 ;
        RECT 217.200 58.200 219.000 60.000 ;
        RECT 220.350 58.800 223.500 60.300 ;
        RECT 227.550 59.700 241.050 60.450 ;
        RECT 227.100 59.550 241.050 59.700 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 154.950 55.950 157.050 58.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 14.700 52.200 15.600 55.950 ;
        RECT 17.100 54.150 18.900 55.950 ;
        RECT 23.100 54.150 24.900 55.950 ;
        RECT 32.100 54.150 33.900 55.950 ;
        RECT 38.100 54.150 39.900 55.950 ;
        RECT 14.700 51.000 18.000 52.200 ;
        RECT 16.200 42.600 18.000 51.000 ;
        RECT 41.700 48.600 42.600 55.950 ;
        RECT 37.500 47.400 42.600 48.600 ;
        RECT 59.400 48.600 60.300 55.950 ;
        RECT 62.100 54.150 63.900 55.950 ;
        RECT 68.100 54.150 69.900 55.950 ;
        RECT 77.100 54.150 78.900 55.950 ;
        RECT 83.100 54.150 84.900 55.950 ;
        RECT 86.400 52.200 87.300 55.950 ;
        RECT 104.100 54.150 105.900 55.950 ;
        RECT 84.000 51.000 87.300 52.200 ;
        RECT 106.950 51.750 108.150 55.950 ;
        RECT 110.100 54.150 111.900 55.950 ;
        RECT 59.400 47.400 64.500 48.600 ;
        RECT 37.500 42.600 39.300 47.400 ;
        RECT 62.700 42.600 64.500 47.400 ;
        RECT 84.000 42.600 85.800 51.000 ;
        RECT 104.400 50.700 108.150 51.750 ;
        RECT 104.400 48.600 105.600 50.700 ;
        RECT 103.800 42.600 105.600 48.600 ;
        RECT 106.800 47.700 114.600 49.050 ;
        RECT 106.800 42.600 108.600 47.700 ;
        RECT 112.800 42.600 114.600 47.700 ;
        RECT 125.400 48.600 126.300 55.950 ;
        RECT 128.100 54.150 129.900 55.950 ;
        RECT 134.100 54.150 135.900 55.950 ;
        RECT 149.100 54.150 150.900 55.950 ;
        RECT 130.950 51.450 133.050 52.050 ;
        RECT 139.950 51.450 142.050 52.050 ;
        RECT 151.950 51.750 153.150 55.950 ;
        RECT 155.100 54.150 156.900 55.950 ;
        RECT 170.100 54.150 171.900 55.950 ;
        RECT 172.950 51.750 174.150 55.950 ;
        RECT 176.100 54.150 177.900 55.950 ;
        RECT 191.100 54.150 192.900 55.950 ;
        RECT 130.950 50.550 142.050 51.450 ;
        RECT 130.950 49.950 133.050 50.550 ;
        RECT 139.950 49.950 142.050 50.550 ;
        RECT 149.400 50.700 153.150 51.750 ;
        RECT 170.400 50.700 174.150 51.750 ;
        RECT 194.850 51.750 196.050 55.950 ;
        RECT 197.100 54.150 198.900 55.950 ;
        RECT 212.400 55.800 214.500 57.900 ;
        RECT 217.200 56.100 219.300 58.200 ;
        RECT 212.700 55.200 214.500 55.800 ;
        RECT 212.700 54.000 219.300 55.200 ;
        RECT 217.200 53.100 219.300 54.000 ;
        RECT 194.850 50.700 198.600 51.750 ;
        RECT 214.650 51.000 216.750 51.600 ;
        RECT 217.650 51.300 219.450 53.100 ;
        RECT 220.350 52.200 221.250 58.800 ;
        RECT 227.100 57.900 228.900 59.550 ;
        RECT 238.950 58.950 241.050 59.550 ;
        RECT 245.400 58.050 246.600 71.400 ;
        RECT 265.800 65.400 267.600 76.500 ;
        RECT 268.800 64.500 270.600 75.600 ;
        RECT 271.800 66.600 273.600 76.500 ;
        RECT 277.800 66.600 279.600 77.400 ;
        RECT 293.400 71.400 295.200 77.400 ;
        RECT 293.700 71.100 295.200 71.400 ;
        RECT 299.400 71.400 301.200 77.400 ;
        RECT 313.800 71.400 315.600 77.400 ;
        RECT 299.400 71.100 300.300 71.400 ;
        RECT 293.700 70.200 300.300 71.100 ;
        RECT 271.800 65.700 279.600 66.600 ;
        RECT 268.800 63.600 273.900 64.500 ;
        RECT 269.100 58.050 270.900 59.850 ;
        RECT 273.000 58.050 273.900 63.600 ;
        RECT 275.100 58.050 276.900 59.850 ;
        RECT 293.100 58.050 294.900 59.850 ;
        RECT 299.400 58.050 300.300 70.200 ;
        RECT 314.700 71.100 315.600 71.400 ;
        RECT 319.800 71.400 321.600 77.400 ;
        RECT 319.800 71.100 321.300 71.400 ;
        RECT 314.700 70.200 321.300 71.100 ;
        RECT 314.700 58.050 315.600 70.200 ;
        RECT 335.400 66.300 337.200 77.400 ;
        RECT 341.400 66.300 343.200 77.400 ;
        RECT 335.400 65.400 343.200 66.300 ;
        RECT 344.400 65.400 346.200 77.400 ;
        RECT 365.400 71.400 367.200 77.400 ;
        RECT 386.400 71.400 388.200 77.400 ;
        RECT 403.800 71.400 405.600 77.400 ;
        RECT 316.950 63.450 319.050 64.050 ;
        RECT 340.950 63.450 343.050 64.050 ;
        RECT 316.950 62.550 343.050 63.450 ;
        RECT 316.950 61.950 319.050 62.550 ;
        RECT 340.950 61.950 343.050 62.550 ;
        RECT 330.000 60.450 334.050 61.050 ;
        RECT 320.100 58.050 321.900 59.850 ;
        RECT 329.550 58.950 334.050 60.450 ;
        RECT 222.300 56.100 224.100 57.900 ;
        RECT 222.150 54.000 224.250 56.100 ;
        RECT 226.950 55.800 229.050 57.900 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 295.950 55.950 298.050 58.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 319.950 55.950 322.050 58.050 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 242.100 54.150 243.900 55.950 ;
        RECT 149.400 48.600 150.600 50.700 ;
        RECT 125.400 47.400 130.500 48.600 ;
        RECT 128.700 42.600 130.500 47.400 ;
        RECT 148.800 42.600 150.600 48.600 ;
        RECT 151.800 47.700 159.600 49.050 ;
        RECT 170.400 48.600 171.600 50.700 ;
        RECT 151.800 42.600 153.600 47.700 ;
        RECT 157.800 42.600 159.600 47.700 ;
        RECT 169.800 42.600 171.600 48.600 ;
        RECT 172.800 47.700 180.600 49.050 ;
        RECT 172.800 42.600 174.600 47.700 ;
        RECT 178.800 42.600 180.600 47.700 ;
        RECT 188.400 47.700 196.200 49.050 ;
        RECT 188.400 42.600 190.200 47.700 ;
        RECT 194.400 42.600 196.200 47.700 ;
        RECT 197.400 48.600 198.600 50.700 ;
        RECT 212.400 49.500 216.750 51.000 ;
        RECT 220.350 50.100 223.500 52.200 ;
        RECT 212.400 48.600 213.900 49.500 ;
        RECT 197.400 42.600 199.200 48.600 ;
        RECT 212.400 42.600 214.200 48.600 ;
        RECT 220.350 48.000 221.400 50.100 ;
        RECT 224.700 49.800 226.800 51.900 ;
        RECT 245.400 50.700 246.600 55.950 ;
        RECT 248.100 54.150 249.900 55.950 ;
        RECT 266.100 54.150 267.900 55.950 ;
        RECT 253.950 51.450 256.050 52.050 ;
        RECT 268.950 51.450 271.050 52.050 ;
        RECT 245.400 49.800 249.600 50.700 ;
        RECT 253.950 50.550 271.050 51.450 ;
        RECT 253.950 49.950 256.050 50.550 ;
        RECT 268.950 49.950 271.050 50.550 ;
        RECT 224.700 48.600 229.200 49.800 ;
        RECT 219.600 42.600 221.400 48.000 ;
        RECT 227.400 42.600 229.200 48.600 ;
        RECT 247.800 42.600 249.600 49.800 ;
        RECT 273.000 48.600 274.050 55.950 ;
        RECT 278.100 54.150 279.900 55.950 ;
        RECT 290.100 54.150 291.900 55.950 ;
        RECT 296.100 54.150 297.900 55.950 ;
        RECT 299.400 52.200 300.300 55.950 ;
        RECT 297.000 51.000 300.300 52.200 ;
        RECT 314.700 52.200 315.600 55.950 ;
        RECT 317.100 54.150 318.900 55.950 ;
        RECT 323.100 54.150 324.900 55.950 ;
        RECT 329.550 54.450 330.450 58.950 ;
        RECT 338.100 58.050 339.900 59.850 ;
        RECT 344.700 58.050 345.600 65.400 ;
        RECT 365.850 58.050 367.050 71.400 ;
        RECT 371.100 58.050 372.900 59.850 ;
        RECT 383.100 58.050 384.900 59.850 ;
        RECT 386.400 58.050 387.600 71.400 ;
        RECT 404.700 71.100 405.600 71.400 ;
        RECT 409.800 71.400 411.600 77.400 ;
        RECT 428.400 71.400 430.200 77.400 ;
        RECT 409.800 71.100 411.300 71.400 ;
        RECT 404.700 70.200 411.300 71.100 ;
        RECT 428.700 71.100 430.200 71.400 ;
        RECT 434.400 71.400 436.200 77.400 ;
        RECT 455.400 71.400 457.200 77.400 ;
        RECT 475.800 71.400 477.600 77.400 ;
        RECT 493.800 71.400 495.600 77.400 ;
        RECT 509.400 71.400 511.200 77.400 ;
        RECT 434.400 71.100 435.300 71.400 ;
        RECT 428.700 70.200 435.300 71.100 ;
        RECT 404.700 58.050 405.600 70.200 ;
        RECT 406.950 63.450 409.050 64.050 ;
        RECT 418.950 63.450 421.050 64.050 ;
        RECT 430.950 63.450 433.050 64.050 ;
        RECT 406.950 62.550 433.050 63.450 ;
        RECT 406.950 61.950 409.050 62.550 ;
        RECT 418.950 61.950 421.050 62.550 ;
        RECT 430.950 61.950 433.050 62.550 ;
        RECT 410.100 58.050 411.900 59.850 ;
        RECT 428.100 58.050 429.900 59.850 ;
        RECT 434.400 58.050 435.300 70.200 ;
        RECT 455.850 58.050 457.050 71.400 ;
        RECT 461.100 58.050 462.900 59.850 ;
        RECT 470.100 58.050 471.900 59.850 ;
        RECT 475.950 58.050 477.150 71.400 ;
        RECT 481.950 60.450 486.000 61.050 ;
        RECT 489.000 60.450 493.050 61.050 ;
        RECT 481.950 58.950 486.450 60.450 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 343.950 55.950 346.050 58.050 ;
        RECT 361.950 55.950 364.050 58.050 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 382.950 55.950 385.050 58.050 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 403.950 55.950 406.050 58.050 ;
        RECT 406.950 55.950 409.050 58.050 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 430.950 55.950 433.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 451.950 55.950 454.050 58.050 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 472.950 55.950 475.050 58.050 ;
        RECT 475.950 55.950 478.050 58.050 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 326.550 54.000 330.450 54.450 ;
        RECT 335.100 54.150 336.900 55.950 ;
        RECT 341.100 54.150 342.900 55.950 ;
        RECT 325.950 53.550 330.450 54.000 ;
        RECT 314.700 51.000 318.000 52.200 ;
        RECT 250.950 45.450 253.050 46.050 ;
        RECT 262.950 45.450 265.050 46.050 ;
        RECT 250.950 44.550 265.050 45.450 ;
        RECT 250.950 43.950 253.050 44.550 ;
        RECT 262.950 43.950 265.050 44.550 ;
        RECT 273.000 42.600 274.800 48.600 ;
        RECT 297.000 42.600 298.800 51.000 ;
        RECT 301.950 48.450 304.050 49.050 ;
        RECT 307.950 48.450 310.050 49.050 ;
        RECT 301.950 47.550 310.050 48.450 ;
        RECT 301.950 46.950 304.050 47.550 ;
        RECT 307.950 46.950 310.050 47.550 ;
        RECT 316.200 42.600 318.000 51.000 ;
        RECT 325.950 49.950 328.050 53.550 ;
        RECT 344.700 48.600 345.600 55.950 ;
        RECT 362.100 54.150 363.900 55.950 ;
        RECT 364.950 51.750 366.150 55.950 ;
        RECT 368.100 54.150 369.900 55.950 ;
        RECT 362.400 50.700 366.150 51.750 ;
        RECT 362.400 48.600 363.600 50.700 ;
        RECT 340.500 47.400 345.600 48.600 ;
        RECT 340.500 42.600 342.300 47.400 ;
        RECT 361.800 42.600 363.600 48.600 ;
        RECT 364.800 47.700 372.600 49.050 ;
        RECT 364.800 42.600 366.600 47.700 ;
        RECT 370.800 42.600 372.600 47.700 ;
        RECT 386.400 45.600 387.600 55.950 ;
        RECT 404.700 52.200 405.600 55.950 ;
        RECT 407.100 54.150 408.900 55.950 ;
        RECT 413.100 54.150 414.900 55.950 ;
        RECT 425.100 54.150 426.900 55.950 ;
        RECT 431.100 54.150 432.900 55.950 ;
        RECT 434.400 52.200 435.300 55.950 ;
        RECT 452.100 54.150 453.900 55.950 ;
        RECT 404.700 51.000 408.000 52.200 ;
        RECT 386.400 42.600 388.200 45.600 ;
        RECT 406.200 42.600 408.000 51.000 ;
        RECT 432.000 51.000 435.300 52.200 ;
        RECT 454.950 51.750 456.150 55.950 ;
        RECT 458.100 54.150 459.900 55.950 ;
        RECT 473.100 54.150 474.900 55.950 ;
        RECT 432.000 42.600 433.800 51.000 ;
        RECT 452.400 50.700 456.150 51.750 ;
        RECT 476.850 51.750 478.050 55.950 ;
        RECT 479.100 54.150 480.900 55.950 ;
        RECT 485.550 55.050 486.450 58.950 ;
        RECT 481.950 53.550 486.450 55.050 ;
        RECT 488.550 58.950 493.050 60.450 ;
        RECT 481.950 52.950 486.000 53.550 ;
        RECT 488.550 52.050 489.450 58.950 ;
        RECT 494.400 58.050 495.600 71.400 ;
        RECT 509.700 71.100 511.200 71.400 ;
        RECT 515.400 71.400 517.200 77.400 ;
        RECT 533.400 71.400 535.200 77.400 ;
        RECT 515.400 71.100 516.300 71.400 ;
        RECT 509.700 70.200 516.300 71.100 ;
        RECT 533.700 71.100 535.200 71.400 ;
        RECT 539.400 71.400 541.200 77.400 ;
        RECT 554.400 71.400 556.200 77.400 ;
        RECT 568.800 71.400 570.600 77.400 ;
        RECT 539.400 71.100 540.300 71.400 ;
        RECT 533.700 70.200 540.300 71.100 ;
        RECT 497.100 58.050 498.900 59.850 ;
        RECT 509.100 58.050 510.900 59.850 ;
        RECT 515.400 58.050 516.300 70.200 ;
        RECT 533.100 58.050 534.900 59.850 ;
        RECT 539.400 58.050 540.300 70.200 ;
        RECT 551.100 58.050 552.900 59.850 ;
        RECT 554.400 58.050 555.600 71.400 ;
        RECT 569.700 71.100 570.600 71.400 ;
        RECT 574.800 71.400 576.600 77.400 ;
        RECT 574.800 71.100 576.300 71.400 ;
        RECT 569.700 70.200 576.300 71.100 ;
        RECT 569.700 58.050 570.600 70.200 ;
        RECT 590.400 66.300 592.200 77.400 ;
        RECT 596.400 66.300 598.200 77.400 ;
        RECT 590.400 65.400 598.200 66.300 ;
        RECT 599.400 65.400 601.200 77.400 ;
        RECT 617.400 71.400 619.200 77.400 ;
        RECT 634.800 71.400 636.600 77.400 ;
        RECT 652.800 76.500 660.600 77.400 ;
        RECT 575.100 58.050 576.900 59.850 ;
        RECT 593.100 58.050 594.900 59.850 ;
        RECT 599.700 58.050 600.600 65.400 ;
        RECT 614.100 58.050 615.900 59.850 ;
        RECT 617.400 58.050 618.600 71.400 ;
        RECT 629.100 58.050 630.900 59.850 ;
        RECT 634.950 58.050 636.150 71.400 ;
        RECT 652.800 65.400 654.600 76.500 ;
        RECT 655.800 64.500 657.600 75.600 ;
        RECT 658.800 66.600 660.600 76.500 ;
        RECT 664.800 66.600 666.600 77.400 ;
        RECT 679.800 71.400 681.600 77.400 ;
        RECT 658.800 65.700 666.600 66.600 ;
        RECT 655.800 63.600 660.900 64.500 ;
        RECT 656.100 58.050 657.900 59.850 ;
        RECT 660.000 58.050 660.900 63.600 ;
        RECT 662.100 58.050 663.900 59.850 ;
        RECT 680.400 58.050 681.600 71.400 ;
        RECT 686.550 65.400 688.350 77.400 ;
        RECT 694.050 71.400 695.850 77.400 ;
        RECT 691.950 69.300 695.850 71.400 ;
        RECT 701.850 70.500 703.650 77.400 ;
        RECT 709.650 71.400 711.450 77.400 ;
        RECT 710.250 70.500 711.450 71.400 ;
        RECT 700.950 69.450 707.550 70.500 ;
        RECT 700.950 68.700 702.750 69.450 ;
        RECT 705.750 68.700 707.550 69.450 ;
        RECT 710.250 68.400 715.050 70.500 ;
        RECT 693.150 66.600 695.850 68.400 ;
        RECT 696.750 67.800 698.550 68.400 ;
        RECT 696.750 66.900 703.050 67.800 ;
        RECT 710.250 67.500 711.450 68.400 ;
        RECT 696.750 66.600 698.550 66.900 ;
        RECT 694.950 65.700 695.850 66.600 ;
        RECT 683.100 58.050 684.900 59.850 ;
        RECT 686.550 58.050 687.750 65.400 ;
        RECT 691.950 64.800 694.050 65.700 ;
        RECT 694.950 64.800 700.050 65.700 ;
        RECT 689.850 63.600 694.050 64.800 ;
        RECT 688.950 61.800 690.750 63.600 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 496.950 55.950 499.050 58.050 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 550.950 55.950 553.050 58.050 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 628.950 55.950 631.050 58.050 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 686.550 57.750 691.050 58.050 ;
        RECT 686.550 55.950 692.850 57.750 ;
        RECT 486.000 51.900 489.450 52.050 ;
        RECT 476.850 50.700 480.600 51.750 ;
        RECT 452.400 48.600 453.600 50.700 ;
        RECT 451.800 42.600 453.600 48.600 ;
        RECT 454.800 47.700 462.600 49.050 ;
        RECT 454.800 42.600 456.600 47.700 ;
        RECT 460.800 42.600 462.600 47.700 ;
        RECT 470.400 47.700 478.200 49.050 ;
        RECT 470.400 42.600 472.200 47.700 ;
        RECT 476.400 42.600 478.200 47.700 ;
        RECT 479.400 48.600 480.600 50.700 ;
        RECT 484.950 50.550 489.450 51.900 ;
        RECT 484.950 49.950 489.000 50.550 ;
        RECT 484.950 49.800 487.050 49.950 ;
        RECT 479.400 42.600 481.200 48.600 ;
        RECT 494.400 45.600 495.600 55.950 ;
        RECT 506.100 54.150 507.900 55.950 ;
        RECT 512.100 54.150 513.900 55.950 ;
        RECT 515.400 52.200 516.300 55.950 ;
        RECT 530.100 54.150 531.900 55.950 ;
        RECT 536.100 54.150 537.900 55.950 ;
        RECT 539.400 52.200 540.300 55.950 ;
        RECT 493.800 42.600 495.600 45.600 ;
        RECT 513.000 51.000 516.300 52.200 ;
        RECT 537.000 51.000 540.300 52.200 ;
        RECT 541.950 51.450 544.050 52.050 ;
        RECT 550.950 51.450 553.050 51.750 ;
        RECT 513.000 42.600 514.800 51.000 ;
        RECT 537.000 42.600 538.800 51.000 ;
        RECT 541.950 50.550 553.050 51.450 ;
        RECT 541.950 49.950 544.050 50.550 ;
        RECT 550.950 49.650 553.050 50.550 ;
        RECT 554.400 45.600 555.600 55.950 ;
        RECT 569.700 52.200 570.600 55.950 ;
        RECT 572.100 54.150 573.900 55.950 ;
        RECT 578.100 54.150 579.900 55.950 ;
        RECT 590.100 54.150 591.900 55.950 ;
        RECT 596.100 54.150 597.900 55.950 ;
        RECT 569.700 51.000 573.000 52.200 ;
        RECT 554.400 42.600 556.200 45.600 ;
        RECT 571.200 42.600 573.000 51.000 ;
        RECT 599.700 48.600 600.600 55.950 ;
        RECT 595.500 47.400 600.600 48.600 ;
        RECT 595.500 42.600 597.300 47.400 ;
        RECT 617.400 45.600 618.600 55.950 ;
        RECT 632.100 54.150 633.900 55.950 ;
        RECT 635.850 51.750 637.050 55.950 ;
        RECT 638.100 54.150 639.900 55.950 ;
        RECT 653.100 54.150 654.900 55.950 ;
        RECT 635.850 50.700 639.600 51.750 ;
        RECT 629.400 47.700 637.200 49.050 ;
        RECT 617.400 42.600 619.200 45.600 ;
        RECT 629.400 42.600 631.200 47.700 ;
        RECT 635.400 42.600 637.200 47.700 ;
        RECT 638.400 48.600 639.600 50.700 ;
        RECT 660.000 48.600 661.050 55.950 ;
        RECT 665.100 54.150 666.900 55.950 ;
        RECT 638.400 42.600 640.200 48.600 ;
        RECT 660.000 42.600 661.800 48.600 ;
        RECT 680.400 45.600 681.600 55.950 ;
        RECT 679.800 42.600 681.600 45.600 ;
        RECT 686.550 48.600 687.750 55.950 ;
        RECT 699.150 52.200 700.050 64.800 ;
        RECT 702.150 64.800 703.050 66.900 ;
        RECT 703.950 66.300 711.450 67.500 ;
        RECT 703.950 65.700 705.750 66.300 ;
        RECT 718.050 65.400 719.850 77.400 ;
        RECT 733.800 71.400 735.600 77.400 ;
        RECT 702.150 64.500 710.550 64.800 ;
        RECT 718.950 64.500 719.850 65.400 ;
        RECT 702.150 63.900 719.850 64.500 ;
        RECT 708.750 63.300 719.850 63.900 ;
        RECT 708.750 63.000 710.550 63.300 ;
        RECT 706.950 56.400 709.050 58.050 ;
        RECT 706.950 55.200 714.900 56.400 ;
        RECT 715.950 55.950 718.050 58.050 ;
        RECT 713.100 54.600 714.900 55.200 ;
        RECT 716.100 54.150 717.900 55.950 ;
        RECT 710.100 53.400 711.900 54.000 ;
        RECT 716.100 53.400 717.000 54.150 ;
        RECT 710.100 52.200 717.000 53.400 ;
        RECT 699.150 51.000 711.150 52.200 ;
        RECT 699.150 50.400 700.950 51.000 ;
        RECT 710.100 49.200 711.150 51.000 ;
        RECT 686.550 42.600 688.350 48.600 ;
        RECT 691.950 47.700 694.050 48.600 ;
        RECT 691.950 46.500 695.700 47.700 ;
        RECT 706.350 47.550 708.150 48.300 ;
        RECT 694.650 45.600 695.700 46.500 ;
        RECT 703.200 46.500 708.150 47.550 ;
        RECT 709.650 47.400 711.450 49.200 ;
        RECT 718.950 48.600 719.850 63.300 ;
        RECT 734.400 58.050 735.600 71.400 ;
        RECT 751.800 76.500 759.600 77.400 ;
        RECT 751.800 65.400 753.600 76.500 ;
        RECT 754.800 64.500 756.600 75.600 ;
        RECT 757.800 66.600 759.600 76.500 ;
        RECT 763.800 66.600 765.600 77.400 ;
        RECT 778.800 71.400 780.600 77.400 ;
        RECT 757.800 65.700 765.600 66.600 ;
        RECT 754.800 63.600 759.900 64.500 ;
        RECT 737.100 58.050 738.900 59.850 ;
        RECT 755.100 58.050 756.900 59.850 ;
        RECT 759.000 58.050 759.900 63.600 ;
        RECT 761.100 58.050 762.900 59.850 ;
        RECT 779.400 58.050 780.600 71.400 ;
        RECT 785.550 65.400 787.350 77.400 ;
        RECT 793.050 71.400 794.850 77.400 ;
        RECT 790.950 69.300 794.850 71.400 ;
        RECT 800.850 70.500 802.650 77.400 ;
        RECT 808.650 71.400 810.450 77.400 ;
        RECT 809.250 70.500 810.450 71.400 ;
        RECT 799.950 69.450 806.550 70.500 ;
        RECT 799.950 68.700 801.750 69.450 ;
        RECT 804.750 68.700 806.550 69.450 ;
        RECT 809.250 68.400 814.050 70.500 ;
        RECT 792.150 66.600 794.850 68.400 ;
        RECT 795.750 67.800 797.550 68.400 ;
        RECT 795.750 66.900 802.050 67.800 ;
        RECT 809.250 67.500 810.450 68.400 ;
        RECT 795.750 66.600 797.550 66.900 ;
        RECT 793.950 65.700 794.850 66.600 ;
        RECT 782.100 58.050 783.900 59.850 ;
        RECT 785.550 58.050 786.750 65.400 ;
        RECT 790.950 64.800 793.050 65.700 ;
        RECT 793.950 64.800 799.050 65.700 ;
        RECT 788.850 63.600 793.050 64.800 ;
        RECT 787.950 61.800 789.750 63.600 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 785.550 57.750 790.050 58.050 ;
        RECT 785.550 55.950 791.850 57.750 ;
        RECT 712.950 46.500 715.050 48.600 ;
        RECT 703.200 45.600 704.250 46.500 ;
        RECT 712.950 45.600 714.000 46.500 ;
        RECT 694.650 42.600 696.450 45.600 ;
        RECT 702.450 42.600 704.250 45.600 ;
        RECT 710.250 44.700 714.000 45.600 ;
        RECT 710.250 42.600 712.050 44.700 ;
        RECT 718.050 42.600 719.850 48.600 ;
        RECT 734.400 45.600 735.600 55.950 ;
        RECT 752.100 54.150 753.900 55.950 ;
        RECT 733.800 42.600 735.600 45.600 ;
        RECT 759.000 48.600 760.050 55.950 ;
        RECT 764.100 54.150 765.900 55.950 ;
        RECT 759.000 42.600 760.800 48.600 ;
        RECT 779.400 45.600 780.600 55.950 ;
        RECT 778.800 42.600 780.600 45.600 ;
        RECT 785.550 48.600 786.750 55.950 ;
        RECT 798.150 52.200 799.050 64.800 ;
        RECT 801.150 64.800 802.050 66.900 ;
        RECT 802.950 66.300 810.450 67.500 ;
        RECT 802.950 65.700 804.750 66.300 ;
        RECT 817.050 65.400 818.850 77.400 ;
        RECT 801.150 64.500 809.550 64.800 ;
        RECT 817.950 64.500 818.850 65.400 ;
        RECT 801.150 63.900 818.850 64.500 ;
        RECT 807.750 63.300 818.850 63.900 ;
        RECT 807.750 63.000 809.550 63.300 ;
        RECT 805.950 56.400 808.050 58.050 ;
        RECT 805.950 55.200 813.900 56.400 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 812.100 54.600 813.900 55.200 ;
        RECT 815.100 54.150 816.900 55.950 ;
        RECT 809.100 53.400 810.900 54.000 ;
        RECT 815.100 53.400 816.000 54.150 ;
        RECT 809.100 52.200 816.000 53.400 ;
        RECT 798.150 51.000 810.150 52.200 ;
        RECT 798.150 50.400 799.950 51.000 ;
        RECT 809.100 49.200 810.150 51.000 ;
        RECT 785.550 42.600 787.350 48.600 ;
        RECT 790.950 47.700 793.050 48.600 ;
        RECT 790.950 46.500 794.700 47.700 ;
        RECT 805.350 47.550 807.150 48.300 ;
        RECT 793.650 45.600 794.700 46.500 ;
        RECT 802.200 46.500 807.150 47.550 ;
        RECT 808.650 47.400 810.450 49.200 ;
        RECT 817.950 48.600 818.850 63.300 ;
        RECT 811.950 46.500 814.050 48.600 ;
        RECT 802.200 45.600 803.250 46.500 ;
        RECT 811.950 45.600 813.000 46.500 ;
        RECT 793.650 42.600 795.450 45.600 ;
        RECT 801.450 42.600 803.250 45.600 ;
        RECT 809.250 44.700 813.000 45.600 ;
        RECT 809.250 42.600 811.050 44.700 ;
        RECT 817.050 42.600 818.850 48.600 ;
        RECT 822.150 65.400 823.950 77.400 ;
        RECT 830.550 71.400 832.350 77.400 ;
        RECT 830.550 70.500 831.750 71.400 ;
        RECT 838.350 70.500 840.150 77.400 ;
        RECT 846.150 71.400 847.950 77.400 ;
        RECT 826.950 68.400 831.750 70.500 ;
        RECT 834.450 69.450 841.050 70.500 ;
        RECT 834.450 68.700 836.250 69.450 ;
        RECT 839.250 68.700 841.050 69.450 ;
        RECT 846.150 69.300 850.050 71.400 ;
        RECT 830.550 67.500 831.750 68.400 ;
        RECT 843.450 67.800 845.250 68.400 ;
        RECT 830.550 66.300 838.050 67.500 ;
        RECT 836.250 65.700 838.050 66.300 ;
        RECT 838.950 66.900 845.250 67.800 ;
        RECT 822.150 64.500 823.050 65.400 ;
        RECT 838.950 64.800 839.850 66.900 ;
        RECT 843.450 66.600 845.250 66.900 ;
        RECT 846.150 66.600 848.850 68.400 ;
        RECT 846.150 65.700 847.050 66.600 ;
        RECT 831.450 64.500 839.850 64.800 ;
        RECT 822.150 63.900 839.850 64.500 ;
        RECT 841.950 64.800 847.050 65.700 ;
        RECT 847.950 64.800 850.050 65.700 ;
        RECT 853.650 65.400 855.450 77.400 ;
        RECT 866.400 71.400 868.200 77.400 ;
        RECT 866.700 71.100 868.200 71.400 ;
        RECT 872.400 71.400 874.200 77.400 ;
        RECT 892.800 71.400 894.600 77.400 ;
        RECT 872.400 71.100 873.300 71.400 ;
        RECT 866.700 70.200 873.300 71.100 ;
        RECT 822.150 63.300 833.250 63.900 ;
        RECT 822.150 48.600 823.050 63.300 ;
        RECT 831.450 63.000 833.250 63.300 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 832.950 56.400 835.050 58.050 ;
        RECT 824.100 54.150 825.900 55.950 ;
        RECT 827.100 55.200 835.050 56.400 ;
        RECT 827.100 54.600 828.900 55.200 ;
        RECT 825.000 53.400 825.900 54.150 ;
        RECT 830.100 53.400 831.900 54.000 ;
        RECT 825.000 52.200 831.900 53.400 ;
        RECT 841.950 52.200 842.850 64.800 ;
        RECT 847.950 63.600 852.150 64.800 ;
        RECT 851.250 61.800 853.050 63.600 ;
        RECT 854.250 58.050 855.450 65.400 ;
        RECT 866.100 58.050 867.900 59.850 ;
        RECT 872.400 58.050 873.300 70.200 ;
        RECT 877.950 63.450 880.050 64.050 ;
        RECT 886.950 63.450 889.050 64.050 ;
        RECT 877.950 62.550 889.050 63.450 ;
        RECT 877.950 61.950 880.050 62.550 ;
        RECT 886.950 61.950 889.050 62.550 ;
        RECT 887.100 58.050 888.900 59.850 ;
        RECT 892.950 58.050 894.150 71.400 ;
        RECT 850.950 57.750 855.450 58.050 ;
        RECT 849.150 55.950 855.450 57.750 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 865.950 55.950 868.050 58.050 ;
        RECT 868.950 55.950 871.050 58.050 ;
        RECT 871.950 55.950 874.050 58.050 ;
        RECT 886.950 55.950 889.050 58.050 ;
        RECT 889.950 55.950 892.050 58.050 ;
        RECT 892.950 55.950 895.050 58.050 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 830.850 51.000 842.850 52.200 ;
        RECT 830.850 49.200 831.900 51.000 ;
        RECT 841.050 50.400 842.850 51.000 ;
        RECT 822.150 42.600 823.950 48.600 ;
        RECT 826.950 46.500 829.050 48.600 ;
        RECT 830.550 47.400 832.350 49.200 ;
        RECT 854.250 48.600 855.450 55.950 ;
        RECT 863.100 54.150 864.900 55.950 ;
        RECT 869.100 54.150 870.900 55.950 ;
        RECT 872.400 52.200 873.300 55.950 ;
        RECT 890.100 54.150 891.900 55.950 ;
        RECT 833.850 47.550 835.650 48.300 ;
        RECT 847.950 47.700 850.050 48.600 ;
        RECT 833.850 46.500 838.800 47.550 ;
        RECT 828.000 45.600 829.050 46.500 ;
        RECT 837.750 45.600 838.800 46.500 ;
        RECT 846.300 46.500 850.050 47.700 ;
        RECT 846.300 45.600 847.350 46.500 ;
        RECT 828.000 44.700 831.750 45.600 ;
        RECT 829.950 42.600 831.750 44.700 ;
        RECT 837.750 42.600 839.550 45.600 ;
        RECT 845.550 42.600 847.350 45.600 ;
        RECT 853.650 42.600 855.450 48.600 ;
        RECT 870.000 51.000 873.300 52.200 ;
        RECT 893.850 51.750 895.050 55.950 ;
        RECT 896.100 54.150 897.900 55.950 ;
        RECT 870.000 42.600 871.800 51.000 ;
        RECT 893.850 50.700 897.600 51.750 ;
        RECT 887.400 47.700 895.200 49.050 ;
        RECT 887.400 42.600 889.200 47.700 ;
        RECT 893.400 42.600 895.200 47.700 ;
        RECT 896.400 48.600 897.600 50.700 ;
        RECT 896.400 42.600 898.200 48.600 ;
        RECT 17.700 33.600 19.500 38.400 ;
        RECT 34.800 35.400 36.600 38.400 ;
        RECT 14.400 32.400 19.500 33.600 ;
        RECT 14.400 25.050 15.300 32.400 ;
        RECT 17.100 25.050 18.900 26.850 ;
        RECT 23.100 25.050 24.900 26.850 ;
        RECT 35.400 25.050 36.600 35.400 ;
        RECT 52.800 32.400 54.600 38.400 ;
        RECT 53.400 30.300 54.600 32.400 ;
        RECT 55.800 33.300 57.600 38.400 ;
        RECT 61.800 33.300 63.600 38.400 ;
        RECT 55.800 31.950 63.600 33.300 ;
        RECT 53.400 29.250 57.150 30.300 ;
        RECT 53.100 25.050 54.900 26.850 ;
        RECT 55.950 25.050 57.150 29.250 ;
        RECT 78.000 30.000 79.800 38.400 ;
        RECT 102.000 30.000 103.800 38.400 ;
        RECT 119.400 33.300 121.200 38.400 ;
        RECT 125.400 33.300 127.200 38.400 ;
        RECT 119.400 31.950 127.200 33.300 ;
        RECT 128.400 32.400 130.200 38.400 ;
        RECT 145.800 35.400 147.600 38.400 ;
        RECT 128.400 30.300 129.600 32.400 ;
        RECT 78.000 28.800 81.300 30.000 ;
        RECT 102.000 28.800 105.300 30.000 ;
        RECT 59.100 25.050 60.900 26.850 ;
        RECT 71.100 25.050 72.900 26.850 ;
        RECT 77.100 25.050 78.900 26.850 ;
        RECT 80.400 25.050 81.300 28.800 ;
        RECT 95.100 25.050 96.900 26.850 ;
        RECT 101.100 25.050 102.900 26.850 ;
        RECT 104.400 25.050 105.300 28.800 ;
        RECT 125.850 29.250 129.600 30.300 ;
        RECT 122.100 25.050 123.900 26.850 ;
        RECT 125.850 25.050 127.050 29.250 ;
        RECT 128.100 25.050 129.900 26.850 ;
        RECT 146.400 25.050 147.600 35.400 ;
        RECT 165.000 30.000 166.800 38.400 ;
        RECT 189.000 30.000 190.800 38.400 ;
        RECT 211.500 33.600 213.300 38.400 ;
        RECT 211.500 32.400 216.600 33.600 ;
        RECT 165.000 28.800 168.300 30.000 ;
        RECT 189.000 28.800 192.300 30.000 ;
        RECT 158.100 25.050 159.900 26.850 ;
        RECT 164.100 25.050 165.900 26.850 ;
        RECT 167.400 25.050 168.300 28.800 ;
        RECT 182.100 25.050 183.900 26.850 ;
        RECT 188.100 25.050 189.900 26.850 ;
        RECT 191.400 25.050 192.300 28.800 ;
        RECT 206.100 25.050 207.900 26.850 ;
        RECT 212.100 25.050 213.900 26.850 ;
        RECT 215.700 25.050 216.600 32.400 ;
        RECT 233.400 31.200 235.200 38.400 ;
        RECT 241.950 36.450 244.050 37.050 ;
        RECT 250.950 36.450 253.050 37.050 ;
        RECT 241.950 35.550 253.050 36.450 ;
        RECT 241.950 34.950 244.050 35.550 ;
        RECT 250.950 34.950 253.050 35.550 ;
        RECT 233.400 30.300 237.600 31.200 ;
        RECT 220.950 27.450 223.050 28.050 ;
        RECT 229.950 27.450 232.050 28.050 ;
        RECT 220.950 26.550 232.050 27.450 ;
        RECT 220.950 25.950 223.050 26.550 ;
        RECT 229.950 25.950 232.050 26.550 ;
        RECT 233.100 25.050 234.900 26.850 ;
        RECT 236.400 25.050 237.600 30.300 ;
        RECT 256.200 30.000 258.000 38.400 ;
        RECT 280.500 33.600 282.300 38.400 ;
        RECT 280.500 32.400 285.600 33.600 ;
        RECT 254.700 28.800 258.000 30.000 ;
        RECT 239.100 25.050 240.900 26.850 ;
        RECT 254.700 25.050 255.600 28.800 ;
        RECT 257.100 25.050 258.900 26.850 ;
        RECT 263.100 25.050 264.900 26.850 ;
        RECT 275.100 25.050 276.900 26.850 ;
        RECT 281.100 25.050 282.900 26.850 ;
        RECT 284.700 25.050 285.600 32.400 ;
        RECT 306.000 30.000 307.800 38.400 ;
        RECT 328.500 33.600 330.300 38.400 ;
        RECT 347.400 35.400 349.200 38.400 ;
        RECT 328.500 32.400 333.600 33.600 ;
        RECT 306.000 28.800 309.300 30.000 ;
        RECT 299.100 25.050 300.900 26.850 ;
        RECT 305.100 25.050 306.900 26.850 ;
        RECT 308.400 25.050 309.300 28.800 ;
        RECT 323.100 25.050 324.900 26.850 ;
        RECT 329.100 25.050 330.900 26.850 ;
        RECT 332.700 25.050 333.600 32.400 ;
        RECT 347.400 25.050 348.600 35.400 ;
        RECT 368.700 33.600 370.500 38.400 ;
        RECT 365.400 32.400 370.500 33.600 ;
        RECT 365.400 25.050 366.300 32.400 ;
        RECT 391.800 31.200 393.600 38.400 ;
        RECT 407.400 33.300 409.200 38.400 ;
        RECT 413.400 33.300 415.200 38.400 ;
        RECT 407.400 31.950 415.200 33.300 ;
        RECT 416.400 32.400 418.200 38.400 ;
        RECT 436.500 33.600 438.300 38.400 ;
        RECT 436.500 32.400 441.600 33.600 ;
        RECT 389.400 30.300 393.600 31.200 ;
        RECT 416.400 30.300 417.600 32.400 ;
        RECT 381.000 27.450 385.050 28.050 ;
        RECT 368.100 25.050 369.900 26.850 ;
        RECT 374.100 25.050 375.900 26.850 ;
        RECT 380.550 25.950 385.050 27.450 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 22.950 22.950 25.050 25.050 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 76.950 22.950 79.050 25.050 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 97.950 22.950 100.050 25.050 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 118.950 22.950 121.050 25.050 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 163.950 22.950 166.050 25.050 ;
        RECT 166.950 22.950 169.050 25.050 ;
        RECT 181.950 22.950 184.050 25.050 ;
        RECT 184.950 22.950 187.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 190.950 22.950 193.050 25.050 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 283.950 22.950 286.050 25.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 304.950 22.950 307.050 25.050 ;
        RECT 307.950 22.950 310.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 331.950 22.950 334.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 367.950 22.950 370.050 25.050 ;
        RECT 370.950 22.950 373.050 25.050 ;
        RECT 373.950 22.950 376.050 25.050 ;
        RECT 14.400 15.600 15.300 22.950 ;
        RECT 20.100 21.150 21.900 22.950 ;
        RECT 13.800 3.600 15.600 15.600 ;
        RECT 16.800 14.700 24.600 15.600 ;
        RECT 16.800 3.600 18.600 14.700 ;
        RECT 22.800 3.600 24.600 14.700 ;
        RECT 35.400 9.600 36.600 22.950 ;
        RECT 38.100 21.150 39.900 22.950 ;
        RECT 56.850 9.600 58.050 22.950 ;
        RECT 62.100 21.150 63.900 22.950 ;
        RECT 74.100 21.150 75.900 22.950 ;
        RECT 80.400 10.800 81.300 22.950 ;
        RECT 98.100 21.150 99.900 22.950 ;
        RECT 85.950 18.450 88.050 19.050 ;
        RECT 100.950 18.450 103.050 19.050 ;
        RECT 85.950 17.550 103.050 18.450 ;
        RECT 85.950 16.950 88.050 17.550 ;
        RECT 100.950 16.950 103.050 17.550 ;
        RECT 104.400 10.800 105.300 22.950 ;
        RECT 119.100 21.150 120.900 22.950 ;
        RECT 74.700 9.900 81.300 10.800 ;
        RECT 74.700 9.600 76.200 9.900 ;
        RECT 34.800 3.600 36.600 9.600 ;
        RECT 56.400 3.600 58.200 9.600 ;
        RECT 74.400 3.600 76.200 9.600 ;
        RECT 80.400 9.600 81.300 9.900 ;
        RECT 98.700 9.900 105.300 10.800 ;
        RECT 98.700 9.600 100.200 9.900 ;
        RECT 80.400 3.600 82.200 9.600 ;
        RECT 98.400 3.600 100.200 9.600 ;
        RECT 104.400 9.600 105.300 9.900 ;
        RECT 124.950 9.600 126.150 22.950 ;
        RECT 146.400 9.600 147.600 22.950 ;
        RECT 149.100 21.150 150.900 22.950 ;
        RECT 161.100 21.150 162.900 22.950 ;
        RECT 148.950 18.450 151.050 19.050 ;
        RECT 163.950 18.450 166.050 19.050 ;
        RECT 148.950 17.550 166.050 18.450 ;
        RECT 148.950 16.950 151.050 17.550 ;
        RECT 163.950 16.950 166.050 17.550 ;
        RECT 167.400 10.800 168.300 22.950 ;
        RECT 185.100 21.150 186.900 22.950 ;
        RECT 172.800 18.000 174.900 19.050 ;
        RECT 175.950 18.450 178.050 19.050 ;
        RECT 187.950 18.450 190.050 19.050 ;
        RECT 172.800 16.950 175.050 18.000 ;
        RECT 175.950 17.550 190.050 18.450 ;
        RECT 175.950 16.950 178.050 17.550 ;
        RECT 187.950 16.950 190.050 17.550 ;
        RECT 172.950 15.450 175.050 16.950 ;
        RECT 184.950 15.450 187.050 15.900 ;
        RECT 172.950 15.000 187.050 15.450 ;
        RECT 173.550 14.550 187.050 15.000 ;
        RECT 184.950 13.800 187.050 14.550 ;
        RECT 191.400 10.800 192.300 22.950 ;
        RECT 209.100 21.150 210.900 22.950 ;
        RECT 215.700 15.600 216.600 22.950 ;
        RECT 161.700 9.900 168.300 10.800 ;
        RECT 161.700 9.600 163.200 9.900 ;
        RECT 104.400 3.600 106.200 9.600 ;
        RECT 124.800 3.600 126.600 9.600 ;
        RECT 145.800 3.600 147.600 9.600 ;
        RECT 161.400 3.600 163.200 9.600 ;
        RECT 167.400 9.600 168.300 9.900 ;
        RECT 185.700 9.900 192.300 10.800 ;
        RECT 185.700 9.600 187.200 9.900 ;
        RECT 167.400 3.600 169.200 9.600 ;
        RECT 185.400 3.600 187.200 9.600 ;
        RECT 191.400 9.600 192.300 9.900 ;
        RECT 206.400 14.700 214.200 15.600 ;
        RECT 191.400 3.600 193.200 9.600 ;
        RECT 206.400 3.600 208.200 14.700 ;
        RECT 212.400 3.600 214.200 14.700 ;
        RECT 215.400 3.600 217.200 15.600 ;
        RECT 236.400 9.600 237.600 22.950 ;
        RECT 254.700 10.800 255.600 22.950 ;
        RECT 260.100 21.150 261.900 22.950 ;
        RECT 278.100 21.150 279.900 22.950 ;
        RECT 284.700 15.600 285.600 22.950 ;
        RECT 302.100 21.150 303.900 22.950 ;
        RECT 275.400 14.700 283.200 15.600 ;
        RECT 254.700 9.900 261.300 10.800 ;
        RECT 254.700 9.600 255.600 9.900 ;
        RECT 235.800 3.600 237.600 9.600 ;
        RECT 253.800 3.600 255.600 9.600 ;
        RECT 259.800 9.600 261.300 9.900 ;
        RECT 259.800 3.600 261.600 9.600 ;
        RECT 275.400 3.600 277.200 14.700 ;
        RECT 281.400 3.600 283.200 14.700 ;
        RECT 284.400 3.600 286.200 15.600 ;
        RECT 308.400 10.800 309.300 22.950 ;
        RECT 313.950 21.450 316.050 22.050 ;
        RECT 319.950 21.450 322.050 22.050 ;
        RECT 313.950 20.550 322.050 21.450 ;
        RECT 326.100 21.150 327.900 22.950 ;
        RECT 313.950 19.950 316.050 20.550 ;
        RECT 319.950 19.950 322.050 20.550 ;
        RECT 310.950 18.450 313.050 19.050 ;
        RECT 328.950 18.450 331.050 19.050 ;
        RECT 310.950 17.550 331.050 18.450 ;
        RECT 310.950 16.950 313.050 17.550 ;
        RECT 328.950 16.950 331.050 17.550 ;
        RECT 332.700 15.600 333.600 22.950 ;
        RECT 344.100 21.150 345.900 22.950 ;
        RECT 302.700 9.900 309.300 10.800 ;
        RECT 302.700 9.600 304.200 9.900 ;
        RECT 302.400 3.600 304.200 9.600 ;
        RECT 308.400 9.600 309.300 9.900 ;
        RECT 323.400 14.700 331.200 15.600 ;
        RECT 308.400 3.600 310.200 9.600 ;
        RECT 323.400 3.600 325.200 14.700 ;
        RECT 329.400 3.600 331.200 14.700 ;
        RECT 332.400 3.600 334.200 15.600 ;
        RECT 347.400 9.600 348.600 22.950 ;
        RECT 365.400 15.600 366.300 22.950 ;
        RECT 371.100 21.150 372.900 22.950 ;
        RECT 380.550 22.050 381.450 25.950 ;
        RECT 386.100 25.050 387.900 26.850 ;
        RECT 389.400 25.050 390.600 30.300 ;
        RECT 413.850 29.250 417.600 30.300 ;
        RECT 424.950 30.450 427.050 31.050 ;
        RECT 436.950 30.450 439.050 31.050 ;
        RECT 424.950 29.550 439.050 30.450 ;
        RECT 392.100 25.050 393.900 26.850 ;
        RECT 410.100 25.050 411.900 26.850 ;
        RECT 413.850 25.050 415.050 29.250 ;
        RECT 424.950 28.950 427.050 29.550 ;
        RECT 436.950 28.950 439.050 29.550 ;
        RECT 416.100 25.050 417.900 26.850 ;
        RECT 431.100 25.050 432.900 26.850 ;
        RECT 437.100 25.050 438.900 26.850 ;
        RECT 440.700 25.050 441.600 32.400 ;
        RECT 459.000 30.000 460.800 38.400 ;
        RECT 478.800 32.400 480.600 38.400 ;
        RECT 479.400 30.300 480.600 32.400 ;
        RECT 481.800 33.300 483.600 38.400 ;
        RECT 487.800 33.300 489.600 38.400 ;
        RECT 506.400 35.400 508.200 38.400 ;
        RECT 512.400 35.400 514.200 38.400 ;
        RECT 507.150 34.500 508.200 35.400 ;
        RECT 513.150 34.500 514.200 35.400 ;
        RECT 507.150 33.600 517.950 34.500 ;
        RECT 481.800 31.950 489.600 33.300 ;
        RECT 459.000 28.800 462.300 30.000 ;
        RECT 479.400 29.250 483.150 30.300 ;
        RECT 442.950 27.450 447.000 28.050 ;
        RECT 442.950 25.950 447.450 27.450 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 415.950 22.950 418.050 25.050 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 376.950 20.550 381.450 22.050 ;
        RECT 376.950 19.950 381.000 20.550 ;
        RECT 347.400 3.600 349.200 9.600 ;
        RECT 364.800 3.600 366.600 15.600 ;
        RECT 367.800 14.700 375.600 15.600 ;
        RECT 367.800 3.600 369.600 14.700 ;
        RECT 373.800 3.600 375.600 14.700 ;
        RECT 389.400 9.600 390.600 22.950 ;
        RECT 407.100 21.150 408.900 22.950 ;
        RECT 412.950 9.600 414.150 22.950 ;
        RECT 434.100 21.150 435.900 22.950 ;
        RECT 440.700 15.600 441.600 22.950 ;
        RECT 446.550 22.050 447.450 25.950 ;
        RECT 452.100 25.050 453.900 26.850 ;
        RECT 458.100 25.050 459.900 26.850 ;
        RECT 461.400 25.050 462.300 28.800 ;
        RECT 479.100 25.050 480.900 26.850 ;
        RECT 481.950 25.050 483.150 29.250 ;
        RECT 485.100 25.050 486.900 26.850 ;
        RECT 509.100 25.200 510.900 27.000 ;
        RECT 516.750 25.200 517.950 33.600 ;
        RECT 536.400 33.300 538.200 38.400 ;
        RECT 542.400 33.300 544.200 38.400 ;
        RECT 536.400 31.950 544.200 33.300 ;
        RECT 545.400 32.400 547.200 38.400 ;
        RECT 563.700 33.600 565.500 38.400 ;
        RECT 560.400 32.400 565.500 33.600 ;
        RECT 583.800 32.400 585.600 38.400 ;
        RECT 591.600 33.000 593.400 38.400 ;
        RECT 545.400 30.300 546.600 32.400 ;
        RECT 542.850 29.250 546.600 30.300 ;
        RECT 451.950 22.950 454.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 502.950 23.100 505.050 25.200 ;
        RECT 508.950 23.100 511.050 25.200 ;
        RECT 511.950 23.100 514.050 25.200 ;
        RECT 516.750 23.100 520.050 25.200 ;
        RECT 539.100 25.050 540.900 26.850 ;
        RECT 542.850 25.050 544.050 29.250 ;
        RECT 545.100 25.050 546.900 26.850 ;
        RECT 560.400 25.050 561.300 32.400 ;
        RECT 583.800 31.200 588.300 32.400 ;
        RECT 586.200 29.100 588.300 31.200 ;
        RECT 591.600 30.900 592.650 33.000 ;
        RECT 598.800 32.400 600.600 38.400 ;
        RECT 599.100 31.500 600.600 32.400 ;
        RECT 589.500 28.800 592.650 30.900 ;
        RECT 596.250 30.000 600.600 31.500 ;
        RECT 611.400 31.200 613.200 38.400 ;
        RECT 634.500 33.600 636.300 38.400 ;
        RECT 656.400 35.400 658.200 38.400 ;
        RECT 634.500 32.400 639.600 33.600 ;
        RECT 611.400 30.300 615.600 31.200 ;
        RECT 563.100 25.050 564.900 26.850 ;
        RECT 569.100 25.050 570.900 26.850 ;
        RECT 446.550 20.550 451.050 22.050 ;
        RECT 455.100 21.150 456.900 22.950 ;
        RECT 447.000 19.950 451.050 20.550 ;
        RECT 431.400 14.700 439.200 15.600 ;
        RECT 389.400 3.600 391.200 9.600 ;
        RECT 412.800 3.600 414.600 9.600 ;
        RECT 418.950 6.450 421.050 7.050 ;
        RECT 424.950 6.450 427.050 7.050 ;
        RECT 418.950 5.550 427.050 6.450 ;
        RECT 418.950 4.950 421.050 5.550 ;
        RECT 424.950 4.950 427.050 5.550 ;
        RECT 431.400 3.600 433.200 14.700 ;
        RECT 437.400 3.600 439.200 14.700 ;
        RECT 440.400 3.600 442.200 15.600 ;
        RECT 461.400 10.800 462.300 22.950 ;
        RECT 455.700 9.900 462.300 10.800 ;
        RECT 455.700 9.600 457.200 9.900 ;
        RECT 455.400 3.600 457.200 9.600 ;
        RECT 461.400 9.600 462.300 9.900 ;
        RECT 482.850 9.600 484.050 22.950 ;
        RECT 488.100 21.150 489.900 22.950 ;
        RECT 503.100 21.300 504.900 23.100 ;
        RECT 512.100 21.300 513.900 23.100 ;
        RECT 516.750 16.800 517.950 23.100 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 544.950 22.950 547.050 25.050 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 568.950 22.950 571.050 25.050 ;
        RECT 583.950 23.100 586.050 25.200 ;
        RECT 588.750 24.900 590.850 27.000 ;
        RECT 588.900 23.100 590.700 24.900 ;
        RECT 536.100 21.150 537.900 22.950 ;
        RECT 516.750 15.600 520.200 16.800 ;
        RECT 500.400 13.500 508.200 14.400 ;
        RECT 461.400 3.600 463.200 9.600 ;
        RECT 482.400 3.600 484.200 9.600 ;
        RECT 500.400 3.600 502.200 13.500 ;
        RECT 506.400 4.500 508.200 13.500 ;
        RECT 509.400 13.200 517.800 14.100 ;
        RECT 509.400 5.400 511.200 13.200 ;
        RECT 512.400 4.500 514.200 12.300 ;
        RECT 506.400 3.600 514.200 4.500 ;
        RECT 516.000 4.500 517.800 13.200 ;
        RECT 519.000 13.200 520.200 15.600 ;
        RECT 519.000 5.400 520.800 13.200 ;
        RECT 522.000 4.500 523.800 13.800 ;
        RECT 541.950 9.600 543.150 22.950 ;
        RECT 560.400 15.600 561.300 22.950 ;
        RECT 566.100 21.150 567.900 22.950 ;
        RECT 574.950 21.450 577.050 22.050 ;
        RECT 584.100 21.450 585.900 23.100 ;
        RECT 591.750 22.200 592.650 28.800 ;
        RECT 593.550 27.900 595.350 29.700 ;
        RECT 596.250 29.400 598.350 30.000 ;
        RECT 593.700 27.000 595.800 27.900 ;
        RECT 593.700 25.800 600.300 27.000 ;
        RECT 598.500 25.200 600.300 25.800 ;
        RECT 598.500 25.050 600.600 25.200 ;
        RECT 611.100 25.050 612.900 26.850 ;
        RECT 614.400 25.050 615.600 30.300 ;
        RECT 619.950 27.450 624.000 28.050 ;
        RECT 617.100 25.050 618.900 26.850 ;
        RECT 619.950 25.950 624.450 27.450 ;
        RECT 593.700 22.800 595.800 24.900 ;
        RECT 598.500 23.100 604.050 25.050 ;
        RECT 600.000 22.950 604.050 23.100 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 574.950 21.300 585.900 21.450 ;
        RECT 574.950 20.550 585.450 21.300 ;
        RECT 589.500 20.700 592.650 22.200 ;
        RECT 594.000 21.000 595.800 22.800 ;
        RECT 574.950 19.950 577.050 20.550 ;
        RECT 589.500 20.100 591.600 20.700 ;
        RECT 586.800 15.600 588.900 16.500 ;
        RECT 516.000 3.600 523.800 4.500 ;
        RECT 541.800 3.600 543.600 9.600 ;
        RECT 559.800 3.600 561.600 15.600 ;
        RECT 562.800 14.700 570.600 15.600 ;
        RECT 562.800 3.600 564.600 14.700 ;
        RECT 568.800 3.600 570.600 14.700 ;
        RECT 583.800 14.400 588.900 15.600 ;
        RECT 589.800 15.600 591.000 20.100 ;
        RECT 592.500 17.700 594.300 19.800 ;
        RECT 592.500 16.800 597.900 17.700 ;
        RECT 595.800 15.900 597.900 16.800 ;
        RECT 589.800 14.700 593.100 15.600 ;
        RECT 595.800 14.700 600.600 15.900 ;
        RECT 583.800 3.600 585.600 14.400 ;
        RECT 591.300 3.600 593.100 14.700 ;
        RECT 598.800 3.600 600.600 14.700 ;
        RECT 614.400 9.600 615.600 22.950 ;
        RECT 623.550 21.450 624.450 25.950 ;
        RECT 629.100 25.050 630.900 26.850 ;
        RECT 635.100 25.050 636.900 26.850 ;
        RECT 638.700 25.050 639.600 32.400 ;
        RECT 656.700 25.050 657.600 35.400 ;
        RECT 671.400 33.300 673.200 38.400 ;
        RECT 677.400 33.300 679.200 38.400 ;
        RECT 671.400 31.950 679.200 33.300 ;
        RECT 680.400 32.400 682.200 38.400 ;
        RECT 695.400 35.400 697.200 38.400 ;
        RECT 680.400 30.300 681.600 32.400 ;
        RECT 695.400 31.500 696.600 35.400 ;
        RECT 701.400 32.400 703.200 38.400 ;
        RECT 695.400 30.600 701.100 31.500 ;
        RECT 677.850 29.250 681.600 30.300 ;
        RECT 699.150 29.700 701.100 30.600 ;
        RECT 666.000 27.450 670.050 28.050 ;
        RECT 665.550 25.950 670.050 27.450 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 637.950 22.950 640.050 25.050 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 623.550 20.550 627.450 21.450 ;
        RECT 632.100 21.150 633.900 22.950 ;
        RECT 626.550 18.450 627.450 20.550 ;
        RECT 631.950 18.450 634.050 19.050 ;
        RECT 626.550 17.550 634.050 18.450 ;
        RECT 631.950 16.950 634.050 17.550 ;
        RECT 638.700 15.600 639.600 22.950 ;
        RECT 653.100 21.150 654.900 22.950 ;
        RECT 656.700 15.600 657.600 22.950 ;
        RECT 659.100 21.150 660.900 22.950 ;
        RECT 665.550 22.050 666.450 25.950 ;
        RECT 674.100 25.050 675.900 26.850 ;
        RECT 677.850 25.050 679.050 29.250 ;
        RECT 680.100 25.050 681.900 26.850 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 673.950 22.950 676.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 694.950 22.950 697.050 25.050 ;
        RECT 661.950 20.550 666.450 22.050 ;
        RECT 671.100 21.150 672.900 22.950 ;
        RECT 661.950 19.950 666.000 20.550 ;
        RECT 613.800 3.600 615.600 9.600 ;
        RECT 629.400 14.700 637.200 15.600 ;
        RECT 629.400 3.600 631.200 14.700 ;
        RECT 635.400 3.600 637.200 14.700 ;
        RECT 638.400 3.600 640.200 15.600 ;
        RECT 656.700 14.400 660.300 15.600 ;
        RECT 658.500 3.600 660.300 14.400 ;
        RECT 676.950 9.600 678.150 22.950 ;
        RECT 695.100 21.150 696.900 22.950 ;
        RECT 699.150 18.300 700.050 29.700 ;
        RECT 702.000 25.050 703.200 32.400 ;
        RECT 700.950 22.950 703.200 25.050 ;
        RECT 699.150 17.400 701.100 18.300 ;
        RECT 695.400 16.500 701.100 17.400 ;
        RECT 695.400 9.600 696.600 16.500 ;
        RECT 702.000 15.600 703.200 22.950 ;
        RECT 676.800 3.600 678.600 9.600 ;
        RECT 695.400 3.600 697.200 9.600 ;
        RECT 701.400 3.600 703.200 15.600 ;
        RECT 708.150 32.400 709.950 38.400 ;
        RECT 715.950 36.300 717.750 38.400 ;
        RECT 714.000 35.400 717.750 36.300 ;
        RECT 723.750 35.400 725.550 38.400 ;
        RECT 731.550 35.400 733.350 38.400 ;
        RECT 714.000 34.500 715.050 35.400 ;
        RECT 723.750 34.500 724.800 35.400 ;
        RECT 712.950 32.400 715.050 34.500 ;
        RECT 708.150 17.700 709.050 32.400 ;
        RECT 716.550 31.800 718.350 33.600 ;
        RECT 719.850 33.450 724.800 34.500 ;
        RECT 732.300 34.500 733.350 35.400 ;
        RECT 719.850 32.700 721.650 33.450 ;
        RECT 732.300 33.300 736.050 34.500 ;
        RECT 733.950 32.400 736.050 33.300 ;
        RECT 739.650 32.400 741.450 38.400 ;
        RECT 716.850 30.000 717.900 31.800 ;
        RECT 727.050 30.000 728.850 30.600 ;
        RECT 716.850 28.800 728.850 30.000 ;
        RECT 711.000 27.600 717.900 28.800 ;
        RECT 711.000 26.850 711.900 27.600 ;
        RECT 716.100 27.000 717.900 27.600 ;
        RECT 710.100 25.050 711.900 26.850 ;
        RECT 713.100 25.800 714.900 26.400 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 713.100 24.600 721.050 25.800 ;
        RECT 718.950 22.950 721.050 24.600 ;
        RECT 717.450 17.700 719.250 18.000 ;
        RECT 708.150 17.100 719.250 17.700 ;
        RECT 708.150 16.500 725.850 17.100 ;
        RECT 708.150 15.600 709.050 16.500 ;
        RECT 717.450 16.200 725.850 16.500 ;
        RECT 708.150 3.600 709.950 15.600 ;
        RECT 722.250 14.700 724.050 15.300 ;
        RECT 716.550 13.500 724.050 14.700 ;
        RECT 724.950 14.100 725.850 16.200 ;
        RECT 727.950 16.200 728.850 28.800 ;
        RECT 740.250 25.050 741.450 32.400 ;
        RECT 752.400 35.400 754.200 38.400 ;
        RECT 752.400 31.500 753.600 35.400 ;
        RECT 758.400 32.400 760.200 38.400 ;
        RECT 752.400 30.600 758.100 31.500 ;
        RECT 756.150 29.700 758.100 30.600 ;
        RECT 735.150 23.250 741.450 25.050 ;
        RECT 736.950 22.950 741.450 23.250 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 737.250 17.400 739.050 19.200 ;
        RECT 733.950 16.200 738.150 17.400 ;
        RECT 727.950 15.300 733.050 16.200 ;
        RECT 733.950 15.300 736.050 16.200 ;
        RECT 740.250 15.600 741.450 22.950 ;
        RECT 752.100 21.150 753.900 22.950 ;
        RECT 756.150 18.300 757.050 29.700 ;
        RECT 759.000 25.050 760.200 32.400 ;
        RECT 757.950 22.950 760.200 25.050 ;
        RECT 756.150 17.400 758.100 18.300 ;
        RECT 732.150 14.400 733.050 15.300 ;
        RECT 729.450 14.100 731.250 14.400 ;
        RECT 716.550 12.600 717.750 13.500 ;
        RECT 724.950 13.200 731.250 14.100 ;
        RECT 729.450 12.600 731.250 13.200 ;
        RECT 732.150 12.600 734.850 14.400 ;
        RECT 712.950 10.500 717.750 12.600 ;
        RECT 720.450 11.550 722.250 12.300 ;
        RECT 725.250 11.550 727.050 12.300 ;
        RECT 720.450 10.500 727.050 11.550 ;
        RECT 716.550 9.600 717.750 10.500 ;
        RECT 716.550 3.600 718.350 9.600 ;
        RECT 724.350 3.600 726.150 10.500 ;
        RECT 732.150 9.600 736.050 11.700 ;
        RECT 732.150 3.600 733.950 9.600 ;
        RECT 739.650 3.600 741.450 15.600 ;
        RECT 752.400 16.500 758.100 17.400 ;
        RECT 752.400 9.600 753.600 16.500 ;
        RECT 759.000 15.600 760.200 22.950 ;
        RECT 752.400 3.600 754.200 9.600 ;
        RECT 758.400 3.600 760.200 15.600 ;
        RECT 765.150 32.400 766.950 38.400 ;
        RECT 772.950 36.300 774.750 38.400 ;
        RECT 771.000 35.400 774.750 36.300 ;
        RECT 780.750 35.400 782.550 38.400 ;
        RECT 788.550 35.400 790.350 38.400 ;
        RECT 771.000 34.500 772.050 35.400 ;
        RECT 780.750 34.500 781.800 35.400 ;
        RECT 769.950 32.400 772.050 34.500 ;
        RECT 765.150 17.700 766.050 32.400 ;
        RECT 773.550 31.800 775.350 33.600 ;
        RECT 776.850 33.450 781.800 34.500 ;
        RECT 789.300 34.500 790.350 35.400 ;
        RECT 776.850 32.700 778.650 33.450 ;
        RECT 789.300 33.300 793.050 34.500 ;
        RECT 790.950 32.400 793.050 33.300 ;
        RECT 796.650 32.400 798.450 38.400 ;
        RECT 773.850 30.000 774.900 31.800 ;
        RECT 784.050 30.000 785.850 30.600 ;
        RECT 773.850 28.800 785.850 30.000 ;
        RECT 768.000 27.600 774.900 28.800 ;
        RECT 768.000 26.850 768.900 27.600 ;
        RECT 773.100 27.000 774.900 27.600 ;
        RECT 767.100 25.050 768.900 26.850 ;
        RECT 770.100 25.800 771.900 26.400 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 770.100 24.600 778.050 25.800 ;
        RECT 775.950 22.950 778.050 24.600 ;
        RECT 774.450 17.700 776.250 18.000 ;
        RECT 765.150 17.100 776.250 17.700 ;
        RECT 765.150 16.500 782.850 17.100 ;
        RECT 765.150 15.600 766.050 16.500 ;
        RECT 774.450 16.200 782.850 16.500 ;
        RECT 765.150 3.600 766.950 15.600 ;
        RECT 779.250 14.700 781.050 15.300 ;
        RECT 773.550 13.500 781.050 14.700 ;
        RECT 781.950 14.100 782.850 16.200 ;
        RECT 784.950 16.200 785.850 28.800 ;
        RECT 797.250 25.050 798.450 32.400 ;
        RECT 806.400 35.400 808.200 38.400 ;
        RECT 806.400 31.500 807.600 35.400 ;
        RECT 812.400 32.400 814.200 38.400 ;
        RECT 806.400 30.600 812.100 31.500 ;
        RECT 810.150 29.700 812.100 30.600 ;
        RECT 792.150 23.250 798.450 25.050 ;
        RECT 793.950 22.950 798.450 23.250 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 794.250 17.400 796.050 19.200 ;
        RECT 790.950 16.200 795.150 17.400 ;
        RECT 784.950 15.300 790.050 16.200 ;
        RECT 790.950 15.300 793.050 16.200 ;
        RECT 797.250 15.600 798.450 22.950 ;
        RECT 806.100 21.150 807.900 22.950 ;
        RECT 810.150 18.300 811.050 29.700 ;
        RECT 813.000 25.050 814.200 32.400 ;
        RECT 827.400 35.400 829.200 38.400 ;
        RECT 827.400 31.500 828.600 35.400 ;
        RECT 833.400 32.400 835.200 38.400 ;
        RECT 827.400 30.600 833.100 31.500 ;
        RECT 831.150 29.700 833.100 30.600 ;
        RECT 811.950 22.950 814.200 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 810.150 17.400 812.100 18.300 ;
        RECT 789.150 14.400 790.050 15.300 ;
        RECT 786.450 14.100 788.250 14.400 ;
        RECT 773.550 12.600 774.750 13.500 ;
        RECT 781.950 13.200 788.250 14.100 ;
        RECT 786.450 12.600 788.250 13.200 ;
        RECT 789.150 12.600 791.850 14.400 ;
        RECT 769.950 10.500 774.750 12.600 ;
        RECT 777.450 11.550 779.250 12.300 ;
        RECT 782.250 11.550 784.050 12.300 ;
        RECT 777.450 10.500 784.050 11.550 ;
        RECT 773.550 9.600 774.750 10.500 ;
        RECT 773.550 3.600 775.350 9.600 ;
        RECT 781.350 3.600 783.150 10.500 ;
        RECT 789.150 9.600 793.050 11.700 ;
        RECT 789.150 3.600 790.950 9.600 ;
        RECT 796.650 3.600 798.450 15.600 ;
        RECT 806.400 16.500 812.100 17.400 ;
        RECT 806.400 9.600 807.600 16.500 ;
        RECT 813.000 15.600 814.200 22.950 ;
        RECT 827.100 21.150 828.900 22.950 ;
        RECT 831.150 18.300 832.050 29.700 ;
        RECT 834.000 25.050 835.200 32.400 ;
        RECT 832.950 22.950 835.200 25.050 ;
        RECT 831.150 17.400 833.100 18.300 ;
        RECT 806.400 3.600 808.200 9.600 ;
        RECT 812.400 3.600 814.200 15.600 ;
        RECT 827.400 16.500 833.100 17.400 ;
        RECT 827.400 9.600 828.600 16.500 ;
        RECT 834.000 15.600 835.200 22.950 ;
        RECT 827.400 3.600 829.200 9.600 ;
        RECT 833.400 3.600 835.200 15.600 ;
        RECT 850.800 32.400 852.600 38.400 ;
        RECT 856.800 35.400 858.600 38.400 ;
        RECT 850.800 25.050 852.000 32.400 ;
        RECT 857.400 31.500 858.600 35.400 ;
        RECT 852.900 30.600 858.600 31.500 ;
        RECT 866.400 35.400 868.200 38.400 ;
        RECT 866.400 31.500 867.600 35.400 ;
        RECT 872.400 32.400 874.200 38.400 ;
        RECT 866.400 30.600 872.100 31.500 ;
        RECT 852.900 29.700 854.850 30.600 ;
        RECT 850.800 22.950 853.050 25.050 ;
        RECT 850.800 15.600 852.000 22.950 ;
        RECT 853.950 18.300 854.850 29.700 ;
        RECT 870.150 29.700 872.100 30.600 ;
        RECT 856.950 22.950 859.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 857.100 21.150 858.900 22.950 ;
        RECT 866.100 21.150 867.900 22.950 ;
        RECT 852.900 17.400 854.850 18.300 ;
        RECT 870.150 18.300 871.050 29.700 ;
        RECT 873.000 25.050 874.200 32.400 ;
        RECT 890.400 31.200 892.200 38.400 ;
        RECT 890.400 30.300 894.600 31.200 ;
        RECT 890.100 25.050 891.900 26.850 ;
        RECT 893.400 25.050 894.600 30.300 ;
        RECT 896.100 25.050 897.900 26.850 ;
        RECT 871.950 22.950 874.200 25.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 892.950 22.950 895.050 25.050 ;
        RECT 895.950 22.950 898.050 25.050 ;
        RECT 870.150 17.400 872.100 18.300 ;
        RECT 852.900 16.500 858.600 17.400 ;
        RECT 850.800 3.600 852.600 15.600 ;
        RECT 857.400 9.600 858.600 16.500 ;
        RECT 856.800 3.600 858.600 9.600 ;
        RECT 866.400 16.500 872.100 17.400 ;
        RECT 866.400 9.600 867.600 16.500 ;
        RECT 873.000 15.600 874.200 22.950 ;
        RECT 866.400 3.600 868.200 9.600 ;
        RECT 872.400 3.600 874.200 15.600 ;
        RECT 893.400 9.600 894.600 22.950 ;
        RECT 895.950 18.450 898.050 19.050 ;
        RECT 910.950 18.450 913.050 19.050 ;
        RECT 895.950 17.550 913.050 18.450 ;
        RECT 895.950 16.950 898.050 17.550 ;
        RECT 910.950 16.950 913.050 17.550 ;
        RECT 892.800 3.600 894.600 9.600 ;
      LAYER metal2 ;
        RECT 664.950 934.950 667.050 937.050 ;
        RECT 847.950 934.950 850.050 937.050 ;
        RECT 43.950 931.950 46.050 934.050 ;
        RECT 97.950 931.950 100.050 934.050 ;
        RECT 136.950 931.950 139.050 934.050 ;
        RECT 652.950 931.950 655.050 934.050 ;
        RECT 13.950 922.950 16.050 925.050 ;
        RECT 37.950 922.950 40.050 925.050 ;
        RECT 14.400 916.050 15.600 922.950 ;
        RECT 25.950 917.100 28.050 919.200 ;
        RECT 31.950 917.100 34.050 919.200 ;
        RECT 13.950 913.950 16.050 916.050 ;
        RECT 16.950 913.950 19.050 916.050 ;
        RECT 17.400 889.050 18.600 913.950 ;
        RECT 26.400 912.600 27.600 917.100 ;
        RECT 32.400 916.050 33.600 917.100 ;
        RECT 38.400 916.050 39.600 922.950 ;
        RECT 44.400 919.050 45.600 931.950 ;
        RECT 76.950 925.950 79.050 928.050 ;
        RECT 58.950 922.950 61.050 925.050 ;
        RECT 43.800 916.950 45.900 919.050 ;
        RECT 46.950 917.100 49.050 919.200 ;
        RECT 52.950 917.100 55.050 919.200 ;
        RECT 31.950 913.950 34.050 916.050 ;
        RECT 34.950 913.950 37.050 916.050 ;
        RECT 37.950 913.950 40.050 916.050 ;
        RECT 40.950 913.950 43.050 916.050 ;
        RECT 35.400 912.900 36.600 913.950 ;
        RECT 41.400 912.900 42.600 913.950 ;
        RECT 47.400 913.050 48.600 917.100 ;
        RECT 53.400 916.050 54.600 917.100 ;
        RECT 59.400 916.050 60.600 922.950 ;
        RECT 77.400 919.200 78.600 925.950 ;
        RECT 88.950 919.950 91.050 922.050 ;
        RECT 76.950 917.100 79.050 919.200 ;
        RECT 77.400 916.050 78.600 917.100 ;
        RECT 52.950 913.950 55.050 916.050 ;
        RECT 55.950 913.950 58.050 916.050 ;
        RECT 58.950 913.950 61.050 916.050 ;
        RECT 61.950 913.950 64.050 916.050 ;
        RECT 76.950 913.950 79.050 916.050 ;
        RECT 79.950 913.950 82.050 916.050 ;
        RECT 26.400 911.400 30.600 912.600 ;
        RECT 16.950 885.000 19.050 889.050 ;
        RECT 17.400 883.050 18.600 885.000 ;
        RECT 22.950 884.100 25.050 886.200 ;
        RECT 29.400 886.050 30.600 911.400 ;
        RECT 34.950 910.800 37.050 912.900 ;
        RECT 40.950 910.800 43.050 912.900 ;
        RECT 46.950 910.950 49.050 913.050 ;
        RECT 41.400 886.200 42.600 910.800 ;
        RECT 56.400 895.050 57.600 913.950 ;
        RECT 62.400 912.900 63.600 913.950 ;
        RECT 61.950 910.800 64.050 912.900 ;
        RECT 70.950 910.800 73.050 912.900 ;
        RECT 55.950 892.950 58.050 895.050 ;
        RECT 23.400 883.050 24.600 884.100 ;
        RECT 28.950 883.950 31.050 886.050 ;
        RECT 31.950 883.950 34.050 886.050 ;
        RECT 40.950 884.100 43.050 886.200 ;
        RECT 49.950 884.100 52.050 886.200 ;
        RECT 58.950 884.100 61.050 889.050 ;
        RECT 64.950 884.100 67.050 886.200 ;
        RECT 13.950 880.950 16.050 883.050 ;
        RECT 16.950 880.950 19.050 883.050 ;
        RECT 19.950 880.950 22.050 883.050 ;
        RECT 22.950 880.950 25.050 883.050 ;
        RECT 25.950 880.950 28.050 883.050 ;
        RECT 14.400 874.050 15.600 880.950 ;
        RECT 13.950 871.950 16.050 874.050 ;
        RECT 14.400 844.050 15.600 871.950 ;
        RECT 13.950 841.950 16.050 844.050 ;
        RECT 10.950 839.100 13.050 841.200 ;
        RECT 11.400 838.050 12.600 839.100 ;
        RECT 10.950 835.950 13.050 838.050 ;
        RECT 13.950 835.950 16.050 838.050 ;
        RECT 4.950 826.950 7.050 829.050 ;
        RECT 1.950 806.100 4.050 808.200 ;
        RECT 2.400 787.050 3.600 806.100 ;
        RECT 1.950 784.950 4.050 787.050 ;
        RECT 5.400 756.900 6.600 826.950 ;
        RECT 14.400 823.050 15.600 835.950 ;
        RECT 20.400 829.050 21.600 880.950 ;
        RECT 26.400 868.050 27.600 880.950 ;
        RECT 28.950 877.950 31.050 880.050 ;
        RECT 29.400 874.050 30.600 877.950 ;
        RECT 28.950 871.950 31.050 874.050 ;
        RECT 25.950 865.950 28.050 868.050 ;
        RECT 22.950 856.950 25.050 859.050 ;
        RECT 19.950 826.950 22.050 829.050 ;
        RECT 13.950 820.950 16.050 823.050 ;
        RECT 19.950 822.600 22.050 823.050 ;
        RECT 23.400 822.600 24.600 856.950 ;
        RECT 32.400 850.050 33.600 883.950 ;
        RECT 41.400 883.050 42.600 884.100 ;
        RECT 37.950 880.950 40.050 883.050 ;
        RECT 40.950 880.950 43.050 883.050 ;
        RECT 43.950 880.950 46.050 883.050 ;
        RECT 38.400 868.050 39.600 880.950 ;
        RECT 44.400 879.900 45.600 880.950 ;
        RECT 43.950 877.800 46.050 879.900 ;
        RECT 37.950 865.950 40.050 868.050 ;
        RECT 44.400 856.050 45.600 877.800 ;
        RECT 50.400 877.050 51.600 884.100 ;
        RECT 59.400 883.050 60.600 884.100 ;
        RECT 65.400 883.050 66.600 884.100 ;
        RECT 55.950 880.950 58.050 883.050 ;
        RECT 58.950 880.950 61.050 883.050 ;
        RECT 61.950 880.950 64.050 883.050 ;
        RECT 64.950 880.950 67.050 883.050 ;
        RECT 49.950 874.950 52.050 877.050 ;
        RECT 56.400 874.050 57.600 880.950 ;
        RECT 62.400 879.900 63.600 880.950 ;
        RECT 61.950 877.800 64.050 879.900 ;
        RECT 58.950 874.950 61.050 877.050 ;
        RECT 55.950 871.950 58.050 874.050 ;
        RECT 43.950 853.950 46.050 856.050 ;
        RECT 31.950 847.950 34.050 850.050 ;
        RECT 40.950 847.950 43.050 850.050 ;
        RECT 25.950 840.600 30.000 841.050 ;
        RECT 25.950 838.950 30.600 840.600 ;
        RECT 34.950 839.100 37.050 841.200 ;
        RECT 29.400 838.050 30.600 838.950 ;
        RECT 35.400 838.050 36.600 839.100 ;
        RECT 28.950 835.950 31.050 838.050 ;
        RECT 31.950 835.950 34.050 838.050 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 32.400 834.900 33.600 835.950 ;
        RECT 31.950 832.800 34.050 834.900 ;
        RECT 19.950 821.400 24.600 822.600 ;
        RECT 19.950 820.950 22.050 821.400 ;
        RECT 7.950 814.950 10.050 817.050 ;
        RECT 8.400 763.200 9.600 814.950 ;
        RECT 20.400 808.200 21.600 820.950 ;
        RECT 28.950 817.950 31.050 820.050 ;
        RECT 19.950 806.100 22.050 808.200 ;
        RECT 20.400 805.050 21.600 806.100 ;
        RECT 13.950 802.950 16.050 805.050 ;
        RECT 19.950 802.950 22.050 805.050 ;
        RECT 22.950 802.950 25.050 805.050 ;
        RECT 14.400 793.050 15.600 802.950 ;
        RECT 23.400 801.000 24.600 802.950 ;
        RECT 22.950 796.950 25.050 801.000 ;
        RECT 29.400 799.050 30.600 817.950 ;
        RECT 37.950 814.950 40.050 817.050 ;
        RECT 31.950 808.950 34.050 811.050 ;
        RECT 32.400 801.900 33.600 808.950 ;
        RECT 38.400 805.050 39.600 814.950 ;
        RECT 41.400 811.050 42.600 847.950 ;
        RECT 43.950 839.100 46.050 841.200 ;
        RECT 49.950 839.100 52.050 841.200 ;
        RECT 55.950 840.000 58.050 844.050 ;
        RECT 59.400 841.050 60.600 874.950 ;
        RECT 71.400 874.050 72.600 910.800 ;
        RECT 80.400 907.050 81.600 913.950 ;
        RECT 89.400 913.050 90.600 919.950 ;
        RECT 98.400 916.050 99.600 931.950 ;
        RECT 112.950 928.950 115.050 931.050 ;
        RECT 109.950 925.950 112.050 928.050 ;
        RECT 103.950 917.100 106.050 919.200 ;
        RECT 110.400 918.600 111.600 925.950 ;
        RECT 113.400 922.050 114.600 928.950 ;
        RECT 130.950 922.950 133.050 925.050 ;
        RECT 112.950 919.950 115.050 922.050 ;
        RECT 110.400 917.400 114.600 918.600 ;
        RECT 118.950 918.000 121.050 922.050 ;
        RECT 127.950 919.950 130.050 922.050 ;
        RECT 104.400 916.050 105.600 917.100 ;
        RECT 113.400 916.050 114.600 917.400 ;
        RECT 119.400 916.050 120.600 918.000 ;
        RECT 94.950 913.950 97.050 916.050 ;
        RECT 97.950 913.950 100.050 916.050 ;
        RECT 100.950 913.950 103.050 916.050 ;
        RECT 103.950 913.950 106.050 916.050 ;
        RECT 112.950 913.950 115.050 916.050 ;
        RECT 115.950 913.950 118.050 916.050 ;
        RECT 118.950 913.950 121.050 916.050 ;
        RECT 121.950 913.950 124.050 916.050 ;
        RECT 88.950 910.950 91.050 913.050 ;
        RECT 95.400 912.900 96.600 913.950 ;
        RECT 101.400 912.900 102.600 913.950 ;
        RECT 116.400 912.900 117.600 913.950 ;
        RECT 122.400 912.900 123.600 913.950 ;
        RECT 94.950 910.800 97.050 912.900 ;
        RECT 100.950 910.800 103.050 912.900 ;
        RECT 115.950 910.800 118.050 912.900 ;
        RECT 121.950 910.800 124.050 912.900 ;
        RECT 116.400 907.050 117.600 910.800 ;
        RECT 128.400 910.050 129.600 919.950 ;
        RECT 131.400 916.050 132.600 922.950 ;
        RECT 137.400 916.050 138.600 931.950 ;
        RECT 214.950 928.950 217.050 931.050 ;
        RECT 298.950 928.950 301.050 931.050 ;
        RECT 310.950 928.950 313.050 931.050 ;
        RECT 334.950 928.950 337.050 931.050 ;
        RECT 163.950 922.950 166.050 925.050 ;
        RECT 178.950 922.950 181.050 925.050 ;
        RECT 205.950 922.950 208.050 925.050 ;
        RECT 142.950 917.100 145.050 919.200 ;
        RECT 151.950 917.100 154.050 919.200 ;
        RECT 143.400 916.050 144.600 917.100 ;
        RECT 130.950 913.950 133.050 916.050 ;
        RECT 136.950 913.950 139.050 916.050 ;
        RECT 139.950 913.950 142.050 916.050 ;
        RECT 142.950 913.950 145.050 916.050 ;
        RECT 145.950 913.950 148.050 916.050 ;
        RECT 140.400 912.900 141.600 913.950 ;
        RECT 139.950 910.800 142.050 912.900 ;
        RECT 127.950 907.950 130.050 910.050 ;
        RECT 79.950 904.950 82.050 907.050 ;
        RECT 94.950 904.950 97.050 907.050 ;
        RECT 115.950 904.950 118.050 907.050 ;
        RECT 88.950 898.950 91.050 901.050 ;
        RECT 73.950 883.950 76.050 886.050 ;
        RECT 82.950 885.000 85.050 889.050 ;
        RECT 70.950 871.950 73.050 874.050 ;
        RECT 70.950 856.950 73.050 859.050 ;
        RECT 44.400 835.050 45.600 839.100 ;
        RECT 50.400 838.050 51.600 839.100 ;
        RECT 56.400 838.050 57.600 840.000 ;
        RECT 58.950 838.950 61.050 841.050 ;
        RECT 64.950 839.100 67.050 844.050 ;
        RECT 65.400 838.050 66.600 839.100 ;
        RECT 71.400 838.050 72.600 856.950 ;
        RECT 74.400 843.600 75.600 883.950 ;
        RECT 83.400 883.050 84.600 885.000 ;
        RECT 89.400 883.050 90.600 898.950 ;
        RECT 95.400 898.050 96.600 904.950 ;
        RECT 118.950 901.950 121.050 904.050 ;
        RECT 119.400 898.050 120.600 901.950 ;
        RECT 128.400 901.050 129.600 907.950 ;
        RECT 146.400 904.050 147.600 913.950 ;
        RECT 145.950 901.950 148.050 904.050 ;
        RECT 127.950 898.950 130.050 901.050 ;
        RECT 152.400 898.050 153.600 917.100 ;
        RECT 164.400 916.050 165.600 922.950 ;
        RECT 169.950 917.100 172.050 919.200 ;
        RECT 170.400 916.050 171.600 917.100 ;
        RECT 160.950 913.950 163.050 916.050 ;
        RECT 163.950 913.950 166.050 916.050 ;
        RECT 166.950 913.950 169.050 916.050 ;
        RECT 169.950 913.950 172.050 916.050 ;
        RECT 95.400 896.400 100.050 898.050 ;
        RECT 96.000 895.950 100.050 896.400 ;
        RECT 118.950 895.950 121.050 898.050 ;
        RECT 151.950 895.950 154.050 898.050 ;
        RECT 94.950 892.950 97.050 895.050 ;
        RECT 79.950 880.950 82.050 883.050 ;
        RECT 82.950 880.950 85.050 883.050 ;
        RECT 85.950 880.950 88.050 883.050 ;
        RECT 88.950 880.950 91.050 883.050 ;
        RECT 80.400 879.900 81.600 880.950 ;
        RECT 86.400 879.900 87.600 880.950 ;
        RECT 79.950 877.800 82.050 879.900 ;
        RECT 85.950 877.800 88.050 879.900 ;
        RECT 91.950 877.800 94.050 879.900 ;
        RECT 92.400 874.050 93.600 877.800 ;
        RECT 82.950 871.950 85.050 874.050 ;
        RECT 91.950 871.950 94.050 874.050 ;
        RECT 74.400 843.000 78.600 843.600 ;
        RECT 74.400 842.400 79.050 843.000 ;
        RECT 76.950 838.950 79.050 842.400 ;
        RECT 79.950 839.100 82.050 841.200 ;
        RECT 49.950 835.950 52.050 838.050 ;
        RECT 52.950 835.950 55.050 838.050 ;
        RECT 55.950 835.950 58.050 838.050 ;
        RECT 64.950 835.950 67.050 838.050 ;
        RECT 67.950 835.950 70.050 838.050 ;
        RECT 70.950 835.950 73.050 838.050 ;
        RECT 73.950 835.950 76.050 838.050 ;
        RECT 43.950 832.950 46.050 835.050 ;
        RECT 53.400 834.900 54.600 835.950 ;
        RECT 44.400 820.050 45.600 832.950 ;
        RECT 52.950 832.800 55.050 834.900 ;
        RECT 58.950 832.950 61.050 835.050 ;
        RECT 59.400 823.050 60.600 832.950 ;
        RECT 68.400 823.050 69.600 835.950 ;
        RECT 74.400 835.050 75.600 835.950 ;
        RECT 74.400 833.400 79.050 835.050 ;
        RECT 75.000 832.950 79.050 833.400 ;
        RECT 80.400 832.050 81.600 839.100 ;
        RECT 83.400 835.050 84.600 871.950 ;
        RECT 91.950 856.950 94.050 859.050 ;
        RECT 85.950 844.950 88.050 847.050 ;
        RECT 82.950 832.950 85.050 835.050 ;
        RECT 70.950 829.950 73.050 832.050 ;
        RECT 79.950 829.950 82.050 832.050 ;
        RECT 52.950 820.950 55.050 823.050 ;
        RECT 58.950 820.950 61.050 823.050 ;
        RECT 67.950 820.950 70.050 823.050 ;
        RECT 43.950 817.950 46.050 820.050 ;
        RECT 43.950 811.950 46.050 814.050 ;
        RECT 40.950 808.950 43.050 811.050 ;
        RECT 44.400 805.050 45.600 811.950 ;
        RECT 37.950 802.950 40.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 43.950 802.950 46.050 805.050 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 41.400 801.900 42.600 802.950 ;
        RECT 31.950 799.800 34.050 801.900 ;
        RECT 40.950 799.800 43.050 801.900 ;
        RECT 28.950 796.950 31.050 799.050 ;
        RECT 47.400 793.050 48.600 802.950 ;
        RECT 13.950 790.950 16.050 793.050 ;
        RECT 46.800 790.950 48.900 793.050 ;
        RECT 49.950 790.950 52.050 793.050 ;
        RECT 28.950 781.950 31.050 784.050 ;
        RECT 13.950 769.950 16.050 772.050 ;
        RECT 7.950 761.100 10.050 763.200 ;
        RECT 14.400 760.050 15.600 769.950 ;
        RECT 19.950 761.100 22.050 763.200 ;
        RECT 20.400 760.050 21.600 761.100 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 22.950 757.950 25.050 760.050 ;
        RECT 4.950 754.800 7.050 756.900 ;
        RECT 17.400 756.000 18.600 757.950 ;
        RECT 23.400 756.900 24.600 757.950 ;
        RECT 16.950 751.950 19.050 756.000 ;
        RECT 22.950 754.800 25.050 756.900 ;
        RECT 25.950 732.600 28.050 733.050 ;
        RECT 29.400 732.600 30.600 781.950 ;
        RECT 50.400 772.050 51.600 790.950 ;
        RECT 53.400 784.050 54.600 820.950 ;
        RECT 61.950 811.950 64.050 814.050 ;
        RECT 62.400 805.050 63.600 811.950 ;
        RECT 58.950 802.950 61.050 805.050 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 64.950 802.950 67.050 805.050 ;
        RECT 59.400 796.050 60.600 802.950 ;
        RECT 61.950 796.950 64.050 799.050 ;
        RECT 58.950 793.950 61.050 796.050 ;
        RECT 52.950 781.950 55.050 784.050 ;
        RECT 49.950 769.950 52.050 772.050 ;
        RECT 37.950 761.100 40.050 763.200 ;
        RECT 43.950 761.100 46.050 763.200 ;
        RECT 38.400 760.050 39.600 761.100 ;
        RECT 44.400 760.050 45.600 761.100 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 43.950 757.950 46.050 760.050 ;
        RECT 35.400 756.900 36.600 757.950 ;
        RECT 34.950 754.800 37.050 756.900 ;
        RECT 41.400 748.050 42.600 757.950 ;
        RECT 40.950 745.950 43.050 748.050 ;
        RECT 25.950 731.400 30.600 732.600 ;
        RECT 25.950 730.950 28.050 731.400 ;
        RECT 16.950 728.100 19.050 730.200 ;
        RECT 17.400 727.050 18.600 728.100 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 19.950 724.950 22.050 727.050 ;
        RECT 14.400 712.050 15.600 724.950 ;
        RECT 20.400 723.000 21.600 724.950 ;
        RECT 19.950 718.950 22.050 723.000 ;
        RECT 22.950 721.950 25.050 724.050 ;
        RECT 13.950 709.950 16.050 712.050 ;
        RECT 1.950 697.950 4.050 700.050 ;
        RECT 2.400 648.600 3.600 697.950 ;
        RECT 10.950 688.950 13.050 691.050 ;
        RECT 11.400 685.200 12.600 688.950 ;
        RECT 23.400 685.200 24.600 721.950 ;
        RECT 26.400 721.050 27.600 730.950 ;
        RECT 34.950 729.000 37.050 733.050 ;
        RECT 35.400 727.050 36.600 729.000 ;
        RECT 40.950 728.100 43.050 730.200 ;
        RECT 41.400 727.050 42.600 728.100 ;
        RECT 46.950 727.950 49.050 730.050 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 37.950 724.950 40.050 727.050 ;
        RECT 40.950 724.950 43.050 727.050 ;
        RECT 25.950 718.950 28.050 721.050 ;
        RECT 4.950 683.100 7.050 685.200 ;
        RECT 10.950 683.100 13.050 685.200 ;
        RECT 16.950 683.100 19.050 685.200 ;
        RECT 22.800 683.100 24.900 685.200 ;
        RECT 26.400 685.050 27.600 718.950 ;
        RECT 32.400 712.050 33.600 724.950 ;
        RECT 38.400 718.050 39.600 724.950 ;
        RECT 47.400 723.900 48.600 727.950 ;
        RECT 46.950 721.800 49.050 723.900 ;
        RECT 50.400 720.600 51.600 769.950 ;
        RECT 52.950 763.950 55.050 766.050 ;
        RECT 53.400 754.050 54.600 763.950 ;
        RECT 62.400 760.050 63.600 796.950 ;
        RECT 65.400 790.050 66.600 802.950 ;
        RECT 71.400 801.600 72.600 829.950 ;
        RECT 82.950 829.800 85.050 831.900 ;
        RECT 83.400 814.050 84.600 829.800 ;
        RECT 82.950 811.950 85.050 814.050 ;
        RECT 76.950 806.100 79.050 808.200 ;
        RECT 77.400 805.050 78.600 806.100 ;
        RECT 83.400 805.050 84.600 811.950 ;
        RECT 86.400 811.050 87.600 844.950 ;
        RECT 92.400 843.600 93.600 856.950 ;
        RECT 95.400 847.050 96.600 892.950 ;
        RECT 161.400 892.050 162.600 913.950 ;
        RECT 167.400 912.900 168.600 913.950 ;
        RECT 166.950 910.800 169.050 912.900 ;
        RECT 179.400 898.050 180.600 922.950 ;
        RECT 184.950 917.100 187.050 919.200 ;
        RECT 199.950 917.100 202.050 919.200 ;
        RECT 185.400 916.050 186.600 917.100 ;
        RECT 200.400 916.050 201.600 917.100 ;
        RECT 206.400 916.050 207.600 922.950 ;
        RECT 184.950 913.950 187.050 916.050 ;
        RECT 187.950 913.950 190.050 916.050 ;
        RECT 199.950 913.950 202.050 916.050 ;
        RECT 202.950 913.950 205.050 916.050 ;
        RECT 205.950 913.950 208.050 916.050 ;
        RECT 208.950 913.950 211.050 916.050 ;
        RECT 188.400 912.000 189.600 913.950 ;
        RECT 187.950 907.950 190.050 912.000 ;
        RECT 199.950 907.950 202.050 910.050 ;
        RECT 178.950 895.950 181.050 898.050 ;
        RECT 148.950 889.950 151.050 892.050 ;
        RECT 160.950 889.950 163.050 892.050 ;
        RECT 109.950 884.100 112.050 886.200 ;
        RECT 110.400 883.050 111.600 884.100 ;
        RECT 121.950 883.950 124.050 886.050 ;
        RECT 133.950 884.100 136.050 886.200 ;
        RECT 139.950 884.100 142.050 886.200 ;
        RECT 106.950 880.950 109.050 883.050 ;
        RECT 109.950 880.950 112.050 883.050 ;
        RECT 115.950 880.950 118.050 883.050 ;
        RECT 107.400 879.000 108.600 880.950 ;
        RECT 106.950 874.950 109.050 879.000 ;
        RECT 116.400 871.050 117.600 880.950 ;
        RECT 106.950 868.950 109.050 871.050 ;
        RECT 115.950 868.950 118.050 871.050 ;
        RECT 94.950 844.950 97.050 847.050 ;
        RECT 92.400 842.400 96.600 843.600 ;
        RECT 95.400 838.050 96.600 842.400 ;
        RECT 100.950 839.100 103.050 841.200 ;
        RECT 101.400 838.050 102.600 839.100 ;
        RECT 91.950 835.950 94.050 838.050 ;
        RECT 94.950 835.950 97.050 838.050 ;
        RECT 97.950 835.950 100.050 838.050 ;
        RECT 100.950 835.950 103.050 838.050 ;
        RECT 92.400 834.900 93.600 835.950 ;
        RECT 91.950 832.800 94.050 834.900 ;
        RECT 98.400 823.050 99.600 835.950 ;
        RECT 107.400 835.050 108.600 868.950 ;
        RECT 122.400 856.050 123.600 883.950 ;
        RECT 134.400 883.050 135.600 884.100 ;
        RECT 140.400 883.050 141.600 884.100 ;
        RECT 130.950 880.950 133.050 883.050 ;
        RECT 133.950 880.950 136.050 883.050 ;
        RECT 136.950 880.950 139.050 883.050 ;
        RECT 139.950 880.950 142.050 883.050 ;
        RECT 121.950 853.950 124.050 856.050 ;
        RECT 127.950 847.950 130.050 850.050 ;
        RECT 118.950 843.600 121.050 847.050 ;
        RECT 116.400 843.000 121.050 843.600 ;
        RECT 116.400 842.400 120.600 843.000 ;
        RECT 116.400 838.050 117.600 842.400 ;
        RECT 121.950 839.100 124.050 841.200 ;
        RECT 122.400 838.050 123.600 839.100 ;
        RECT 128.400 838.050 129.600 847.950 ;
        RECT 112.950 835.950 115.050 838.050 ;
        RECT 115.950 835.950 118.050 838.050 ;
        RECT 118.950 835.950 121.050 838.050 ;
        RECT 121.950 835.950 124.050 838.050 ;
        RECT 127.950 835.950 130.050 838.050 ;
        RECT 106.950 832.950 109.050 835.050 ;
        RECT 113.400 834.900 114.600 835.950 ;
        RECT 119.400 834.900 120.600 835.950 ;
        RECT 112.950 832.800 115.050 834.900 ;
        RECT 118.950 832.800 121.050 834.900 ;
        RECT 131.400 829.050 132.600 880.950 ;
        RECT 137.400 879.000 138.600 880.950 ;
        RECT 136.950 874.950 139.050 879.000 ;
        RECT 136.950 839.100 139.050 841.200 ;
        RECT 137.400 838.050 138.600 839.100 ;
        RECT 136.950 835.950 139.050 838.050 ;
        RECT 139.950 835.950 142.050 838.050 ;
        RECT 140.400 829.050 141.600 835.950 ;
        RECT 130.950 826.950 133.050 829.050 ;
        RECT 139.950 826.950 142.050 829.050 ;
        RECT 97.950 820.950 100.050 823.050 ;
        RECT 149.400 817.050 150.600 889.950 ;
        RECT 157.950 884.100 160.050 886.200 ;
        RECT 169.950 884.100 172.050 886.200 ;
        RECT 173.400 884.400 180.600 885.600 ;
        RECT 184.950 885.000 187.050 889.050 ;
        RECT 158.400 883.050 159.600 884.100 ;
        RECT 154.950 880.950 157.050 883.050 ;
        RECT 157.950 880.950 160.050 883.050 ;
        RECT 163.950 880.950 166.050 883.050 ;
        RECT 155.400 879.000 156.600 880.950 ;
        RECT 154.950 874.950 157.050 879.000 ;
        RECT 164.400 853.050 165.600 880.950 ;
        RECT 163.950 850.950 166.050 853.050 ;
        RECT 154.950 844.950 157.050 847.050 ;
        RECT 155.400 838.050 156.600 844.950 ;
        RECT 164.400 838.050 165.600 850.950 ;
        RECT 170.400 844.050 171.600 884.100 ;
        RECT 173.400 853.050 174.600 884.400 ;
        RECT 179.400 883.050 180.600 884.400 ;
        RECT 185.400 883.050 186.600 885.000 ;
        RECT 193.950 884.100 196.050 886.200 ;
        RECT 194.400 883.050 195.600 884.100 ;
        RECT 200.400 883.050 201.600 907.950 ;
        RECT 203.400 901.050 204.600 913.950 ;
        RECT 209.400 904.050 210.600 913.950 ;
        RECT 215.400 912.900 216.600 928.950 ;
        RECT 247.950 922.950 250.050 925.050 ;
        RECT 265.950 922.950 268.050 925.050 ;
        RECT 280.950 922.950 283.050 925.050 ;
        RECT 220.950 917.100 223.050 919.200 ;
        RECT 226.950 917.100 229.050 919.200 ;
        RECT 235.950 917.100 238.050 919.200 ;
        RECT 221.400 916.050 222.600 917.100 ;
        RECT 227.400 916.050 228.600 917.100 ;
        RECT 220.950 913.950 223.050 916.050 ;
        RECT 223.950 913.950 226.050 916.050 ;
        RECT 226.950 913.950 229.050 916.050 ;
        RECT 229.950 913.950 232.050 916.050 ;
        RECT 224.400 912.900 225.600 913.950 ;
        RECT 214.950 910.800 217.050 912.900 ;
        RECT 223.950 910.800 226.050 912.900 ;
        RECT 223.950 904.950 226.050 907.050 ;
        RECT 208.950 901.950 211.050 904.050 ;
        RECT 202.950 898.950 205.050 901.050 ;
        RECT 209.400 892.050 210.600 901.950 ;
        RECT 211.950 895.950 214.050 898.050 ;
        RECT 208.950 889.950 211.050 892.050 ;
        RECT 208.950 884.100 211.050 886.200 ;
        RECT 178.950 880.950 181.050 883.050 ;
        RECT 181.950 880.950 184.050 883.050 ;
        RECT 184.950 880.950 187.050 883.050 ;
        RECT 193.950 880.950 196.050 883.050 ;
        RECT 196.950 880.950 199.050 883.050 ;
        RECT 199.950 880.950 202.050 883.050 ;
        RECT 202.950 880.950 205.050 883.050 ;
        RECT 182.400 879.900 183.600 880.950 ;
        RECT 197.400 879.900 198.600 880.950 ;
        RECT 181.950 877.800 184.050 879.900 ;
        RECT 196.950 877.800 199.050 879.900 ;
        RECT 203.400 874.050 204.600 880.950 ;
        RECT 205.950 874.950 208.050 877.050 ;
        RECT 187.950 871.950 190.050 874.050 ;
        RECT 202.950 871.950 205.050 874.050 ;
        RECT 172.950 850.950 175.050 853.050 ;
        RECT 169.950 841.950 172.050 844.050 ;
        RECT 154.950 835.950 157.050 838.050 ;
        RECT 160.950 835.950 163.050 838.050 ;
        RECT 163.950 835.950 166.050 838.050 ;
        RECT 161.400 834.900 162.600 835.950 ;
        RECT 170.400 835.050 171.600 841.950 ;
        RECT 173.400 841.200 174.600 850.950 ;
        RECT 188.400 850.050 189.600 871.950 ;
        RECT 190.950 865.950 193.050 868.050 ;
        RECT 187.950 847.950 190.050 850.050 ;
        RECT 172.950 839.100 175.050 841.200 ;
        RECT 178.950 839.100 181.050 841.200 ;
        RECT 184.950 840.000 187.050 844.050 ;
        RECT 188.400 841.050 189.600 847.950 ;
        RECT 160.950 832.800 163.050 834.900 ;
        RECT 169.950 832.950 172.050 835.050 ;
        RECT 148.950 814.950 151.050 817.050 ;
        RECT 112.950 811.950 115.050 814.050 ;
        RECT 124.950 811.950 127.050 814.050 ;
        RECT 136.950 811.950 139.050 814.050 ;
        RECT 85.950 808.950 88.050 811.050 ;
        RECT 91.950 808.950 94.050 811.050 ;
        RECT 76.950 802.950 79.050 805.050 ;
        RECT 79.950 802.950 82.050 805.050 ;
        RECT 82.950 802.950 85.050 805.050 ;
        RECT 85.950 802.950 88.050 805.050 ;
        RECT 71.400 800.400 75.600 801.600 ;
        RECT 64.950 787.950 67.050 790.050 ;
        RECT 67.950 769.950 70.050 772.050 ;
        RECT 68.400 760.050 69.600 769.950 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 64.950 757.950 67.050 760.050 ;
        RECT 67.950 757.950 70.050 760.050 ;
        RECT 52.950 751.950 55.050 754.050 ;
        RECT 59.400 736.050 60.600 757.950 ;
        RECT 65.400 748.050 66.600 757.950 ;
        RECT 74.400 751.050 75.600 800.400 ;
        RECT 80.400 793.050 81.600 802.950 ;
        RECT 86.400 801.900 87.600 802.950 ;
        RECT 92.400 801.900 93.600 808.950 ;
        RECT 100.950 807.000 103.050 811.050 ;
        RECT 101.400 805.050 102.600 807.000 ;
        RECT 106.950 806.100 109.050 808.200 ;
        RECT 107.400 805.050 108.600 806.100 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 100.950 802.950 103.050 805.050 ;
        RECT 103.950 802.950 106.050 805.050 ;
        RECT 106.950 802.950 109.050 805.050 ;
        RECT 98.400 801.900 99.600 802.950 ;
        RECT 85.950 799.800 88.050 801.900 ;
        RECT 91.950 799.800 94.050 801.900 ;
        RECT 97.950 799.800 100.050 801.900 ;
        RECT 104.400 796.050 105.600 802.950 ;
        RECT 113.400 801.900 114.600 811.950 ;
        RECT 115.950 805.950 118.050 808.050 ;
        RECT 112.950 799.800 115.050 801.900 ;
        RECT 103.950 793.950 106.050 796.050 ;
        RECT 79.950 790.950 82.050 793.050 ;
        RECT 82.950 784.950 85.050 787.050 ;
        RECT 76.950 778.950 79.050 781.050 ;
        RECT 77.400 763.200 78.600 778.950 ;
        RECT 83.400 772.050 84.600 784.950 ;
        RECT 104.400 781.050 105.600 793.950 ;
        RECT 103.950 778.950 106.050 781.050 ;
        RECT 116.400 775.050 117.600 805.950 ;
        RECT 125.400 805.050 126.600 811.950 ;
        RECT 130.950 806.100 133.050 808.200 ;
        RECT 131.400 805.050 132.600 806.100 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 127.950 802.950 130.050 805.050 ;
        RECT 130.950 802.950 133.050 805.050 ;
        RECT 122.400 801.000 123.600 802.950 ;
        RECT 121.950 796.950 124.050 801.000 ;
        RECT 128.400 796.050 129.600 802.950 ;
        RECT 127.950 793.950 130.050 796.050 ;
        RECT 115.950 772.950 118.050 775.050 ;
        RECT 82.950 769.950 85.050 772.050 ;
        RECT 76.950 761.100 79.050 763.200 ;
        RECT 73.950 748.950 76.050 751.050 ;
        RECT 64.950 745.950 67.050 748.050 ;
        RECT 77.400 745.050 78.600 761.100 ;
        RECT 83.400 760.050 84.600 769.950 ;
        RECT 100.950 762.000 103.050 766.050 ;
        RECT 101.400 760.050 102.600 762.000 ;
        RECT 106.950 761.100 109.050 763.200 ;
        RECT 112.950 761.100 115.050 763.200 ;
        RECT 107.400 760.050 108.600 761.100 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 85.950 757.950 88.050 760.050 ;
        RECT 97.950 757.950 100.050 760.050 ;
        RECT 100.950 757.950 103.050 760.050 ;
        RECT 103.950 757.950 106.050 760.050 ;
        RECT 106.950 757.950 109.050 760.050 ;
        RECT 86.400 745.050 87.600 757.950 ;
        RECT 94.950 748.950 97.050 751.050 ;
        RECT 61.950 742.950 64.050 745.050 ;
        RECT 76.950 742.950 79.050 745.050 ;
        RECT 85.950 742.950 88.050 745.050 ;
        RECT 58.950 733.950 61.050 736.050 ;
        RECT 55.950 728.100 58.050 730.200 ;
        RECT 56.400 727.050 57.600 728.100 ;
        RECT 62.400 727.050 63.600 742.950 ;
        RECT 73.950 733.950 76.050 736.050 ;
        RECT 70.950 728.100 73.050 730.200 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 58.950 724.950 61.050 727.050 ;
        RECT 61.950 724.950 64.050 727.050 ;
        RECT 64.950 724.950 67.050 727.050 ;
        RECT 59.400 723.900 60.600 724.950 ;
        RECT 65.400 723.900 66.600 724.950 ;
        RECT 58.950 721.800 61.050 723.900 ;
        RECT 64.950 721.800 67.050 723.900 ;
        RECT 47.400 719.400 51.600 720.600 ;
        RECT 37.950 715.950 40.050 718.050 ;
        RECT 28.950 709.950 31.050 712.050 ;
        RECT 31.950 709.950 34.050 712.050 ;
        RECT 5.400 651.600 6.600 683.100 ;
        RECT 11.400 682.050 12.600 683.100 ;
        RECT 17.400 682.050 18.600 683.100 ;
        RECT 10.950 679.950 13.050 682.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 14.400 670.050 15.600 679.950 ;
        RECT 13.950 667.950 16.050 670.050 ;
        RECT 7.950 651.600 10.050 652.200 ;
        RECT 5.400 650.400 10.050 651.600 ;
        RECT 7.950 650.100 10.050 650.400 ;
        RECT 13.950 650.100 16.050 652.200 ;
        RECT 23.400 652.050 24.600 683.100 ;
        RECT 25.950 682.950 28.050 685.050 ;
        RECT 29.400 682.050 30.600 709.950 ;
        RECT 34.950 688.950 37.050 691.050 ;
        RECT 35.400 682.050 36.600 688.950 ;
        RECT 43.950 682.950 46.050 685.050 ;
        RECT 28.950 679.950 31.050 682.050 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 37.950 679.950 40.050 682.050 ;
        RECT 32.400 678.900 33.600 679.950 ;
        RECT 31.950 676.800 34.050 678.900 ;
        RECT 25.950 670.950 28.050 673.050 ;
        RECT 22.950 651.600 25.050 652.050 ;
        RECT 20.400 650.400 25.050 651.600 ;
        RECT 2.400 647.400 6.600 648.600 ;
        RECT 1.950 589.950 4.050 592.050 ;
        RECT 2.400 544.050 3.600 589.950 ;
        RECT 1.950 541.950 4.050 544.050 ;
        RECT 2.400 403.050 3.600 541.950 ;
        RECT 5.400 517.050 6.600 647.400 ;
        RECT 8.400 601.050 9.600 650.100 ;
        RECT 14.400 649.050 15.600 650.100 ;
        RECT 20.400 649.050 21.600 650.400 ;
        RECT 22.950 649.950 25.050 650.400 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 17.400 645.900 18.600 646.950 ;
        RECT 26.400 646.050 27.600 670.950 ;
        RECT 34.950 655.950 37.050 658.050 ;
        RECT 35.400 649.050 36.600 655.950 ;
        RECT 38.400 655.050 39.600 679.950 ;
        RECT 44.400 673.050 45.600 682.950 ;
        RECT 47.400 679.050 48.600 719.400 ;
        RECT 49.950 715.950 52.050 718.050 ;
        RECT 50.400 709.050 51.600 715.950 ;
        RECT 49.950 706.950 52.050 709.050 ;
        RECT 46.950 676.950 49.050 679.050 ;
        RECT 43.950 670.950 46.050 673.050 ;
        RECT 44.400 655.050 45.600 670.950 ;
        RECT 37.950 652.950 40.050 655.050 ;
        RECT 43.950 652.950 46.050 655.050 ;
        RECT 40.950 650.100 43.050 652.200 ;
        RECT 46.800 650.100 48.900 652.200 ;
        RECT 50.400 652.050 51.600 706.950 ;
        RECT 59.400 688.200 60.600 721.800 ;
        RECT 71.400 703.050 72.600 728.100 ;
        RECT 70.950 700.950 73.050 703.050 ;
        RECT 74.400 694.050 75.600 733.950 ;
        RECT 82.950 729.000 85.050 733.050 ;
        RECT 83.400 727.050 84.600 729.000 ;
        RECT 88.950 728.100 91.050 730.200 ;
        RECT 89.400 727.050 90.600 728.100 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 80.400 712.050 81.600 724.950 ;
        RECT 82.950 718.950 85.050 721.050 ;
        RECT 79.950 709.950 82.050 712.050 ;
        RECT 73.950 691.950 76.050 694.050 ;
        RECT 58.950 686.100 61.050 688.200 ;
        RECT 70.950 685.950 73.050 688.050 ;
        RECT 58.950 682.950 61.050 685.050 ;
        RECT 64.950 683.100 67.050 685.200 ;
        RECT 59.400 682.050 60.600 682.950 ;
        RECT 65.400 682.050 66.600 683.100 ;
        RECT 55.950 679.950 58.050 682.050 ;
        RECT 58.950 679.950 61.050 682.050 ;
        RECT 61.950 679.950 64.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 56.400 678.900 57.600 679.950 ;
        RECT 55.950 676.800 58.050 678.900 ;
        RECT 62.400 670.050 63.600 679.950 ;
        RECT 61.950 667.950 64.050 670.050 ;
        RECT 55.950 655.950 58.050 658.050 ;
        RECT 41.400 649.050 42.600 650.100 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 37.950 646.950 40.050 649.050 ;
        RECT 40.950 646.950 43.050 649.050 ;
        RECT 16.950 643.800 19.050 645.900 ;
        RECT 25.950 643.950 28.050 646.050 ;
        RECT 32.400 645.900 33.600 646.950 ;
        RECT 31.950 643.800 34.050 645.900 ;
        RECT 16.950 610.950 19.050 613.050 ;
        RECT 17.400 604.050 18.600 610.950 ;
        RECT 38.400 610.050 39.600 646.950 ;
        RECT 47.400 613.050 48.600 650.100 ;
        RECT 49.950 649.950 52.050 652.050 ;
        RECT 56.400 649.050 57.600 655.950 ;
        RECT 67.950 652.950 70.050 655.050 ;
        RECT 63.000 651.600 67.050 652.050 ;
        RECT 62.400 649.950 67.050 651.600 ;
        RECT 62.400 649.050 63.600 649.950 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 55.950 646.950 58.050 649.050 ;
        RECT 58.950 646.950 61.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 53.400 645.900 54.600 646.950 ;
        RECT 52.950 643.800 55.050 645.900 ;
        RECT 59.400 645.000 60.600 646.950 ;
        RECT 58.950 640.950 61.050 645.000 ;
        RECT 64.950 643.950 67.050 646.050 ;
        RECT 65.400 636.600 66.600 643.950 ;
        RECT 68.400 640.050 69.600 652.950 ;
        RECT 71.400 651.600 72.600 685.950 ;
        RECT 83.400 685.200 84.600 718.950 ;
        RECT 86.400 709.050 87.600 724.950 ;
        RECT 85.950 706.950 88.050 709.050 ;
        RECT 91.950 700.950 94.050 703.050 ;
        RECT 76.950 683.100 79.050 685.200 ;
        RECT 82.950 683.100 85.050 685.200 ;
        RECT 77.400 682.050 78.600 683.100 ;
        RECT 83.400 682.050 84.600 683.100 ;
        RECT 92.400 682.050 93.600 700.950 ;
        RECT 76.950 679.950 79.050 682.050 ;
        RECT 79.950 679.950 82.050 682.050 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 85.950 679.950 88.050 682.050 ;
        RECT 91.950 679.950 94.050 682.050 ;
        RECT 80.400 678.900 81.600 679.950 ;
        RECT 79.950 676.800 82.050 678.900 ;
        RECT 80.400 670.050 81.600 676.800 ;
        RECT 86.400 670.050 87.600 679.950 ;
        RECT 95.400 676.050 96.600 748.950 ;
        RECT 98.400 724.050 99.600 757.950 ;
        RECT 104.400 756.000 105.600 757.950 ;
        RECT 103.950 751.950 106.050 756.000 ;
        RECT 113.400 745.050 114.600 761.100 ;
        RECT 116.400 754.050 117.600 772.950 ;
        RECT 137.400 765.600 138.600 811.950 ;
        RECT 161.400 811.050 162.600 832.800 ;
        RECT 173.400 832.050 174.600 839.100 ;
        RECT 179.400 838.050 180.600 839.100 ;
        RECT 185.400 838.050 186.600 840.000 ;
        RECT 187.950 838.950 190.050 841.050 ;
        RECT 178.950 835.950 181.050 838.050 ;
        RECT 181.950 835.950 184.050 838.050 ;
        RECT 184.950 835.950 187.050 838.050 ;
        RECT 182.400 834.900 183.600 835.950 ;
        RECT 181.950 832.800 184.050 834.900 ;
        RECT 163.950 829.950 166.050 832.050 ;
        RECT 172.950 829.950 175.050 832.050 ;
        RECT 160.950 808.950 163.050 811.050 ;
        RECT 139.950 806.100 142.050 808.200 ;
        RECT 145.950 806.100 148.050 808.200 ;
        RECT 151.950 806.100 154.050 808.200 ;
        RECT 140.400 787.050 141.600 806.100 ;
        RECT 146.400 805.050 147.600 806.100 ;
        RECT 152.400 805.050 153.600 806.100 ;
        RECT 160.950 805.800 163.050 807.900 ;
        RECT 145.950 802.950 148.050 805.050 ;
        RECT 148.950 802.950 151.050 805.050 ;
        RECT 151.950 802.950 154.050 805.050 ;
        RECT 154.950 802.950 157.050 805.050 ;
        RECT 149.400 801.900 150.600 802.950 ;
        RECT 148.950 799.800 151.050 801.900 ;
        RECT 155.400 796.050 156.600 802.950 ;
        RECT 161.400 796.050 162.600 805.800 ;
        RECT 145.950 793.950 148.050 796.050 ;
        RECT 154.950 793.950 157.050 796.050 ;
        RECT 160.950 793.950 163.050 796.050 ;
        RECT 139.950 784.950 142.050 787.050 ;
        RECT 146.400 775.050 147.600 793.950 ;
        RECT 164.400 781.050 165.600 829.950 ;
        RECT 166.950 814.950 169.050 817.050 ;
        RECT 167.400 799.050 168.600 814.950 ;
        RECT 175.950 811.950 178.050 814.050 ;
        RECT 176.400 805.050 177.600 811.950 ;
        RECT 191.400 808.200 192.600 865.950 ;
        RECT 196.950 839.100 199.050 841.200 ;
        RECT 206.400 840.600 207.600 874.950 ;
        RECT 203.400 839.400 207.600 840.600 ;
        RECT 197.400 838.050 198.600 839.100 ;
        RECT 203.400 838.050 204.600 839.400 ;
        RECT 196.950 835.950 199.050 838.050 ;
        RECT 199.950 835.950 202.050 838.050 ;
        RECT 202.950 835.950 205.050 838.050 ;
        RECT 200.400 829.050 201.600 835.950 ;
        RECT 209.400 829.050 210.600 884.100 ;
        RECT 212.400 880.050 213.600 895.950 ;
        RECT 224.400 883.050 225.600 904.950 ;
        RECT 220.950 880.950 223.050 883.050 ;
        RECT 223.950 880.950 226.050 883.050 ;
        RECT 211.950 877.950 214.050 880.050 ;
        RECT 221.400 879.900 222.600 880.950 ;
        RECT 220.950 877.800 223.050 879.900 ;
        RECT 230.400 868.050 231.600 913.950 ;
        RECT 236.400 901.050 237.600 917.100 ;
        RECT 248.400 916.050 249.600 922.950 ;
        RECT 259.950 918.600 262.050 919.200 ;
        RECT 254.400 917.400 262.050 918.600 ;
        RECT 254.400 916.050 255.600 917.400 ;
        RECT 259.950 917.100 262.050 917.400 ;
        RECT 244.950 913.950 247.050 916.050 ;
        RECT 247.950 913.950 250.050 916.050 ;
        RECT 250.950 913.950 253.050 916.050 ;
        RECT 253.950 913.950 256.050 916.050 ;
        RECT 235.950 898.950 238.050 901.050 ;
        RECT 245.400 892.050 246.600 913.950 ;
        RECT 251.400 912.900 252.600 913.950 ;
        RECT 250.950 910.800 253.050 912.900 ;
        RECT 256.950 910.800 259.050 912.900 ;
        RECT 244.950 889.950 247.050 892.050 ;
        RECT 232.950 884.100 235.050 886.200 ;
        RECT 241.950 884.100 244.050 886.200 ;
        RECT 250.950 884.100 253.050 886.200 ;
        RECT 233.400 874.050 234.600 884.100 ;
        RECT 242.400 883.050 243.600 884.100 ;
        RECT 251.400 883.050 252.600 884.100 ;
        RECT 257.400 883.050 258.600 910.800 ;
        RECT 260.400 904.050 261.600 917.100 ;
        RECT 266.400 916.050 267.600 922.950 ;
        RECT 271.950 917.100 274.050 919.200 ;
        RECT 272.400 916.050 273.600 917.100 ;
        RECT 265.950 913.950 268.050 916.050 ;
        RECT 268.950 913.950 271.050 916.050 ;
        RECT 271.950 913.950 274.050 916.050 ;
        RECT 274.950 913.950 277.050 916.050 ;
        RECT 269.400 912.900 270.600 913.950 ;
        RECT 268.950 910.800 271.050 912.900 ;
        RECT 275.400 907.050 276.600 913.950 ;
        RECT 274.950 904.950 277.050 907.050 ;
        RECT 259.950 901.950 262.050 904.050 ;
        RECT 281.400 895.050 282.600 922.950 ;
        RECT 286.950 917.100 289.050 919.200 ;
        RECT 292.950 917.100 295.050 919.200 ;
        RECT 287.400 912.900 288.600 917.100 ;
        RECT 293.400 916.050 294.600 917.100 ;
        RECT 299.400 916.050 300.600 928.950 ;
        RECT 304.950 925.950 307.050 928.050 ;
        RECT 292.950 913.950 295.050 916.050 ;
        RECT 295.950 913.950 298.050 916.050 ;
        RECT 298.950 913.950 301.050 916.050 ;
        RECT 286.950 910.800 289.050 912.900 ;
        RECT 296.400 912.000 297.600 913.950 ;
        RECT 265.950 892.950 268.050 895.050 ;
        RECT 280.950 892.950 283.050 895.050 ;
        RECT 238.950 880.950 241.050 883.050 ;
        RECT 241.950 880.950 244.050 883.050 ;
        RECT 250.950 880.950 253.050 883.050 ;
        RECT 253.950 880.950 256.050 883.050 ;
        RECT 256.950 880.950 259.050 883.050 ;
        RECT 259.950 880.950 262.050 883.050 ;
        RECT 239.400 879.900 240.600 880.950 ;
        RECT 254.400 879.900 255.600 880.950 ;
        RECT 238.950 877.800 241.050 879.900 ;
        RECT 253.950 877.800 256.050 879.900 ;
        RECT 260.400 879.600 261.600 880.950 ;
        RECT 260.400 878.400 264.600 879.600 ;
        RECT 232.950 871.950 235.050 874.050 ;
        RECT 229.950 865.950 232.050 868.050 ;
        RECT 233.400 858.600 234.600 871.950 ;
        RECT 259.950 859.950 262.050 862.050 ;
        RECT 230.400 857.400 234.600 858.600 ;
        RECT 220.950 839.100 223.050 841.200 ;
        RECT 221.400 838.050 222.600 839.100 ;
        RECT 217.950 835.950 220.050 838.050 ;
        RECT 220.950 835.950 223.050 838.050 ;
        RECT 223.950 835.950 226.050 838.050 ;
        RECT 199.950 826.950 202.050 829.050 ;
        RECT 208.950 826.950 211.050 829.050 ;
        RECT 218.400 826.050 219.600 835.950 ;
        RECT 224.400 829.050 225.600 835.950 ;
        RECT 230.400 835.050 231.600 857.400 ;
        RECT 235.950 839.100 238.050 841.200 ;
        RECT 241.950 840.000 244.050 844.050 ;
        RECT 236.400 838.050 237.600 839.100 ;
        RECT 242.400 838.050 243.600 840.000 ;
        RECT 247.950 838.950 250.050 841.050 ;
        RECT 235.950 835.950 238.050 838.050 ;
        RECT 238.950 835.950 241.050 838.050 ;
        RECT 241.950 835.950 244.050 838.050 ;
        RECT 229.950 832.950 232.050 835.050 ;
        RECT 239.400 834.900 240.600 835.950 ;
        RECT 248.400 834.900 249.600 838.950 ;
        RECT 260.400 838.050 261.600 859.950 ;
        RECT 263.400 859.050 264.600 878.400 ;
        RECT 262.950 856.950 265.050 859.050 ;
        RECT 266.400 853.050 267.600 892.950 ;
        RECT 283.950 889.950 286.050 892.050 ;
        RECT 271.950 884.100 274.050 886.200 ;
        RECT 280.950 884.100 283.050 886.200 ;
        RECT 272.400 883.050 273.600 884.100 ;
        RECT 271.950 880.950 274.050 883.050 ;
        RECT 274.950 880.950 277.050 883.050 ;
        RECT 268.950 877.950 271.050 880.050 ;
        RECT 275.400 879.900 276.600 880.950 ;
        RECT 269.400 862.050 270.600 877.950 ;
        RECT 274.950 877.800 277.050 879.900 ;
        RECT 281.400 874.050 282.600 884.100 ;
        RECT 280.950 871.950 283.050 874.050 ;
        RECT 268.950 859.950 271.050 862.050 ;
        RECT 284.400 858.600 285.600 889.950 ;
        RECT 287.400 868.050 288.600 910.800 ;
        RECT 295.950 907.950 298.050 912.000 ;
        RECT 305.400 910.050 306.600 925.950 ;
        RECT 311.400 916.050 312.600 928.950 ;
        RECT 316.950 917.100 319.050 919.200 ;
        RECT 325.950 917.100 328.050 919.200 ;
        RECT 317.400 916.050 318.600 917.100 ;
        RECT 310.950 913.950 313.050 916.050 ;
        RECT 313.950 913.950 316.050 916.050 ;
        RECT 316.950 913.950 319.050 916.050 ;
        RECT 319.950 913.950 322.050 916.050 ;
        RECT 314.400 912.900 315.600 913.950 ;
        RECT 313.950 910.800 316.050 912.900 ;
        RECT 304.950 907.950 307.050 910.050 ;
        RECT 292.950 901.950 295.050 904.050 ;
        RECT 293.400 883.050 294.600 901.950 ;
        RECT 307.950 898.950 310.050 901.050 ;
        RECT 298.950 884.100 301.050 886.200 ;
        RECT 299.400 883.050 300.600 884.100 ;
        RECT 292.950 880.950 295.050 883.050 ;
        RECT 295.950 880.950 298.050 883.050 ;
        RECT 298.950 880.950 301.050 883.050 ;
        RECT 301.950 880.950 304.050 883.050 ;
        RECT 296.400 879.900 297.600 880.950 ;
        RECT 302.400 879.900 303.600 880.950 ;
        RECT 295.950 877.800 298.050 879.900 ;
        RECT 301.950 877.800 304.050 879.900 ;
        RECT 308.400 877.050 309.600 898.950 ;
        RECT 320.400 895.050 321.600 913.950 ;
        RECT 326.400 913.050 327.600 917.100 ;
        RECT 335.400 916.050 336.600 928.950 ;
        RECT 337.950 925.950 340.050 928.050 ;
        RECT 355.950 925.950 358.050 928.050 ;
        RECT 370.950 925.950 373.050 928.050 ;
        RECT 463.950 925.950 466.050 928.050 ;
        RECT 505.950 925.950 508.050 928.050 ;
        RECT 338.400 922.050 339.600 925.950 ;
        RECT 340.950 922.050 343.050 922.200 ;
        RECT 338.400 920.550 343.050 922.050 ;
        RECT 339.000 920.100 343.050 920.550 ;
        RECT 339.000 919.950 342.000 920.100 ;
        RECT 340.950 916.950 343.050 919.050 ;
        RECT 349.950 918.000 352.050 922.050 ;
        RECT 341.400 916.050 342.600 916.950 ;
        RECT 350.400 916.050 351.600 918.000 ;
        RECT 356.400 916.050 357.600 925.950 ;
        RECT 367.950 917.100 370.050 919.200 ;
        RECT 334.950 913.950 337.050 916.050 ;
        RECT 337.950 913.950 340.050 916.050 ;
        RECT 340.950 913.950 343.050 916.050 ;
        RECT 349.950 913.950 352.050 916.050 ;
        RECT 352.950 913.950 355.050 916.050 ;
        RECT 355.950 913.950 358.050 916.050 ;
        RECT 358.950 913.950 361.050 916.050 ;
        RECT 325.950 910.950 328.050 913.050 ;
        RECT 338.400 912.900 339.600 913.950 ;
        RECT 353.400 912.900 354.600 913.950 ;
        RECT 337.950 910.800 340.050 912.900 ;
        RECT 352.950 910.800 355.050 912.900 ;
        RECT 319.950 892.950 322.050 895.050 ;
        RECT 316.950 888.600 319.050 892.050 ;
        RECT 319.950 888.600 322.050 889.050 ;
        RECT 316.950 888.000 322.050 888.600 ;
        RECT 317.400 887.400 322.050 888.000 ;
        RECT 319.950 886.950 322.050 887.400 ;
        RECT 320.400 883.050 321.600 886.950 ;
        RECT 328.950 885.600 331.050 889.050 ;
        RECT 328.950 885.000 333.600 885.600 ;
        RECT 329.400 884.400 333.600 885.000 ;
        RECT 332.400 883.050 333.600 884.400 ;
        RECT 337.950 884.100 340.050 886.200 ;
        RECT 352.950 884.100 355.050 886.200 ;
        RECT 359.400 885.600 360.600 913.950 ;
        RECT 364.950 892.950 367.050 895.050 ;
        RECT 359.400 884.400 363.600 885.600 ;
        RECT 338.400 883.050 339.600 884.100 ;
        RECT 353.400 883.050 354.600 884.100 ;
        RECT 316.950 880.950 319.050 883.050 ;
        RECT 319.950 880.950 322.050 883.050 ;
        RECT 331.950 880.950 334.050 883.050 ;
        RECT 334.950 880.950 337.050 883.050 ;
        RECT 337.950 880.950 340.050 883.050 ;
        RECT 340.950 880.950 343.050 883.050 ;
        RECT 352.950 880.950 355.050 883.050 ;
        RECT 355.950 880.950 358.050 883.050 ;
        RECT 317.400 879.900 318.600 880.950 ;
        RECT 316.950 877.800 319.050 879.900 ;
        RECT 307.950 874.950 310.050 877.050 ;
        RECT 286.950 865.950 289.050 868.050 ;
        RECT 335.400 862.050 336.600 880.950 ;
        RECT 341.400 874.050 342.600 880.950 ;
        RECT 356.400 879.900 357.600 880.950 ;
        RECT 355.950 877.800 358.050 879.900 ;
        RECT 340.950 871.950 343.050 874.050 ;
        RECT 334.950 859.950 337.050 862.050 ;
        RECT 362.400 859.050 363.600 884.400 ;
        RECT 286.950 858.600 289.050 859.050 ;
        RECT 284.400 857.400 289.050 858.600 ;
        RECT 286.950 856.950 289.050 857.400 ;
        RECT 361.950 856.950 364.050 859.050 ;
        RECT 265.950 850.950 268.050 853.050 ;
        RECT 268.950 841.950 271.050 844.050 ;
        RECT 256.950 835.950 259.050 838.050 ;
        RECT 259.950 835.950 262.050 838.050 ;
        RECT 262.950 835.950 265.050 838.050 ;
        RECT 257.400 834.900 258.600 835.950 ;
        RECT 238.950 832.800 241.050 834.900 ;
        RECT 247.950 832.800 250.050 834.900 ;
        RECT 256.950 832.800 259.050 834.900 ;
        RECT 223.950 826.950 226.050 829.050 ;
        RECT 217.950 823.950 220.050 826.050 ;
        RECT 244.950 823.950 247.050 829.050 ;
        RECT 253.950 826.950 256.050 829.050 ;
        RECT 218.400 820.050 219.600 823.950 ;
        RECT 254.400 823.050 255.600 826.950 ;
        RECT 256.950 823.950 259.050 829.050 ;
        RECT 253.950 820.950 256.050 823.050 ;
        RECT 202.950 817.950 205.050 820.050 ;
        RECT 217.800 817.950 219.900 820.050 ;
        RECT 190.950 806.100 193.050 808.200 ;
        RECT 196.950 806.100 199.050 808.200 ;
        RECT 191.400 805.050 192.600 806.100 ;
        RECT 197.400 805.050 198.600 806.100 ;
        RECT 172.950 802.950 175.050 805.050 ;
        RECT 175.950 802.950 178.050 805.050 ;
        RECT 178.950 802.950 181.050 805.050 ;
        RECT 187.950 802.950 190.050 805.050 ;
        RECT 190.950 802.950 193.050 805.050 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 169.950 799.950 172.050 802.050 ;
        RECT 173.400 801.000 174.600 802.950 ;
        RECT 179.400 801.900 180.600 802.950 ;
        RECT 166.950 796.950 169.050 799.050 ;
        RECT 170.400 787.050 171.600 799.950 ;
        RECT 172.950 796.950 175.050 801.000 ;
        RECT 178.950 799.800 181.050 801.900 ;
        RECT 173.400 793.050 174.600 796.950 ;
        RECT 188.400 793.050 189.600 802.950 ;
        RECT 194.400 796.050 195.600 802.950 ;
        RECT 193.950 793.950 196.050 796.050 ;
        RECT 172.950 790.950 175.050 793.050 ;
        RECT 187.950 790.950 190.050 793.050 ;
        RECT 169.950 784.950 172.050 787.050 ;
        RECT 184.950 784.950 187.050 787.050 ;
        RECT 163.950 778.950 166.050 781.050 ;
        RECT 175.950 778.950 178.050 781.050 ;
        RECT 145.950 772.950 148.050 775.050 ;
        RECT 163.950 772.950 166.050 775.050 ;
        RECT 137.400 764.400 141.600 765.600 ;
        RECT 121.950 761.100 124.050 763.200 ;
        RECT 122.400 760.050 123.600 761.100 ;
        RECT 130.950 760.950 133.050 763.050 ;
        RECT 121.950 757.950 124.050 760.050 ;
        RECT 124.950 757.950 127.050 760.050 ;
        RECT 125.400 756.900 126.600 757.950 ;
        RECT 124.950 754.800 127.050 756.900 ;
        RECT 131.400 754.050 132.600 760.950 ;
        RECT 140.400 760.050 141.600 764.400 ;
        RECT 146.400 760.050 147.600 772.950 ;
        RECT 164.400 763.200 165.600 772.950 ;
        RECT 172.950 766.950 175.050 769.050 ;
        RECT 152.400 761.400 159.600 762.600 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 139.950 757.950 142.050 760.050 ;
        RECT 142.950 757.950 145.050 760.050 ;
        RECT 145.950 757.950 148.050 760.050 ;
        RECT 115.950 751.950 118.050 754.050 ;
        RECT 130.950 751.950 133.050 754.050 ;
        RECT 112.950 742.950 115.050 745.050 ;
        RECT 118.800 742.950 120.900 745.050 ;
        RECT 121.950 742.950 124.050 745.050 ;
        RECT 103.950 729.000 106.050 733.050 ;
        RECT 104.400 727.050 105.600 729.000 ;
        RECT 109.950 728.100 112.050 730.200 ;
        RECT 110.400 727.050 111.600 728.100 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 97.950 721.950 100.050 724.050 ;
        RECT 107.400 718.050 108.600 724.950 ;
        RECT 106.950 715.950 109.050 718.050 ;
        RECT 109.950 709.950 112.050 712.050 ;
        RECT 110.400 688.050 111.600 709.950 ;
        RECT 113.400 709.050 114.600 724.950 ;
        RECT 112.950 706.950 115.050 709.050 ;
        RECT 115.950 703.950 118.050 706.050 ;
        RECT 116.400 700.050 117.600 703.950 ;
        RECT 115.950 697.950 118.050 700.050 ;
        RECT 109.950 685.950 112.050 688.050 ;
        RECT 100.950 683.100 103.050 685.200 ;
        RECT 106.950 683.100 109.050 685.200 ;
        RECT 101.400 682.050 102.600 683.100 ;
        RECT 107.400 682.050 108.600 683.100 ;
        RECT 115.950 682.950 118.050 685.050 ;
        RECT 100.950 679.950 103.050 682.050 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 97.950 676.950 100.050 679.050 ;
        RECT 104.400 678.900 105.600 679.950 ;
        RECT 88.950 673.950 91.050 676.050 ;
        RECT 94.950 673.950 97.050 676.050 ;
        RECT 79.950 667.950 82.050 670.050 ;
        RECT 85.950 667.950 88.050 670.050 ;
        RECT 71.400 650.400 75.600 651.600 ;
        RECT 74.400 649.050 75.600 650.400 ;
        RECT 79.950 650.100 82.050 652.200 ;
        RECT 80.400 649.050 81.600 650.100 ;
        RECT 73.950 646.950 76.050 649.050 ;
        RECT 76.950 646.950 79.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 70.950 643.950 73.050 646.050 ;
        RECT 67.950 637.950 70.050 640.050 ;
        RECT 65.400 635.400 69.600 636.600 ;
        RECT 46.950 610.950 49.050 613.050 ;
        RECT 58.950 610.950 61.050 613.050 ;
        RECT 22.950 605.100 25.050 607.200 ;
        RECT 28.950 605.100 31.050 610.050 ;
        RECT 37.950 607.950 40.050 610.050 ;
        RECT 34.950 605.100 37.050 607.200 ;
        RECT 40.950 606.000 43.050 610.050 ;
        RECT 23.400 604.050 24.600 605.100 ;
        RECT 13.950 601.950 16.050 604.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 19.950 601.950 22.050 604.050 ;
        RECT 22.950 601.950 25.050 604.050 ;
        RECT 7.950 598.950 10.050 601.050 ;
        RECT 14.400 600.900 15.600 601.950 ;
        RECT 13.950 598.800 16.050 600.900 ;
        RECT 20.400 600.000 21.600 601.950 ;
        RECT 19.950 595.950 22.050 600.000 ;
        RECT 16.950 586.950 19.050 589.050 ;
        RECT 7.950 574.950 10.050 577.050 ;
        RECT 8.400 567.900 9.600 574.950 ;
        RECT 17.400 571.050 18.600 586.950 ;
        RECT 22.950 583.950 25.050 586.050 ;
        RECT 23.400 571.050 24.600 583.950 ;
        RECT 29.400 574.050 30.600 605.100 ;
        RECT 35.400 604.050 36.600 605.100 ;
        RECT 41.400 604.050 42.600 606.000 ;
        RECT 49.950 604.950 52.050 607.050 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 43.950 601.950 46.050 604.050 ;
        RECT 31.950 598.950 34.050 601.050 ;
        RECT 28.950 571.950 31.050 574.050 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 19.950 568.950 22.050 571.050 ;
        RECT 22.950 568.950 25.050 571.050 ;
        RECT 25.950 568.950 28.050 571.050 ;
        RECT 14.400 567.900 15.600 568.950 ;
        RECT 7.950 565.800 10.050 567.900 ;
        RECT 13.950 565.800 16.050 567.900 ;
        RECT 20.400 532.050 21.600 568.950 ;
        RECT 26.400 562.050 27.600 568.950 ;
        RECT 25.950 559.950 28.050 562.050 ;
        RECT 28.950 538.950 31.050 541.050 ;
        RECT 7.950 529.950 10.050 532.050 ;
        RECT 19.950 529.950 22.050 532.050 ;
        RECT 8.400 522.750 9.600 529.950 ;
        RECT 19.950 526.800 22.050 528.900 ;
        RECT 20.400 525.900 21.600 526.800 ;
        RECT 29.400 525.900 30.600 538.950 ;
        RECT 32.400 528.600 33.600 598.950 ;
        RECT 38.400 598.050 39.600 601.950 ;
        RECT 37.950 595.950 40.050 598.050 ;
        RECT 38.400 577.050 39.600 595.950 ;
        RECT 40.950 583.950 43.050 586.050 ;
        RECT 37.950 574.950 40.050 577.050 ;
        RECT 41.400 571.050 42.600 583.950 ;
        RECT 44.400 574.050 45.600 601.950 ;
        RECT 50.400 589.050 51.600 604.950 ;
        RECT 59.400 604.050 60.600 610.950 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 58.950 601.950 61.050 604.050 ;
        RECT 61.950 601.950 64.050 604.050 ;
        RECT 49.950 586.950 52.050 589.050 ;
        RECT 56.400 583.050 57.600 601.950 ;
        RECT 62.400 592.050 63.600 601.950 ;
        RECT 68.400 601.050 69.600 635.400 ;
        RECT 67.950 598.950 70.050 601.050 ;
        RECT 71.400 595.050 72.600 643.950 ;
        RECT 73.950 640.950 76.050 643.050 ;
        RECT 74.400 613.050 75.600 640.950 ;
        RECT 77.400 640.050 78.600 646.950 ;
        RECT 83.400 645.000 84.600 646.950 ;
        RECT 82.950 640.950 85.050 645.000 ;
        RECT 76.950 637.950 79.050 640.050 ;
        RECT 89.400 637.050 90.600 673.950 ;
        RECT 98.400 661.050 99.600 676.950 ;
        RECT 103.950 676.800 106.050 678.900 ;
        RECT 91.950 658.950 94.050 661.050 ;
        RECT 97.950 658.950 100.050 661.050 ;
        RECT 92.400 643.050 93.600 658.950 ;
        RECT 110.400 655.050 111.600 679.950 ;
        RECT 116.400 675.600 117.600 682.950 ;
        RECT 119.400 679.050 120.600 742.950 ;
        RECT 122.400 724.050 123.600 742.950 ;
        RECT 131.400 732.600 132.600 751.950 ;
        RECT 137.400 748.050 138.600 757.950 ;
        RECT 136.950 745.950 139.050 748.050 ;
        RECT 143.400 745.050 144.600 757.950 ;
        RECT 148.950 751.950 151.050 754.050 ;
        RECT 142.950 742.950 145.050 745.050 ;
        RECT 131.400 731.400 135.600 732.600 ;
        RECT 127.950 728.100 130.050 730.200 ;
        RECT 128.400 727.050 129.600 728.100 ;
        RECT 134.400 727.050 135.600 731.400 ;
        RECT 149.400 727.050 150.600 751.950 ;
        RECT 152.400 742.050 153.600 761.400 ;
        RECT 158.400 760.050 159.600 761.400 ;
        RECT 163.950 761.100 166.050 763.200 ;
        RECT 164.400 760.050 165.600 761.100 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 163.950 757.950 166.050 760.050 ;
        RECT 166.950 757.950 169.050 760.050 ;
        RECT 161.400 748.050 162.600 757.950 ;
        RECT 160.950 745.950 163.050 748.050 ;
        RECT 151.950 739.950 154.050 742.050 ;
        RECT 152.400 733.050 153.600 739.950 ;
        RECT 151.950 730.950 154.050 733.050 ;
        RECT 155.400 728.400 162.600 729.600 ;
        RECT 155.400 727.050 156.600 728.400 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 130.950 724.950 133.050 727.050 ;
        RECT 133.950 724.950 136.050 727.050 ;
        RECT 136.950 724.950 139.050 727.050 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 148.950 724.950 151.050 727.050 ;
        RECT 151.950 724.950 154.050 727.050 ;
        RECT 154.950 724.950 157.050 727.050 ;
        RECT 121.950 721.950 124.050 724.050 ;
        RECT 131.400 723.900 132.600 724.950 ;
        RECT 122.400 685.050 123.600 721.950 ;
        RECT 130.950 721.800 133.050 723.900 ;
        RECT 137.400 723.000 138.600 724.950 ;
        RECT 146.400 723.900 147.600 724.950 ;
        RECT 152.400 723.900 153.600 724.950 ;
        RECT 136.950 718.950 139.050 723.000 ;
        RECT 145.950 721.800 148.050 723.900 ;
        RECT 151.950 718.950 154.050 723.900 ;
        RECT 130.950 715.950 133.050 718.050 ;
        RECT 131.400 697.050 132.600 715.950 ;
        RECT 157.950 706.950 160.050 709.050 ;
        RECT 130.950 694.950 133.050 697.050 ;
        RECT 145.950 691.950 148.050 694.050 ;
        RECT 127.800 687.300 129.900 689.400 ;
        RECT 137.400 688.500 139.500 690.600 ;
        RECT 121.950 682.950 124.050 685.050 ;
        RECT 125.400 682.050 126.600 684.600 ;
        RECT 125.400 679.950 127.500 682.050 ;
        RECT 118.950 676.950 121.050 679.050 ;
        RECT 121.950 676.950 124.050 679.050 ;
        RECT 128.700 678.300 129.600 687.300 ;
        RECT 131.100 683.700 133.200 685.800 ;
        RECT 134.400 684.900 135.600 687.450 ;
        RECT 132.300 681.300 133.200 683.700 ;
        RECT 134.100 682.800 136.200 684.900 ;
        RECT 138.000 681.300 139.050 688.500 ;
        RECT 132.300 680.100 139.050 681.300 ;
        RECT 135.150 678.300 137.250 679.200 ;
        RECT 128.700 677.100 137.250 678.300 ;
        RECT 113.400 674.400 117.600 675.600 ;
        RECT 109.950 652.950 112.050 655.050 ;
        RECT 100.950 650.100 103.050 652.200 ;
        RECT 101.400 649.050 102.600 650.100 ;
        RECT 97.950 646.950 100.050 649.050 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 106.950 646.950 109.050 649.050 ;
        RECT 91.950 640.950 94.050 643.050 ;
        RECT 88.950 634.950 91.050 637.050 ;
        RECT 98.400 631.050 99.600 646.950 ;
        RECT 103.950 643.950 106.050 646.050 ;
        RECT 97.950 628.950 100.050 631.050 ;
        RECT 104.400 622.050 105.600 643.950 ;
        RECT 107.400 637.050 108.600 646.950 ;
        RECT 113.400 637.050 114.600 674.400 ;
        RECT 122.400 673.050 123.600 676.950 ;
        RECT 130.200 675.300 132.300 677.100 ;
        RECT 134.100 676.050 136.200 676.200 ;
        RECT 133.950 674.100 136.200 676.050 ;
        RECT 138.150 674.700 139.050 680.100 ;
        RECT 139.950 679.950 142.050 682.050 ;
        RECT 140.400 677.400 141.600 679.950 ;
        RECT 133.950 673.950 136.050 674.100 ;
        RECT 121.950 670.950 124.050 673.050 ;
        RECT 127.950 670.950 130.050 673.050 ;
        RECT 134.400 671.550 135.600 673.950 ;
        RECT 137.400 672.600 139.500 674.700 ;
        RECT 115.950 667.950 118.050 670.050 ;
        RECT 116.400 643.050 117.600 667.950 ;
        RECT 128.400 658.050 129.600 670.950 ;
        RECT 146.400 664.050 147.600 691.950 ;
        RECT 154.950 688.950 157.050 691.050 ;
        RECT 155.400 685.050 156.600 688.950 ;
        RECT 158.400 687.600 159.600 706.950 ;
        RECT 161.400 691.050 162.600 728.400 ;
        RECT 163.950 728.100 166.050 730.200 ;
        RECT 167.400 730.050 168.600 757.950 ;
        RECT 173.400 757.050 174.600 766.950 ;
        RECT 172.950 754.950 175.050 757.050 ;
        RECT 176.400 748.050 177.600 778.950 ;
        RECT 185.400 760.050 186.600 784.950 ;
        RECT 203.400 769.050 204.600 817.950 ;
        RECT 220.950 816.600 223.050 820.050 ;
        RECT 218.400 816.000 223.050 816.600 ;
        RECT 218.400 815.400 222.600 816.000 ;
        RECT 214.650 809.400 216.750 811.500 ;
        RECT 208.950 805.950 211.050 808.050 ;
        RECT 209.400 778.050 210.600 805.950 ;
        RECT 212.400 803.100 214.500 805.200 ;
        RECT 212.400 800.550 213.600 803.100 ;
        RECT 215.400 796.800 216.300 809.400 ;
        RECT 218.400 807.900 219.600 815.400 ;
        RECT 221.400 810.900 222.600 813.450 ;
        RECT 221.400 808.800 223.500 810.900 ;
        RECT 224.700 809.100 226.800 811.200 ;
        RECT 217.200 807.000 219.600 807.900 ;
        RECT 217.200 805.800 224.250 807.000 ;
        RECT 222.150 804.900 224.250 805.800 ;
        RECT 217.200 804.000 219.300 804.900 ;
        RECT 225.150 804.000 226.050 809.100 ;
        RECT 227.400 805.200 228.600 807.600 ;
        RECT 232.950 805.950 235.050 808.050 ;
        RECT 244.950 806.100 247.050 808.200 ;
        RECT 217.200 803.100 226.050 804.000 ;
        RECT 226.950 803.100 229.050 805.200 ;
        RECT 217.200 802.800 219.300 803.100 ;
        RECT 221.400 800.100 223.500 802.200 ;
        RECT 215.100 794.700 217.200 796.800 ;
        RECT 221.400 790.050 222.600 800.100 ;
        RECT 225.150 796.500 226.050 803.100 ;
        RECT 233.400 802.050 234.600 805.950 ;
        RECT 245.400 805.050 246.600 806.100 ;
        RECT 241.950 802.950 244.050 805.050 ;
        RECT 244.950 802.950 247.050 805.050 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 232.950 799.950 235.050 802.050 ;
        RECT 224.100 794.400 226.200 796.500 ;
        RECT 220.950 787.950 223.050 790.050 ;
        RECT 235.950 787.950 238.050 790.050 ;
        RECT 223.950 784.950 226.050 787.050 ;
        RECT 208.950 775.950 211.050 778.050 ;
        RECT 205.950 772.950 208.050 775.050 ;
        RECT 217.950 772.950 220.050 775.050 ;
        RECT 202.950 766.950 205.050 769.050 ;
        RECT 193.950 763.950 196.050 766.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 182.400 757.050 183.600 757.950 ;
        RECT 178.950 755.400 183.600 757.050 ;
        RECT 188.400 756.000 189.600 757.950 ;
        RECT 178.950 754.950 183.000 755.400 ;
        RECT 181.950 751.950 184.050 754.050 ;
        RECT 187.950 751.950 190.050 756.000 ;
        RECT 194.400 754.050 195.600 763.950 ;
        RECT 199.950 762.000 202.050 766.050 ;
        RECT 200.400 760.050 201.600 762.000 ;
        RECT 206.400 760.050 207.600 772.950 ;
        RECT 218.400 763.200 219.600 772.950 ;
        RECT 220.950 763.950 223.050 766.050 ;
        RECT 211.950 761.100 214.050 763.200 ;
        RECT 217.950 761.100 220.050 763.200 ;
        RECT 212.400 760.050 213.600 761.100 ;
        RECT 199.950 757.950 202.050 760.050 ;
        RECT 202.950 757.950 205.050 760.050 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 203.400 756.900 204.600 757.950 ;
        RECT 202.950 754.800 205.050 756.900 ;
        RECT 209.400 756.000 210.600 757.950 ;
        RECT 193.950 751.950 196.050 754.050 ;
        RECT 199.950 751.950 202.050 754.050 ;
        RECT 175.950 745.950 178.050 748.050 ;
        RECT 164.400 715.050 165.600 728.100 ;
        RECT 166.950 727.950 169.050 730.050 ;
        RECT 169.950 728.100 172.050 730.200 ;
        RECT 170.400 727.050 171.600 728.100 ;
        RECT 178.950 727.950 181.050 730.050 ;
        RECT 169.950 724.950 172.050 727.050 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 173.400 723.900 174.600 724.950 ;
        RECT 172.950 721.800 175.050 723.900 ;
        RECT 163.950 712.950 166.050 715.050 ;
        RECT 179.400 706.050 180.600 727.950 ;
        RECT 178.950 703.950 181.050 706.050 ;
        RECT 182.400 700.050 183.600 751.950 ;
        RECT 190.950 739.950 193.050 742.050 ;
        RECT 191.400 727.050 192.600 739.950 ;
        RECT 196.950 736.950 199.050 739.050 ;
        RECT 197.400 730.050 198.600 736.950 ;
        RECT 196.950 727.950 199.050 730.050 ;
        RECT 187.950 724.950 190.050 727.050 ;
        RECT 190.950 724.950 193.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 188.400 718.050 189.600 724.950 ;
        RECT 187.950 715.950 190.050 718.050 ;
        RECT 194.400 706.050 195.600 724.950 ;
        RECT 200.400 721.050 201.600 751.950 ;
        RECT 203.400 730.200 204.600 754.800 ;
        RECT 208.950 751.950 211.050 756.000 ;
        RECT 218.400 742.050 219.600 761.100 ;
        RECT 221.400 754.050 222.600 763.950 ;
        RECT 220.950 751.950 223.050 754.050 ;
        RECT 217.950 739.950 220.050 742.050 ;
        RECT 202.950 728.100 205.050 730.200 ;
        RECT 211.950 728.100 214.050 730.200 ;
        RECT 199.950 718.950 202.050 721.050 ;
        RECT 203.400 712.050 204.600 728.100 ;
        RECT 212.400 727.050 213.600 728.100 ;
        RECT 208.950 724.950 211.050 727.050 ;
        RECT 211.950 724.950 214.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 209.400 718.050 210.600 724.950 ;
        RECT 218.400 721.050 219.600 724.950 ;
        RECT 217.950 718.950 220.050 721.050 ;
        RECT 208.950 715.950 211.050 718.050 ;
        RECT 202.950 709.950 205.050 712.050 ;
        RECT 209.400 709.050 210.600 715.950 ;
        RECT 202.950 706.800 205.050 708.900 ;
        RECT 208.950 706.950 211.050 709.050 ;
        RECT 193.950 703.950 196.050 706.050 ;
        RECT 181.950 697.950 184.050 700.050 ;
        RECT 193.950 697.950 196.050 700.050 ;
        RECT 172.950 694.950 175.050 697.050 ;
        RECT 160.950 688.950 163.050 691.050 ;
        RECT 158.400 686.400 162.600 687.600 ;
        RECT 154.950 682.950 157.050 685.050 ;
        RECT 161.400 682.050 162.600 686.400 ;
        RECT 169.950 685.950 172.050 688.050 ;
        RECT 148.950 679.950 151.050 682.050 ;
        RECT 157.950 679.950 160.050 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 145.950 661.950 148.050 664.050 ;
        RECT 149.400 661.050 150.600 679.950 ;
        RECT 154.950 676.950 157.050 679.050 ;
        RECT 127.950 655.950 130.050 658.050 ;
        RECT 130.950 657.000 133.050 661.050 ;
        RECT 142.950 658.950 145.050 661.050 ;
        RECT 148.950 658.950 151.050 661.050 ;
        RECT 118.950 652.950 121.050 655.050 ;
        RECT 124.650 653.400 126.750 655.500 ;
        RECT 115.950 640.950 118.050 643.050 ;
        RECT 106.950 634.950 109.050 637.050 ;
        RECT 112.950 634.950 115.050 637.050 ;
        RECT 115.950 628.950 118.050 631.050 ;
        RECT 103.950 619.950 106.050 622.050 ;
        RECT 73.950 610.950 76.050 613.050 ;
        RECT 112.950 610.950 115.050 613.050 ;
        RECT 73.950 605.100 76.050 607.200 ;
        RECT 79.950 605.100 82.050 607.200 ;
        RECT 85.950 605.100 88.050 607.200 ;
        RECT 100.950 605.100 103.050 607.200 ;
        RECT 70.950 592.950 73.050 595.050 ;
        RECT 74.400 592.050 75.600 605.100 ;
        RECT 80.400 604.050 81.600 605.100 ;
        RECT 86.400 604.050 87.600 605.100 ;
        RECT 101.400 604.050 102.600 605.100 ;
        RECT 79.950 601.950 82.050 604.050 ;
        RECT 82.950 601.950 85.050 604.050 ;
        RECT 85.950 601.950 88.050 604.050 ;
        RECT 88.950 601.950 91.050 604.050 ;
        RECT 97.950 601.950 100.050 604.050 ;
        RECT 100.950 601.950 103.050 604.050 ;
        RECT 103.950 601.950 106.050 604.050 ;
        RECT 76.950 595.950 79.050 601.050 ;
        RECT 83.400 600.900 84.600 601.950 ;
        RECT 82.950 598.800 85.050 600.900 ;
        RECT 61.950 589.950 64.050 592.050 ;
        RECT 73.950 589.950 76.050 592.050 ;
        RECT 55.950 580.950 58.050 583.050 ;
        RECT 76.950 580.950 79.050 583.050 ;
        RECT 43.950 571.950 46.050 574.050 ;
        RECT 52.950 571.950 55.050 574.050 ;
        RECT 61.950 573.000 64.050 577.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 40.950 568.950 43.050 571.050 ;
        RECT 46.950 568.950 49.050 571.050 ;
        RECT 38.400 567.900 39.600 568.950 ;
        RECT 37.950 565.800 40.050 567.900 ;
        RECT 47.400 562.050 48.600 568.950 ;
        RECT 46.950 559.950 49.050 562.050 ;
        RECT 49.950 541.950 52.050 544.050 ;
        RECT 40.950 535.950 43.050 538.050 ;
        RECT 34.950 528.600 37.050 529.050 ;
        RECT 32.400 527.400 37.050 528.600 ;
        RECT 34.950 526.950 37.050 527.400 ;
        RECT 13.950 523.800 16.050 525.900 ;
        RECT 19.950 523.800 22.050 525.900 ;
        RECT 22.950 523.800 25.050 525.900 ;
        RECT 28.950 523.800 31.050 525.900 ;
        RECT 7.950 520.650 10.050 522.750 ;
        RECT 10.950 520.950 13.050 523.050 ;
        RECT 14.400 522.750 15.600 523.800 ;
        RECT 4.950 514.950 7.050 517.050 ;
        RECT 11.400 496.200 12.600 520.950 ;
        RECT 13.950 520.650 16.050 522.750 ;
        RECT 23.400 522.600 24.600 523.800 ;
        RECT 23.400 521.400 27.600 522.600 ;
        RECT 23.400 521.250 24.600 521.400 ;
        RECT 22.950 517.950 25.050 520.050 ;
        RECT 16.950 508.950 19.050 511.050 ;
        RECT 4.950 493.950 7.050 496.050 ;
        RECT 10.950 494.100 13.050 496.200 ;
        RECT 5.400 444.900 6.600 493.950 ;
        RECT 11.400 493.050 12.600 494.100 ;
        RECT 17.400 493.050 18.600 508.950 ;
        RECT 23.400 496.050 24.600 517.950 ;
        RECT 22.950 493.950 25.050 496.050 ;
        RECT 10.950 490.950 13.050 493.050 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 19.950 490.950 22.050 493.050 ;
        RECT 14.400 489.900 15.600 490.950 ;
        RECT 13.950 487.800 16.050 489.900 ;
        RECT 14.400 448.050 15.600 487.800 ;
        RECT 20.400 484.050 21.600 490.950 ;
        RECT 19.950 481.950 22.050 484.050 ;
        RECT 26.400 483.600 27.600 521.400 ;
        RECT 35.400 520.050 36.600 526.950 ;
        RECT 34.950 517.950 37.050 520.050 ;
        RECT 28.950 496.950 31.050 499.050 ;
        RECT 29.400 486.600 30.600 496.950 ;
        RECT 34.950 495.000 37.050 499.050 ;
        RECT 41.400 496.200 42.600 535.950 ;
        RECT 50.400 526.050 51.600 541.950 ;
        RECT 53.400 538.050 54.600 571.950 ;
        RECT 62.400 571.050 63.600 573.000 ;
        RECT 58.950 568.950 61.050 571.050 ;
        RECT 61.950 568.950 64.050 571.050 ;
        RECT 64.950 568.950 67.050 571.050 ;
        RECT 59.400 567.900 60.600 568.950 ;
        RECT 58.950 565.800 61.050 567.900 ;
        RECT 55.950 562.950 58.050 565.050 ;
        RECT 52.950 535.950 55.050 538.050 ;
        RECT 56.400 526.050 57.600 562.950 ;
        RECT 65.400 544.050 66.600 568.950 ;
        RECT 77.400 567.900 78.600 580.950 ;
        RECT 89.400 577.050 90.600 601.950 ;
        RECT 88.950 574.950 91.050 577.050 ;
        RECT 94.950 574.950 97.050 577.050 ;
        RECT 85.950 572.100 88.050 574.200 ;
        RECT 86.400 571.050 87.600 572.100 ;
        RECT 82.950 568.950 85.050 571.050 ;
        RECT 85.950 568.950 88.050 571.050 ;
        RECT 88.950 568.950 91.050 571.050 ;
        RECT 83.400 567.900 84.600 568.950 ;
        RECT 76.950 565.800 79.050 567.900 ;
        RECT 82.950 565.800 85.050 567.900 ;
        RECT 89.400 559.050 90.600 568.950 ;
        RECT 91.950 565.950 94.050 568.050 ;
        RECT 88.950 556.950 91.050 559.050 ;
        RECT 64.950 541.950 67.050 544.050 ;
        RECT 92.400 532.050 93.600 565.950 ;
        RECT 64.950 527.100 67.050 529.200 ;
        RECT 73.950 527.100 76.050 532.050 ;
        RECT 79.950 528.000 82.050 532.050 ;
        RECT 88.950 528.000 91.050 532.050 ;
        RECT 91.950 529.950 94.050 532.050 ;
        RECT 95.400 529.200 96.600 574.950 ;
        RECT 98.400 574.050 99.600 601.950 ;
        RECT 104.400 600.600 105.600 601.950 ;
        RECT 104.400 600.000 108.600 600.600 ;
        RECT 104.400 599.400 109.050 600.000 ;
        RECT 106.950 597.600 109.050 599.400 ;
        RECT 106.950 596.400 111.600 597.600 ;
        RECT 106.950 595.950 109.050 596.400 ;
        RECT 100.950 592.950 103.050 595.050 ;
        RECT 101.400 589.050 102.600 592.950 ;
        RECT 103.950 589.950 106.050 592.050 ;
        RECT 100.950 586.950 103.050 589.050 ;
        RECT 97.950 571.950 100.050 574.050 ;
        RECT 104.400 571.050 105.600 589.950 ;
        RECT 110.400 574.050 111.600 596.400 ;
        RECT 113.400 588.600 114.600 610.950 ;
        RECT 116.400 604.050 117.600 628.950 ;
        RECT 119.400 628.050 120.600 652.950 ;
        RECT 122.400 647.100 124.500 649.200 ;
        RECT 122.400 645.900 123.600 647.100 ;
        RECT 121.950 643.800 124.050 645.900 ;
        RECT 125.400 640.800 126.300 653.400 ;
        RECT 128.400 651.900 129.600 655.950 ;
        RECT 131.400 654.900 132.600 657.000 ;
        RECT 131.400 652.800 133.500 654.900 ;
        RECT 134.700 653.100 136.800 655.200 ;
        RECT 127.200 651.000 129.600 651.900 ;
        RECT 127.200 649.800 134.250 651.000 ;
        RECT 132.150 648.900 134.250 649.800 ;
        RECT 127.200 648.000 129.300 648.900 ;
        RECT 135.150 648.000 136.050 653.100 ;
        RECT 137.400 649.200 138.600 651.600 ;
        RECT 127.200 647.100 136.050 648.000 ;
        RECT 136.950 647.100 139.050 649.200 ;
        RECT 127.200 646.800 129.300 647.100 ;
        RECT 131.400 644.100 133.500 646.200 ;
        RECT 131.400 641.550 132.600 644.100 ;
        RECT 125.100 638.700 127.200 640.800 ;
        RECT 135.150 640.500 136.050 647.100 ;
        RECT 143.400 646.050 144.600 658.950 ;
        RECT 149.400 649.050 150.600 658.950 ;
        RECT 155.400 649.050 156.600 676.950 ;
        RECT 158.400 673.050 159.600 679.950 ;
        RECT 164.400 678.900 165.600 679.950 ;
        RECT 163.950 676.800 166.050 678.900 ;
        RECT 157.950 670.950 160.050 673.050 ;
        RECT 170.400 664.050 171.600 685.950 ;
        RECT 173.400 670.050 174.600 694.950 ;
        RECT 181.950 684.000 184.050 688.050 ;
        RECT 182.400 682.050 183.600 684.000 ;
        RECT 187.950 683.100 190.050 685.200 ;
        RECT 194.400 685.050 195.600 697.950 ;
        RECT 188.400 682.050 189.600 683.100 ;
        RECT 193.950 682.950 196.050 685.050 ;
        RECT 196.950 683.100 199.050 685.200 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 682.050 ;
        RECT 184.950 679.950 187.050 682.050 ;
        RECT 187.950 679.950 190.050 682.050 ;
        RECT 190.950 679.950 193.050 682.050 ;
        RECT 179.400 678.900 180.600 679.950 ;
        RECT 185.400 678.900 186.600 679.950 ;
        RECT 175.800 676.800 177.900 678.900 ;
        RECT 178.950 676.800 181.050 678.900 ;
        RECT 184.950 676.800 187.050 678.900 ;
        RECT 172.950 667.950 175.050 670.050 ;
        RECT 176.400 667.050 177.600 676.800 ;
        RECT 184.950 670.950 187.050 673.050 ;
        RECT 175.950 664.950 178.050 667.050 ;
        RECT 166.800 661.950 168.900 664.050 ;
        RECT 169.950 661.950 172.050 664.050 ;
        RECT 163.950 652.950 166.050 655.050 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 151.950 646.950 154.050 649.050 ;
        RECT 154.950 646.950 157.050 649.050 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 142.950 643.950 145.050 646.050 ;
        RECT 152.400 645.900 153.600 646.950 ;
        RECT 158.400 645.900 159.600 646.950 ;
        RECT 164.400 645.900 165.600 652.950 ;
        RECT 151.950 643.800 154.050 645.900 ;
        RECT 157.950 643.800 160.050 645.900 ;
        RECT 163.950 643.800 166.050 645.900 ;
        RECT 139.950 640.950 142.050 643.050 ;
        RECT 134.100 638.400 136.200 640.500 ;
        RECT 118.950 625.950 121.050 628.050 ;
        RECT 136.950 625.950 139.050 628.050 ;
        RECT 133.950 619.950 136.050 622.050 ;
        RECT 119.100 610.200 121.200 612.300 ;
        RECT 128.100 610.500 130.200 612.600 ;
        RECT 115.950 603.900 118.050 604.050 ;
        RECT 115.950 601.950 118.500 603.900 ;
        RECT 116.400 601.800 118.500 601.950 ;
        RECT 119.400 597.600 120.300 610.200 ;
        RECT 125.400 606.900 126.600 609.450 ;
        RECT 125.400 604.800 127.500 606.900 ;
        RECT 121.200 603.900 123.300 604.200 ;
        RECT 129.150 603.900 130.050 610.500 ;
        RECT 134.400 607.050 135.600 619.950 ;
        RECT 133.950 604.950 136.050 607.050 ;
        RECT 121.200 603.000 130.050 603.900 ;
        RECT 121.200 602.100 123.300 603.000 ;
        RECT 126.150 601.200 128.250 602.100 ;
        RECT 121.200 600.000 128.250 601.200 ;
        RECT 121.200 599.100 123.600 600.000 ;
        RECT 118.650 595.500 120.750 597.600 ;
        RECT 122.400 592.050 123.600 599.100 ;
        RECT 125.400 596.100 127.500 598.200 ;
        RECT 129.150 597.900 130.050 603.000 ;
        RECT 130.950 601.800 133.050 603.900 ;
        RECT 131.400 599.400 132.600 601.800 ;
        RECT 121.950 589.950 124.050 592.050 ;
        RECT 113.400 587.400 117.600 588.600 ;
        RECT 112.950 583.950 115.050 586.050 ;
        RECT 109.950 571.950 112.050 574.050 ;
        RECT 100.950 568.950 103.050 571.050 ;
        RECT 103.950 568.950 106.050 571.050 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 101.400 567.900 102.600 568.950 ;
        RECT 107.400 567.900 108.600 568.950 ;
        RECT 113.400 567.900 114.600 583.950 ;
        RECT 116.400 574.050 117.600 587.400 ;
        RECT 125.400 583.050 126.600 596.100 ;
        RECT 128.700 595.800 130.800 597.900 ;
        RECT 130.950 589.950 133.050 592.050 ;
        RECT 127.950 586.950 130.050 589.050 ;
        RECT 124.950 580.950 127.050 583.050 ;
        RECT 115.950 571.950 118.050 574.050 ;
        RECT 121.950 573.000 124.050 577.050 ;
        RECT 128.400 574.050 129.600 586.950 ;
        RECT 122.400 571.050 123.600 573.000 ;
        RECT 127.950 571.950 130.050 574.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 121.950 568.950 124.050 571.050 ;
        RECT 124.950 568.950 127.050 571.050 ;
        RECT 100.950 565.800 103.050 567.900 ;
        RECT 101.400 559.050 102.600 565.800 ;
        RECT 106.950 562.950 109.050 567.900 ;
        RECT 112.950 565.800 115.050 567.900 ;
        RECT 115.950 565.950 118.050 568.050 ;
        RECT 119.400 567.900 120.600 568.950 ;
        RECT 100.950 556.950 103.050 559.050 ;
        RECT 103.950 547.950 106.050 550.050 ;
        RECT 100.950 532.950 103.050 535.050 ;
        RECT 49.950 523.950 52.050 526.050 ;
        RECT 52.950 523.950 55.050 526.050 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 53.400 522.900 54.600 523.950 ;
        RECT 65.400 523.050 66.600 527.100 ;
        RECT 74.400 526.050 75.600 527.100 ;
        RECT 80.400 526.050 81.600 528.000 ;
        RECT 89.400 526.050 90.600 528.000 ;
        RECT 94.950 527.100 97.050 529.200 ;
        RECT 101.400 529.050 102.600 532.950 ;
        RECT 95.400 526.050 96.600 527.100 ;
        RECT 100.950 526.950 103.050 529.050 ;
        RECT 70.950 523.950 73.050 526.050 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 52.950 520.800 55.050 522.900 ;
        RECT 64.950 520.950 67.050 523.050 ;
        RECT 55.950 502.950 58.050 505.050 ;
        RECT 71.400 504.600 72.600 523.950 ;
        RECT 77.400 522.900 78.600 523.950 ;
        RECT 76.950 520.800 79.050 522.900 ;
        RECT 92.400 519.600 93.600 523.950 ;
        RECT 98.400 522.000 99.600 523.950 ;
        RECT 92.400 518.400 96.600 519.600 ;
        RECT 88.950 514.950 91.050 517.050 ;
        RECT 95.400 516.600 96.600 518.400 ;
        RECT 97.950 517.950 100.050 522.000 ;
        RECT 100.950 520.950 103.050 523.050 ;
        RECT 101.400 516.600 102.600 520.950 ;
        RECT 95.400 515.400 102.600 516.600 ;
        RECT 68.400 503.400 72.600 504.600 ;
        RECT 56.400 496.200 57.600 502.950 ;
        RECT 61.950 499.950 64.050 502.050 ;
        RECT 35.400 493.050 36.600 495.000 ;
        RECT 40.950 494.100 43.050 496.200 ;
        RECT 55.950 494.100 58.050 496.200 ;
        RECT 41.400 493.050 42.600 494.100 ;
        RECT 56.400 493.050 57.600 494.100 ;
        RECT 62.400 493.050 63.600 499.950 ;
        RECT 68.400 493.050 69.600 503.400 ;
        RECT 79.950 502.950 82.050 505.050 ;
        RECT 70.950 499.950 73.050 502.050 ;
        RECT 34.950 490.950 37.050 493.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 55.950 490.950 58.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 61.950 490.950 64.050 493.050 ;
        RECT 67.950 490.950 70.050 493.050 ;
        RECT 29.400 485.400 33.600 486.600 ;
        RECT 28.950 483.600 31.050 484.050 ;
        RECT 26.400 482.400 31.050 483.600 ;
        RECT 28.950 481.950 31.050 482.400 ;
        RECT 25.950 466.950 28.050 469.050 ;
        RECT 26.400 451.200 27.600 466.950 ;
        RECT 19.950 449.100 22.050 451.200 ;
        RECT 25.950 449.100 28.050 451.200 ;
        RECT 20.400 448.050 21.600 449.100 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 11.400 444.900 12.600 445.950 ;
        RECT 17.400 444.900 18.600 445.950 ;
        RECT 4.950 442.800 7.050 444.900 ;
        RECT 10.950 442.800 13.050 444.900 ;
        RECT 16.950 442.800 19.050 444.900 ;
        RECT 19.950 433.950 22.050 436.050 ;
        RECT 7.950 415.950 10.050 418.050 ;
        RECT 13.950 416.100 16.050 418.200 ;
        RECT 1.950 400.950 4.050 403.050 ;
        RECT 8.400 391.050 9.600 415.950 ;
        RECT 14.400 415.050 15.600 416.100 ;
        RECT 20.400 415.050 21.600 433.950 ;
        RECT 26.400 424.050 27.600 449.100 ;
        RECT 25.950 421.950 28.050 424.050 ;
        RECT 13.950 412.950 16.050 415.050 ;
        RECT 16.950 412.950 19.050 415.050 ;
        RECT 19.950 412.950 22.050 415.050 ;
        RECT 22.950 412.950 25.050 415.050 ;
        RECT 17.400 411.000 18.600 412.950 ;
        RECT 23.400 411.900 24.600 412.950 ;
        RECT 16.950 406.950 19.050 411.000 ;
        RECT 22.950 409.800 25.050 411.900 ;
        RECT 29.400 411.600 30.600 481.950 ;
        RECT 32.400 451.200 33.600 485.400 ;
        RECT 38.400 484.050 39.600 490.950 ;
        RECT 44.400 489.900 45.600 490.950 ;
        RECT 53.400 489.900 54.600 490.950 ;
        RECT 59.400 489.900 60.600 490.950 ;
        RECT 43.950 487.800 46.050 489.900 ;
        RECT 52.950 487.800 55.050 489.900 ;
        RECT 58.950 487.800 61.050 489.900 ;
        RECT 37.950 481.950 40.050 484.050 ;
        RECT 46.950 472.950 49.050 475.050 ;
        RECT 31.950 449.100 34.050 451.200 ;
        RECT 40.950 449.100 43.050 454.050 ;
        RECT 41.400 448.050 42.600 449.100 ;
        RECT 47.400 448.050 48.600 472.950 ;
        RECT 59.400 469.050 60.600 487.800 ;
        RECT 68.400 487.050 69.600 490.950 ;
        RECT 67.950 484.950 70.050 487.050 ;
        RECT 71.400 478.050 72.600 499.950 ;
        RECT 80.400 493.050 81.600 502.950 ;
        RECT 85.950 494.100 88.050 496.200 ;
        RECT 89.400 496.050 90.600 514.950 ;
        RECT 104.400 514.050 105.600 547.950 ;
        RECT 112.950 538.950 115.050 541.050 ;
        RECT 113.400 531.600 114.600 538.950 ;
        RECT 116.400 535.050 117.600 565.950 ;
        RECT 118.950 565.800 121.050 567.900 ;
        RECT 125.400 562.050 126.600 568.950 ;
        RECT 127.950 565.950 130.050 568.050 ;
        RECT 124.950 559.950 127.050 562.050 ;
        RECT 115.950 532.950 118.050 535.050 ;
        RECT 113.400 530.400 117.600 531.600 ;
        RECT 109.950 527.100 112.050 529.200 ;
        RECT 110.400 526.050 111.600 527.100 ;
        RECT 116.400 526.050 117.600 530.400 ;
        RECT 124.950 527.100 127.050 529.200 ;
        RECT 109.950 523.950 112.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 94.950 511.950 97.050 514.050 ;
        RECT 103.800 511.950 105.900 514.050 ;
        RECT 106.950 511.950 109.050 514.050 ;
        RECT 91.950 499.950 94.050 502.050 ;
        RECT 86.400 493.050 87.600 494.100 ;
        RECT 88.950 493.950 91.050 496.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 77.400 489.000 78.600 490.950 ;
        RECT 83.400 489.900 84.600 490.950 ;
        RECT 76.950 484.950 79.050 489.000 ;
        RECT 82.950 487.800 85.050 489.900 ;
        RECT 88.950 487.950 91.050 490.050 ;
        RECT 92.400 489.900 93.600 499.950 ;
        RECT 89.400 484.050 90.600 487.950 ;
        RECT 91.950 487.800 94.050 489.900 ;
        RECT 95.400 489.600 96.600 511.950 ;
        RECT 107.400 502.050 108.600 511.950 ;
        RECT 113.400 511.050 114.600 523.950 ;
        RECT 119.400 522.900 120.600 523.950 ;
        RECT 125.400 523.050 126.600 527.100 ;
        RECT 118.950 520.800 121.050 522.900 ;
        RECT 124.950 520.950 127.050 523.050 ;
        RECT 128.400 520.050 129.600 565.950 ;
        RECT 131.400 550.050 132.600 589.950 ;
        RECT 133.950 577.950 136.050 580.050 ;
        RECT 134.400 574.050 135.600 577.950 ;
        RECT 137.400 574.050 138.600 625.950 ;
        RECT 140.400 576.600 141.600 640.950 ;
        RECT 160.950 634.950 163.050 637.050 ;
        RECT 161.400 616.050 162.600 634.950 ;
        RECT 167.400 628.050 168.600 661.950 ;
        RECT 185.400 661.050 186.600 670.950 ;
        RECT 191.400 661.050 192.600 679.950 ;
        RECT 197.400 679.050 198.600 683.100 ;
        RECT 203.400 682.050 204.600 706.800 ;
        RECT 208.950 694.950 211.050 697.050 ;
        RECT 209.400 682.050 210.600 694.950 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 196.950 676.950 199.050 679.050 ;
        RECT 199.950 676.950 202.050 679.050 ;
        RECT 206.400 678.900 207.600 679.950 ;
        RECT 218.400 679.050 219.600 718.950 ;
        RECT 224.400 703.050 225.600 784.950 ;
        RECT 229.950 778.950 232.050 781.050 ;
        RECT 230.400 766.050 231.600 778.950 ;
        RECT 229.950 762.000 232.050 766.050 ;
        RECT 230.400 760.050 231.600 762.000 ;
        RECT 236.400 760.050 237.600 787.950 ;
        RECT 242.400 775.050 243.600 802.950 ;
        RECT 248.400 787.050 249.600 802.950 ;
        RECT 254.400 801.600 255.600 820.950 ;
        RECT 263.400 814.050 264.600 835.950 ;
        RECT 269.400 814.050 270.600 841.950 ;
        RECT 274.950 839.100 277.050 841.200 ;
        RECT 280.950 839.100 283.050 841.200 ;
        RECT 275.400 838.050 276.600 839.100 ;
        RECT 281.400 838.050 282.600 839.100 ;
        RECT 274.950 835.950 277.050 838.050 ;
        RECT 277.950 835.950 280.050 838.050 ;
        RECT 280.950 835.950 283.050 838.050 ;
        RECT 278.400 834.900 279.600 835.950 ;
        RECT 287.400 835.050 288.600 856.950 ;
        RECT 289.950 853.950 292.050 856.050 ;
        RECT 290.400 841.200 291.600 853.950 ;
        RECT 298.950 850.950 301.050 853.050 ;
        RECT 292.950 841.950 295.050 844.050 ;
        RECT 289.950 839.100 292.050 841.200 ;
        RECT 277.950 832.800 280.050 834.900 ;
        RECT 286.950 832.950 289.050 835.050 ;
        RECT 290.400 826.050 291.600 839.100 ;
        RECT 293.400 832.050 294.600 841.950 ;
        RECT 299.400 838.050 300.600 850.950 ;
        RECT 365.400 850.050 366.600 892.950 ;
        RECT 368.400 886.050 369.600 917.100 ;
        RECT 371.400 912.600 372.600 925.950 ;
        RECT 415.950 922.950 418.050 925.050 ;
        RECT 427.950 922.950 430.050 925.050 ;
        RECT 379.950 918.000 382.050 922.050 ;
        RECT 397.950 921.600 402.000 922.050 ;
        RECT 397.950 919.950 402.600 921.600 ;
        RECT 380.400 916.050 381.600 918.000 ;
        RECT 385.950 917.100 388.050 919.200 ;
        RECT 386.400 916.050 387.600 917.100 ;
        RECT 401.400 916.050 402.600 919.950 ;
        RECT 416.400 919.200 417.600 922.950 ;
        RECT 409.950 917.100 412.050 919.200 ;
        RECT 415.950 917.100 418.050 919.200 ;
        RECT 421.950 917.100 424.050 919.200 ;
        RECT 410.400 916.050 411.600 917.100 ;
        RECT 376.950 913.950 379.050 916.050 ;
        RECT 379.950 913.950 382.050 916.050 ;
        RECT 382.950 913.950 385.050 916.050 ;
        RECT 385.950 913.950 388.050 916.050 ;
        RECT 400.950 913.950 403.050 916.050 ;
        RECT 406.950 913.950 409.050 916.050 ;
        RECT 409.950 913.950 412.050 916.050 ;
        RECT 377.400 912.900 378.600 913.950 ;
        RECT 371.400 911.400 375.600 912.600 ;
        RECT 367.950 883.950 370.050 886.050 ;
        RECT 374.400 883.050 375.600 911.400 ;
        RECT 376.950 910.800 379.050 912.900 ;
        RECT 383.400 892.050 384.600 913.950 ;
        RECT 407.400 912.900 408.600 913.950 ;
        RECT 406.950 910.800 409.050 912.900 ;
        RECT 416.400 912.600 417.600 917.100 ;
        RECT 422.400 916.050 423.600 917.100 ;
        RECT 428.400 916.050 429.600 922.950 ;
        RECT 442.950 917.100 445.050 919.200 ;
        RECT 443.400 916.050 444.600 917.100 ;
        RECT 454.950 916.950 457.050 919.050 ;
        RECT 421.950 913.950 424.050 916.050 ;
        RECT 424.950 913.950 427.050 916.050 ;
        RECT 427.950 913.950 430.050 916.050 ;
        RECT 442.950 913.950 445.050 916.050 ;
        RECT 445.950 913.950 448.050 916.050 ;
        RECT 416.400 911.400 420.600 912.600 ;
        RECT 407.400 907.050 408.600 910.800 ;
        RECT 406.950 904.950 409.050 907.050 ;
        RECT 412.950 904.950 415.050 907.050 ;
        RECT 382.950 889.950 385.050 892.050 ;
        RECT 394.950 889.950 397.050 892.050 ;
        RECT 379.950 884.100 382.050 886.200 ;
        RECT 385.950 884.100 388.050 886.200 ;
        RECT 380.400 883.050 381.600 884.100 ;
        RECT 370.950 880.950 373.050 883.050 ;
        RECT 373.950 880.950 376.050 883.050 ;
        RECT 376.950 880.950 379.050 883.050 ;
        RECT 379.950 880.950 382.050 883.050 ;
        RECT 371.400 879.900 372.600 880.950 ;
        RECT 370.950 877.800 373.050 879.900 ;
        RECT 377.400 874.050 378.600 880.950 ;
        RECT 386.400 877.050 387.600 884.100 ;
        RECT 395.400 883.050 396.600 889.950 ;
        RECT 400.950 884.100 403.050 886.200 ;
        RECT 401.400 883.050 402.600 884.100 ;
        RECT 406.950 883.950 409.050 886.050 ;
        RECT 391.950 880.950 394.050 883.050 ;
        RECT 394.950 880.950 397.050 883.050 ;
        RECT 397.950 880.950 400.050 883.050 ;
        RECT 400.950 880.950 403.050 883.050 ;
        RECT 392.400 879.900 393.600 880.950 ;
        RECT 398.400 879.900 399.600 880.950 ;
        RECT 391.950 877.800 394.050 879.900 ;
        RECT 385.950 874.950 388.050 877.050 ;
        RECT 397.950 874.950 400.050 879.900 ;
        RECT 376.950 871.950 379.050 874.050 ;
        RECT 364.950 847.950 367.050 850.050 ;
        RECT 403.950 847.950 406.050 850.050 ;
        RECT 388.950 844.950 391.050 847.050 ;
        RECT 307.950 839.100 310.050 841.200 ;
        RECT 319.950 839.100 322.050 844.050 ;
        RECT 325.950 839.100 328.050 841.200 ;
        RECT 331.950 839.100 334.050 844.050 ;
        RECT 334.950 841.950 337.050 844.050 ;
        RECT 337.950 841.950 340.050 844.050 ;
        RECT 308.400 838.050 309.600 839.100 ;
        RECT 320.400 838.050 321.600 839.100 ;
        RECT 326.400 838.050 327.600 839.100 ;
        RECT 298.950 835.950 301.050 838.050 ;
        RECT 301.950 835.950 304.050 838.050 ;
        RECT 307.950 835.950 310.050 838.050 ;
        RECT 319.950 835.950 322.050 838.050 ;
        RECT 322.950 835.950 325.050 838.050 ;
        RECT 325.950 835.950 328.050 838.050 ;
        RECT 328.950 835.950 331.050 838.050 ;
        RECT 292.950 829.950 295.050 832.050 ;
        RECT 283.950 823.950 289.050 826.050 ;
        RECT 289.950 823.950 292.050 826.050 ;
        RECT 295.950 823.950 298.050 826.050 ;
        RECT 296.400 820.050 297.600 823.950 ;
        RECT 292.800 817.950 294.900 820.050 ;
        RECT 295.950 817.950 298.050 820.050 ;
        RECT 262.950 811.950 265.050 814.050 ;
        RECT 268.950 811.950 271.050 814.050 ;
        RECT 262.950 806.100 265.050 808.200 ;
        RECT 263.400 805.050 264.600 806.100 ;
        RECT 269.400 805.050 270.600 811.950 ;
        RECT 274.950 806.100 277.050 808.200 ;
        RECT 280.950 806.100 283.050 808.200 ;
        RECT 286.950 806.100 289.050 808.200 ;
        RECT 275.400 805.050 276.600 806.100 ;
        RECT 262.950 802.950 265.050 805.050 ;
        RECT 265.950 802.950 268.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 274.950 802.950 277.050 805.050 ;
        RECT 251.400 800.400 255.600 801.600 ;
        RECT 247.950 784.950 250.050 787.050 ;
        RECT 241.950 772.950 244.050 775.050 ;
        RECT 241.950 761.100 244.050 763.200 ;
        RECT 247.950 761.100 250.050 763.200 ;
        RECT 242.400 760.050 243.600 761.100 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 233.400 754.050 234.600 757.950 ;
        RECT 239.400 756.900 240.600 757.950 ;
        RECT 238.950 754.800 241.050 756.900 ;
        RECT 232.950 751.950 235.050 754.050 ;
        RECT 233.400 736.050 234.600 751.950 ;
        RECT 235.950 748.950 238.050 751.050 ;
        RECT 232.950 733.950 235.050 736.050 ;
        RECT 236.400 732.600 237.600 748.950 ;
        RECT 239.400 748.050 240.600 754.800 ;
        RECT 238.950 745.950 241.050 748.050 ;
        RECT 248.400 739.050 249.600 761.100 ;
        RECT 251.400 751.050 252.600 800.400 ;
        RECT 266.400 790.050 267.600 802.950 ;
        RECT 268.950 796.950 271.050 799.050 ;
        RECT 265.950 787.950 268.050 790.050 ;
        RECT 262.950 766.950 265.050 769.050 ;
        RECT 263.400 763.200 264.600 766.950 ;
        RECT 253.950 762.600 258.000 763.050 ;
        RECT 253.950 760.950 258.600 762.600 ;
        RECT 262.950 761.100 265.050 763.200 ;
        RECT 257.400 760.050 258.600 760.950 ;
        RECT 263.400 760.050 264.600 761.100 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 253.950 754.950 256.050 757.050 ;
        RECT 260.400 756.900 261.600 757.950 ;
        RECT 250.950 748.950 253.050 751.050 ;
        RECT 247.950 736.950 250.050 739.050 ;
        RECT 254.400 736.050 255.600 754.950 ;
        RECT 259.950 754.800 262.050 756.900 ;
        RECT 265.950 754.950 268.050 757.050 ;
        RECT 262.950 748.950 265.050 751.050 ;
        RECT 259.950 742.950 262.050 745.050 ;
        RECT 256.950 739.950 259.050 742.050 ;
        RECT 253.950 733.950 256.050 736.050 ;
        RECT 233.400 731.400 237.600 732.600 ;
        RECT 233.400 727.050 234.600 731.400 ;
        RECT 238.950 727.950 241.050 730.050 ;
        RECT 247.950 728.100 250.050 730.200 ;
        RECT 229.950 724.950 232.050 727.050 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 230.400 723.900 231.600 724.950 ;
        RECT 229.950 721.800 232.050 723.900 ;
        RECT 239.400 715.050 240.600 727.950 ;
        RECT 248.400 727.050 249.600 728.100 ;
        RECT 244.950 724.950 247.050 727.050 ;
        RECT 247.950 724.950 250.050 727.050 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 245.400 718.050 246.600 724.950 ;
        RECT 244.950 715.950 247.050 718.050 ;
        RECT 232.950 712.950 235.050 715.050 ;
        RECT 238.950 712.950 241.050 715.050 ;
        RECT 223.950 700.950 226.050 703.050 ;
        RECT 233.400 685.200 234.600 712.950 ;
        RECT 251.400 703.050 252.600 724.950 ;
        RECT 257.400 724.050 258.600 739.950 ;
        RECT 256.950 721.950 259.050 724.050 ;
        RECT 241.950 700.950 244.050 703.050 ;
        RECT 250.950 700.950 253.050 703.050 ;
        RECT 238.950 694.950 241.050 697.050 ;
        RECT 226.950 683.100 229.050 685.200 ;
        RECT 232.950 683.100 235.050 685.200 ;
        RECT 227.400 682.050 228.600 683.100 ;
        RECT 233.400 682.050 234.600 683.100 ;
        RECT 223.950 679.950 226.050 682.050 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 197.400 667.050 198.600 676.950 ;
        RECT 200.400 667.050 201.600 676.950 ;
        RECT 205.950 676.800 208.050 678.900 ;
        RECT 211.950 675.600 214.050 679.050 ;
        RECT 217.950 676.950 220.050 679.050 ;
        RECT 220.950 676.950 223.050 679.050 ;
        RECT 209.400 675.000 214.050 675.600 ;
        RECT 209.400 674.400 213.600 675.000 ;
        RECT 196.800 664.950 198.900 667.050 ;
        RECT 199.950 664.950 202.050 667.050 ;
        RECT 184.950 658.950 187.050 661.050 ;
        RECT 190.950 658.950 193.050 661.050 ;
        RECT 172.950 654.600 175.050 655.050 ;
        RECT 178.950 654.600 181.050 655.050 ;
        RECT 172.950 653.400 181.050 654.600 ;
        RECT 172.950 652.950 175.050 653.400 ;
        RECT 178.950 652.950 181.050 653.400 ;
        RECT 175.950 650.100 178.050 652.200 ;
        RECT 176.400 649.050 177.600 650.100 ;
        RECT 172.950 646.950 175.050 649.050 ;
        RECT 175.950 646.950 178.050 649.050 ;
        RECT 178.950 646.950 181.050 649.050 ;
        RECT 173.400 645.600 174.600 646.950 ;
        RECT 170.400 644.400 174.600 645.600 ;
        RECT 170.400 634.050 171.600 644.400 ;
        RECT 172.950 637.950 175.050 640.050 ;
        RECT 169.950 631.950 172.050 634.050 ;
        RECT 166.950 625.950 169.050 628.050 ;
        RECT 170.400 624.600 171.600 631.950 ;
        RECT 167.400 623.400 171.600 624.600 ;
        RECT 163.950 619.950 166.050 622.050 ;
        RECT 160.950 613.950 163.050 616.050 ;
        RECT 145.800 609.300 147.900 611.400 ;
        RECT 155.400 610.500 157.500 612.600 ;
        RECT 143.400 604.050 144.600 606.600 ;
        RECT 143.400 603.900 145.500 604.050 ;
        RECT 142.950 601.950 145.500 603.900 ;
        RECT 142.950 601.800 145.050 601.950 ;
        RECT 146.700 600.300 147.600 609.300 ;
        RECT 149.100 605.700 151.200 607.800 ;
        RECT 152.400 606.900 153.600 609.450 ;
        RECT 150.300 603.300 151.200 605.700 ;
        RECT 152.100 604.800 154.200 606.900 ;
        RECT 156.000 603.300 157.050 610.500 ;
        RECT 164.400 604.050 165.600 619.950 ;
        RECT 150.300 602.100 157.050 603.300 ;
        RECT 153.150 600.300 155.250 601.200 ;
        RECT 146.700 599.100 155.250 600.300 ;
        RECT 148.200 597.300 150.300 599.100 ;
        RECT 152.100 598.050 154.200 598.200 ;
        RECT 151.950 596.100 154.200 598.050 ;
        RECT 156.150 596.700 157.050 602.100 ;
        RECT 157.950 601.950 160.050 604.050 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 158.400 599.400 159.600 601.950 ;
        RECT 151.950 595.950 154.050 596.100 ;
        RECT 152.400 593.550 153.600 595.950 ;
        RECT 155.400 594.600 157.500 596.700 ;
        RECT 148.950 589.950 151.050 592.050 ;
        RECT 140.400 575.400 144.600 576.600 ;
        RECT 143.400 574.200 144.600 575.400 ;
        RECT 133.950 571.950 136.050 574.050 ;
        RECT 136.950 571.950 139.050 574.050 ;
        RECT 142.950 572.100 145.050 574.200 ;
        RECT 134.400 567.900 135.600 571.950 ;
        RECT 143.400 571.050 144.600 572.100 ;
        RECT 149.400 571.050 150.600 589.950 ;
        RECT 167.400 586.050 168.600 623.400 ;
        RECT 173.400 604.050 174.600 637.950 ;
        RECT 179.400 631.050 180.600 646.950 ;
        RECT 181.950 643.950 184.050 646.050 ;
        RECT 178.950 628.950 181.050 631.050 ;
        RECT 182.400 622.050 183.600 643.950 ;
        RECT 185.400 637.050 186.600 658.950 ;
        RECT 199.950 651.000 202.050 655.050 ;
        RECT 200.400 649.050 201.600 651.000 ;
        RECT 209.400 649.050 210.600 674.400 ;
        RECT 221.400 673.050 222.600 676.950 ;
        RECT 220.950 670.950 223.050 673.050 ;
        RECT 217.950 669.600 220.050 670.050 ;
        RECT 224.400 669.600 225.600 679.950 ;
        RECT 230.400 678.900 231.600 679.950 ;
        RECT 229.950 676.800 232.050 678.900 ;
        RECT 217.950 668.400 225.600 669.600 ;
        RECT 217.950 667.950 220.050 668.400 ;
        RECT 211.950 664.950 214.050 667.050 ;
        RECT 212.400 649.050 213.600 664.950 ;
        RECT 223.950 655.950 226.050 658.050 ;
        RECT 235.950 655.950 238.050 658.050 ;
        RECT 220.200 653.100 222.300 655.200 ;
        RECT 224.400 654.900 225.600 655.950 ;
        RECT 218.400 649.200 219.600 651.600 ;
        RECT 190.950 646.950 193.050 649.050 ;
        RECT 196.950 646.950 199.050 649.050 ;
        RECT 199.950 646.950 202.050 649.050 ;
        RECT 202.950 646.950 205.050 649.050 ;
        RECT 208.800 646.950 210.900 649.050 ;
        RECT 211.950 646.950 214.050 649.050 ;
        RECT 217.950 647.100 220.050 649.200 ;
        RECT 220.950 648.000 221.850 653.100 ;
        RECT 223.500 652.800 225.600 654.900 ;
        RECT 230.250 653.400 232.350 655.500 ;
        RECT 227.700 651.000 229.800 651.900 ;
        RECT 222.750 649.800 229.800 651.000 ;
        RECT 222.750 648.900 224.850 649.800 ;
        RECT 227.700 648.000 229.800 648.900 ;
        RECT 220.950 647.100 229.800 648.000 ;
        RECT 184.950 634.950 187.050 637.050 ;
        RECT 191.400 630.600 192.600 646.950 ;
        RECT 197.400 645.000 198.600 646.950 ;
        RECT 203.400 645.000 204.600 646.950 ;
        RECT 196.950 640.950 199.050 645.000 ;
        RECT 202.950 640.950 205.050 645.000 ;
        RECT 214.950 643.800 217.050 645.900 ;
        RECT 193.950 630.600 196.050 631.050 ;
        RECT 191.400 629.400 196.050 630.600 ;
        RECT 193.950 628.950 196.050 629.400 ;
        RECT 181.950 619.950 184.050 622.050 ;
        RECT 187.950 613.950 190.050 616.050 ;
        RECT 178.950 605.100 181.050 607.200 ;
        RECT 179.400 604.050 180.600 605.100 ;
        RECT 172.950 601.950 175.050 604.050 ;
        RECT 175.950 601.950 178.050 604.050 ;
        RECT 178.950 601.950 181.050 604.050 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 176.400 597.600 177.600 601.950 ;
        RECT 173.400 596.400 177.600 597.600 ;
        RECT 154.950 583.950 157.050 586.050 ;
        RECT 166.950 583.950 169.050 586.050 ;
        RECT 139.950 568.950 142.050 571.050 ;
        RECT 142.950 568.950 145.050 571.050 ;
        RECT 145.950 568.950 148.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 140.400 567.900 141.600 568.950 ;
        RECT 133.950 565.800 136.050 567.900 ;
        RECT 139.950 565.800 142.050 567.900 ;
        RECT 146.400 567.000 147.600 568.950 ;
        RECT 136.950 562.950 139.050 565.050 ;
        RECT 145.950 562.950 148.050 567.000 ;
        RECT 133.950 556.950 136.050 559.050 ;
        RECT 130.950 547.950 133.050 550.050 ;
        RECT 134.400 546.600 135.600 556.950 ;
        RECT 131.400 545.400 135.600 546.600 ;
        RECT 127.950 517.950 130.050 520.050 ;
        RECT 131.400 517.050 132.600 545.400 ;
        RECT 137.400 529.200 138.600 562.950 ;
        RECT 155.400 559.050 156.600 583.950 ;
        RECT 173.400 580.050 174.600 596.400 ;
        RECT 178.950 589.950 181.050 592.050 ;
        RECT 175.950 583.950 178.050 586.050 ;
        RECT 172.950 577.950 175.050 580.050 ;
        RECT 163.950 572.100 166.050 574.200 ;
        RECT 169.950 572.100 172.050 574.200 ;
        RECT 164.400 571.050 165.600 572.100 ;
        RECT 170.400 571.050 171.600 572.100 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 163.950 568.950 166.050 571.050 ;
        RECT 166.950 568.950 169.050 571.050 ;
        RECT 169.950 568.950 172.050 571.050 ;
        RECT 161.400 568.050 162.600 568.950 ;
        RECT 157.950 566.400 162.600 568.050 ;
        RECT 157.950 565.950 162.000 566.400 ;
        RECT 167.400 565.050 168.600 568.950 ;
        RECT 176.400 565.050 177.600 583.950 ;
        RECT 166.950 562.950 169.050 565.050 ;
        RECT 175.950 562.950 178.050 565.050 ;
        RECT 154.950 556.950 157.050 559.050 ;
        RECT 148.950 550.950 151.050 553.050 ;
        RECT 142.950 538.950 145.050 541.050 ;
        RECT 143.400 535.050 144.600 538.950 ;
        RECT 142.950 532.950 145.050 535.050 ;
        RECT 136.950 527.100 139.050 529.200 ;
        RECT 137.400 526.050 138.600 527.100 ;
        RECT 143.400 526.050 144.600 532.950 ;
        RECT 149.400 529.050 150.600 550.950 ;
        RECT 160.950 538.950 163.050 541.050 ;
        RECT 151.950 532.950 154.050 535.050 ;
        RECT 148.950 526.950 151.050 529.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 133.950 520.950 136.050 523.050 ;
        RECT 140.400 522.900 141.600 523.950 ;
        RECT 130.950 514.950 133.050 517.050 ;
        RECT 134.400 514.050 135.600 520.950 ;
        RECT 139.950 520.800 142.050 522.900 ;
        RECT 146.400 522.000 147.600 523.950 ;
        RECT 145.950 517.950 148.050 522.000 ;
        RECT 136.950 514.950 139.050 517.050 ;
        RECT 133.950 511.950 136.050 514.050 ;
        RECT 112.950 508.950 115.050 511.050 ;
        RECT 127.950 508.950 130.050 511.050 ;
        RECT 113.400 505.050 114.600 508.950 ;
        RECT 112.950 502.950 115.050 505.050 ;
        RECT 106.950 499.950 109.050 502.050 ;
        RECT 97.950 495.600 102.000 496.050 ;
        RECT 97.950 493.950 102.600 495.600 ;
        RECT 106.950 494.100 109.050 496.200 ;
        RECT 113.400 496.050 114.600 502.950 ;
        RECT 101.400 493.050 102.600 493.950 ;
        RECT 107.400 493.050 108.600 494.100 ;
        RECT 112.950 493.950 115.050 496.050 ;
        RECT 115.950 494.100 118.050 496.200 ;
        RECT 121.950 494.100 124.050 496.200 ;
        RECT 100.950 490.950 103.050 493.050 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 104.400 489.900 105.600 490.950 ;
        RECT 110.400 490.050 111.600 490.950 ;
        RECT 95.400 488.400 99.600 489.600 ;
        RECT 94.950 484.950 97.050 487.050 ;
        RECT 88.950 481.950 91.050 484.050 ;
        RECT 70.950 475.950 73.050 478.050 ;
        RECT 64.950 472.950 67.050 475.050 ;
        RECT 58.950 466.950 61.050 469.050 ;
        RECT 52.950 451.950 55.050 454.050 ;
        RECT 37.950 445.950 40.050 448.050 ;
        RECT 40.950 445.950 43.050 448.050 ;
        RECT 43.950 445.950 46.050 448.050 ;
        RECT 46.950 445.950 49.050 448.050 ;
        RECT 38.400 430.050 39.600 445.950 ;
        RECT 44.400 444.900 45.600 445.950 ;
        RECT 43.950 442.800 46.050 444.900 ;
        RECT 40.950 433.950 43.050 436.050 ;
        RECT 31.950 427.950 34.050 430.050 ;
        RECT 37.950 427.950 40.050 430.050 ;
        RECT 32.400 418.050 33.600 427.950 ;
        RECT 41.400 420.600 42.600 433.950 ;
        RECT 49.950 421.950 52.050 424.050 ;
        RECT 38.400 419.400 42.600 420.600 ;
        RECT 31.950 415.950 34.050 418.050 ;
        RECT 38.400 415.050 39.600 419.400 ;
        RECT 43.950 416.100 46.050 418.200 ;
        RECT 44.400 415.050 45.600 416.100 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 37.950 412.950 40.050 415.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 43.950 412.950 46.050 415.050 ;
        RECT 35.400 411.900 36.600 412.950 ;
        RECT 26.400 410.400 30.600 411.600 ;
        RECT 22.950 400.950 25.050 403.050 ;
        RECT 7.950 388.950 10.050 391.050 ;
        RECT 1.950 385.950 4.050 388.050 ;
        RECT 2.400 37.050 3.600 385.950 ;
        RECT 4.950 376.950 7.050 379.050 ;
        RECT 5.400 358.050 6.600 376.950 ;
        RECT 10.950 371.100 13.050 373.200 ;
        RECT 19.950 371.100 22.050 373.200 ;
        RECT 23.400 373.050 24.600 400.950 ;
        RECT 11.400 370.050 12.600 371.100 ;
        RECT 20.400 370.050 21.600 371.100 ;
        RECT 22.950 370.950 25.050 373.050 ;
        RECT 10.950 367.950 13.050 370.050 ;
        RECT 13.950 367.950 16.050 370.050 ;
        RECT 19.950 367.950 22.050 370.050 ;
        RECT 7.950 361.950 10.050 364.050 ;
        RECT 4.950 355.950 7.050 358.050 ;
        RECT 4.950 277.950 7.050 280.050 ;
        RECT 5.400 181.050 6.600 277.950 ;
        RECT 8.400 271.050 9.600 361.950 ;
        RECT 14.400 358.050 15.600 367.950 ;
        RECT 16.950 364.950 19.050 367.050 ;
        RECT 13.950 355.950 16.050 358.050 ;
        RECT 17.400 352.050 18.600 364.950 ;
        RECT 26.400 364.050 27.600 410.400 ;
        RECT 34.950 409.800 37.050 411.900 ;
        RECT 31.950 394.950 34.050 397.050 ;
        RECT 32.400 379.050 33.600 394.950 ;
        RECT 41.400 385.050 42.600 412.950 ;
        RECT 46.950 406.950 49.050 409.050 ;
        RECT 43.950 400.950 46.050 403.050 ;
        RECT 40.950 382.950 43.050 385.050 ;
        RECT 37.950 379.950 40.050 382.050 ;
        RECT 31.950 376.950 34.050 379.050 ;
        RECT 32.400 370.050 33.600 376.950 ;
        RECT 38.400 373.200 39.600 379.950 ;
        RECT 37.950 371.100 40.050 373.200 ;
        RECT 38.400 370.050 39.600 371.100 ;
        RECT 31.950 367.950 34.050 370.050 ;
        RECT 34.950 367.950 37.050 370.050 ;
        RECT 37.950 367.950 40.050 370.050 ;
        RECT 25.800 361.950 27.900 364.050 ;
        RECT 28.950 361.950 31.050 367.050 ;
        RECT 10.950 349.950 13.050 352.050 ;
        RECT 16.950 349.950 19.050 352.050 ;
        RECT 28.950 349.950 31.050 352.050 ;
        RECT 11.400 340.050 12.600 349.950 ;
        RECT 16.950 343.950 19.050 346.050 ;
        RECT 10.950 337.950 13.050 340.050 ;
        RECT 17.400 337.050 18.600 343.950 ;
        RECT 22.950 338.100 25.050 340.200 ;
        RECT 23.400 337.050 24.600 338.100 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 16.950 334.950 19.050 337.050 ;
        RECT 19.950 334.950 22.050 337.050 ;
        RECT 22.950 334.950 25.050 337.050 ;
        RECT 14.400 333.900 15.600 334.950 ;
        RECT 13.950 331.800 16.050 333.900 ;
        RECT 13.950 328.650 16.050 330.750 ;
        RECT 14.400 304.050 15.600 328.650 ;
        RECT 20.400 319.050 21.600 334.950 ;
        RECT 25.950 331.950 28.050 334.050 ;
        RECT 29.400 333.600 30.600 349.950 ;
        RECT 35.400 340.200 36.600 367.950 ;
        RECT 44.400 358.050 45.600 400.950 ;
        RECT 37.950 355.950 40.050 358.050 ;
        RECT 43.950 355.950 46.050 358.050 ;
        RECT 38.400 346.050 39.600 355.950 ;
        RECT 43.950 349.950 46.050 352.050 ;
        RECT 37.950 343.950 40.050 346.050 ;
        RECT 39.000 342.600 43.050 343.050 ;
        RECT 38.400 340.950 43.050 342.600 ;
        RECT 34.950 339.600 37.050 340.200 ;
        RECT 32.400 339.000 37.050 339.600 ;
        RECT 31.950 338.400 37.050 339.000 ;
        RECT 31.950 334.950 34.050 338.400 ;
        RECT 34.950 338.100 37.050 338.400 ;
        RECT 38.400 337.050 39.600 340.950 ;
        RECT 44.400 337.050 45.600 349.950 ;
        RECT 47.400 343.050 48.600 406.950 ;
        RECT 50.400 403.050 51.600 421.950 ;
        RECT 53.400 409.050 54.600 451.950 ;
        RECT 58.950 450.000 61.050 454.050 ;
        RECT 59.400 448.050 60.600 450.000 ;
        RECT 65.400 448.050 66.600 472.950 ;
        RECT 73.950 457.950 76.050 460.050 ;
        RECT 58.950 445.950 61.050 448.050 ;
        RECT 61.950 445.950 64.050 448.050 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 67.950 445.950 70.050 448.050 ;
        RECT 62.400 444.900 63.600 445.950 ;
        RECT 68.400 444.900 69.600 445.950 ;
        RECT 74.400 445.050 75.600 457.950 ;
        RECT 76.950 449.100 79.050 451.200 ;
        RECT 82.950 449.100 85.050 451.200 ;
        RECT 88.950 450.000 91.050 454.050 ;
        RECT 95.400 451.050 96.600 484.950 ;
        RECT 61.950 442.800 64.050 444.900 ;
        RECT 67.950 442.800 70.050 444.900 ;
        RECT 73.950 442.950 76.050 445.050 ;
        RECT 58.950 430.950 61.050 433.050 ;
        RECT 59.400 415.050 60.600 430.950 ;
        RECT 77.400 430.050 78.600 449.100 ;
        RECT 83.400 448.050 84.600 449.100 ;
        RECT 89.400 448.050 90.600 450.000 ;
        RECT 94.950 448.950 97.050 451.050 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 91.950 445.950 94.050 448.050 ;
        RECT 86.400 444.900 87.600 445.950 ;
        RECT 85.950 442.800 88.050 444.900 ;
        RECT 86.400 436.050 87.600 442.800 ;
        RECT 92.400 439.050 93.600 445.950 ;
        RECT 94.950 439.950 97.050 442.050 ;
        RECT 91.950 436.950 94.050 439.050 ;
        RECT 85.950 433.950 88.050 436.050 ;
        RECT 76.950 427.950 79.050 430.050 ;
        RECT 82.950 424.950 85.050 427.050 ;
        RECT 73.950 421.950 76.050 424.050 ;
        RECT 64.950 416.100 67.050 418.200 ;
        RECT 65.400 415.050 66.600 416.100 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 61.950 412.950 64.050 415.050 ;
        RECT 64.950 412.950 67.050 415.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 62.400 411.900 63.600 412.950 ;
        RECT 52.950 406.950 55.050 409.050 ;
        RECT 61.950 406.950 64.050 411.900 ;
        RECT 68.400 411.600 69.600 412.950 ;
        RECT 74.400 411.900 75.600 421.950 ;
        RECT 83.400 418.200 84.600 424.950 ;
        RECT 82.950 416.100 85.050 418.200 ;
        RECT 88.950 416.100 91.050 418.200 ;
        RECT 83.400 415.050 84.600 416.100 ;
        RECT 89.400 415.050 90.600 416.100 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 82.950 412.950 85.050 415.050 ;
        RECT 85.950 412.950 88.050 415.050 ;
        RECT 88.950 412.950 91.050 415.050 ;
        RECT 73.950 411.600 76.050 411.900 ;
        RECT 68.400 410.400 76.050 411.600 ;
        RECT 80.400 411.000 81.600 412.950 ;
        RECT 86.400 411.900 87.600 412.950 ;
        RECT 73.950 409.800 76.050 410.400 ;
        RECT 79.950 406.950 82.050 411.000 ;
        RECT 85.950 409.800 88.050 411.900 ;
        RECT 76.950 403.950 79.050 406.050 ;
        RECT 49.950 400.950 52.050 403.050 ;
        RECT 77.400 391.050 78.600 403.950 ;
        RECT 76.950 388.950 79.050 391.050 ;
        RECT 95.400 385.050 96.600 439.950 ;
        RECT 98.400 394.050 99.600 488.400 ;
        RECT 103.950 487.800 106.050 489.900 ;
        RECT 110.400 488.400 115.050 490.050 ;
        RECT 111.000 487.950 115.050 488.400 ;
        RECT 106.950 484.950 109.050 487.050 ;
        RECT 107.400 478.050 108.600 484.950 ;
        RECT 106.950 475.950 109.050 478.050 ;
        RECT 116.400 475.050 117.600 494.100 ;
        RECT 122.400 493.050 123.600 494.100 ;
        RECT 128.400 493.050 129.600 508.950 ;
        RECT 134.400 496.050 135.600 511.950 ;
        RECT 133.950 493.950 136.050 496.050 ;
        RECT 121.950 490.950 124.050 493.050 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 127.950 490.950 130.050 493.050 ;
        RECT 130.950 490.950 133.050 493.050 ;
        RECT 125.400 489.000 126.600 490.950 ;
        RECT 131.400 489.900 132.600 490.950 ;
        RECT 124.950 484.950 127.050 489.000 ;
        RECT 130.950 487.800 133.050 489.900 ;
        RECT 137.400 481.050 138.600 514.950 ;
        RECT 152.400 511.050 153.600 532.950 ;
        RECT 161.400 526.050 162.600 538.950 ;
        RECT 167.400 535.050 168.600 562.950 ;
        RECT 172.950 556.950 175.050 559.050 ;
        RECT 166.950 532.950 169.050 535.050 ;
        RECT 167.400 526.050 168.600 532.950 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 166.950 523.950 169.050 526.050 ;
        RECT 158.400 522.600 159.600 523.950 ;
        RECT 155.400 522.000 159.600 522.600 ;
        RECT 154.950 521.400 159.600 522.000 ;
        RECT 154.950 517.950 157.050 521.400 ;
        RECT 164.400 517.050 165.600 523.950 ;
        RECT 163.950 514.950 166.050 517.050 ;
        RECT 173.400 511.050 174.600 556.950 ;
        RECT 175.950 538.950 178.050 541.050 ;
        RECT 151.950 508.950 154.050 511.050 ;
        RECT 172.950 508.950 175.050 511.050 ;
        RECT 148.950 502.950 151.050 505.050 ;
        RECT 154.950 502.950 157.050 505.050 ;
        RECT 166.950 502.950 169.050 505.050 ;
        RECT 172.950 502.950 175.050 505.050 ;
        RECT 149.400 493.050 150.600 502.950 ;
        RECT 155.400 493.050 156.600 502.950 ;
        RECT 167.400 499.050 168.600 502.950 ;
        RECT 173.400 499.050 174.600 502.950 ;
        RECT 166.950 496.950 169.050 499.050 ;
        RECT 172.950 496.950 175.050 499.050 ;
        RECT 173.400 493.050 174.600 496.950 ;
        RECT 176.400 496.050 177.600 538.950 ;
        RECT 179.400 535.050 180.600 589.950 ;
        RECT 182.400 567.900 183.600 601.950 ;
        RECT 188.400 595.050 189.600 613.950 ;
        RECT 190.950 605.100 193.050 607.200 ;
        RECT 187.950 592.950 190.050 595.050 ;
        RECT 184.950 589.950 187.050 592.050 ;
        RECT 185.400 574.050 186.600 589.950 ;
        RECT 191.400 586.050 192.600 605.100 ;
        RECT 194.400 601.050 195.600 628.950 ;
        RECT 199.950 625.950 202.050 628.050 ;
        RECT 200.400 610.050 201.600 625.950 ;
        RECT 215.400 616.050 216.600 643.800 ;
        RECT 220.950 640.500 221.850 647.100 ;
        RECT 227.700 646.800 229.800 647.100 ;
        RECT 223.500 644.100 225.600 646.200 ;
        RECT 224.400 641.550 225.600 644.100 ;
        RECT 230.700 640.800 231.600 653.400 ;
        RECT 232.500 647.100 234.600 649.200 ;
        RECT 236.400 649.050 237.600 655.950 ;
        RECT 233.400 645.000 234.600 647.100 ;
        RECT 235.950 646.950 238.050 649.050 ;
        RECT 232.950 640.950 235.050 645.000 ;
        RECT 220.800 638.400 222.900 640.500 ;
        RECT 229.800 638.700 231.900 640.800 ;
        RECT 220.950 634.950 223.050 637.050 ;
        RECT 205.950 613.950 208.050 616.050 ;
        RECT 214.950 613.950 217.050 616.050 ;
        RECT 199.950 607.950 202.050 610.050 ;
        RECT 200.400 604.050 201.600 607.950 ;
        RECT 206.400 604.050 207.600 613.950 ;
        RECT 214.950 607.950 217.050 610.050 ;
        RECT 211.950 604.950 214.050 607.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 202.950 601.950 205.050 604.050 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 193.950 598.950 196.050 601.050 ;
        RECT 190.950 583.950 193.050 586.050 ;
        RECT 190.950 577.950 193.050 580.050 ;
        RECT 184.950 571.950 187.050 574.050 ;
        RECT 191.400 571.050 192.600 577.950 ;
        RECT 196.950 572.100 199.050 574.200 ;
        RECT 203.400 574.050 204.600 601.950 ;
        RECT 208.950 592.950 211.050 595.050 ;
        RECT 209.400 576.600 210.600 592.950 ;
        RECT 212.400 592.050 213.600 604.950 ;
        RECT 211.950 589.950 214.050 592.050 ;
        RECT 215.400 583.050 216.600 607.950 ;
        RECT 221.400 607.200 222.600 634.950 ;
        RECT 239.400 634.050 240.600 694.950 ;
        RECT 242.400 634.050 243.600 700.950 ;
        RECT 260.400 700.050 261.600 742.950 ;
        RECT 259.950 697.950 262.050 700.050 ;
        RECT 256.950 691.950 259.050 694.050 ;
        RECT 257.400 685.200 258.600 691.950 ;
        RECT 250.950 683.100 253.050 685.200 ;
        RECT 256.950 683.100 259.050 685.200 ;
        RECT 251.400 682.050 252.600 683.100 ;
        RECT 257.400 682.050 258.600 683.100 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 248.400 664.050 249.600 679.950 ;
        RECT 254.400 678.000 255.600 679.950 ;
        RECT 253.950 670.950 256.050 678.000 ;
        RECT 259.950 673.950 262.050 676.050 ;
        RECT 247.950 661.950 250.050 664.050 ;
        RECT 250.950 658.950 253.050 661.050 ;
        RECT 251.400 649.050 252.600 658.950 ;
        RECT 247.950 646.950 250.050 649.050 ;
        RECT 250.950 646.950 253.050 649.050 ;
        RECT 253.950 646.950 256.050 649.050 ;
        RECT 244.950 643.950 247.050 646.050 ;
        RECT 238.800 631.950 240.900 634.050 ;
        RECT 241.950 631.950 244.050 634.050 ;
        RECT 238.950 628.800 241.050 630.900 ;
        RECT 235.950 625.950 238.050 628.050 ;
        RECT 229.950 622.950 232.050 625.050 ;
        RECT 220.950 605.100 223.050 607.200 ;
        RECT 221.400 604.050 222.600 605.100 ;
        RECT 230.400 604.050 231.600 622.950 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 223.950 601.950 226.050 604.050 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 224.400 600.900 225.600 601.950 ;
        RECT 223.950 598.800 226.050 600.900 ;
        RECT 232.950 598.950 235.050 601.050 ;
        RECT 217.950 592.950 220.050 595.050 ;
        RECT 214.950 580.950 217.050 583.050 ;
        RECT 209.400 575.400 213.600 576.600 ;
        RECT 197.400 571.050 198.600 572.100 ;
        RECT 202.950 571.950 205.050 574.050 ;
        RECT 212.400 571.050 213.600 575.400 ;
        RECT 218.400 571.050 219.600 592.950 ;
        RECT 224.400 577.050 225.600 598.800 ;
        RECT 229.950 580.950 232.050 583.050 ;
        RECT 226.950 577.950 229.050 580.050 ;
        RECT 223.950 574.950 226.050 577.050 ;
        RECT 223.950 571.800 226.050 573.900 ;
        RECT 187.950 568.950 190.050 571.050 ;
        RECT 190.950 568.950 193.050 571.050 ;
        RECT 193.950 568.950 196.050 571.050 ;
        RECT 196.950 568.950 199.050 571.050 ;
        RECT 181.950 565.800 184.050 567.900 ;
        RECT 184.950 565.950 187.050 568.050 ;
        RECT 188.400 567.900 189.600 568.950 ;
        RECT 194.400 567.900 195.600 568.950 ;
        RECT 202.950 568.800 205.050 570.900 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 217.950 568.950 220.050 571.050 ;
        RECT 185.400 541.050 186.600 565.950 ;
        RECT 187.950 565.800 190.050 567.900 ;
        RECT 193.950 565.800 196.050 567.900 ;
        RECT 199.950 565.950 202.050 568.050 ;
        RECT 188.400 547.050 189.600 565.800 ;
        RECT 187.950 544.950 190.050 547.050 ;
        RECT 184.950 538.950 187.050 541.050 ;
        RECT 200.400 535.050 201.600 565.950 ;
        RECT 203.400 562.050 204.600 568.800 ;
        RECT 205.950 565.950 208.050 568.050 ;
        RECT 202.950 559.950 205.050 562.050 ;
        RECT 206.400 538.050 207.600 565.950 ;
        RECT 209.400 562.050 210.600 568.950 ;
        RECT 215.400 567.900 216.600 568.950 ;
        RECT 214.950 565.800 217.050 567.900 ;
        RECT 208.950 559.950 211.050 562.050 ;
        RECT 205.950 535.950 208.050 538.050 ;
        RECT 178.950 532.950 181.050 535.050 ;
        RECT 187.950 532.950 190.050 535.050 ;
        RECT 193.950 532.950 196.050 535.050 ;
        RECT 199.950 532.950 202.050 535.050 ;
        RECT 188.400 529.200 189.600 532.950 ;
        RECT 187.950 527.100 190.050 529.200 ;
        RECT 188.400 526.050 189.600 527.100 ;
        RECT 194.400 526.050 195.600 532.950 ;
        RECT 208.950 527.100 211.050 529.200 ;
        RECT 214.950 527.100 217.050 529.200 ;
        RECT 224.400 528.600 225.600 571.800 ;
        RECT 227.400 567.900 228.600 577.950 ;
        RECT 226.950 565.800 229.050 567.900 ;
        RECT 230.400 562.050 231.600 580.950 ;
        RECT 233.400 574.050 234.600 598.950 ;
        RECT 236.400 595.050 237.600 625.950 ;
        RECT 239.400 607.050 240.600 628.800 ;
        RECT 245.400 615.600 246.600 643.950 ;
        RECT 248.400 619.050 249.600 646.950 ;
        RECT 250.950 637.950 253.050 640.050 ;
        RECT 247.950 616.950 250.050 619.050 ;
        RECT 245.400 614.400 249.600 615.600 ;
        RECT 238.950 604.950 241.050 607.050 ;
        RECT 244.950 605.100 247.050 607.200 ;
        RECT 248.400 607.050 249.600 614.400 ;
        RECT 245.400 604.050 246.600 605.100 ;
        RECT 247.950 604.950 250.050 607.050 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 238.950 598.950 241.050 601.050 ;
        RECT 235.950 592.950 238.050 595.050 ;
        RECT 239.400 592.050 240.600 598.950 ;
        RECT 242.400 597.600 243.600 601.950 ;
        RECT 251.400 600.600 252.600 637.950 ;
        RECT 254.400 637.050 255.600 646.950 ;
        RECT 256.950 643.950 259.050 646.050 ;
        RECT 253.950 634.950 256.050 637.050 ;
        RECT 257.400 633.600 258.600 643.950 ;
        RECT 260.400 640.050 261.600 673.950 ;
        RECT 263.400 673.050 264.600 748.950 ;
        RECT 266.400 748.050 267.600 754.950 ;
        RECT 269.400 754.050 270.600 796.950 ;
        RECT 272.400 796.050 273.600 802.950 ;
        RECT 281.400 799.050 282.600 806.100 ;
        RECT 287.400 805.050 288.600 806.100 ;
        RECT 293.400 805.050 294.600 817.950 ;
        RECT 302.400 817.050 303.600 835.950 ;
        RECT 323.400 834.900 324.600 835.950 ;
        RECT 322.950 832.800 325.050 834.900 ;
        RECT 316.950 829.950 319.050 832.050 ;
        RECT 301.950 814.950 304.050 817.050 ;
        RECT 301.950 806.100 304.050 808.200 ;
        RECT 307.950 806.100 310.050 808.200 ;
        RECT 286.950 802.950 289.050 805.050 ;
        RECT 289.950 802.950 292.050 805.050 ;
        RECT 292.950 802.950 295.050 805.050 ;
        RECT 295.950 802.950 298.050 805.050 ;
        RECT 280.950 796.950 283.050 799.050 ;
        RECT 290.400 796.050 291.600 802.950 ;
        RECT 296.400 801.000 297.600 802.950 ;
        RECT 295.950 796.950 298.050 801.000 ;
        RECT 271.950 793.950 274.050 796.050 ;
        RECT 289.950 793.950 292.050 796.050 ;
        RECT 272.400 763.050 273.600 793.950 ;
        RECT 290.400 787.050 291.600 793.950 ;
        RECT 302.400 790.050 303.600 806.100 ;
        RECT 308.400 805.050 309.600 806.100 ;
        RECT 307.950 802.950 310.050 805.050 ;
        RECT 310.950 802.950 313.050 805.050 ;
        RECT 311.400 799.050 312.600 802.950 ;
        RECT 307.950 797.400 312.600 799.050 ;
        RECT 307.950 796.950 312.000 797.400 ;
        RECT 310.950 793.950 313.050 796.050 ;
        RECT 301.950 787.950 304.050 790.050 ;
        RECT 307.950 787.950 310.050 790.050 ;
        RECT 286.800 784.950 288.900 787.050 ;
        RECT 289.950 784.950 292.050 787.050 ;
        RECT 287.400 781.050 288.600 784.950 ;
        RECT 301.950 781.950 304.050 784.050 ;
        RECT 280.950 778.950 283.050 781.050 ;
        RECT 286.950 778.950 289.050 781.050 ;
        RECT 271.800 760.950 273.900 763.050 ;
        RECT 274.950 761.100 277.050 763.200 ;
        RECT 275.400 760.050 276.600 761.100 ;
        RECT 281.400 760.050 282.600 778.950 ;
        RECT 286.950 761.100 289.050 763.200 ;
        RECT 292.950 761.100 295.050 763.200 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 278.400 756.000 279.600 757.950 ;
        RECT 268.950 751.950 271.050 754.050 ;
        RECT 277.950 751.950 280.050 756.000 ;
        RECT 283.950 754.950 286.050 757.050 ;
        RECT 265.950 745.950 268.050 748.050 ;
        RECT 271.950 733.950 274.050 736.050 ;
        RECT 272.400 730.200 273.600 733.950 ;
        RECT 271.950 728.100 274.050 730.200 ;
        RECT 272.400 727.050 273.600 728.100 ;
        RECT 268.950 724.950 271.050 727.050 ;
        RECT 271.950 724.950 274.050 727.050 ;
        RECT 277.950 724.950 280.050 727.050 ;
        RECT 269.400 711.600 270.600 724.950 ;
        RECT 278.400 723.900 279.600 724.950 ;
        RECT 277.950 721.800 280.050 723.900 ;
        RECT 280.950 717.600 283.050 718.050 ;
        RECT 284.400 717.600 285.600 754.950 ;
        RECT 287.400 754.050 288.600 761.100 ;
        RECT 293.400 760.050 294.600 761.100 ;
        RECT 302.400 760.050 303.600 781.950 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 301.950 757.950 304.050 760.050 ;
        RECT 286.950 751.950 289.050 754.050 ;
        RECT 292.950 751.950 295.050 754.050 ;
        RECT 293.400 727.050 294.600 751.950 ;
        RECT 296.400 748.050 297.600 757.950 ;
        RECT 308.400 757.050 309.600 787.950 ;
        RECT 311.400 784.050 312.600 793.950 ;
        RECT 317.400 790.050 318.600 829.950 ;
        RECT 322.950 826.950 325.050 829.050 ;
        RECT 319.950 823.950 322.050 826.050 ;
        RECT 316.950 787.950 319.050 790.050 ;
        RECT 310.950 781.950 313.050 784.050 ;
        RECT 320.400 778.050 321.600 823.950 ;
        RECT 323.400 796.050 324.600 826.950 ;
        RECT 329.400 826.050 330.600 835.950 ;
        RECT 335.400 829.050 336.600 841.950 ;
        RECT 338.400 835.050 339.600 841.950 ;
        RECT 343.950 840.000 346.050 844.050 ;
        RECT 358.950 841.950 361.050 844.050 ;
        RECT 344.400 838.050 345.600 840.000 ;
        RECT 349.950 839.100 352.050 841.200 ;
        RECT 350.400 838.050 351.600 839.100 ;
        RECT 343.950 835.950 346.050 838.050 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 349.950 835.950 352.050 838.050 ;
        RECT 352.950 835.950 355.050 838.050 ;
        RECT 337.950 832.950 340.050 835.050 ;
        RECT 340.950 832.950 343.050 835.050 ;
        RECT 347.400 834.000 348.600 835.950 ;
        RECT 341.400 829.050 342.600 832.950 ;
        RECT 346.950 829.950 349.050 834.000 ;
        RECT 353.400 829.050 354.600 835.950 ;
        RECT 359.400 832.050 360.600 841.950 ;
        RECT 367.950 839.100 370.050 841.200 ;
        RECT 373.950 840.000 376.050 844.050 ;
        RECT 382.950 841.950 385.050 844.050 ;
        RECT 368.400 838.050 369.600 839.100 ;
        RECT 374.400 838.050 375.600 840.000 ;
        RECT 379.950 839.100 382.050 841.200 ;
        RECT 364.950 835.950 367.050 838.050 ;
        RECT 367.950 835.950 370.050 838.050 ;
        RECT 370.950 835.950 373.050 838.050 ;
        RECT 373.950 835.950 376.050 838.050 ;
        RECT 358.950 829.950 361.050 832.050 ;
        RECT 334.950 826.950 337.050 829.050 ;
        RECT 340.950 826.950 343.050 829.050 ;
        RECT 346.950 826.800 349.050 828.900 ;
        RECT 352.950 826.950 355.050 829.050 ;
        RECT 328.950 823.950 331.050 826.050 ;
        RECT 337.950 823.950 340.050 826.050 ;
        RECT 331.950 814.950 334.050 817.050 ;
        RECT 332.400 805.050 333.600 814.950 ;
        RECT 338.400 805.050 339.600 823.950 ;
        RECT 347.400 820.050 348.600 826.800 ;
        RECT 358.950 823.950 361.050 826.050 ;
        RECT 346.950 817.950 349.050 820.050 ;
        RECT 340.950 811.950 343.050 814.050 ;
        RECT 341.400 808.050 342.600 811.950 ;
        RECT 347.400 808.200 348.600 817.950 ;
        RECT 359.400 816.600 360.600 823.950 ;
        RECT 365.400 823.050 366.600 835.950 ;
        RECT 364.950 820.950 367.050 823.050 ;
        RECT 359.400 815.400 363.600 816.600 ;
        RECT 352.950 811.950 355.050 814.050 ;
        RECT 340.950 805.950 343.050 808.050 ;
        RECT 346.950 806.100 349.050 808.200 ;
        RECT 347.400 805.050 348.600 806.100 ;
        RECT 353.400 805.050 354.600 811.950 ;
        RECT 328.950 802.950 331.050 805.050 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 334.950 802.950 337.050 805.050 ;
        RECT 337.950 802.950 340.050 805.050 ;
        RECT 346.950 802.950 349.050 805.050 ;
        RECT 349.950 802.950 352.050 805.050 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 355.950 802.950 358.050 805.050 ;
        RECT 322.950 793.950 325.050 796.050 ;
        RECT 329.400 787.050 330.600 802.950 ;
        RECT 335.400 790.050 336.600 802.950 ;
        RECT 343.950 799.950 346.050 802.050 ;
        RECT 340.950 790.950 343.050 793.050 ;
        RECT 334.950 787.950 337.050 790.050 ;
        RECT 328.950 784.950 331.050 787.050 ;
        RECT 322.950 778.950 325.050 781.050 ;
        RECT 310.950 775.950 313.050 778.050 ;
        RECT 319.950 775.950 322.050 778.050 ;
        RECT 307.950 754.950 310.050 757.050 ;
        RECT 304.950 748.950 307.050 751.050 ;
        RECT 295.950 745.950 298.050 748.050 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 292.950 724.950 295.050 727.050 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 286.950 721.800 289.050 723.900 ;
        RECT 290.400 723.000 291.600 724.950 ;
        RECT 296.400 723.900 297.600 724.950 ;
        RECT 295.950 723.600 298.050 723.900 ;
        RECT 280.950 716.400 285.600 717.600 ;
        RECT 280.950 715.950 283.050 716.400 ;
        RECT 269.400 710.400 273.600 711.600 ;
        RECT 268.950 706.950 271.050 709.050 ;
        RECT 269.400 682.050 270.600 706.950 ;
        RECT 272.400 706.050 273.600 710.400 ;
        RECT 271.950 703.950 274.050 706.050 ;
        RECT 274.950 683.100 277.050 685.200 ;
        RECT 281.400 685.050 282.600 715.950 ;
        RECT 287.400 694.050 288.600 721.800 ;
        RECT 289.950 718.950 292.050 723.000 ;
        RECT 295.950 722.400 300.600 723.600 ;
        RECT 295.950 721.800 298.050 722.400 ;
        RECT 290.400 703.050 291.600 718.950 ;
        RECT 299.400 718.050 300.600 722.400 ;
        RECT 298.950 715.950 301.050 718.050 ;
        RECT 298.950 709.950 301.050 712.050 ;
        RECT 289.950 700.950 292.050 703.050 ;
        RECT 283.800 691.950 285.900 694.050 ;
        RECT 286.950 691.950 289.050 694.050 ;
        RECT 275.400 682.050 276.600 683.100 ;
        RECT 280.950 682.950 283.050 685.050 ;
        RECT 268.950 679.950 271.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 274.950 679.950 277.050 682.050 ;
        RECT 277.950 679.950 280.050 682.050 ;
        RECT 265.950 673.950 268.050 679.050 ;
        RECT 272.400 678.900 273.600 679.950 ;
        RECT 271.950 676.800 274.050 678.900 ;
        RECT 278.400 673.050 279.600 679.950 ;
        RECT 284.400 679.050 285.600 691.950 ;
        RECT 292.950 683.100 295.050 685.200 ;
        RECT 293.400 682.050 294.600 683.100 ;
        RECT 299.400 682.050 300.600 709.950 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 295.950 679.950 298.050 682.050 ;
        RECT 298.950 679.950 301.050 682.050 ;
        RECT 283.950 676.950 286.050 679.050 ;
        RECT 283.950 673.800 286.050 675.900 ;
        RECT 262.950 670.950 265.050 673.050 ;
        RECT 277.950 670.950 280.050 673.050 ;
        RECT 277.950 661.950 280.050 664.050 ;
        RECT 271.950 655.950 274.050 658.050 ;
        RECT 265.950 650.100 268.050 652.200 ;
        RECT 266.400 649.050 267.600 650.100 ;
        RECT 272.400 649.050 273.600 655.950 ;
        RECT 278.400 649.050 279.600 661.950 ;
        RECT 280.950 658.950 283.050 661.050 ;
        RECT 281.400 652.050 282.600 658.950 ;
        RECT 280.950 649.950 283.050 652.050 ;
        RECT 265.950 646.950 268.050 649.050 ;
        RECT 268.950 646.950 271.050 649.050 ;
        RECT 271.950 646.950 274.050 649.050 ;
        RECT 274.950 646.950 277.050 649.050 ;
        RECT 277.950 646.950 280.050 649.050 ;
        RECT 259.950 637.950 262.050 640.050 ;
        RECT 259.950 634.800 262.050 636.900 ;
        RECT 248.400 599.400 252.600 600.600 ;
        RECT 254.400 632.400 258.600 633.600 ;
        RECT 242.400 596.400 246.600 597.600 ;
        RECT 241.950 592.950 244.050 595.050 ;
        RECT 238.950 589.950 241.050 592.050 ;
        RECT 238.950 583.950 241.050 586.050 ;
        RECT 232.950 571.950 235.050 574.050 ;
        RECT 239.400 571.050 240.600 583.950 ;
        RECT 242.400 577.050 243.600 592.950 ;
        RECT 245.400 586.050 246.600 596.400 ;
        RECT 244.950 583.950 247.050 586.050 ;
        RECT 244.950 577.950 247.050 580.050 ;
        RECT 241.950 574.950 244.050 577.050 ;
        RECT 245.400 574.050 246.600 577.950 ;
        RECT 244.950 571.950 247.050 574.050 ;
        RECT 235.950 568.950 238.050 571.050 ;
        RECT 238.950 568.950 241.050 571.050 ;
        RECT 241.950 568.950 244.050 571.050 ;
        RECT 232.950 565.950 235.050 568.050 ;
        RECT 236.400 567.900 237.600 568.950 ;
        RECT 229.950 559.950 232.050 562.050 ;
        RECT 229.950 550.950 232.050 553.050 ;
        RECT 221.400 527.400 225.600 528.600 ;
        RECT 209.400 526.050 210.600 527.100 ;
        RECT 215.400 526.050 216.600 527.100 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 187.950 523.950 190.050 526.050 ;
        RECT 190.950 523.950 193.050 526.050 ;
        RECT 193.950 523.950 196.050 526.050 ;
        RECT 205.950 523.950 208.050 526.050 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 211.950 523.950 214.050 526.050 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 185.400 507.600 186.600 523.950 ;
        RECT 191.400 517.050 192.600 523.950 ;
        RECT 190.950 514.950 193.050 517.050 ;
        RECT 206.400 513.600 207.600 523.950 ;
        RECT 212.400 517.050 213.600 523.950 ;
        RECT 217.950 520.950 220.050 523.050 ;
        RECT 218.400 517.050 219.600 520.950 ;
        RECT 211.950 514.950 214.050 517.050 ;
        RECT 217.950 514.950 220.050 517.050 ;
        RECT 206.400 512.400 210.600 513.600 ;
        RECT 205.950 508.950 208.050 511.050 ;
        RECT 185.400 506.400 189.600 507.600 ;
        RECT 184.950 502.950 187.050 505.050 ;
        RECT 175.950 493.950 178.050 496.050 ;
        RECT 145.950 490.950 148.050 493.050 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 157.950 490.950 160.050 493.050 ;
        RECT 169.950 490.950 172.050 493.050 ;
        RECT 172.950 490.950 175.050 493.050 ;
        RECT 178.950 490.950 181.050 493.050 ;
        RECT 146.400 489.900 147.600 490.950 ;
        RECT 145.950 487.800 148.050 489.900 ;
        RECT 124.950 478.950 127.050 481.050 ;
        RECT 136.950 478.950 139.050 481.050 ;
        RECT 115.950 472.950 118.050 475.050 ;
        RECT 118.950 460.950 121.050 463.050 ;
        RECT 112.950 457.950 115.050 460.050 ;
        RECT 100.950 448.950 103.050 451.050 ;
        RECT 106.950 450.000 109.050 454.050 ;
        RECT 101.400 439.050 102.600 448.950 ;
        RECT 107.400 448.050 108.600 450.000 ;
        RECT 113.400 448.050 114.600 457.950 ;
        RECT 119.400 451.050 120.600 460.950 ;
        RECT 118.800 448.950 120.900 451.050 ;
        RECT 121.950 449.100 124.050 451.200 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 100.950 436.950 103.050 439.050 ;
        RECT 110.400 427.050 111.600 445.950 ;
        RECT 116.400 445.050 117.600 445.950 ;
        RECT 116.400 443.400 121.050 445.050 ;
        RECT 117.000 442.950 121.050 443.400 ;
        RECT 122.400 442.050 123.600 449.100 ;
        RECT 121.950 439.950 124.050 442.050 ;
        RECT 121.950 430.950 124.050 433.050 ;
        RECT 109.950 424.950 112.050 427.050 ;
        RECT 100.950 415.950 103.050 418.050 ;
        RECT 109.950 416.100 112.050 418.200 ;
        RECT 115.950 417.000 118.050 421.050 ;
        RECT 101.400 400.050 102.600 415.950 ;
        RECT 110.400 415.050 111.600 416.100 ;
        RECT 116.400 415.050 117.600 417.000 ;
        RECT 106.950 412.950 109.050 415.050 ;
        RECT 109.950 412.950 112.050 415.050 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 115.950 412.950 118.050 415.050 ;
        RECT 100.950 397.950 103.050 400.050 ;
        RECT 97.950 391.950 100.050 394.050 ;
        RECT 107.400 388.050 108.600 412.950 ;
        RECT 113.400 411.900 114.600 412.950 ;
        RECT 112.950 409.800 115.050 411.900 ;
        RECT 122.400 394.050 123.600 430.950 ;
        RECT 125.400 418.050 126.600 478.950 ;
        RECT 152.400 469.050 153.600 490.950 ;
        RECT 158.400 484.050 159.600 490.950 ;
        RECT 170.400 489.900 171.600 490.950 ;
        RECT 169.950 487.800 172.050 489.900 ;
        RECT 179.400 489.000 180.600 490.950 ;
        RECT 157.950 481.950 160.050 484.050 ;
        RECT 178.950 481.950 181.050 489.000 ;
        RECT 181.950 487.950 184.050 490.050 ;
        RECT 185.400 489.600 186.600 502.950 ;
        RECT 188.400 502.050 189.600 506.400 ;
        RECT 187.950 499.950 190.050 502.050 ;
        RECT 193.950 494.100 196.050 496.200 ;
        RECT 194.400 493.050 195.600 494.100 ;
        RECT 202.950 493.950 205.050 496.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 191.400 489.600 192.600 490.950 ;
        RECT 197.400 489.900 198.600 490.950 ;
        RECT 185.400 488.400 192.600 489.600 ;
        RECT 142.950 466.950 145.050 469.050 ;
        RECT 151.950 466.950 154.050 469.050 ;
        RECT 136.950 454.950 139.050 457.050 ;
        RECT 130.950 449.100 133.050 451.200 ;
        RECT 131.400 448.050 132.600 449.100 ;
        RECT 137.400 448.050 138.600 454.950 ;
        RECT 143.400 451.050 144.600 466.950 ;
        RECT 151.950 460.950 154.050 463.050 ;
        RECT 142.950 448.950 145.050 451.050 ;
        RECT 152.400 448.050 153.600 460.950 ;
        RECT 163.950 451.950 166.050 454.050 ;
        RECT 159.000 450.600 163.050 451.050 ;
        RECT 158.400 448.950 163.050 450.600 ;
        RECT 158.400 448.050 159.600 448.950 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 133.950 445.950 136.050 448.050 ;
        RECT 136.950 445.950 139.050 448.050 ;
        RECT 139.950 445.950 142.050 448.050 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 151.950 445.950 154.050 448.050 ;
        RECT 154.950 445.950 157.050 448.050 ;
        RECT 157.950 445.950 160.050 448.050 ;
        RECT 127.950 439.950 130.050 445.050 ;
        RECT 134.400 433.050 135.600 445.950 ;
        RECT 140.400 444.900 141.600 445.950 ;
        RECT 139.950 439.950 142.050 444.900 ;
        RECT 149.400 444.600 150.600 445.950 ;
        RECT 155.400 444.900 156.600 445.950 ;
        RECT 164.400 445.050 165.600 451.950 ;
        RECT 169.950 449.100 172.050 451.200 ;
        RECT 175.950 449.100 178.050 451.200 ;
        RECT 182.400 450.600 183.600 487.950 ;
        RECT 190.950 484.950 196.050 487.050 ;
        RECT 196.950 484.950 199.050 489.900 ;
        RECT 187.950 478.950 190.050 481.050 ;
        RECT 182.400 449.400 186.600 450.600 ;
        RECT 170.400 448.050 171.600 449.100 ;
        RECT 176.400 448.050 177.600 449.100 ;
        RECT 169.950 445.950 172.050 448.050 ;
        RECT 172.950 445.950 175.050 448.050 ;
        RECT 175.950 445.950 178.050 448.050 ;
        RECT 178.950 445.950 181.050 448.050 ;
        RECT 146.400 443.400 150.600 444.600 ;
        RECT 133.950 430.950 136.050 433.050 ;
        RECT 124.950 415.950 127.050 418.050 ;
        RECT 127.950 417.000 130.050 421.050 ;
        RECT 128.400 415.050 129.600 417.000 ;
        RECT 134.400 415.050 135.600 430.950 ;
        RECT 146.400 424.050 147.600 443.400 ;
        RECT 154.950 442.800 157.050 444.900 ;
        RECT 160.950 442.950 163.050 445.050 ;
        RECT 163.950 442.950 166.050 445.050 ;
        RECT 161.400 439.050 162.600 442.950 ;
        RECT 163.950 439.800 166.050 441.900 ;
        RECT 160.950 436.950 163.050 439.050 ;
        RECT 157.950 424.950 160.050 427.050 ;
        RECT 145.950 421.950 148.050 424.050 ;
        RECT 146.400 418.050 147.600 421.950 ;
        RECT 142.950 415.950 145.050 418.050 ;
        RECT 145.950 415.950 148.050 418.050 ;
        RECT 148.950 416.100 151.050 418.200 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 133.950 412.950 136.050 415.050 ;
        RECT 136.950 412.950 139.050 415.050 ;
        RECT 124.950 409.950 127.050 412.050 ;
        RECT 131.400 411.000 132.600 412.950 ;
        RECT 109.950 391.950 112.050 394.050 ;
        RECT 121.950 391.950 124.050 394.050 ;
        RECT 106.950 385.950 109.050 388.050 ;
        RECT 70.950 382.950 73.050 385.050 ;
        RECT 94.950 382.950 97.050 385.050 ;
        RECT 58.950 376.950 61.050 379.050 ;
        RECT 52.950 371.100 55.050 373.200 ;
        RECT 53.400 370.050 54.600 371.100 ;
        RECT 59.400 370.050 60.600 376.950 ;
        RECT 67.950 370.950 70.050 373.050 ;
        RECT 52.950 367.950 55.050 370.050 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 58.950 367.950 61.050 370.050 ;
        RECT 61.950 367.950 64.050 370.050 ;
        RECT 56.400 363.600 57.600 367.950 ;
        RECT 62.400 366.000 63.600 367.950 ;
        RECT 53.400 362.400 57.600 363.600 ;
        RECT 53.400 352.050 54.600 362.400 ;
        RECT 61.950 361.950 64.050 366.000 ;
        RECT 52.950 349.950 55.050 352.050 ;
        RECT 58.950 349.950 61.050 352.050 ;
        RECT 55.950 343.950 58.050 346.050 ;
        RECT 46.950 340.950 49.050 343.050 ;
        RECT 52.950 340.950 55.050 343.050 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 46.950 334.950 49.050 337.050 ;
        RECT 29.400 332.400 33.600 333.600 ;
        RECT 19.950 316.950 22.050 319.050 ;
        RECT 13.950 301.950 16.050 304.050 ;
        RECT 16.950 293.100 19.050 295.200 ;
        RECT 26.400 295.050 27.600 331.950 ;
        RECT 32.400 322.050 33.600 332.400 ;
        RECT 34.950 331.800 37.050 333.900 ;
        RECT 35.400 328.050 36.600 331.800 ;
        RECT 34.950 325.950 37.050 328.050 ;
        RECT 31.950 319.950 34.050 322.050 ;
        RECT 41.400 319.050 42.600 334.950 ;
        RECT 47.400 333.900 48.600 334.950 ;
        RECT 46.950 331.800 49.050 333.900 ;
        RECT 43.950 328.950 46.050 331.050 ;
        RECT 28.950 316.950 31.050 319.050 ;
        RECT 40.950 316.950 43.050 319.050 ;
        RECT 25.950 294.600 28.050 295.050 ;
        RECT 23.400 293.400 28.050 294.600 ;
        RECT 17.400 292.050 18.600 293.100 ;
        RECT 23.400 292.050 24.600 293.400 ;
        RECT 25.950 292.950 28.050 293.400 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 22.950 289.950 25.050 292.050 ;
        RECT 14.400 280.050 15.600 289.950 ;
        RECT 16.950 283.950 19.050 286.050 ;
        RECT 13.950 277.950 16.050 280.050 ;
        RECT 17.400 277.050 18.600 283.950 ;
        RECT 20.400 280.050 21.600 289.950 ;
        RECT 25.950 286.950 28.050 289.050 ;
        RECT 19.950 277.950 22.050 280.050 ;
        RECT 16.950 274.950 19.050 277.050 ;
        RECT 7.950 268.950 10.050 271.050 ;
        RECT 7.950 259.950 10.050 262.050 ;
        RECT 16.950 260.100 19.050 262.200 ;
        RECT 22.950 260.100 25.050 262.200 ;
        RECT 26.400 262.050 27.600 286.950 ;
        RECT 29.400 286.050 30.600 316.950 ;
        RECT 44.400 310.050 45.600 328.950 ;
        RECT 49.950 325.950 52.050 328.050 ;
        RECT 43.950 307.950 46.050 310.050 ;
        RECT 43.950 301.950 46.050 304.050 ;
        RECT 44.400 295.200 45.600 301.950 ;
        RECT 37.950 293.100 40.050 295.200 ;
        RECT 43.950 293.100 46.050 295.200 ;
        RECT 38.400 292.050 39.600 293.100 ;
        RECT 44.400 292.050 45.600 293.100 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 43.950 289.950 46.050 292.050 ;
        RECT 31.950 286.950 34.050 289.050 ;
        RECT 28.950 283.950 31.050 286.050 ;
        RECT 4.950 178.950 7.050 181.050 ;
        RECT 4.950 151.950 7.050 154.050 ;
        RECT 5.400 109.050 6.600 151.950 ;
        RECT 8.400 151.050 9.600 259.950 ;
        RECT 17.400 259.050 18.600 260.100 ;
        RECT 23.400 259.050 24.600 260.100 ;
        RECT 25.950 259.950 28.050 262.050 ;
        RECT 13.950 256.950 16.050 259.050 ;
        RECT 16.950 256.950 19.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 22.950 256.950 25.050 259.050 ;
        RECT 14.400 238.050 15.600 256.950 ;
        RECT 20.400 255.900 21.600 256.950 ;
        RECT 29.400 255.900 30.600 283.950 ;
        RECT 32.400 262.050 33.600 286.950 ;
        RECT 35.400 271.050 36.600 289.950 ;
        RECT 41.400 277.050 42.600 289.950 ;
        RECT 46.950 286.950 49.050 289.050 ;
        RECT 40.950 274.950 43.050 277.050 ;
        RECT 34.950 268.950 37.050 271.050 ;
        RECT 37.950 265.950 40.050 268.050 ;
        RECT 31.950 259.950 34.050 262.050 ;
        RECT 38.400 259.050 39.600 265.950 ;
        RECT 47.400 265.050 48.600 286.950 ;
        RECT 50.400 280.050 51.600 325.950 ;
        RECT 53.400 295.050 54.600 340.950 ;
        RECT 56.400 333.900 57.600 343.950 ;
        RECT 59.400 340.050 60.600 349.950 ;
        RECT 68.400 343.050 69.600 370.950 ;
        RECT 71.400 366.600 72.600 382.950 ;
        RECT 106.950 382.800 109.050 384.900 ;
        RECT 76.950 371.100 79.050 373.200 ;
        RECT 94.950 371.100 97.050 373.200 ;
        RECT 100.950 371.100 103.050 373.200 ;
        RECT 77.400 370.050 78.600 371.100 ;
        RECT 95.400 370.050 96.600 371.100 ;
        RECT 101.400 370.050 102.600 371.100 ;
        RECT 76.950 367.950 79.050 370.050 ;
        RECT 79.950 367.950 82.050 370.050 ;
        RECT 85.950 367.950 88.050 370.050 ;
        RECT 91.950 367.950 94.050 370.050 ;
        RECT 94.950 367.950 97.050 370.050 ;
        RECT 97.950 367.950 100.050 370.050 ;
        RECT 100.950 367.950 103.050 370.050 ;
        RECT 71.400 365.400 75.600 366.600 ;
        RECT 70.950 355.950 73.050 358.050 ;
        RECT 67.950 340.950 70.050 343.050 ;
        RECT 58.950 337.950 61.050 340.050 ;
        RECT 64.950 338.100 67.050 340.200 ;
        RECT 65.400 337.050 66.600 338.100 ;
        RECT 71.400 337.050 72.600 355.950 ;
        RECT 74.400 340.050 75.600 365.400 ;
        RECT 80.400 358.050 81.600 367.950 ;
        RECT 79.950 355.950 82.050 358.050 ;
        RECT 86.400 352.050 87.600 367.950 ;
        RECT 92.400 358.050 93.600 367.950 ;
        RECT 98.400 364.050 99.600 367.950 ;
        RECT 103.950 364.950 106.050 367.050 ;
        RECT 98.400 362.400 103.050 364.050 ;
        RECT 99.000 361.950 103.050 362.400 ;
        RECT 91.950 355.950 94.050 358.050 ;
        RECT 85.950 349.950 88.050 352.050 ;
        RECT 76.950 340.950 79.050 343.050 ;
        RECT 73.950 337.950 76.050 340.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 64.950 334.950 67.050 337.050 ;
        RECT 67.950 334.950 70.050 337.050 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 62.400 333.900 63.600 334.950 ;
        RECT 55.950 331.800 58.050 333.900 ;
        RECT 61.950 331.800 64.050 333.900 ;
        RECT 64.950 328.950 67.050 331.050 ;
        RECT 52.950 292.950 55.050 295.050 ;
        RECT 58.950 294.000 61.050 298.050 ;
        RECT 65.400 295.200 66.600 328.950 ;
        RECT 68.400 325.050 69.600 334.950 ;
        RECT 77.400 333.900 78.600 340.950 ;
        RECT 86.400 337.050 87.600 349.950 ;
        RECT 100.950 340.950 103.050 343.050 ;
        RECT 91.950 338.100 94.050 340.200 ;
        RECT 92.400 337.050 93.600 338.100 ;
        RECT 97.950 337.950 100.050 340.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 88.950 334.950 91.050 337.050 ;
        RECT 91.950 334.950 94.050 337.050 ;
        RECT 76.950 331.800 79.050 333.900 ;
        RECT 79.950 331.950 82.050 334.050 ;
        RECT 83.400 333.900 84.600 334.950 ;
        RECT 67.950 322.950 70.050 325.050 ;
        RECT 80.400 304.050 81.600 331.950 ;
        RECT 82.950 331.800 85.050 333.900 ;
        RECT 89.400 328.050 90.600 334.950 ;
        RECT 88.950 325.950 91.050 328.050 ;
        RECT 89.400 319.050 90.600 325.950 ;
        RECT 88.950 316.950 91.050 319.050 ;
        RECT 88.950 307.950 91.050 310.050 ;
        RECT 79.950 301.950 82.050 304.050 ;
        RECT 59.400 292.050 60.600 294.000 ;
        RECT 64.950 293.100 67.050 295.200 ;
        RECT 73.950 294.000 76.050 298.050 ;
        RECT 65.400 292.050 66.600 293.100 ;
        RECT 74.400 292.050 75.600 294.000 ;
        RECT 79.950 293.100 82.050 295.200 ;
        RECT 80.400 292.050 81.600 293.100 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 61.950 289.950 64.050 292.050 ;
        RECT 64.950 289.950 67.050 292.050 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 52.950 286.950 55.050 289.050 ;
        RECT 56.400 288.000 57.600 289.950 ;
        RECT 62.400 288.900 63.600 289.950 ;
        RECT 77.400 288.900 78.600 289.950 ;
        RECT 49.950 277.950 52.050 280.050 ;
        RECT 46.950 262.950 49.050 265.050 ;
        RECT 43.950 260.100 46.050 262.200 ;
        RECT 44.400 259.050 45.600 260.100 ;
        RECT 49.950 259.950 52.050 262.050 ;
        RECT 34.950 256.950 37.050 259.050 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 35.400 256.050 36.600 256.950 ;
        RECT 19.950 253.800 22.050 255.900 ;
        RECT 28.950 253.800 31.050 255.900 ;
        RECT 31.950 254.400 36.600 256.050 ;
        RECT 41.400 255.900 42.600 256.950 ;
        RECT 31.950 253.950 36.000 254.400 ;
        RECT 40.950 253.800 43.050 255.900 ;
        RECT 13.950 235.950 16.050 238.050 ;
        RECT 50.400 235.050 51.600 259.950 ;
        RECT 22.950 232.950 25.050 235.050 ;
        RECT 49.950 232.950 52.050 235.050 ;
        RECT 16.950 226.950 19.050 229.050 ;
        RECT 17.400 214.050 18.600 226.950 ;
        RECT 23.400 214.050 24.600 232.950 ;
        RECT 31.950 226.950 34.050 229.050 ;
        RECT 32.400 214.050 33.600 226.950 ;
        RECT 37.950 223.950 40.050 226.050 ;
        RECT 46.950 223.950 49.050 226.050 ;
        RECT 38.400 214.050 39.600 223.950 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 19.950 211.950 22.050 214.050 ;
        RECT 22.950 211.950 25.050 214.050 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 14.400 187.050 15.600 211.950 ;
        RECT 20.400 205.050 21.600 211.950 ;
        RECT 35.400 210.900 36.600 211.950 ;
        RECT 34.950 208.800 37.050 210.900 ;
        RECT 19.950 202.950 22.050 205.050 ;
        RECT 16.950 196.950 19.050 199.050 ;
        RECT 13.950 184.950 16.050 187.050 ;
        RECT 17.400 181.050 18.600 196.950 ;
        RECT 41.400 190.050 42.600 211.950 ;
        RECT 47.400 205.050 48.600 223.950 ;
        RECT 50.400 210.900 51.600 232.950 ;
        RECT 49.950 208.800 52.050 210.900 ;
        RECT 46.950 202.950 49.050 205.050 ;
        RECT 46.950 199.800 49.050 201.900 ;
        RECT 28.950 187.950 31.050 190.050 ;
        RECT 40.950 187.950 43.050 190.050 ;
        RECT 22.950 182.100 25.050 184.200 ;
        RECT 23.400 181.050 24.600 182.100 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 22.950 178.950 25.050 181.050 ;
        RECT 10.950 175.950 13.050 178.050 ;
        RECT 14.400 177.900 15.600 178.950 ;
        RECT 20.400 177.900 21.600 178.950 ;
        RECT 29.400 177.900 30.600 187.950 ;
        RECT 37.950 182.100 40.050 184.200 ;
        RECT 38.400 181.050 39.600 182.100 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 35.400 177.900 36.600 178.950 ;
        RECT 7.950 148.950 10.050 151.050 ;
        RECT 11.400 142.050 12.600 175.950 ;
        RECT 13.950 175.800 16.050 177.900 ;
        RECT 19.950 175.800 22.050 177.900 ;
        RECT 28.950 175.800 31.050 177.900 ;
        RECT 34.950 175.800 37.050 177.900 ;
        RECT 41.400 177.600 42.600 178.950 ;
        RECT 47.400 177.600 48.600 199.800 ;
        RECT 53.400 199.050 54.600 286.950 ;
        RECT 55.950 283.950 58.050 288.000 ;
        RECT 61.950 286.800 64.050 288.900 ;
        RECT 76.950 286.800 79.050 288.900 ;
        RECT 83.400 283.050 84.600 289.950 ;
        RECT 89.400 288.900 90.600 307.950 ;
        RECT 91.950 301.950 94.050 304.050 ;
        RECT 88.950 286.800 91.050 288.900 ;
        RECT 82.950 280.950 85.050 283.050 ;
        RECT 64.950 274.950 67.050 277.050 ;
        RECT 55.950 261.600 60.000 262.050 ;
        RECT 55.950 259.950 60.600 261.600 ;
        RECT 59.400 259.050 60.600 259.950 ;
        RECT 65.400 259.050 66.600 274.950 ;
        RECT 83.400 265.050 84.600 280.950 ;
        RECT 73.950 262.950 76.050 265.050 ;
        RECT 82.950 262.950 85.050 265.050 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 67.950 256.950 70.050 259.050 ;
        RECT 55.950 253.950 58.050 256.050 ;
        RECT 62.400 255.900 63.600 256.950 ;
        RECT 68.400 255.900 69.600 256.950 ;
        RECT 74.400 255.900 75.600 262.950 ;
        RECT 85.950 260.100 88.050 262.200 ;
        RECT 86.400 259.050 87.600 260.100 ;
        RECT 82.950 256.950 85.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 56.400 247.050 57.600 253.950 ;
        RECT 61.950 253.800 64.050 255.900 ;
        RECT 67.950 253.800 70.050 255.900 ;
        RECT 73.950 253.800 76.050 255.900 ;
        RECT 55.950 244.950 58.050 247.050 ;
        RECT 58.950 238.950 61.050 241.050 ;
        RECT 59.400 214.050 60.600 238.950 ;
        RECT 62.400 238.050 63.600 253.800 ;
        RECT 64.950 250.950 67.050 253.050 ;
        RECT 61.950 235.950 64.050 238.050 ;
        RECT 65.400 229.050 66.600 250.950 ;
        RECT 70.950 232.950 73.050 235.050 ;
        RECT 64.950 226.950 67.050 229.050 ;
        RECT 64.950 215.100 67.050 217.200 ;
        RECT 65.400 214.050 66.600 215.100 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 52.950 196.950 55.050 199.050 ;
        RECT 62.400 184.200 63.600 211.950 ;
        RECT 71.400 202.050 72.600 232.950 ;
        RECT 83.400 220.050 84.600 256.950 ;
        RECT 88.950 253.950 91.050 256.050 ;
        RECT 89.400 241.050 90.600 253.950 ;
        RECT 88.950 238.950 91.050 241.050 ;
        RECT 82.950 217.950 85.050 220.050 ;
        RECT 76.950 215.100 79.050 217.200 ;
        RECT 77.400 214.050 78.600 215.100 ;
        RECT 83.400 214.050 84.600 217.950 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 79.950 211.950 82.050 214.050 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 70.950 199.950 73.050 202.050 ;
        RECT 73.950 193.950 76.050 196.050 ;
        RECT 49.950 181.950 52.050 184.050 ;
        RECT 55.950 182.100 58.050 184.200 ;
        RECT 61.950 182.100 64.050 184.200 ;
        RECT 41.400 176.400 48.600 177.600 ;
        RECT 14.400 160.050 15.600 175.800 ;
        RECT 13.950 157.950 16.050 160.050 ;
        RECT 22.950 148.950 25.050 151.050 ;
        RECT 10.950 141.600 13.050 142.050 ;
        RECT 8.400 140.400 13.050 141.600 ;
        RECT 8.400 130.050 9.600 140.400 ;
        RECT 10.950 139.950 13.050 140.400 ;
        RECT 16.950 138.000 19.050 142.050 ;
        RECT 17.400 136.050 18.600 138.000 ;
        RECT 23.400 136.050 24.600 148.950 ;
        RECT 29.400 139.050 30.600 175.800 ;
        RECT 46.950 148.950 49.050 151.050 ;
        RECT 28.950 136.950 31.050 139.050 ;
        RECT 31.950 138.000 34.050 142.050 ;
        RECT 37.950 139.950 40.050 145.050 ;
        RECT 32.400 136.050 33.600 138.000 ;
        RECT 38.400 136.050 39.600 139.950 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 22.950 133.950 25.050 136.050 ;
        RECT 31.950 133.950 34.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 7.950 127.950 10.050 130.050 ;
        RECT 7.950 112.950 10.050 115.050 ;
        RECT 4.950 106.950 7.050 109.050 ;
        RECT 5.400 94.050 6.600 106.950 ;
        RECT 8.400 99.900 9.600 112.950 ;
        RECT 14.400 109.050 15.600 133.950 ;
        RECT 20.400 132.000 21.600 133.950 ;
        RECT 19.950 127.950 22.050 132.000 ;
        RECT 25.950 130.950 28.050 133.050 ;
        RECT 35.400 132.900 36.600 133.950 ;
        RECT 16.950 109.950 19.050 112.050 ;
        RECT 13.950 106.950 16.050 109.050 ;
        RECT 17.400 103.050 18.600 109.950 ;
        RECT 26.400 106.200 27.600 130.950 ;
        RECT 34.950 130.800 37.050 132.900 ;
        RECT 41.400 118.050 42.600 133.950 ;
        RECT 47.400 132.900 48.600 148.950 ;
        RECT 46.950 130.800 49.050 132.900 ;
        RECT 40.950 115.950 43.050 118.050 ;
        RECT 28.950 109.950 31.050 112.050 ;
        RECT 25.950 105.600 28.050 106.200 ;
        RECT 23.400 104.400 28.050 105.600 ;
        RECT 23.400 103.050 24.600 104.400 ;
        RECT 25.950 104.100 28.050 104.400 ;
        RECT 13.950 100.950 16.050 103.050 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 19.950 100.950 22.050 103.050 ;
        RECT 22.950 100.950 25.050 103.050 ;
        RECT 14.400 99.900 15.600 100.950 ;
        RECT 7.950 97.800 10.050 99.900 ;
        RECT 13.950 97.800 16.050 99.900 ;
        RECT 20.400 94.050 21.600 100.950 ;
        RECT 4.950 91.950 7.050 94.050 ;
        RECT 19.950 91.950 22.050 94.050 ;
        RECT 16.950 70.950 19.050 73.050 ;
        RECT 17.400 58.050 18.600 70.950 ;
        RECT 22.950 60.000 25.050 64.050 ;
        RECT 29.400 61.050 30.600 109.950 ;
        RECT 41.400 108.600 42.600 115.950 ;
        RECT 41.400 107.400 45.600 108.600 ;
        RECT 32.400 104.400 39.600 105.600 ;
        RECT 32.400 64.050 33.600 104.400 ;
        RECT 38.400 103.050 39.600 104.400 ;
        RECT 44.400 103.050 45.600 107.400 ;
        RECT 50.400 105.600 51.600 181.950 ;
        RECT 56.400 181.050 57.600 182.100 ;
        RECT 62.400 181.050 63.600 182.100 ;
        RECT 74.400 181.050 75.600 193.950 ;
        RECT 80.400 193.050 81.600 211.950 ;
        RECT 92.400 211.050 93.600 301.950 ;
        RECT 94.950 295.050 97.050 298.050 ;
        RECT 98.400 295.200 99.600 337.950 ;
        RECT 101.400 298.050 102.600 340.950 ;
        RECT 104.400 340.050 105.600 364.950 ;
        RECT 107.400 364.050 108.600 382.800 ;
        RECT 106.950 361.950 109.050 364.050 ;
        RECT 106.950 355.950 109.050 358.050 ;
        RECT 103.950 337.950 106.050 340.050 ;
        RECT 107.400 337.050 108.600 355.950 ;
        RECT 110.400 355.050 111.600 391.950 ;
        RECT 125.400 385.050 126.600 409.950 ;
        RECT 130.950 406.950 133.050 411.000 ;
        RECT 137.400 406.050 138.600 412.950 ;
        RECT 143.400 409.050 144.600 415.950 ;
        RECT 149.400 415.050 150.600 416.100 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 142.950 406.950 145.050 409.050 ;
        RECT 145.950 406.950 148.050 412.050 ;
        RECT 152.400 411.900 153.600 412.950 ;
        RECT 151.950 409.800 154.050 411.900 ;
        RECT 136.950 403.950 139.050 406.050 ;
        RECT 137.400 403.050 138.600 403.950 ;
        RECT 137.400 401.400 142.050 403.050 ;
        RECT 138.000 400.950 142.050 401.400 ;
        RECT 145.950 400.950 151.050 403.050 ;
        RECT 130.950 388.950 133.050 391.050 ;
        RECT 124.950 382.950 127.050 385.050 ;
        RECT 112.950 376.950 115.050 379.050 ;
        RECT 121.950 376.950 124.050 379.050 ;
        RECT 113.400 361.050 114.600 376.950 ;
        RECT 122.400 370.050 123.600 376.950 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 124.950 367.950 127.050 370.050 ;
        RECT 112.950 358.950 115.050 361.050 ;
        RECT 119.400 355.050 120.600 367.950 ;
        RECT 109.950 352.950 112.050 355.050 ;
        RECT 118.950 352.950 121.050 355.050 ;
        RECT 125.400 346.050 126.600 367.950 ;
        RECT 127.950 358.950 130.050 361.050 ;
        RECT 124.950 343.950 127.050 346.050 ;
        RECT 112.950 339.000 115.050 343.050 ;
        RECT 124.950 340.800 127.050 342.900 ;
        RECT 113.400 337.050 114.600 339.000 ;
        RECT 106.950 334.950 109.050 337.050 ;
        RECT 109.950 334.950 112.050 337.050 ;
        RECT 112.950 334.950 115.050 337.050 ;
        RECT 115.950 334.950 118.050 337.050 ;
        RECT 103.950 331.950 106.050 334.050 ;
        RECT 104.400 328.050 105.600 331.950 ;
        RECT 110.400 328.050 111.600 334.950 ;
        RECT 116.400 333.900 117.600 334.950 ;
        RECT 125.400 334.050 126.600 340.800 ;
        RECT 115.950 331.800 118.050 333.900 ;
        RECT 124.950 331.950 127.050 334.050 ;
        RECT 103.950 325.950 106.050 328.050 ;
        RECT 109.950 325.950 112.050 328.050 ;
        RECT 116.400 322.050 117.600 331.800 ;
        RECT 128.400 328.050 129.600 358.950 ;
        RECT 131.400 343.050 132.600 388.950 ;
        RECT 145.950 382.950 148.050 385.050 ;
        RECT 133.950 379.950 136.050 382.050 ;
        RECT 134.400 361.050 135.600 379.950 ;
        RECT 139.950 376.950 142.050 379.050 ;
        RECT 140.400 370.050 141.600 376.950 ;
        RECT 146.400 370.050 147.600 382.950 ;
        RECT 154.950 379.950 157.050 382.050 ;
        RECT 151.950 371.100 154.050 373.200 ;
        RECT 155.400 373.050 156.600 379.950 ;
        RECT 158.400 373.200 159.600 424.950 ;
        RECT 161.400 403.050 162.600 436.950 ;
        RECT 164.400 418.050 165.600 439.800 ;
        RECT 173.400 433.050 174.600 445.950 ;
        RECT 179.400 444.900 180.600 445.950 ;
        RECT 178.950 442.800 181.050 444.900 ;
        RECT 185.400 435.600 186.600 449.400 ;
        RECT 182.400 434.400 186.600 435.600 ;
        RECT 169.950 430.950 172.050 433.050 ;
        RECT 172.950 430.950 175.050 433.050 ;
        RECT 163.950 415.950 166.050 418.050 ;
        RECT 170.400 415.050 171.600 430.950 ;
        RECT 175.950 417.000 178.050 421.050 ;
        RECT 176.400 415.050 177.600 417.000 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 172.950 412.950 175.050 415.050 ;
        RECT 175.950 412.950 178.050 415.050 ;
        RECT 167.400 411.900 168.600 412.950 ;
        RECT 166.950 409.800 169.050 411.900 ;
        RECT 160.950 400.950 163.050 403.050 ;
        RECT 167.400 382.050 168.600 409.800 ;
        RECT 173.400 403.050 174.600 412.950 ;
        RECT 172.950 400.950 175.050 403.050 ;
        RECT 166.950 379.950 169.050 382.050 ;
        RECT 163.950 376.950 166.050 379.050 ;
        RECT 169.950 376.950 172.050 379.050 ;
        RECT 175.950 376.950 178.050 382.050 ;
        RECT 139.950 367.950 142.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 145.950 367.950 148.050 370.050 ;
        RECT 133.950 358.950 136.050 361.050 ;
        RECT 143.400 352.050 144.600 367.950 ;
        RECT 152.400 364.050 153.600 371.100 ;
        RECT 154.950 370.950 157.050 373.050 ;
        RECT 157.950 371.100 160.050 373.200 ;
        RECT 158.400 370.050 159.600 371.100 ;
        RECT 164.400 370.050 165.600 376.950 ;
        RECT 157.950 367.950 160.050 370.050 ;
        RECT 160.950 367.950 163.050 370.050 ;
        RECT 163.950 367.950 166.050 370.050 ;
        RECT 154.950 364.950 157.050 367.050 ;
        RECT 145.950 361.950 148.050 364.050 ;
        RECT 151.950 361.950 154.050 364.050 ;
        RECT 136.950 349.950 139.050 352.050 ;
        RECT 142.950 349.950 145.050 352.050 ;
        RECT 130.950 340.950 133.050 343.050 ;
        RECT 137.400 337.050 138.600 349.950 ;
        RECT 142.950 346.800 145.050 348.900 ;
        RECT 133.950 334.950 136.050 337.050 ;
        RECT 136.950 334.950 139.050 337.050 ;
        RECT 130.950 331.950 133.050 334.050 ;
        RECT 134.400 333.900 135.600 334.950 ;
        RECT 127.950 325.950 130.050 328.050 ;
        RECT 115.950 319.950 118.050 322.050 ;
        RECT 103.950 301.950 106.050 304.050 ;
        RECT 115.950 303.600 120.000 304.050 ;
        RECT 115.950 303.000 120.600 303.600 ;
        RECT 115.950 301.950 121.050 303.000 ;
        RECT 100.950 295.950 103.050 298.050 ;
        RECT 94.800 294.000 97.050 295.050 ;
        RECT 94.800 292.950 96.900 294.000 ;
        RECT 97.950 293.100 100.050 295.200 ;
        RECT 98.400 292.050 99.600 293.100 ;
        RECT 104.400 292.050 105.600 301.950 ;
        RECT 118.950 298.950 121.050 301.950 ;
        RECT 131.400 298.050 132.600 331.950 ;
        RECT 133.950 331.800 136.050 333.900 ;
        RECT 139.950 331.950 142.050 334.050 ;
        RECT 133.950 304.950 136.050 307.050 ;
        RECT 115.950 295.950 118.050 298.050 ;
        RECT 130.950 295.950 133.050 298.050 ;
        RECT 112.950 292.950 115.050 295.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 100.950 289.950 103.050 292.050 ;
        RECT 103.950 289.950 106.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 94.950 286.950 97.050 289.050 ;
        RECT 101.400 288.900 102.600 289.950 ;
        RECT 95.400 262.050 96.600 286.950 ;
        RECT 100.950 286.800 103.050 288.900 ;
        RECT 107.400 277.050 108.600 289.950 ;
        RECT 106.950 274.950 109.050 277.050 ;
        RECT 106.950 268.950 109.050 271.050 ;
        RECT 94.950 259.950 97.050 262.050 ;
        RECT 100.950 260.100 103.050 262.200 ;
        RECT 101.400 259.050 102.600 260.100 ;
        RECT 107.400 259.050 108.600 268.950 ;
        RECT 113.400 262.200 114.600 292.950 ;
        RECT 116.400 283.050 117.600 295.950 ;
        RECT 121.950 293.100 124.050 295.200 ;
        RECT 127.950 293.100 130.050 295.200 ;
        RECT 134.400 295.050 135.600 304.950 ;
        RECT 136.950 298.950 139.050 301.050 ;
        RECT 122.400 292.050 123.600 293.100 ;
        RECT 128.400 292.050 129.600 293.100 ;
        RECT 133.950 292.950 136.050 295.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 124.950 289.950 127.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 118.950 286.950 121.050 289.050 ;
        RECT 115.950 280.950 118.050 283.050 ;
        RECT 119.400 265.050 120.600 286.950 ;
        RECT 125.400 283.050 126.600 289.950 ;
        RECT 131.400 288.900 132.600 289.950 ;
        RECT 137.400 289.050 138.600 298.950 ;
        RECT 130.950 286.800 133.050 288.900 ;
        RECT 133.950 286.950 136.050 289.050 ;
        RECT 136.950 286.950 139.050 289.050 ;
        RECT 127.950 283.950 130.050 286.050 ;
        RECT 124.950 280.950 127.050 283.050 ;
        RECT 128.400 274.050 129.600 283.950 ;
        RECT 127.950 271.950 130.050 274.050 ;
        RECT 118.950 262.950 121.050 265.050 ;
        RECT 130.950 262.950 133.050 265.050 ;
        RECT 112.950 260.100 115.050 262.200 ;
        RECT 121.950 260.100 124.050 262.200 ;
        RECT 122.400 259.050 123.600 260.100 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 98.400 255.900 99.600 256.950 ;
        RECT 97.950 253.800 100.050 255.900 ;
        RECT 104.400 247.050 105.600 256.950 ;
        RECT 110.400 255.900 111.600 256.950 ;
        RECT 109.950 253.800 112.050 255.900 ;
        RECT 119.400 255.000 120.600 256.950 ;
        RECT 112.950 250.950 115.050 253.050 ;
        RECT 118.950 250.950 121.050 255.000 ;
        RECT 103.950 244.950 106.050 247.050 ;
        RECT 106.950 222.600 109.050 223.050 ;
        RECT 95.400 221.400 109.050 222.600 ;
        RECT 95.400 217.200 96.600 221.400 ;
        RECT 106.950 220.950 109.050 221.400 ;
        RECT 94.950 215.100 97.050 217.200 ;
        RECT 97.950 216.000 100.050 220.050 ;
        RECT 103.950 216.000 106.050 220.050 ;
        RECT 98.400 214.050 99.600 216.000 ;
        RECT 104.400 214.050 105.600 216.000 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 85.950 208.950 88.050 211.050 ;
        RECT 91.950 208.950 94.050 211.050 ;
        RECT 79.950 190.950 82.050 193.050 ;
        RECT 82.950 184.950 85.050 187.050 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 73.950 178.950 76.050 181.050 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 59.400 172.050 60.600 178.950 ;
        RECT 58.950 169.950 61.050 172.050 ;
        RECT 65.400 163.050 66.600 178.950 ;
        RECT 70.950 175.950 73.050 178.050 ;
        RECT 77.400 177.900 78.600 178.950 ;
        RECT 64.950 160.950 67.050 163.050 ;
        RECT 58.950 157.950 61.050 160.050 ;
        RECT 59.400 142.050 60.600 157.950 ;
        RECT 61.950 151.950 64.050 154.050 ;
        RECT 58.950 139.950 61.050 142.050 ;
        RECT 55.950 137.100 58.050 139.200 ;
        RECT 56.400 136.050 57.600 137.100 ;
        RECT 62.400 136.050 63.600 151.950 ;
        RECT 55.950 133.950 58.050 136.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 52.950 130.950 55.050 133.050 ;
        RECT 53.400 118.050 54.600 130.950 ;
        RECT 52.950 115.950 55.050 118.050 ;
        RECT 59.400 115.050 60.600 133.950 ;
        RECT 65.400 127.050 66.600 133.950 ;
        RECT 71.400 132.900 72.600 175.950 ;
        RECT 76.950 175.800 79.050 177.900 ;
        RECT 77.400 136.050 78.600 175.800 ;
        RECT 83.400 172.050 84.600 184.950 ;
        RECT 86.400 175.050 87.600 208.950 ;
        RECT 101.400 207.600 102.600 211.950 ;
        RECT 98.400 206.400 102.600 207.600 ;
        RECT 94.950 187.950 97.050 190.050 ;
        RECT 95.400 181.050 96.600 187.950 ;
        RECT 98.400 187.050 99.600 206.400 ;
        RECT 103.950 205.050 106.050 208.050 ;
        RECT 107.400 205.050 108.600 211.950 ;
        RECT 100.950 204.000 106.050 205.050 ;
        RECT 100.950 203.400 105.600 204.000 ;
        RECT 100.950 202.950 105.000 203.400 ;
        RECT 106.950 202.950 109.050 205.050 ;
        RECT 100.950 199.800 103.050 201.900 ;
        RECT 97.950 184.950 100.050 187.050 ;
        RECT 101.400 181.050 102.600 199.800 ;
        RECT 113.400 193.050 114.600 250.950 ;
        RECT 125.400 235.050 126.600 256.950 ;
        RECT 131.400 255.900 132.600 262.950 ;
        RECT 130.950 253.800 133.050 255.900 ;
        RECT 124.950 232.950 127.050 235.050 ;
        RECT 121.950 220.950 124.050 223.050 ;
        RECT 122.400 214.050 123.600 220.950 ;
        RECT 130.950 217.950 133.050 220.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 121.950 211.950 124.050 214.050 ;
        RECT 124.950 211.950 127.050 214.050 ;
        RECT 119.400 205.050 120.600 211.950 ;
        RECT 125.400 210.900 126.600 211.950 ;
        RECT 131.400 210.900 132.600 217.950 ;
        RECT 124.950 208.800 127.050 210.900 ;
        RECT 130.950 208.800 133.050 210.900 ;
        RECT 134.400 207.600 135.600 286.950 ;
        RECT 136.950 268.950 139.050 271.050 ;
        RECT 137.400 223.050 138.600 268.950 ;
        RECT 140.400 262.050 141.600 331.950 ;
        RECT 143.400 295.200 144.600 346.800 ;
        RECT 146.400 334.050 147.600 361.950 ;
        RECT 155.400 349.050 156.600 364.950 ;
        RECT 157.950 361.950 160.050 364.050 ;
        RECT 154.950 346.950 157.050 349.050 ;
        RECT 158.400 340.200 159.600 361.950 ;
        RECT 161.400 355.050 162.600 367.950 ;
        RECT 170.400 361.050 171.600 376.950 ;
        RECT 178.950 372.000 181.050 376.050 ;
        RECT 182.400 373.050 183.600 434.400 ;
        RECT 184.950 430.950 187.050 433.050 ;
        RECT 185.400 373.050 186.600 430.950 ;
        RECT 188.400 427.050 189.600 478.950 ;
        RECT 203.400 475.050 204.600 493.950 ;
        RECT 202.950 472.950 205.050 475.050 ;
        RECT 206.400 471.600 207.600 508.950 ;
        RECT 203.400 470.400 207.600 471.600 ;
        RECT 196.950 449.100 199.050 451.200 ;
        RECT 197.400 448.050 198.600 449.100 ;
        RECT 193.950 445.950 196.050 448.050 ;
        RECT 196.950 445.950 199.050 448.050 ;
        RECT 194.400 439.050 195.600 445.950 ;
        RECT 199.950 442.950 202.050 445.050 ;
        RECT 193.950 436.950 196.050 439.050 ;
        RECT 200.400 433.050 201.600 442.950 ;
        RECT 203.400 441.600 204.600 470.400 ;
        RECT 205.950 457.950 208.050 460.050 ;
        RECT 206.400 445.050 207.600 457.950 ;
        RECT 205.950 442.950 208.050 445.050 ;
        RECT 203.400 440.400 207.600 441.600 ;
        RECT 199.950 430.950 202.050 433.050 ;
        RECT 187.950 424.950 190.050 427.050 ;
        RECT 199.950 421.950 202.050 424.050 ;
        RECT 193.950 416.100 196.050 421.050 ;
        RECT 194.400 415.050 195.600 416.100 ;
        RECT 200.400 415.050 201.600 421.950 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 193.950 412.950 196.050 415.050 ;
        RECT 196.950 412.950 199.050 415.050 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 191.400 394.050 192.600 412.950 ;
        RECT 190.950 391.950 193.050 394.050 ;
        RECT 197.400 391.050 198.600 412.950 ;
        RECT 196.950 388.950 199.050 391.050 ;
        RECT 206.400 385.050 207.600 440.400 ;
        RECT 209.400 439.050 210.600 512.400 ;
        RECT 221.400 511.050 222.600 527.400 ;
        RECT 230.400 526.050 231.600 550.950 ;
        RECT 233.400 541.050 234.600 565.950 ;
        RECT 235.950 565.800 238.050 567.900 ;
        RECT 242.400 556.050 243.600 568.950 ;
        RECT 244.950 565.950 247.050 568.050 ;
        RECT 241.950 553.950 244.050 556.050 ;
        RECT 232.950 538.950 235.050 541.050 ;
        RECT 241.950 538.950 244.050 541.050 ;
        RECT 232.950 532.950 235.050 537.900 ;
        RECT 235.950 532.950 238.050 535.050 ;
        RECT 236.400 529.200 237.600 532.950 ;
        RECT 235.950 527.100 238.050 529.200 ;
        RECT 236.400 526.050 237.600 527.100 ;
        RECT 226.950 523.950 229.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 220.950 508.950 223.050 511.050 ;
        RECT 214.950 494.100 217.050 496.200 ;
        RECT 220.950 494.100 223.050 496.200 ;
        RECT 227.400 496.050 228.600 523.950 ;
        RECT 233.400 522.900 234.600 523.950 ;
        RECT 232.950 520.800 235.050 522.900 ;
        RECT 242.400 508.050 243.600 538.950 ;
        RECT 245.400 529.050 246.600 565.950 ;
        RECT 248.400 550.050 249.600 599.400 ;
        RECT 254.400 586.050 255.600 632.400 ;
        RECT 256.950 613.950 259.050 616.050 ;
        RECT 253.950 585.600 256.050 586.050 ;
        RECT 251.400 584.400 256.050 585.600 ;
        RECT 251.400 574.050 252.600 584.400 ;
        RECT 253.950 583.950 256.050 584.400 ;
        RECT 253.950 577.950 256.050 580.050 ;
        RECT 250.950 571.950 253.050 574.050 ;
        RECT 254.400 571.050 255.600 577.950 ;
        RECT 257.400 577.050 258.600 613.950 ;
        RECT 260.400 610.050 261.600 634.800 ;
        RECT 269.400 613.050 270.600 646.950 ;
        RECT 275.400 645.900 276.600 646.950 ;
        RECT 274.950 643.800 277.050 645.900 ;
        RECT 284.400 637.050 285.600 673.800 ;
        RECT 286.950 670.950 289.050 673.050 ;
        RECT 283.950 634.950 286.050 637.050 ;
        RECT 268.950 610.950 271.050 613.050 ;
        RECT 287.400 610.200 288.600 670.950 ;
        RECT 296.400 664.050 297.600 679.950 ;
        RECT 298.950 673.950 301.050 676.050 ;
        RECT 295.950 661.950 298.050 664.050 ;
        RECT 299.400 655.050 300.600 673.950 ;
        RECT 305.400 672.600 306.600 748.950 ;
        RECT 311.400 736.050 312.600 775.950 ;
        RECT 316.950 766.950 319.050 769.050 ;
        RECT 317.400 760.050 318.600 766.950 ;
        RECT 323.400 763.200 324.600 778.950 ;
        RECT 328.950 775.950 331.050 778.050 ;
        RECT 322.950 761.100 325.050 763.200 ;
        RECT 323.400 760.050 324.600 761.100 ;
        RECT 316.950 757.950 319.050 760.050 ;
        RECT 319.950 757.950 322.050 760.050 ;
        RECT 322.950 757.950 325.050 760.050 ;
        RECT 320.400 748.050 321.600 757.950 ;
        RECT 329.400 751.050 330.600 775.950 ;
        RECT 341.400 760.050 342.600 790.950 ;
        RECT 344.400 787.050 345.600 799.950 ;
        RECT 346.950 796.950 349.050 799.050 ;
        RECT 343.950 784.950 346.050 787.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 340.950 757.950 343.050 760.050 ;
        RECT 328.950 748.950 331.050 751.050 ;
        RECT 338.400 748.050 339.600 757.950 ;
        RECT 343.950 754.950 346.050 757.050 ;
        RECT 319.950 745.950 322.050 748.050 ;
        RECT 337.950 745.950 340.050 748.050 ;
        RECT 344.400 745.050 345.600 754.950 ;
        RECT 343.950 742.950 346.050 745.050 ;
        RECT 310.950 733.950 313.050 736.050 ;
        RECT 322.950 733.950 325.050 736.050 ;
        RECT 313.950 729.000 316.050 733.050 ;
        RECT 319.950 730.950 322.050 733.050 ;
        RECT 314.400 727.050 315.600 729.000 ;
        RECT 310.950 724.950 313.050 727.050 ;
        RECT 313.950 724.950 316.050 727.050 ;
        RECT 311.400 723.900 312.600 724.950 ;
        RECT 310.950 721.800 313.050 723.900 ;
        RECT 316.950 715.950 319.050 718.050 ;
        RECT 317.400 709.050 318.600 715.950 ;
        RECT 320.400 715.050 321.600 730.950 ;
        RECT 319.950 712.950 322.050 715.050 ;
        RECT 316.950 706.950 319.050 709.050 ;
        RECT 313.950 703.950 316.050 706.050 ;
        RECT 307.950 683.100 310.050 685.200 ;
        RECT 308.400 676.050 309.600 683.100 ;
        RECT 314.400 682.050 315.600 703.950 ;
        RECT 323.400 688.050 324.600 733.950 ;
        RECT 347.400 732.600 348.600 796.950 ;
        RECT 350.400 796.050 351.600 802.950 ;
        RECT 356.400 801.000 357.600 802.950 ;
        RECT 362.400 802.050 363.600 815.400 ;
        RECT 371.400 810.600 372.600 835.950 ;
        RECT 380.400 811.050 381.600 839.100 ;
        RECT 371.400 809.400 375.600 810.600 ;
        RECT 374.400 808.200 375.600 809.400 ;
        RECT 379.950 808.950 382.050 811.050 ;
        RECT 373.950 806.100 376.050 808.200 ;
        RECT 383.400 807.600 384.600 841.950 ;
        RECT 389.400 838.050 390.600 844.950 ;
        RECT 397.950 839.100 400.050 841.200 ;
        RECT 398.400 838.050 399.600 839.100 ;
        RECT 388.950 835.950 391.050 838.050 ;
        RECT 391.950 835.950 394.050 838.050 ;
        RECT 397.950 835.950 400.050 838.050 ;
        RECT 392.400 826.050 393.600 835.950 ;
        RECT 400.950 832.950 403.050 835.050 ;
        RECT 391.950 823.950 394.050 826.050 ;
        RECT 397.950 817.950 400.050 820.050 ;
        RECT 388.950 811.950 391.050 814.050 ;
        RECT 380.400 806.400 387.600 807.600 ;
        RECT 374.400 805.050 375.600 806.100 ;
        RECT 380.400 805.050 381.600 806.400 ;
        RECT 370.950 802.950 373.050 805.050 ;
        RECT 373.950 802.950 376.050 805.050 ;
        RECT 376.950 802.950 379.050 805.050 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 355.950 796.950 358.050 801.000 ;
        RECT 361.950 799.950 364.050 802.050 ;
        RECT 367.950 799.950 370.050 802.050 ;
        RECT 349.950 793.950 352.050 796.050 ;
        RECT 364.950 793.950 367.050 796.050 ;
        RECT 349.950 784.950 352.050 787.050 ;
        RECT 350.400 760.050 351.600 784.950 ;
        RECT 352.950 763.950 355.050 766.050 ;
        RECT 349.950 757.950 352.050 760.050 ;
        RECT 350.400 733.050 351.600 757.950 ;
        RECT 353.400 754.050 354.600 763.950 ;
        RECT 358.950 762.000 361.050 766.050 ;
        RECT 365.400 763.050 366.600 793.950 ;
        RECT 359.400 760.050 360.600 762.000 ;
        RECT 364.950 760.950 367.050 763.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 361.950 757.950 364.050 760.050 ;
        RECT 362.400 756.000 363.600 757.950 ;
        RECT 368.400 756.900 369.600 799.950 ;
        RECT 371.400 793.050 372.600 802.950 ;
        RECT 377.400 799.050 378.600 802.950 ;
        RECT 376.950 796.950 379.050 799.050 ;
        RECT 370.950 790.950 373.050 793.050 ;
        RECT 377.400 775.050 378.600 796.950 ;
        RECT 386.400 796.050 387.600 806.400 ;
        RECT 382.950 793.950 385.050 796.050 ;
        RECT 385.950 793.950 388.050 796.050 ;
        RECT 383.400 790.050 384.600 793.950 ;
        RECT 382.800 787.950 384.900 790.050 ;
        RECT 385.950 787.950 388.050 790.050 ;
        RECT 376.950 772.950 379.050 775.050 ;
        RECT 386.400 769.050 387.600 787.950 ;
        RECT 389.400 778.050 390.600 811.950 ;
        RECT 391.950 805.950 394.050 811.050 ;
        RECT 398.400 805.050 399.600 817.950 ;
        RECT 401.400 811.050 402.600 832.950 ;
        RECT 400.950 808.950 403.050 811.050 ;
        RECT 404.400 808.050 405.600 847.950 ;
        RECT 407.400 814.050 408.600 883.950 ;
        RECT 413.400 883.050 414.600 904.950 ;
        RECT 419.400 889.050 420.600 911.400 ;
        RECT 425.400 892.050 426.600 913.950 ;
        RECT 424.950 889.950 427.050 892.050 ;
        RECT 433.950 889.950 436.050 892.050 ;
        RECT 418.950 885.000 421.050 889.050 ;
        RECT 427.950 886.950 430.050 889.050 ;
        RECT 419.400 883.050 420.600 885.000 ;
        RECT 412.950 880.950 415.050 883.050 ;
        RECT 415.950 880.950 418.050 883.050 ;
        RECT 418.950 880.950 421.050 883.050 ;
        RECT 416.400 879.900 417.600 880.950 ;
        RECT 415.950 877.800 418.050 879.900 ;
        RECT 428.400 871.050 429.600 886.950 ;
        RECT 434.400 883.050 435.600 889.950 ;
        RECT 446.400 889.050 447.600 913.950 ;
        RECT 455.400 912.900 456.600 916.950 ;
        RECT 464.400 916.050 465.600 925.950 ;
        RECT 493.950 919.950 496.050 922.050 ;
        RECT 460.950 913.950 463.050 916.050 ;
        RECT 463.950 913.950 466.050 916.050 ;
        RECT 481.950 913.950 484.050 916.050 ;
        RECT 461.400 912.900 462.600 913.950 ;
        RECT 482.400 912.900 483.600 913.950 ;
        RECT 494.400 913.050 495.600 919.950 ;
        RECT 499.950 918.000 502.050 922.050 ;
        RECT 500.400 916.050 501.600 918.000 ;
        RECT 506.400 916.050 507.600 925.950 ;
        RECT 556.950 922.950 559.050 925.050 ;
        RECT 571.950 922.950 574.050 925.050 ;
        RECT 583.950 922.950 586.050 925.050 ;
        RECT 601.950 922.950 604.050 925.050 ;
        RECT 643.950 922.950 646.050 925.050 ;
        RECT 517.950 917.100 520.050 919.200 ;
        RECT 523.950 917.100 526.050 919.200 ;
        RECT 535.950 917.100 538.050 919.200 ;
        RECT 541.950 917.100 544.050 919.200 ;
        RECT 547.950 917.100 550.050 919.200 ;
        RECT 499.950 913.950 502.050 916.050 ;
        RECT 502.950 913.950 505.050 916.050 ;
        RECT 505.950 913.950 508.050 916.050 ;
        RECT 508.950 913.950 511.050 916.050 ;
        RECT 454.950 910.800 457.050 912.900 ;
        RECT 460.950 910.800 463.050 912.900 ;
        RECT 481.950 912.600 484.050 912.900 ;
        RECT 481.950 911.400 486.600 912.600 ;
        RECT 481.950 910.800 484.050 911.400 ;
        RECT 448.950 904.950 451.050 907.050 ;
        RECT 445.950 886.950 448.050 889.050 ;
        RECT 433.950 880.950 436.050 883.050 ;
        RECT 436.950 880.950 439.050 883.050 ;
        RECT 430.950 877.800 433.050 879.900 ;
        RECT 409.950 868.950 412.050 871.050 ;
        RECT 427.950 868.950 430.050 871.050 ;
        RECT 410.400 841.050 411.600 868.950 ;
        RECT 424.950 856.950 427.050 859.050 ;
        RECT 412.950 844.950 415.050 847.050 ;
        RECT 409.950 838.950 412.050 841.050 ;
        RECT 413.400 838.050 414.600 844.950 ;
        RECT 418.950 839.100 421.050 841.200 ;
        RECT 419.400 838.050 420.600 839.100 ;
        RECT 412.950 835.950 415.050 838.050 ;
        RECT 415.950 835.950 418.050 838.050 ;
        RECT 418.950 835.950 421.050 838.050 ;
        RECT 416.400 834.900 417.600 835.950 ;
        RECT 415.950 832.800 418.050 834.900 ;
        RECT 418.950 829.950 421.050 832.050 ;
        RECT 406.950 811.950 409.050 814.050 ;
        RECT 403.950 805.950 406.050 808.050 ;
        RECT 406.950 806.100 409.050 808.200 ;
        RECT 412.950 806.100 415.050 808.200 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 400.950 802.950 403.050 805.050 ;
        RECT 391.950 799.950 394.050 802.050 ;
        RECT 395.400 801.900 396.600 802.950 ;
        RECT 401.400 801.900 402.600 802.950 ;
        RECT 392.400 790.050 393.600 799.950 ;
        RECT 394.950 799.800 397.050 801.900 ;
        RECT 400.950 799.800 403.050 801.900 ;
        RECT 403.950 799.950 406.050 802.050 ;
        RECT 394.950 793.950 400.050 796.050 ;
        RECT 391.950 787.950 394.050 790.050 ;
        RECT 391.950 778.950 394.050 781.050 ;
        RECT 388.950 775.950 391.050 778.050 ;
        RECT 376.950 766.950 379.050 769.050 ;
        RECT 385.950 768.600 388.050 769.050 ;
        RECT 385.950 767.400 390.600 768.600 ;
        RECT 385.950 766.950 388.050 767.400 ;
        RECT 377.400 760.050 378.600 766.950 ;
        RECT 382.950 761.100 385.050 763.200 ;
        RECT 389.400 763.050 390.600 767.400 ;
        RECT 392.400 766.050 393.600 778.950 ;
        RECT 401.400 775.050 402.600 799.800 ;
        RECT 400.950 772.950 403.050 775.050 ;
        RECT 404.400 769.050 405.600 799.950 ;
        RECT 407.400 781.050 408.600 806.100 ;
        RECT 413.400 805.050 414.600 806.100 ;
        RECT 419.400 805.050 420.600 829.950 ;
        RECT 425.400 808.050 426.600 856.950 ;
        RECT 427.950 853.950 430.050 856.050 ;
        RECT 428.400 820.050 429.600 853.950 ;
        RECT 431.400 832.050 432.600 877.800 ;
        RECT 437.400 874.050 438.600 880.950 ;
        RECT 446.400 880.050 447.600 886.950 ;
        RECT 449.400 883.050 450.600 904.950 ;
        RECT 454.950 884.100 457.050 886.200 ;
        RECT 472.950 885.000 475.050 889.050 ;
        RECT 455.400 883.050 456.600 884.100 ;
        RECT 473.400 883.050 474.600 885.000 ;
        RECT 478.950 884.100 481.050 886.200 ;
        RECT 479.400 883.050 480.600 884.100 ;
        RECT 448.950 880.950 451.050 883.050 ;
        RECT 454.950 880.950 457.050 883.050 ;
        RECT 469.950 880.950 472.050 883.050 ;
        RECT 472.950 880.950 475.050 883.050 ;
        RECT 475.950 880.950 478.050 883.050 ;
        RECT 478.950 880.950 481.050 883.050 ;
        RECT 445.950 877.950 448.050 880.050 ;
        RECT 451.950 877.950 454.050 880.050 ;
        RECT 470.400 879.900 471.600 880.950 ;
        RECT 476.400 879.900 477.600 880.950 ;
        RECT 436.950 871.950 439.050 874.050 ;
        RECT 452.400 856.050 453.600 877.950 ;
        RECT 469.950 877.800 472.050 879.900 ;
        RECT 475.950 877.800 478.050 879.900 ;
        RECT 436.950 853.950 439.050 856.050 ;
        RECT 451.950 853.950 454.050 856.050 ;
        RECT 437.400 838.050 438.600 853.950 ;
        RECT 442.950 839.100 445.050 841.200 ;
        RECT 448.950 839.100 451.050 844.050 ;
        RECT 443.400 838.050 444.600 839.100 ;
        RECT 436.950 835.950 439.050 838.050 ;
        RECT 439.950 835.950 442.050 838.050 ;
        RECT 442.950 835.950 445.050 838.050 ;
        RECT 430.950 829.950 433.050 832.050 ;
        RECT 440.400 826.050 441.600 835.950 ;
        RECT 442.950 829.950 445.050 832.050 ;
        RECT 439.950 823.950 442.050 826.050 ;
        RECT 428.400 818.400 433.050 820.050 ;
        RECT 429.000 817.950 433.050 818.400 ;
        RECT 427.950 814.950 430.050 817.050 ;
        RECT 424.950 805.950 427.050 808.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 415.950 802.950 418.050 805.050 ;
        RECT 418.950 802.950 421.050 805.050 ;
        RECT 421.950 802.950 424.050 805.050 ;
        RECT 416.400 801.000 417.600 802.950 ;
        RECT 422.400 801.900 423.600 802.950 ;
        RECT 415.950 796.950 418.050 801.000 ;
        RECT 421.950 799.800 424.050 801.900 ;
        RECT 424.950 799.950 427.050 802.050 ;
        RECT 428.400 801.900 429.600 814.950 ;
        RECT 433.950 806.100 436.050 808.200 ;
        RECT 434.400 805.050 435.600 806.100 ;
        RECT 433.950 802.950 436.050 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 415.950 781.950 418.050 784.050 ;
        RECT 406.950 778.950 409.050 781.050 ;
        RECT 412.950 775.950 415.050 778.050 ;
        RECT 394.950 766.950 397.050 769.050 ;
        RECT 403.950 766.950 406.050 769.050 ;
        RECT 391.950 763.950 394.050 766.050 ;
        RECT 383.400 760.050 384.600 761.100 ;
        RECT 388.950 760.950 391.050 763.050 ;
        RECT 391.950 760.800 394.050 762.900 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 379.950 757.950 382.050 760.050 ;
        RECT 382.950 757.950 385.050 760.050 ;
        RECT 385.950 757.950 388.050 760.050 ;
        RECT 352.950 751.950 355.050 754.050 ;
        RECT 361.950 751.950 364.050 756.000 ;
        RECT 367.950 754.800 370.050 756.900 ;
        RECT 370.950 754.950 373.050 757.050 ;
        RECT 374.400 756.900 375.600 757.950 ;
        RECT 362.400 748.050 363.600 751.950 ;
        RECT 361.950 745.950 364.050 748.050 ;
        RECT 358.950 736.950 361.050 739.050 ;
        RECT 352.950 733.950 355.050 736.050 ;
        RECT 344.400 731.400 348.600 732.600 ;
        RECT 331.950 728.100 334.050 730.200 ;
        RECT 332.400 727.050 333.600 728.100 ;
        RECT 340.950 727.950 343.050 730.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 331.950 724.950 334.050 727.050 ;
        RECT 334.950 724.950 337.050 727.050 ;
        RECT 329.400 723.900 330.600 724.950 ;
        RECT 335.400 723.900 336.600 724.950 ;
        RECT 328.950 721.800 331.050 723.900 ;
        RECT 334.950 721.800 337.050 723.900 ;
        RECT 341.400 721.050 342.600 727.950 ;
        RECT 344.400 723.900 345.600 731.400 ;
        RECT 349.950 730.950 352.050 733.050 ;
        RECT 353.400 727.050 354.600 733.950 ;
        RECT 359.400 727.050 360.600 736.950 ;
        RECT 364.950 733.950 367.050 736.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 352.950 724.950 355.050 727.050 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 343.950 721.800 346.050 723.900 ;
        RECT 350.400 723.000 351.600 724.950 ;
        RECT 356.400 723.000 357.600 724.950 ;
        RECT 340.950 718.950 343.050 721.050 ;
        RECT 337.950 709.950 340.050 712.050 ;
        RECT 328.950 700.950 331.050 703.050 ;
        RECT 322.950 685.950 325.050 688.050 ;
        RECT 319.950 683.100 322.050 685.200 ;
        RECT 320.400 682.050 321.600 683.100 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 316.950 679.950 319.050 682.050 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 322.950 679.950 325.050 682.050 ;
        RECT 317.400 678.900 318.600 679.950 ;
        RECT 316.950 676.800 319.050 678.900 ;
        RECT 307.950 673.950 310.050 676.050 ;
        RECT 305.400 671.400 309.600 672.600 ;
        RECT 298.950 651.600 301.050 655.050 ;
        RECT 296.400 651.000 301.050 651.600 ;
        RECT 296.400 650.400 300.600 651.000 ;
        RECT 296.400 649.050 297.600 650.400 ;
        RECT 292.950 646.950 295.050 649.050 ;
        RECT 295.950 646.950 298.050 649.050 ;
        RECT 301.950 646.950 304.050 649.050 ;
        RECT 259.950 607.950 262.050 610.050 ;
        RECT 265.950 606.000 268.050 610.050 ;
        RECT 277.950 607.950 280.050 610.050 ;
        RECT 266.400 604.050 267.600 606.000 ;
        RECT 271.950 605.100 274.050 607.200 ;
        RECT 272.400 604.050 273.600 605.100 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 265.950 601.950 268.050 604.050 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 259.950 598.950 262.050 601.050 ;
        RECT 260.400 585.600 261.600 598.950 ;
        RECT 263.400 589.050 264.600 601.950 ;
        RECT 269.400 600.900 270.600 601.950 ;
        RECT 268.950 598.800 271.050 600.900 ;
        RECT 274.950 598.950 277.050 601.050 ;
        RECT 265.950 597.600 270.000 598.050 ;
        RECT 265.950 597.000 270.600 597.600 ;
        RECT 265.950 595.950 271.050 597.000 ;
        RECT 268.950 592.950 271.050 595.950 ;
        RECT 275.400 595.050 276.600 598.950 ;
        RECT 274.950 592.950 277.050 595.050 ;
        RECT 265.950 589.950 268.050 592.050 ;
        RECT 262.950 586.950 265.050 589.050 ;
        RECT 260.400 585.000 264.600 585.600 ;
        RECT 260.400 584.400 265.050 585.000 ;
        RECT 262.950 580.950 265.050 584.400 ;
        RECT 259.950 577.950 262.050 580.050 ;
        RECT 256.950 574.950 259.050 577.050 ;
        RECT 260.400 571.050 261.600 577.950 ;
        RECT 266.400 574.050 267.600 589.950 ;
        RECT 275.400 576.600 276.600 592.950 ;
        RECT 278.400 592.050 279.600 607.950 ;
        RECT 280.950 604.950 283.050 610.050 ;
        RECT 286.950 608.100 289.050 610.200 ;
        RECT 293.400 610.050 294.600 646.950 ;
        RECT 302.400 645.000 303.600 646.950 ;
        RECT 295.950 640.950 298.050 643.050 ;
        RECT 301.950 640.950 304.050 645.000 ;
        RECT 296.400 631.050 297.600 640.950 ;
        RECT 298.950 631.950 301.050 634.050 ;
        RECT 295.950 628.950 298.050 631.050 ;
        RECT 292.950 607.950 295.050 610.050 ;
        RECT 286.950 604.950 289.050 607.050 ;
        RECT 287.400 604.050 288.600 604.950 ;
        RECT 283.950 601.950 286.050 604.050 ;
        RECT 286.950 601.950 289.050 604.050 ;
        RECT 284.400 600.900 285.600 601.950 ;
        RECT 283.950 598.800 286.050 600.900 ;
        RECT 293.400 600.600 294.600 607.950 ;
        RECT 295.950 605.100 298.050 607.200 ;
        RECT 299.400 607.050 300.600 631.950 ;
        RECT 308.400 619.050 309.600 671.400 ;
        RECT 310.950 670.950 313.050 673.050 ;
        RECT 311.400 643.050 312.600 670.950 ;
        RECT 323.400 670.050 324.600 679.950 ;
        RECT 325.950 676.950 328.050 679.050 ;
        RECT 326.400 673.050 327.600 676.950 ;
        RECT 329.400 676.050 330.600 700.950 ;
        RECT 331.950 685.950 334.050 688.050 ;
        RECT 328.950 673.950 331.050 676.050 ;
        RECT 325.800 670.950 327.900 673.050 ;
        RECT 328.950 670.800 331.050 672.900 ;
        RECT 322.950 667.950 325.050 670.050 ;
        RECT 319.950 658.950 322.050 661.050 ;
        RECT 320.400 649.050 321.600 658.950 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 317.400 643.050 318.600 646.950 ;
        RECT 310.950 640.950 313.050 643.050 ;
        RECT 316.950 640.950 319.050 643.050 ;
        RECT 313.950 634.950 316.050 637.050 ;
        RECT 317.400 636.600 318.600 640.950 ;
        RECT 317.400 635.400 321.600 636.600 ;
        RECT 307.950 616.950 310.050 619.050 ;
        RECT 290.400 599.400 294.600 600.600 ;
        RECT 277.950 589.950 280.050 592.050 ;
        RECT 283.950 580.950 286.050 583.050 ;
        RECT 277.950 577.950 280.050 580.050 ;
        RECT 272.400 575.400 276.600 576.600 ;
        RECT 265.950 571.950 268.050 574.050 ;
        RECT 272.400 571.050 273.600 575.400 ;
        RECT 278.400 571.050 279.600 577.950 ;
        RECT 284.400 574.050 285.600 580.950 ;
        RECT 286.950 577.950 289.050 580.050 ;
        RECT 283.950 571.950 286.050 574.050 ;
        RECT 253.950 568.950 256.050 571.050 ;
        RECT 256.950 568.950 259.050 571.050 ;
        RECT 259.950 568.950 262.050 571.050 ;
        RECT 262.950 568.950 265.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 277.950 568.950 280.050 571.050 ;
        RECT 280.950 568.950 283.050 571.050 ;
        RECT 257.400 567.900 258.600 568.950 ;
        RECT 250.950 565.800 253.050 567.900 ;
        RECT 256.950 565.800 259.050 567.900 ;
        RECT 263.400 567.000 264.600 568.950 ;
        RECT 251.400 562.050 252.600 565.800 ;
        RECT 255.000 564.750 258.000 565.050 ;
        RECT 253.950 562.950 259.050 564.750 ;
        RECT 262.950 562.950 265.050 567.000 ;
        RECT 265.950 565.950 268.050 568.050 ;
        RECT 275.400 567.900 276.600 568.950 ;
        RECT 281.400 568.050 282.600 568.950 ;
        RECT 253.950 562.650 256.050 562.950 ;
        RECT 256.950 562.650 259.050 562.950 ;
        RECT 250.950 559.950 253.050 562.050 ;
        RECT 262.950 559.800 265.050 561.900 ;
        RECT 247.950 547.950 250.050 550.050 ;
        RECT 256.950 547.950 259.050 550.050 ;
        RECT 247.950 544.800 250.050 546.900 ;
        RECT 248.400 535.050 249.600 544.800 ;
        RECT 247.950 532.950 250.050 535.050 ;
        RECT 257.400 532.050 258.600 547.950 ;
        RECT 259.950 541.950 262.050 544.050 ;
        RECT 260.400 538.050 261.600 541.950 ;
        RECT 263.400 541.050 264.600 559.800 ;
        RECT 266.400 559.050 267.600 565.950 ;
        RECT 274.950 565.800 277.050 567.900 ;
        RECT 281.400 566.400 286.050 568.050 ;
        RECT 282.000 565.950 286.050 566.400 ;
        RECT 275.400 564.600 276.600 565.800 ;
        RECT 287.400 565.050 288.600 577.950 ;
        RECT 290.400 577.050 291.600 599.400 ;
        RECT 292.950 595.950 295.050 598.050 ;
        RECT 289.950 574.950 292.050 577.050 ;
        RECT 293.400 574.050 294.600 595.950 ;
        RECT 296.400 595.050 297.600 605.100 ;
        RECT 298.950 604.950 301.050 607.050 ;
        RECT 301.950 606.000 304.050 610.050 ;
        RECT 302.400 604.050 303.600 606.000 ;
        RECT 307.950 605.100 310.050 607.200 ;
        RECT 308.400 604.050 309.600 605.100 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 304.950 601.950 307.050 604.050 ;
        RECT 307.950 601.950 310.050 604.050 ;
        RECT 295.950 592.950 298.050 595.050 ;
        RECT 305.400 592.050 306.600 601.950 ;
        RECT 314.400 601.050 315.600 634.950 ;
        RECT 320.400 627.600 321.600 635.400 ;
        RECT 323.400 630.600 324.600 646.950 ;
        RECT 329.400 637.050 330.600 670.800 ;
        RECT 328.950 634.950 331.050 637.050 ;
        RECT 323.400 629.400 327.600 630.600 ;
        RECT 320.400 626.400 324.600 627.600 ;
        RECT 316.950 616.950 319.050 619.050 ;
        RECT 310.950 598.950 313.050 601.050 ;
        RECT 313.950 598.950 316.050 601.050 ;
        RECT 304.950 589.950 307.050 592.050 ;
        RECT 301.950 577.950 304.050 580.050 ;
        RECT 289.950 571.800 292.050 573.900 ;
        RECT 292.950 571.950 295.050 574.050 ;
        RECT 295.950 572.100 298.050 574.200 ;
        RECT 275.400 563.400 279.600 564.600 ;
        RECT 268.950 559.950 271.050 562.050 ;
        RECT 274.950 559.950 277.050 562.050 ;
        RECT 265.950 556.950 268.050 559.050 ;
        RECT 269.400 556.050 270.600 559.950 ;
        RECT 275.400 556.050 276.600 559.950 ;
        RECT 278.400 558.600 279.600 563.400 ;
        RECT 286.950 562.950 289.050 565.050 ;
        RECT 278.400 557.400 282.600 558.600 ;
        RECT 268.950 553.950 271.050 556.050 ;
        RECT 274.950 553.950 277.050 556.050 ;
        RECT 271.950 550.950 274.050 553.050 ;
        RECT 262.950 538.950 265.050 541.050 ;
        RECT 259.950 535.950 262.050 538.050 ;
        RECT 256.950 529.950 259.050 532.050 ;
        RECT 244.950 526.950 247.050 529.050 ;
        RECT 250.950 527.100 253.050 529.200 ;
        RECT 251.400 526.050 252.600 527.100 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 250.950 523.950 253.050 526.050 ;
        RECT 244.950 520.950 247.050 523.050 ;
        RECT 248.400 522.900 249.600 523.950 ;
        RECT 229.950 505.950 232.050 508.050 ;
        RECT 241.950 505.950 244.050 508.050 ;
        RECT 215.400 493.050 216.600 494.100 ;
        RECT 221.400 493.050 222.600 494.100 ;
        RECT 226.950 493.950 229.050 496.050 ;
        RECT 214.950 490.950 217.050 493.050 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 220.950 490.950 223.050 493.050 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 211.950 469.950 214.050 472.050 ;
        RECT 212.400 451.050 213.600 469.950 ;
        RECT 218.400 469.050 219.600 490.950 ;
        RECT 224.400 489.900 225.600 490.950 ;
        RECT 223.950 487.800 226.050 489.900 ;
        RECT 223.950 478.950 226.050 481.050 ;
        RECT 217.950 466.950 220.050 469.050 ;
        RECT 224.400 451.200 225.600 478.950 ;
        RECT 211.950 448.950 214.050 451.050 ;
        RECT 217.950 449.100 220.050 451.200 ;
        RECT 223.950 449.100 226.050 451.200 ;
        RECT 218.400 448.050 219.600 449.100 ;
        RECT 224.400 448.050 225.600 449.100 ;
        RECT 214.950 445.950 217.050 448.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 220.950 445.950 223.050 448.050 ;
        RECT 223.950 445.950 226.050 448.050 ;
        RECT 215.400 444.900 216.600 445.950 ;
        RECT 214.950 442.800 217.050 444.900 ;
        RECT 221.400 439.050 222.600 445.950 ;
        RECT 226.950 442.950 229.050 445.050 ;
        RECT 208.950 436.950 211.050 439.050 ;
        RECT 220.950 438.600 223.050 439.050 ;
        RECT 220.950 437.400 225.600 438.600 ;
        RECT 220.950 436.950 223.050 437.400 ;
        RECT 224.400 421.050 225.600 437.400 ;
        RECT 227.400 421.050 228.600 442.950 ;
        RECT 214.950 416.100 217.050 418.200 ;
        RECT 220.950 417.000 223.050 421.050 ;
        RECT 223.950 418.950 226.050 421.050 ;
        RECT 226.950 418.950 229.050 421.050 ;
        RECT 230.400 420.600 231.600 505.950 ;
        RECT 232.950 499.950 235.050 502.050 ;
        RECT 241.950 499.950 244.050 502.050 ;
        RECT 233.400 496.050 234.600 499.950 ;
        RECT 242.400 496.050 243.600 499.950 ;
        RECT 232.950 493.950 235.050 496.050 ;
        RECT 240.000 495.600 244.050 496.050 ;
        RECT 239.400 493.950 244.050 495.600 ;
        RECT 239.400 493.050 240.600 493.950 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 232.950 487.950 235.050 490.050 ;
        RECT 236.400 489.900 237.600 490.950 ;
        RECT 233.400 442.050 234.600 487.950 ;
        RECT 235.950 487.800 238.050 489.900 ;
        RECT 245.400 472.050 246.600 520.950 ;
        RECT 247.950 520.800 250.050 522.900 ;
        RECT 248.400 517.050 249.600 520.800 ;
        RECT 257.400 520.050 258.600 529.950 ;
        RECT 260.400 526.050 261.600 535.950 ;
        RECT 265.950 527.100 268.050 529.200 ;
        RECT 266.400 526.050 267.600 527.100 ;
        RECT 272.400 526.050 273.600 550.950 ;
        RECT 281.400 550.050 282.600 557.400 ;
        RECT 280.950 547.950 283.050 550.050 ;
        RECT 277.950 532.950 280.050 538.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 268.950 523.950 271.050 526.050 ;
        RECT 271.950 523.950 274.050 526.050 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 256.950 517.950 259.050 520.050 ;
        RECT 260.400 517.050 261.600 523.950 ;
        RECT 265.950 517.950 268.050 520.050 ;
        RECT 247.950 514.950 250.050 517.050 ;
        RECT 259.950 514.950 262.050 517.050 ;
        RECT 248.400 499.050 249.600 514.950 ;
        RECT 262.950 499.950 265.050 502.050 ;
        RECT 247.950 496.950 250.050 499.050 ;
        RECT 247.950 493.800 250.050 495.900 ;
        RECT 256.950 495.000 259.050 499.050 ;
        RECT 248.400 481.050 249.600 493.800 ;
        RECT 257.400 493.050 258.600 495.000 ;
        RECT 263.400 493.050 264.600 499.950 ;
        RECT 266.400 496.050 267.600 517.950 ;
        RECT 269.400 517.050 270.600 523.950 ;
        RECT 275.400 522.900 276.600 523.950 ;
        RECT 274.950 520.800 277.050 522.900 ;
        RECT 275.400 519.600 276.600 520.800 ;
        RECT 272.400 518.400 276.600 519.600 ;
        RECT 268.950 514.950 271.050 517.050 ;
        RECT 268.950 496.950 271.050 499.050 ;
        RECT 265.950 493.950 268.050 496.050 ;
        RECT 253.950 490.950 256.050 493.050 ;
        RECT 256.950 490.950 259.050 493.050 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 262.950 490.950 265.050 493.050 ;
        RECT 250.950 489.600 253.050 490.050 ;
        RECT 254.400 489.600 255.600 490.950 ;
        RECT 250.950 488.400 255.600 489.600 ;
        RECT 250.950 487.950 253.050 488.400 ;
        RECT 247.950 478.950 250.050 481.050 ;
        RECT 251.400 478.050 252.600 487.950 ;
        RECT 253.950 484.950 256.050 487.050 ;
        RECT 250.950 475.950 253.050 478.050 ;
        RECT 254.400 472.050 255.600 484.950 ;
        RECT 256.950 481.950 259.050 484.050 ;
        RECT 244.950 469.950 247.050 472.050 ;
        RECT 253.950 469.950 256.050 472.050 ;
        RECT 257.400 469.050 258.600 481.950 ;
        RECT 260.400 481.050 261.600 490.950 ;
        RECT 265.950 487.950 268.050 490.050 ;
        RECT 259.950 478.950 262.050 481.050 ;
        RECT 256.950 466.950 259.050 469.050 ;
        RECT 250.950 463.950 253.050 466.050 ;
        RECT 241.950 460.950 244.050 463.050 ;
        RECT 242.400 457.050 243.600 460.950 ;
        RECT 251.400 460.050 252.600 463.950 ;
        RECT 262.950 460.950 265.050 463.050 ;
        RECT 250.800 457.950 252.900 460.050 ;
        RECT 253.950 457.950 256.050 460.050 ;
        RECT 241.950 454.950 244.050 457.050 ;
        RECT 242.400 448.050 243.600 454.950 ;
        RECT 247.950 450.000 250.050 454.050 ;
        RECT 254.400 451.050 255.600 457.950 ;
        RECT 248.400 448.050 249.600 450.000 ;
        RECT 253.950 448.950 256.050 451.050 ;
        RECT 256.950 450.000 259.050 454.050 ;
        RECT 257.400 448.050 258.600 450.000 ;
        RECT 263.400 448.050 264.600 460.950 ;
        RECT 266.400 460.050 267.600 487.950 ;
        RECT 269.400 481.050 270.600 496.950 ;
        RECT 268.950 478.950 271.050 481.050 ;
        RECT 265.950 457.950 268.050 460.050 ;
        RECT 272.400 454.050 273.600 518.400 ;
        RECT 281.400 517.050 282.600 547.950 ;
        RECT 283.950 538.950 286.050 541.050 ;
        RECT 284.400 529.050 285.600 538.950 ;
        RECT 290.400 538.050 291.600 571.800 ;
        RECT 296.400 571.050 297.600 572.100 ;
        RECT 302.400 571.050 303.600 577.950 ;
        RECT 295.950 568.950 298.050 571.050 ;
        RECT 298.950 568.950 301.050 571.050 ;
        RECT 301.950 568.950 304.050 571.050 ;
        RECT 304.950 568.950 307.050 571.050 ;
        RECT 292.950 565.950 295.050 568.050 ;
        RECT 299.400 567.900 300.600 568.950 ;
        RECT 293.400 556.050 294.600 565.950 ;
        RECT 298.950 565.800 301.050 567.900 ;
        RECT 305.400 567.000 306.600 568.950 ;
        RECT 304.950 562.950 307.050 567.000 ;
        RECT 307.950 565.950 310.050 568.050 ;
        RECT 292.950 553.950 295.050 556.050 ;
        RECT 295.950 544.950 298.050 547.050 ;
        RECT 292.950 541.950 295.050 544.050 ;
        RECT 286.950 535.950 289.050 538.050 ;
        RECT 289.950 535.950 292.050 538.050 ;
        RECT 283.950 526.950 286.050 529.050 ;
        RECT 287.400 528.600 288.600 535.950 ;
        RECT 293.400 532.050 294.600 541.950 ;
        RECT 292.950 529.950 295.050 532.050 ;
        RECT 287.400 527.400 291.600 528.600 ;
        RECT 290.400 526.050 291.600 527.400 ;
        RECT 296.400 526.050 297.600 544.950 ;
        RECT 308.400 529.050 309.600 565.950 ;
        RECT 311.400 565.050 312.600 598.950 ;
        RECT 313.950 592.950 316.050 595.050 ;
        RECT 314.400 565.050 315.600 592.950 ;
        RECT 310.950 562.950 313.050 565.050 ;
        RECT 313.950 562.950 316.050 565.050 ;
        RECT 317.400 559.050 318.600 616.950 ;
        RECT 319.950 604.950 322.050 610.050 ;
        RECT 323.400 607.200 324.600 626.400 ;
        RECT 326.400 619.050 327.600 629.400 ;
        RECT 325.950 616.950 328.050 619.050 ;
        RECT 332.400 610.050 333.600 685.950 ;
        RECT 338.400 682.050 339.600 709.950 ;
        RECT 344.400 694.050 345.600 721.800 ;
        RECT 349.950 718.950 352.050 723.000 ;
        RECT 355.950 718.950 358.050 723.000 ;
        RECT 361.950 721.950 364.050 724.050 ;
        RECT 358.950 709.950 361.050 712.050 ;
        RECT 352.950 703.950 355.050 706.050 ;
        RECT 349.950 697.950 352.050 700.050 ;
        RECT 343.950 691.950 346.050 694.050 ;
        RECT 337.950 679.950 340.050 682.050 ;
        RECT 343.950 679.950 346.050 682.050 ;
        RECT 344.400 673.050 345.600 679.950 ;
        RECT 343.950 670.950 346.050 673.050 ;
        RECT 343.950 661.950 346.050 664.050 ;
        RECT 344.400 649.050 345.600 661.950 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 343.950 646.950 346.050 649.050 ;
        RECT 338.400 622.050 339.600 646.950 ;
        RECT 337.950 619.950 340.050 622.050 ;
        RECT 337.950 616.800 340.050 618.900 ;
        RECT 331.950 607.950 334.050 610.050 ;
        RECT 322.950 605.100 325.050 607.200 ;
        RECT 323.400 604.050 324.600 605.100 ;
        RECT 331.950 604.800 334.050 606.900 ;
        RECT 322.950 601.950 325.050 604.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 326.400 600.600 327.600 601.950 ;
        RECT 326.400 599.400 330.600 600.600 ;
        RECT 319.950 592.950 322.050 595.050 ;
        RECT 320.400 574.050 321.600 592.950 ;
        RECT 325.950 580.950 328.050 583.050 ;
        RECT 319.950 571.950 322.050 574.050 ;
        RECT 326.400 571.050 327.600 580.950 ;
        RECT 329.400 574.050 330.600 599.400 ;
        RECT 332.400 577.050 333.600 604.800 ;
        RECT 338.400 604.050 339.600 616.800 ;
        RECT 350.400 613.050 351.600 697.950 ;
        RECT 353.400 685.200 354.600 703.950 ;
        RECT 359.400 700.050 360.600 709.950 ;
        RECT 362.400 706.050 363.600 721.950 ;
        RECT 365.400 709.050 366.600 733.950 ;
        RECT 364.950 706.950 367.050 709.050 ;
        RECT 361.950 703.950 364.050 706.050 ;
        RECT 358.950 697.950 361.050 700.050 ;
        RECT 364.950 691.950 367.050 694.050 ;
        RECT 355.950 688.950 358.050 691.050 ;
        RECT 352.950 683.100 355.050 685.200 ;
        RECT 356.400 682.050 357.600 688.950 ;
        RECT 365.400 685.050 366.600 691.950 ;
        RECT 364.950 682.950 367.050 685.050 ;
        RECT 368.400 682.050 369.600 754.800 ;
        RECT 371.400 739.050 372.600 754.950 ;
        RECT 373.950 754.800 376.050 756.900 ;
        RECT 380.400 739.050 381.600 757.950 ;
        RECT 386.400 756.900 387.600 757.950 ;
        RECT 385.950 754.800 388.050 756.900 ;
        RECT 370.950 736.950 373.050 739.050 ;
        RECT 376.800 736.950 378.900 739.050 ;
        RECT 379.950 736.950 382.050 739.050 ;
        RECT 388.950 736.950 391.050 739.050 ;
        RECT 373.650 731.400 375.750 733.500 ;
        RECT 371.400 725.100 373.500 727.200 ;
        RECT 371.400 722.550 372.600 725.100 ;
        RECT 374.400 718.800 375.300 731.400 ;
        RECT 377.400 729.900 378.600 736.950 ;
        RECT 380.400 732.900 381.600 735.450 ;
        RECT 380.400 730.800 382.500 732.900 ;
        RECT 383.700 731.100 385.800 733.200 ;
        RECT 389.400 733.050 390.600 736.950 ;
        RECT 392.400 736.050 393.600 760.800 ;
        RECT 391.950 733.950 394.050 736.050 ;
        RECT 376.200 729.000 378.600 729.900 ;
        RECT 376.200 727.800 383.250 729.000 ;
        RECT 381.150 726.900 383.250 727.800 ;
        RECT 376.200 726.000 378.300 726.900 ;
        RECT 384.150 726.000 385.050 731.100 ;
        RECT 388.950 730.950 391.050 733.050 ;
        RECT 391.950 730.800 394.050 732.900 ;
        RECT 386.400 727.200 387.600 729.600 ;
        RECT 376.200 725.100 385.050 726.000 ;
        RECT 385.950 725.100 388.050 727.200 ;
        RECT 376.200 724.800 378.300 725.100 ;
        RECT 380.400 722.100 382.500 724.200 ;
        RECT 374.100 716.700 376.200 718.800 ;
        RECT 380.400 715.050 381.600 722.100 ;
        RECT 384.150 718.500 385.050 725.100 ;
        RECT 392.400 724.050 393.600 730.800 ;
        RECT 391.950 718.950 394.050 724.050 ;
        RECT 383.100 716.400 385.200 718.500 ;
        RECT 379.950 712.950 382.050 715.050 ;
        RECT 380.400 691.050 381.600 712.950 ;
        RECT 376.500 688.500 378.600 690.600 ;
        RECT 379.950 688.950 382.050 691.050 ;
        RECT 355.950 679.950 358.050 682.050 ;
        RECT 361.950 679.950 364.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 373.950 679.950 376.050 682.050 ;
        RECT 376.950 681.300 378.000 688.500 ;
        RECT 380.400 684.900 381.600 687.450 ;
        RECT 386.100 687.300 388.200 689.400 ;
        RECT 391.950 688.950 394.050 691.050 ;
        RECT 379.800 682.800 381.900 684.900 ;
        RECT 382.800 683.700 384.900 685.800 ;
        RECT 382.800 681.300 383.700 683.700 ;
        RECT 376.950 680.100 383.700 681.300 ;
        RECT 362.400 678.600 363.600 679.950 ;
        RECT 362.400 677.400 366.600 678.600 ;
        RECT 352.950 673.950 355.050 676.050 ;
        RECT 353.400 652.050 354.600 673.950 ;
        RECT 365.400 666.600 366.600 677.400 ;
        RECT 368.400 670.050 369.600 679.950 ;
        RECT 374.400 677.400 375.600 679.950 ;
        RECT 376.950 674.700 377.850 680.100 ;
        RECT 378.750 678.300 380.850 679.200 ;
        RECT 386.400 678.300 387.300 687.300 ;
        RECT 389.400 682.050 390.600 684.600 ;
        RECT 392.400 682.050 393.600 688.950 ;
        RECT 388.500 679.950 390.600 682.050 ;
        RECT 391.950 679.950 394.050 682.050 ;
        RECT 378.750 677.100 387.300 678.300 ;
        RECT 376.500 672.600 378.600 674.700 ;
        RECT 379.800 674.100 381.900 676.200 ;
        RECT 383.700 675.300 385.800 677.100 ;
        RECT 367.950 667.950 370.050 670.050 ;
        RECT 370.950 666.600 373.050 667.050 ;
        RECT 365.400 665.400 373.050 666.600 ;
        RECT 370.950 664.950 373.050 665.400 ;
        RECT 380.400 664.050 381.600 674.100 ;
        RECT 364.950 661.950 367.050 664.050 ;
        RECT 373.950 661.950 376.050 664.050 ;
        RECT 379.950 661.950 382.050 664.050 ;
        RECT 361.950 658.950 364.050 661.050 ;
        RECT 362.400 652.050 363.600 658.950 ;
        RECT 365.400 655.050 366.600 661.950 ;
        RECT 367.950 655.950 370.050 658.050 ;
        RECT 364.950 652.950 367.050 655.050 ;
        RECT 368.400 652.050 369.600 655.950 ;
        RECT 352.950 649.950 355.050 652.050 ;
        RECT 361.950 649.950 364.050 652.050 ;
        RECT 367.950 651.600 370.050 652.050 ;
        RECT 365.400 650.400 370.050 651.600 ;
        RECT 353.400 645.600 354.600 649.950 ;
        RECT 365.400 649.050 366.600 650.400 ;
        RECT 367.950 649.950 370.050 650.400 ;
        RECT 374.400 649.050 375.600 661.950 ;
        RECT 395.400 661.050 396.600 766.950 ;
        RECT 403.950 761.100 406.050 763.200 ;
        RECT 404.400 760.050 405.600 761.100 ;
        RECT 400.950 757.950 403.050 760.050 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 406.950 757.950 409.050 760.050 ;
        RECT 401.400 757.050 402.600 757.950 ;
        RECT 397.950 755.400 402.600 757.050 ;
        RECT 407.400 756.900 408.600 757.950 ;
        RECT 397.950 754.950 402.000 755.400 ;
        RECT 406.950 754.800 409.050 756.900 ;
        RECT 409.950 754.950 412.050 757.050 ;
        RECT 400.950 732.600 405.000 733.050 ;
        RECT 400.950 730.950 405.600 732.600 ;
        RECT 404.400 727.050 405.600 730.950 ;
        RECT 410.400 730.050 411.600 754.950 ;
        RECT 413.400 732.600 414.600 775.950 ;
        RECT 416.400 757.050 417.600 781.950 ;
        RECT 425.400 766.050 426.600 799.950 ;
        RECT 427.800 799.800 429.900 801.900 ;
        RECT 430.950 798.600 433.050 802.050 ;
        RECT 437.400 801.000 438.600 802.950 ;
        RECT 443.400 802.050 444.600 829.950 ;
        RECT 449.400 828.600 450.600 839.100 ;
        RECT 452.400 829.050 453.600 853.950 ;
        RECT 457.950 840.000 460.050 844.050 ;
        RECT 476.400 841.200 477.600 877.800 ;
        RECT 478.950 871.950 481.050 874.050 ;
        RECT 458.400 838.050 459.600 840.000 ;
        RECT 475.950 839.100 478.050 841.200 ;
        RECT 479.400 838.050 480.600 871.950 ;
        RECT 485.400 871.050 486.600 911.400 ;
        RECT 493.950 910.950 496.050 913.050 ;
        RECT 503.400 892.050 504.600 913.950 ;
        RECT 509.400 907.050 510.600 913.950 ;
        RECT 518.400 907.050 519.600 917.100 ;
        RECT 524.400 916.050 525.600 917.100 ;
        RECT 523.950 913.950 526.050 916.050 ;
        RECT 526.950 913.950 529.050 916.050 ;
        RECT 508.950 904.950 511.050 907.050 ;
        RECT 517.950 904.950 520.050 907.050 ;
        RECT 523.950 895.950 526.050 898.050 ;
        RECT 490.950 889.950 493.050 892.050 ;
        RECT 502.950 889.950 505.050 892.050 ;
        RECT 484.950 868.950 487.050 871.050 ;
        RECT 491.400 868.050 492.600 889.950 ;
        RECT 499.950 884.100 502.050 886.200 ;
        RECT 505.950 884.100 508.050 886.200 ;
        RECT 517.950 884.100 520.050 886.200 ;
        RECT 500.400 883.050 501.600 884.100 ;
        RECT 506.400 883.050 507.600 884.100 ;
        RECT 518.400 883.050 519.600 884.100 ;
        RECT 524.400 883.050 525.600 895.950 ;
        RECT 527.400 889.050 528.600 913.950 ;
        RECT 532.950 898.950 535.050 901.050 ;
        RECT 526.950 886.950 529.050 889.050 ;
        RECT 496.950 880.950 499.050 883.050 ;
        RECT 499.950 880.950 502.050 883.050 ;
        RECT 502.950 880.950 505.050 883.050 ;
        RECT 505.950 880.950 508.050 883.050 ;
        RECT 508.950 880.950 511.050 883.050 ;
        RECT 517.950 880.950 520.050 883.050 ;
        RECT 520.950 880.950 523.050 883.050 ;
        RECT 523.950 880.950 526.050 883.050 ;
        RECT 526.950 880.950 529.050 883.050 ;
        RECT 497.400 879.900 498.600 880.950 ;
        RECT 503.400 879.900 504.600 880.950 ;
        RECT 496.950 877.800 499.050 879.900 ;
        RECT 502.950 877.800 505.050 879.900 ;
        RECT 502.950 874.650 505.050 876.750 ;
        RECT 490.950 865.950 493.050 868.050 ;
        RECT 499.950 859.950 502.050 862.050 ;
        RECT 500.400 841.200 501.600 859.950 ;
        RECT 503.400 850.050 504.600 874.650 ;
        RECT 509.400 874.050 510.600 880.950 ;
        RECT 508.950 871.950 511.050 874.050 ;
        RECT 511.950 868.950 514.050 871.050 ;
        RECT 505.950 856.950 508.050 859.050 ;
        RECT 502.950 847.950 505.050 850.050 ;
        RECT 490.950 838.950 493.050 841.050 ;
        RECT 499.950 839.100 502.050 841.200 ;
        RECT 457.950 835.950 460.050 838.050 ;
        RECT 460.950 835.950 463.050 838.050 ;
        RECT 478.950 835.950 481.050 838.050 ;
        RECT 481.950 835.950 484.050 838.050 ;
        RECT 446.400 827.400 450.600 828.600 ;
        RECT 446.400 808.050 447.600 827.400 ;
        RECT 451.950 826.950 454.050 829.050 ;
        RECT 457.950 826.950 460.050 829.050 ;
        RECT 448.950 817.950 451.050 820.050 ;
        RECT 454.950 817.950 457.050 820.050 ;
        RECT 445.950 805.950 448.050 808.050 ;
        RECT 449.400 805.050 450.600 817.950 ;
        RECT 455.400 808.050 456.600 817.950 ;
        RECT 454.950 805.950 457.050 808.050 ;
        RECT 448.950 802.950 451.050 805.050 ;
        RECT 451.950 802.950 454.050 805.050 ;
        RECT 430.950 798.000 435.600 798.600 ;
        RECT 431.400 797.400 435.600 798.000 ;
        RECT 430.950 790.950 433.050 793.050 ;
        RECT 424.950 763.950 427.050 766.050 ;
        RECT 421.950 761.100 424.050 763.200 ;
        RECT 422.400 760.050 423.600 761.100 ;
        RECT 431.400 760.050 432.600 790.950 ;
        RECT 434.400 790.050 435.600 797.400 ;
        RECT 436.950 796.950 439.050 801.000 ;
        RECT 442.950 799.950 445.050 802.050 ;
        RECT 445.950 799.950 448.050 802.050 ;
        RECT 433.950 787.950 436.050 790.050 ;
        RECT 439.950 787.950 442.050 790.050 ;
        RECT 436.950 778.950 439.050 781.050 ;
        RECT 421.950 757.950 424.050 760.050 ;
        RECT 424.950 757.950 427.050 760.050 ;
        RECT 430.950 757.950 433.050 760.050 ;
        RECT 415.950 754.950 418.050 757.050 ;
        RECT 421.950 751.950 424.050 754.050 ;
        RECT 418.950 733.950 421.050 736.050 ;
        RECT 413.400 731.400 417.600 732.600 ;
        RECT 409.950 727.950 412.050 730.050 ;
        RECT 412.950 727.950 415.050 730.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 403.950 724.950 406.050 727.050 ;
        RECT 406.950 724.950 409.050 727.050 ;
        RECT 401.400 723.900 402.600 724.950 ;
        RECT 407.400 723.900 408.600 724.950 ;
        RECT 400.950 721.800 403.050 723.900 ;
        RECT 406.950 721.800 409.050 723.900 ;
        RECT 409.950 721.950 412.050 724.050 ;
        RECT 413.400 723.900 414.600 727.950 ;
        RECT 403.950 697.950 406.050 700.050 ;
        RECT 397.950 688.950 400.050 691.050 ;
        RECT 398.400 667.050 399.600 688.950 ;
        RECT 404.400 682.050 405.600 697.950 ;
        RECT 410.400 697.050 411.600 721.950 ;
        RECT 412.950 721.800 415.050 723.900 ;
        RECT 409.950 694.950 412.050 697.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 397.950 664.950 400.050 667.050 ;
        RECT 403.950 664.950 406.050 667.050 ;
        RECT 394.950 658.950 397.050 661.050 ;
        RECT 382.500 654.300 384.600 656.400 ;
        RECT 386.400 654.900 387.600 657.450 ;
        RECT 380.400 649.050 381.600 651.600 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 373.950 646.950 376.050 649.050 ;
        RECT 379.950 646.950 382.050 649.050 ;
        RECT 382.950 648.900 383.850 654.300 ;
        RECT 385.800 652.800 387.900 654.900 ;
        RECT 389.700 651.900 391.800 653.700 ;
        RECT 384.750 650.700 393.300 651.900 ;
        RECT 384.750 649.800 386.850 650.700 ;
        RECT 382.950 647.700 389.700 648.900 ;
        RECT 353.400 644.400 357.600 645.600 ;
        RECT 356.400 634.050 357.600 644.400 ;
        RECT 355.950 631.950 358.050 634.050 ;
        RECT 343.950 610.950 346.050 613.050 ;
        RECT 349.950 610.950 352.050 613.050 ;
        RECT 344.400 604.050 345.600 610.950 ;
        RECT 349.950 606.600 352.050 607.200 ;
        RECT 352.950 606.600 355.050 610.050 ;
        RECT 349.950 606.000 355.050 606.600 ;
        RECT 349.950 605.400 354.600 606.000 ;
        RECT 349.950 605.100 352.050 605.400 ;
        RECT 350.400 604.050 351.600 605.100 ;
        RECT 337.950 601.950 340.050 604.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 343.950 601.950 346.050 604.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 334.950 586.950 337.050 589.050 ;
        RECT 331.950 574.950 334.050 577.050 ;
        RECT 335.400 574.050 336.600 586.950 ;
        RECT 341.400 583.050 342.600 601.950 ;
        RECT 347.400 597.600 348.600 601.950 ;
        RECT 352.950 598.950 355.050 601.050 ;
        RECT 349.950 597.600 352.050 598.050 ;
        RECT 347.400 596.400 352.050 597.600 ;
        RECT 349.950 595.950 352.050 596.400 ;
        RECT 340.950 580.950 343.050 583.050 ;
        RECT 337.950 574.950 340.050 577.050 ;
        RECT 328.950 571.950 331.050 574.050 ;
        RECT 334.950 571.950 337.050 574.050 ;
        RECT 322.950 568.950 325.050 571.050 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 323.400 567.000 324.600 568.950 ;
        RECT 332.400 567.900 333.600 568.950 ;
        RECT 328.800 567.000 330.900 567.900 ;
        RECT 319.950 562.950 322.050 565.050 ;
        RECT 322.950 562.950 325.050 567.000 ;
        RECT 328.800 565.800 331.050 567.000 ;
        RECT 331.950 565.800 334.050 567.900 ;
        RECT 328.950 565.050 331.050 565.800 ;
        RECT 328.950 564.750 333.000 565.050 ;
        RECT 328.950 564.000 334.050 564.750 ;
        RECT 329.400 563.400 334.050 564.000 ;
        RECT 330.000 562.950 334.050 563.400 ;
        RECT 313.800 556.950 315.900 559.050 ;
        RECT 316.950 556.950 319.050 559.050 ;
        RECT 304.950 526.950 307.050 529.050 ;
        RECT 307.950 526.950 310.050 529.050 ;
        RECT 283.950 523.800 286.050 525.900 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 292.950 523.950 295.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 274.950 514.950 277.050 517.050 ;
        RECT 280.950 514.950 283.050 517.050 ;
        RECT 275.400 496.050 276.600 514.950 ;
        RECT 284.400 508.050 285.600 523.800 ;
        RECT 293.400 522.900 294.600 523.950 ;
        RECT 292.950 520.800 295.050 522.900 ;
        RECT 289.950 511.950 292.050 514.050 ;
        RECT 283.950 505.950 286.050 508.050 ;
        RECT 280.950 502.950 283.050 505.050 ;
        RECT 274.950 493.950 277.050 496.050 ;
        RECT 281.400 493.050 282.600 502.950 ;
        RECT 286.950 494.100 289.050 496.200 ;
        RECT 290.400 496.050 291.600 511.950 ;
        RECT 299.400 508.050 300.600 523.950 ;
        RECT 305.400 514.050 306.600 526.950 ;
        RECT 314.400 526.050 315.600 556.950 ;
        RECT 320.400 556.050 321.600 562.950 ;
        RECT 331.950 562.650 334.050 562.950 ;
        RECT 319.950 553.950 322.050 556.050 ;
        RECT 322.950 547.950 325.050 550.050 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 307.950 517.950 310.050 523.050 ;
        RECT 304.950 511.950 307.050 514.050 ;
        RECT 301.950 508.950 304.050 511.050 ;
        RECT 298.950 505.950 301.050 508.050 ;
        RECT 302.400 505.050 303.600 508.950 ;
        RECT 301.950 502.950 304.050 505.050 ;
        RECT 301.950 499.800 304.050 501.900 ;
        RECT 302.400 496.200 303.600 499.800 ;
        RECT 308.400 499.050 309.600 517.950 ;
        RECT 311.400 511.050 312.600 523.950 ;
        RECT 317.400 522.000 318.600 523.950 ;
        RECT 316.950 517.950 319.050 522.000 ;
        RECT 319.950 520.950 322.050 523.050 ;
        RECT 320.400 517.050 321.600 520.950 ;
        RECT 319.950 514.950 322.050 517.050 ;
        RECT 310.950 508.950 313.050 511.050 ;
        RECT 323.400 499.050 324.600 547.950 ;
        RECT 328.950 535.950 331.050 538.050 ;
        RECT 329.400 526.050 330.600 535.950 ;
        RECT 338.400 531.600 339.600 574.950 ;
        RECT 341.400 568.050 342.600 580.950 ;
        RECT 350.400 574.050 351.600 595.950 ;
        RECT 353.400 574.200 354.600 598.950 ;
        RECT 356.400 598.050 357.600 631.950 ;
        RECT 359.400 610.050 360.600 646.950 ;
        RECT 361.950 643.950 364.050 646.050 ;
        RECT 358.950 607.950 361.050 610.050 ;
        RECT 362.400 606.600 363.600 643.950 ;
        RECT 374.400 640.050 375.600 646.950 ;
        RECT 376.950 640.950 379.050 643.050 ;
        RECT 373.950 637.950 376.050 640.050 ;
        RECT 364.950 619.950 367.050 622.050 ;
        RECT 359.400 605.400 363.600 606.600 ;
        RECT 355.950 595.950 358.050 598.050 ;
        RECT 349.800 571.950 351.900 574.050 ;
        RECT 352.950 572.100 355.050 574.200 ;
        RECT 353.400 571.050 354.600 572.100 ;
        RECT 346.950 568.950 349.050 571.050 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 340.950 565.950 343.050 568.050 ;
        RECT 347.400 567.900 348.600 568.950 ;
        RECT 341.400 538.050 342.600 565.950 ;
        RECT 346.800 565.800 348.900 567.900 ;
        RECT 349.950 565.950 352.050 568.050 ;
        RECT 350.400 562.050 351.600 565.950 ;
        RECT 355.950 562.950 358.050 565.050 ;
        RECT 343.950 559.950 346.050 562.050 ;
        RECT 349.950 559.950 352.050 562.050 ;
        RECT 340.950 535.950 343.050 538.050 ;
        RECT 338.400 530.400 342.600 531.600 ;
        RECT 334.950 527.100 337.050 529.200 ;
        RECT 335.400 526.050 336.600 527.100 ;
        RECT 341.400 526.050 342.600 530.400 ;
        RECT 344.400 529.050 345.600 559.950 ;
        RECT 346.950 556.950 349.050 559.050 ;
        RECT 343.950 526.950 346.050 529.050 ;
        RECT 328.950 523.950 331.050 526.050 ;
        RECT 331.950 523.950 334.050 526.050 ;
        RECT 334.950 523.950 337.050 526.050 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 332.400 519.600 333.600 523.950 ;
        RECT 338.400 522.000 339.600 523.950 ;
        RECT 332.400 518.400 336.600 519.600 ;
        RECT 335.400 513.600 336.600 518.400 ;
        RECT 337.950 514.950 340.050 522.000 ;
        RECT 343.950 520.950 346.050 523.050 ;
        RECT 340.950 513.600 343.050 514.050 ;
        RECT 344.400 513.600 345.600 520.950 ;
        RECT 335.400 512.400 345.600 513.600 ;
        RECT 340.950 511.950 343.050 512.400 ;
        RECT 331.950 508.950 334.050 511.050 ;
        RECT 337.950 508.950 340.050 511.050 ;
        RECT 328.950 499.950 331.050 502.050 ;
        RECT 307.950 496.950 310.050 499.050 ;
        RECT 322.950 496.950 325.050 499.050 ;
        RECT 287.400 493.050 288.600 494.100 ;
        RECT 289.950 493.950 292.050 496.050 ;
        RECT 292.950 494.100 295.050 496.200 ;
        RECT 301.950 494.100 304.050 496.200 ;
        RECT 319.950 494.100 322.050 496.200 ;
        RECT 277.950 490.950 280.050 493.050 ;
        RECT 280.950 490.950 283.050 493.050 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 286.950 490.950 289.050 493.050 ;
        RECT 274.950 487.950 277.050 490.050 ;
        RECT 271.950 451.950 274.050 454.050 ;
        RECT 271.950 448.800 274.050 450.900 ;
        RECT 238.950 445.950 241.050 448.050 ;
        RECT 241.950 445.950 244.050 448.050 ;
        RECT 244.950 445.950 247.050 448.050 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 265.950 445.950 268.050 448.050 ;
        RECT 235.950 442.950 238.050 445.050 ;
        RECT 232.950 439.950 235.050 442.050 ;
        RECT 232.950 430.950 235.050 433.050 ;
        RECT 233.400 424.050 234.600 430.950 ;
        RECT 232.950 421.950 235.050 424.050 ;
        RECT 230.400 419.400 234.600 420.600 ;
        RECT 215.400 415.050 216.600 416.100 ;
        RECT 221.400 415.050 222.600 417.000 ;
        RECT 229.950 415.950 232.050 418.050 ;
        RECT 211.950 412.950 214.050 415.050 ;
        RECT 214.950 412.950 217.050 415.050 ;
        RECT 217.950 412.950 220.050 415.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 212.400 403.050 213.600 412.950 ;
        RECT 218.400 406.050 219.600 412.950 ;
        RECT 224.400 411.900 225.600 412.950 ;
        RECT 230.400 412.050 231.600 415.950 ;
        RECT 223.950 409.800 226.050 411.900 ;
        RECT 229.950 409.950 232.050 412.050 ;
        RECT 229.950 406.800 232.050 408.900 ;
        RECT 217.950 403.950 220.050 406.050 ;
        RECT 211.950 400.950 214.050 403.050 ;
        RECT 208.950 385.950 211.050 388.050 ;
        RECT 205.950 382.950 208.050 385.050 ;
        RECT 179.400 370.050 180.600 372.000 ;
        RECT 181.950 370.950 184.050 373.050 ;
        RECT 184.950 370.950 187.050 373.050 ;
        RECT 187.950 370.950 190.050 376.050 ;
        RECT 196.950 371.100 199.050 373.200 ;
        RECT 202.950 372.000 205.050 376.050 ;
        RECT 197.400 370.050 198.600 371.100 ;
        RECT 203.400 370.050 204.600 372.000 ;
        RECT 175.950 367.950 178.050 370.050 ;
        RECT 178.950 367.950 181.050 370.050 ;
        RECT 163.950 358.950 166.050 361.050 ;
        RECT 169.950 358.950 172.050 361.050 ;
        RECT 164.400 355.050 165.600 358.950 ;
        RECT 166.950 355.950 169.050 358.050 ;
        RECT 172.950 355.950 175.050 358.050 ;
        RECT 160.800 352.950 162.900 355.050 ;
        RECT 163.950 352.950 166.050 355.050 ;
        RECT 151.950 338.100 154.050 340.200 ;
        RECT 157.950 338.100 160.050 340.200 ;
        RECT 152.400 337.050 153.600 338.100 ;
        RECT 158.400 337.050 159.600 338.100 ;
        RECT 151.950 334.950 154.050 337.050 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 145.950 331.950 148.050 334.050 ;
        RECT 155.400 333.000 156.600 334.950 ;
        RECT 154.950 328.950 157.050 333.000 ;
        RECT 155.400 310.050 156.600 328.950 ;
        RECT 161.400 328.050 162.600 334.950 ;
        RECT 160.950 325.950 163.050 328.050 ;
        RECT 167.400 325.050 168.600 355.950 ;
        RECT 173.400 348.600 174.600 355.950 ;
        RECT 176.400 349.050 177.600 367.950 ;
        RECT 184.950 367.800 187.050 369.900 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 199.950 367.950 202.050 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 185.400 358.050 186.600 367.800 ;
        RECT 194.400 367.050 195.600 367.950 ;
        RECT 190.950 365.400 195.600 367.050 ;
        RECT 200.400 366.900 201.600 367.950 ;
        RECT 190.950 364.950 195.000 365.400 ;
        RECT 199.950 364.800 202.050 366.900 ;
        RECT 205.950 364.950 208.050 367.050 ;
        RECT 206.400 361.050 207.600 364.950 ;
        RECT 205.950 358.950 208.050 361.050 ;
        RECT 184.950 355.950 187.050 358.050 ;
        RECT 199.950 349.950 202.050 352.050 ;
        RECT 170.400 347.400 174.600 348.600 ;
        RECT 170.400 340.050 171.600 347.400 ;
        RECT 175.950 346.950 178.050 349.050 ;
        RECT 190.950 346.950 193.050 349.050 ;
        RECT 172.950 345.600 175.050 346.050 ;
        RECT 178.950 345.600 181.050 346.050 ;
        RECT 172.950 344.400 181.050 345.600 ;
        RECT 172.950 343.950 175.050 344.400 ;
        RECT 178.950 343.950 181.050 344.400 ;
        RECT 169.950 337.950 172.050 340.050 ;
        RECT 175.950 338.100 178.050 340.200 ;
        RECT 181.950 338.100 184.050 340.200 ;
        RECT 176.400 337.050 177.600 338.100 ;
        RECT 182.400 337.050 183.600 338.100 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 175.950 334.950 178.050 337.050 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 173.400 328.050 174.600 334.950 ;
        RECT 172.950 325.950 175.050 328.050 ;
        RECT 179.400 325.050 180.600 334.950 ;
        RECT 185.400 333.900 186.600 334.950 ;
        RECT 191.400 333.900 192.600 346.950 ;
        RECT 200.400 340.200 201.600 349.950 ;
        RECT 199.950 338.100 202.050 340.200 ;
        RECT 200.400 337.050 201.600 338.100 ;
        RECT 206.400 337.050 207.600 358.950 ;
        RECT 209.400 352.050 210.600 385.950 ;
        RECT 211.950 376.950 214.050 379.050 ;
        RECT 208.950 349.950 211.050 352.050 ;
        RECT 212.400 349.050 213.600 376.950 ;
        RECT 214.950 373.950 217.050 376.050 ;
        RECT 211.950 346.950 214.050 349.050 ;
        RECT 215.400 343.050 216.600 373.950 ;
        RECT 223.950 372.000 226.050 376.050 ;
        RECT 224.400 370.050 225.600 372.000 ;
        RECT 230.400 370.050 231.600 406.800 ;
        RECT 233.400 388.050 234.600 419.400 ;
        RECT 236.400 418.050 237.600 442.950 ;
        RECT 239.400 424.050 240.600 445.950 ;
        RECT 245.400 444.000 246.600 445.950 ;
        RECT 244.950 439.950 247.050 444.000 ;
        RECT 253.950 442.950 256.050 445.050 ;
        RECT 250.950 433.950 253.050 436.050 ;
        RECT 244.950 430.950 247.050 433.050 ;
        RECT 241.950 427.950 244.050 430.050 ;
        RECT 238.950 421.950 241.050 424.050 ;
        RECT 238.950 420.600 241.050 420.900 ;
        RECT 242.400 420.600 243.600 427.950 ;
        RECT 245.400 424.050 246.600 430.950 ;
        RECT 247.950 424.950 250.050 427.050 ;
        RECT 244.950 421.950 247.050 424.050 ;
        RECT 238.950 419.400 243.600 420.600 ;
        RECT 238.950 418.800 241.050 419.400 ;
        RECT 235.950 415.950 238.050 418.050 ;
        RECT 239.400 415.050 240.600 418.800 ;
        RECT 238.950 412.950 241.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 235.950 408.600 238.050 412.050 ;
        RECT 242.400 411.900 243.600 412.950 ;
        RECT 241.950 409.800 244.050 411.900 ;
        RECT 244.950 409.950 247.050 412.050 ;
        RECT 235.950 408.000 240.600 408.600 ;
        RECT 236.400 407.400 240.600 408.000 ;
        RECT 232.950 385.950 235.050 388.050 ;
        RECT 235.950 382.950 238.050 385.050 ;
        RECT 220.950 367.950 223.050 370.050 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 226.950 367.950 229.050 370.050 ;
        RECT 229.950 367.950 232.050 370.050 ;
        RECT 221.400 355.050 222.600 367.950 ;
        RECT 227.400 366.000 228.600 367.950 ;
        RECT 226.950 361.950 229.050 366.000 ;
        RECT 220.950 352.950 223.050 355.050 ;
        RECT 232.950 352.950 235.050 355.050 ;
        RECT 217.950 349.950 220.050 352.050 ;
        RECT 214.950 340.950 217.050 343.050 ;
        RECT 218.400 339.600 219.600 349.950 ;
        RECT 215.400 338.400 219.600 339.600 ;
        RECT 223.950 339.000 226.050 343.050 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 197.400 333.900 198.600 334.950 ;
        RECT 184.950 331.800 187.050 333.900 ;
        RECT 190.950 331.800 193.050 333.900 ;
        RECT 196.950 331.800 199.050 333.900 ;
        RECT 191.400 325.050 192.600 331.800 ;
        RECT 197.400 328.050 198.600 331.800 ;
        RECT 196.950 325.950 199.050 328.050 ;
        RECT 166.950 322.950 169.050 325.050 ;
        RECT 178.950 322.950 181.050 325.050 ;
        RECT 190.950 322.950 193.050 325.050 ;
        RECT 196.950 316.950 199.050 319.050 ;
        RECT 154.950 307.950 157.050 310.050 ;
        RECT 148.950 298.950 151.050 301.050 ;
        RECT 142.950 293.100 145.050 295.200 ;
        RECT 149.400 292.050 150.600 298.950 ;
        RECT 197.400 298.050 198.600 316.950 ;
        RECT 203.400 307.050 204.600 334.950 ;
        RECT 205.950 328.950 208.050 331.050 ;
        RECT 202.950 304.950 205.050 307.050 ;
        RECT 154.950 293.100 157.050 298.050 ;
        RECT 160.950 295.950 163.050 298.050 ;
        RECT 155.400 292.050 156.600 293.100 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 146.400 288.900 147.600 289.950 ;
        RECT 152.400 288.900 153.600 289.950 ;
        RECT 145.950 286.800 148.050 288.900 ;
        RECT 151.950 286.800 154.050 288.900 ;
        RECT 152.400 285.600 153.600 286.800 ;
        RECT 149.400 284.400 153.600 285.600 ;
        RECT 142.950 268.950 145.050 271.050 ;
        RECT 139.950 259.950 142.050 262.050 ;
        RECT 143.400 259.050 144.600 268.950 ;
        RECT 149.400 262.200 150.600 284.400 ;
        RECT 161.400 283.050 162.600 295.950 ;
        RECT 166.950 293.100 169.050 295.200 ;
        RECT 172.950 294.000 175.050 298.050 ;
        RECT 196.950 295.950 199.050 298.050 ;
        RECT 167.400 292.050 168.600 293.100 ;
        RECT 173.400 292.050 174.600 294.000 ;
        RECT 184.950 293.100 187.050 295.200 ;
        RECT 190.950 293.100 193.050 295.200 ;
        RECT 166.950 289.950 169.050 292.050 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 170.400 285.600 171.600 289.950 ;
        RECT 176.400 288.900 177.600 289.950 ;
        RECT 175.950 286.800 178.050 288.900 ;
        RECT 170.400 284.400 174.600 285.600 ;
        RECT 160.950 280.950 163.050 283.050 ;
        RECT 169.950 280.950 172.050 283.050 ;
        RECT 160.950 271.950 163.050 274.050 ;
        RECT 148.950 260.100 151.050 262.200 ;
        RECT 149.400 259.050 150.600 260.100 ;
        RECT 161.400 259.050 162.600 271.950 ;
        RECT 142.950 256.950 145.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 160.950 256.950 163.050 259.050 ;
        RECT 163.950 256.950 166.050 259.050 ;
        RECT 146.400 255.900 147.600 256.950 ;
        RECT 145.950 253.800 148.050 255.900 ;
        RECT 152.400 255.000 153.600 256.950 ;
        RECT 164.400 255.900 165.600 256.950 ;
        RECT 151.950 250.950 154.050 255.000 ;
        RECT 163.950 253.800 166.050 255.900 ;
        RECT 170.400 253.050 171.600 280.950 ;
        RECT 173.400 270.600 174.600 284.400 ;
        RECT 185.400 273.600 186.600 293.100 ;
        RECT 191.400 292.050 192.600 293.100 ;
        RECT 197.400 292.050 198.600 295.950 ;
        RECT 203.400 295.050 204.600 304.950 ;
        RECT 202.950 292.950 205.050 295.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 199.950 289.950 202.050 292.050 ;
        RECT 187.950 273.600 190.050 274.050 ;
        RECT 185.400 272.400 190.050 273.600 ;
        RECT 187.950 271.950 190.050 272.400 ;
        RECT 173.400 269.400 177.600 270.600 ;
        RECT 172.950 265.950 175.050 268.050 ;
        RECT 169.950 250.950 172.050 253.050 ;
        RECT 148.950 238.950 151.050 241.050 ;
        RECT 154.950 238.950 157.050 241.050 ;
        RECT 149.400 235.050 150.600 238.950 ;
        RECT 148.950 232.950 151.050 235.050 ;
        RECT 136.950 220.950 139.050 223.050 ;
        RECT 142.950 216.000 145.050 220.050 ;
        RECT 143.400 214.050 144.600 216.000 ;
        RECT 149.400 214.050 150.600 232.950 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 142.950 211.950 145.050 214.050 ;
        RECT 145.950 211.950 148.050 214.050 ;
        RECT 148.950 211.950 151.050 214.050 ;
        RECT 131.400 206.400 135.600 207.600 ;
        RECT 118.950 202.950 121.050 205.050 ;
        RECT 127.950 193.950 130.050 196.050 ;
        RECT 106.950 190.950 109.050 193.050 ;
        RECT 112.950 190.950 115.050 193.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 92.400 177.900 93.600 178.950 ;
        RECT 98.400 177.900 99.600 178.950 ;
        RECT 107.400 177.900 108.600 190.950 ;
        RECT 121.950 187.950 124.050 190.050 ;
        RECT 109.950 181.950 112.050 184.050 ;
        RECT 115.950 182.100 118.050 184.200 ;
        RECT 91.950 175.800 94.050 177.900 ;
        RECT 97.950 175.800 100.050 177.900 ;
        RECT 106.950 175.800 109.050 177.900 ;
        RECT 85.950 172.950 88.050 175.050 ;
        RECT 91.950 172.650 94.050 174.750 ;
        RECT 82.950 169.950 85.050 172.050 ;
        RECT 83.400 136.050 84.600 169.950 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 80.400 132.900 81.600 133.950 ;
        RECT 86.400 132.900 87.600 133.950 ;
        RECT 70.950 130.800 73.050 132.900 ;
        RECT 79.950 130.800 82.050 132.900 ;
        RECT 85.950 130.800 88.050 132.900 ;
        RECT 92.400 127.050 93.600 172.650 ;
        RECT 97.950 169.950 100.050 172.050 ;
        RECT 94.950 139.950 97.050 142.050 ;
        RECT 64.950 124.950 67.050 127.050 ;
        RECT 91.950 124.950 94.050 127.050 ;
        RECT 77.400 116.400 84.600 117.600 ;
        RECT 58.950 112.950 61.050 115.050 ;
        RECT 50.400 104.400 54.600 105.600 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 43.950 100.950 46.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 41.400 88.050 42.600 100.950 ;
        RECT 47.400 99.900 48.600 100.950 ;
        RECT 53.400 99.900 54.600 104.400 ;
        RECT 58.950 104.100 61.050 106.200 ;
        RECT 64.950 104.100 67.050 106.200 ;
        RECT 59.400 103.050 60.600 104.100 ;
        RECT 65.400 103.050 66.600 104.100 ;
        RECT 73.950 103.950 76.050 106.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 46.950 97.800 49.050 99.900 ;
        RECT 52.950 97.800 55.050 99.900 ;
        RECT 62.400 99.000 63.600 100.950 ;
        RECT 53.400 94.050 54.600 97.800 ;
        RECT 61.950 94.950 64.050 99.000 ;
        RECT 68.400 94.050 69.600 100.950 ;
        RECT 52.950 91.950 55.050 94.050 ;
        RECT 67.950 91.950 70.050 94.050 ;
        RECT 40.950 85.950 43.050 88.050 ;
        RECT 61.950 73.950 64.050 76.050 ;
        RECT 37.950 70.950 40.050 73.050 ;
        RECT 31.950 61.950 34.050 64.050 ;
        RECT 28.950 60.600 31.050 61.050 ;
        RECT 23.400 58.050 24.600 60.000 ;
        RECT 28.950 59.400 33.600 60.600 ;
        RECT 28.950 58.950 31.050 59.400 ;
        RECT 32.400 58.050 33.600 59.400 ;
        RECT 38.400 58.050 39.600 70.950 ;
        RECT 46.950 61.950 49.050 64.050 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 31.950 55.950 34.050 58.050 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 14.400 43.050 15.600 55.950 ;
        RECT 20.400 54.900 21.600 55.950 ;
        RECT 19.950 52.800 22.050 54.900 ;
        RECT 35.400 49.050 36.600 55.950 ;
        RECT 34.950 46.950 37.050 49.050 ;
        RECT 13.950 40.950 16.050 43.050 ;
        RECT 19.950 40.950 22.050 43.050 ;
        RECT 1.950 34.950 4.050 37.050 ;
        RECT 13.950 34.950 16.050 37.050 ;
        RECT 14.400 25.050 15.600 34.950 ;
        RECT 20.400 25.050 21.600 40.950 ;
        RECT 41.400 37.050 42.600 55.950 ;
        RECT 47.400 49.050 48.600 61.950 ;
        RECT 62.400 58.050 63.600 73.950 ;
        RECT 74.400 67.050 75.600 103.950 ;
        RECT 67.950 60.000 70.050 64.050 ;
        RECT 73.950 61.950 76.050 67.050 ;
        RECT 77.400 61.200 78.600 116.400 ;
        RECT 79.950 112.950 82.050 115.050 ;
        RECT 80.400 106.050 81.600 112.950 ;
        RECT 83.400 112.050 84.600 116.400 ;
        RECT 85.950 115.950 88.050 118.050 ;
        RECT 82.950 109.950 85.050 112.050 ;
        RECT 79.950 103.950 82.050 106.050 ;
        RECT 86.400 103.050 87.600 115.950 ;
        RECT 91.950 109.950 94.050 112.050 ;
        RECT 92.400 103.050 93.600 109.950 ;
        RECT 95.400 106.050 96.600 139.950 ;
        RECT 94.950 103.950 97.050 106.050 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 83.400 99.900 84.600 100.950 ;
        RECT 82.950 97.800 85.050 99.900 ;
        RECT 89.400 99.000 90.600 100.950 ;
        RECT 88.950 94.950 91.050 99.000 ;
        RECT 89.400 88.050 90.600 94.950 ;
        RECT 88.950 85.950 91.050 88.050 ;
        RECT 82.950 73.950 85.050 76.050 ;
        RECT 68.400 58.050 69.600 60.000 ;
        RECT 76.950 59.100 79.050 61.200 ;
        RECT 77.400 58.050 78.600 59.100 ;
        RECT 83.400 58.050 84.600 73.950 ;
        RECT 91.950 64.950 94.050 67.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 59.400 49.050 60.600 55.950 ;
        RECT 65.400 54.900 66.600 55.950 ;
        RECT 64.950 52.800 67.050 54.900 ;
        RECT 46.950 46.950 49.050 49.050 ;
        RECT 58.950 46.950 61.050 49.050 ;
        RECT 40.950 34.950 43.050 37.050 ;
        RECT 37.950 31.950 40.050 34.050 ;
        RECT 38.400 25.050 39.600 31.950 ;
        RECT 41.400 28.050 42.600 34.950 ;
        RECT 59.400 31.050 60.600 46.950 ;
        RECT 80.400 46.050 81.600 55.950 ;
        RECT 86.400 54.900 87.600 55.950 ;
        RECT 85.950 52.800 88.050 54.900 ;
        RECT 79.950 43.950 82.050 46.050 ;
        RECT 73.950 40.950 76.050 43.050 ;
        RECT 61.950 34.950 64.050 37.050 ;
        RECT 58.950 28.950 61.050 31.050 ;
        RECT 62.400 28.200 63.600 34.950 ;
        RECT 40.950 25.950 43.050 28.050 ;
        RECT 46.950 25.950 49.050 28.050 ;
        RECT 55.950 26.100 58.050 28.200 ;
        RECT 61.950 26.100 64.050 28.200 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 22.950 22.950 25.050 25.050 ;
        RECT 34.950 22.950 37.050 25.050 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 17.400 21.900 18.600 22.950 ;
        RECT 23.400 21.900 24.600 22.950 ;
        RECT 35.400 21.900 36.600 22.950 ;
        RECT 16.950 19.800 19.050 21.900 ;
        RECT 22.950 19.800 25.050 21.900 ;
        RECT 34.950 19.800 37.050 21.900 ;
        RECT 47.400 10.050 48.600 25.950 ;
        RECT 56.400 25.050 57.600 26.100 ;
        RECT 62.400 25.050 63.600 26.100 ;
        RECT 74.400 25.050 75.600 40.950 ;
        RECT 79.950 37.950 82.050 40.050 ;
        RECT 80.400 25.050 81.600 37.950 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 76.950 22.950 79.050 25.050 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 53.400 21.900 54.600 22.950 ;
        RECT 59.400 21.900 60.600 22.950 ;
        RECT 52.950 16.950 55.050 21.900 ;
        RECT 58.950 19.800 61.050 21.900 ;
        RECT 71.400 21.000 72.600 22.950 ;
        RECT 77.400 21.000 78.600 22.950 ;
        RECT 70.950 16.950 73.050 21.000 ;
        RECT 76.950 16.950 79.050 21.000 ;
        RECT 86.400 19.050 87.600 52.800 ;
        RECT 92.400 46.050 93.600 64.950 ;
        RECT 94.950 59.100 97.050 61.200 ;
        RECT 95.400 55.050 96.600 59.100 ;
        RECT 94.950 52.950 97.050 55.050 ;
        RECT 98.400 52.050 99.600 169.950 ;
        RECT 103.950 137.100 106.050 139.200 ;
        RECT 104.400 136.050 105.600 137.100 ;
        RECT 110.400 136.050 111.600 181.950 ;
        RECT 116.400 181.050 117.600 182.100 ;
        RECT 122.400 181.050 123.600 187.950 ;
        RECT 128.400 184.050 129.600 193.950 ;
        RECT 127.950 181.950 130.050 184.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 119.400 177.900 120.600 178.950 ;
        RECT 125.400 177.900 126.600 178.950 ;
        RECT 118.950 175.800 121.050 177.900 ;
        RECT 124.950 175.800 127.050 177.900 ;
        RECT 125.400 163.050 126.600 175.800 ;
        RECT 131.400 172.050 132.600 206.400 ;
        RECT 140.400 205.050 141.600 211.950 ;
        RECT 142.950 205.950 145.050 208.050 ;
        RECT 139.950 202.950 142.050 205.050 ;
        RECT 136.950 182.100 139.050 184.200 ;
        RECT 137.400 181.050 138.600 182.100 ;
        RECT 143.400 181.050 144.600 205.950 ;
        RECT 146.400 190.050 147.600 211.950 ;
        RECT 151.950 199.950 154.050 202.050 ;
        RECT 145.950 187.950 148.050 190.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 142.950 178.950 145.050 181.050 ;
        RECT 145.950 178.950 148.050 181.050 ;
        RECT 140.400 177.000 141.600 178.950 ;
        RECT 139.950 172.950 142.050 177.000 ;
        RECT 130.950 169.950 133.050 172.050 ;
        RECT 124.950 160.950 127.050 163.050 ;
        RECT 115.950 142.950 118.050 145.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 107.400 115.050 108.600 133.950 ;
        RECT 116.400 133.050 117.600 142.950 ;
        RECT 127.950 138.000 130.050 142.050 ;
        RECT 128.400 136.050 129.600 138.000 ;
        RECT 133.950 137.100 136.050 139.200 ;
        RECT 134.400 136.050 135.600 137.100 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 115.950 130.950 118.050 133.050 ;
        RECT 125.400 132.900 126.600 133.950 ;
        RECT 124.950 130.800 127.050 132.900 ;
        RECT 131.400 127.050 132.600 133.950 ;
        RECT 140.400 132.900 141.600 172.950 ;
        RECT 146.400 157.050 147.600 178.950 ;
        RECT 148.950 175.950 151.050 178.050 ;
        RECT 145.950 156.600 148.050 157.050 ;
        RECT 143.400 155.400 148.050 156.600 ;
        RECT 139.950 130.800 142.050 132.900 ;
        RECT 121.950 124.950 124.050 127.050 ;
        RECT 130.950 124.950 133.050 127.050 ;
        RECT 118.950 115.950 121.050 118.050 ;
        RECT 106.950 112.950 109.050 115.050 ;
        RECT 112.950 109.950 115.050 112.050 ;
        RECT 100.950 103.950 103.050 106.050 ;
        RECT 101.400 97.050 102.600 103.950 ;
        RECT 113.400 103.050 114.600 109.950 ;
        RECT 119.400 103.050 120.600 115.950 ;
        RECT 122.400 106.050 123.600 124.950 ;
        RECT 140.400 118.050 141.600 130.800 ;
        RECT 143.400 130.050 144.600 155.400 ;
        RECT 145.950 154.950 148.050 155.400 ;
        RECT 149.400 151.050 150.600 175.950 ;
        RECT 152.400 175.050 153.600 199.950 ;
        RECT 155.400 196.050 156.600 238.950 ;
        RECT 160.950 226.950 163.050 229.050 ;
        RECT 157.950 220.950 160.050 223.050 ;
        RECT 158.400 208.050 159.600 220.950 ;
        RECT 157.950 205.950 160.050 208.050 ;
        RECT 161.400 199.050 162.600 226.950 ;
        RECT 173.400 223.050 174.600 265.950 ;
        RECT 176.400 229.050 177.600 269.400 ;
        RECT 181.950 265.950 184.050 268.050 ;
        RECT 182.400 259.050 183.600 265.950 ;
        RECT 188.400 259.050 189.600 271.950 ;
        RECT 194.400 262.050 195.600 289.950 ;
        RECT 200.400 288.900 201.600 289.950 ;
        RECT 199.950 286.800 202.050 288.900 ;
        RECT 206.400 283.050 207.600 328.950 ;
        RECT 209.400 325.050 210.600 334.950 ;
        RECT 215.400 331.050 216.600 338.400 ;
        RECT 224.400 337.050 225.600 339.000 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 221.400 333.900 222.600 334.950 ;
        RECT 227.400 333.900 228.600 334.950 ;
        RECT 233.400 334.050 234.600 352.950 ;
        RECT 220.950 331.800 223.050 333.900 ;
        RECT 226.800 331.800 228.900 333.900 ;
        RECT 229.950 331.950 232.050 334.050 ;
        RECT 232.950 331.950 235.050 334.050 ;
        RECT 214.950 328.950 217.050 331.050 ;
        RECT 208.950 322.950 211.050 325.050 ;
        RECT 211.950 307.950 214.050 310.050 ;
        RECT 212.400 292.050 213.600 307.950 ;
        RECT 217.950 304.950 220.050 307.050 ;
        RECT 218.400 292.050 219.600 304.950 ;
        RECT 221.400 301.050 222.600 331.800 ;
        RECT 230.400 322.050 231.600 331.950 ;
        RECT 229.950 319.950 232.050 322.050 ;
        RECT 236.400 310.050 237.600 382.950 ;
        RECT 239.400 382.050 240.600 407.400 ;
        RECT 245.400 397.050 246.600 409.950 ;
        RECT 248.400 406.050 249.600 424.950 ;
        RECT 251.400 409.050 252.600 433.950 ;
        RECT 254.400 412.050 255.600 442.950 ;
        RECT 256.950 439.950 259.050 442.050 ;
        RECT 257.400 424.050 258.600 439.950 ;
        RECT 260.400 439.050 261.600 445.950 ;
        RECT 259.950 436.950 262.050 439.050 ;
        RECT 256.950 421.950 259.050 424.050 ;
        RECT 266.400 421.050 267.600 445.950 ;
        RECT 272.400 442.050 273.600 448.800 ;
        RECT 271.950 439.950 274.050 442.050 ;
        RECT 275.400 436.050 276.600 487.950 ;
        RECT 278.400 472.050 279.600 490.950 ;
        RECT 284.400 489.900 285.600 490.950 ;
        RECT 283.950 487.800 286.050 489.900 ;
        RECT 289.950 487.950 292.050 490.050 ;
        RECT 293.400 489.600 294.600 494.100 ;
        RECT 302.400 493.050 303.600 494.100 ;
        RECT 320.400 493.050 321.600 494.100 ;
        RECT 298.950 490.950 301.050 493.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 307.950 490.950 310.050 493.050 ;
        RECT 316.950 490.950 319.050 493.050 ;
        RECT 319.950 490.950 322.050 493.050 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 299.400 489.900 300.600 490.950 ;
        RECT 293.400 488.400 297.600 489.600 ;
        RECT 277.950 469.950 280.050 472.050 ;
        RECT 277.950 463.950 280.050 466.050 ;
        RECT 286.950 463.950 289.050 466.050 ;
        RECT 278.400 451.050 279.600 463.950 ;
        RECT 283.950 454.950 286.050 457.050 ;
        RECT 277.950 448.950 280.050 451.050 ;
        RECT 284.400 448.050 285.600 454.950 ;
        RECT 287.400 454.050 288.600 463.950 ;
        RECT 290.400 457.050 291.600 487.950 ;
        RECT 292.950 466.950 295.050 469.050 ;
        RECT 289.950 454.950 292.050 457.050 ;
        RECT 287.400 453.900 291.000 454.050 ;
        RECT 287.400 452.250 292.050 453.900 ;
        RECT 288.000 451.950 292.050 452.250 ;
        RECT 289.950 451.800 292.050 451.950 ;
        RECT 293.400 451.050 294.600 466.950 ;
        RECT 289.950 448.950 292.050 451.050 ;
        RECT 292.950 448.950 295.050 451.050 ;
        RECT 290.400 448.050 291.600 448.950 ;
        RECT 280.950 445.950 283.050 448.050 ;
        RECT 283.950 445.950 286.050 448.050 ;
        RECT 286.950 445.950 289.050 448.050 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 274.950 433.950 277.050 436.050 ;
        RECT 281.400 433.050 282.600 445.950 ;
        RECT 287.400 444.900 288.600 445.950 ;
        RECT 286.950 442.800 289.050 444.900 ;
        RECT 296.400 444.600 297.600 488.400 ;
        RECT 298.950 487.800 301.050 489.900 ;
        RECT 308.400 489.000 309.600 490.950 ;
        RECT 301.950 484.950 304.050 487.050 ;
        RECT 307.950 484.950 310.050 489.000 ;
        RECT 310.950 486.600 313.050 490.050 ;
        RECT 317.400 487.050 318.600 490.950 ;
        RECT 310.950 486.000 315.600 486.600 ;
        RECT 311.400 485.400 315.600 486.000 ;
        RECT 317.400 485.400 322.050 487.050 ;
        RECT 302.400 475.050 303.600 484.950 ;
        RECT 310.950 481.950 313.050 484.050 ;
        RECT 307.950 478.950 310.050 481.050 ;
        RECT 301.950 472.950 304.050 475.050 ;
        RECT 298.950 454.950 301.050 457.050 ;
        RECT 293.400 443.400 297.600 444.600 ;
        RECT 293.400 442.050 294.600 443.400 ;
        RECT 292.950 439.950 295.050 442.050 ;
        RECT 295.950 439.950 298.050 442.050 ;
        RECT 280.950 430.950 283.050 433.050 ;
        RECT 266.400 419.400 271.050 421.050 ;
        RECT 267.000 418.950 271.050 419.400 ;
        RECT 256.950 417.600 261.000 418.050 ;
        RECT 256.950 415.950 261.600 417.600 ;
        RECT 265.950 416.100 268.050 418.200 ;
        RECT 274.950 416.100 277.050 418.200 ;
        RECT 286.950 417.000 289.050 421.050 ;
        RECT 260.400 415.050 261.600 415.950 ;
        RECT 266.400 415.050 267.600 416.100 ;
        RECT 259.950 412.950 262.050 415.050 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 263.400 411.900 264.600 412.950 ;
        RECT 269.400 411.900 270.600 412.950 ;
        RECT 250.950 406.950 253.050 409.050 ;
        RECT 259.800 406.950 261.900 409.050 ;
        RECT 262.950 406.950 265.050 411.900 ;
        RECT 268.950 409.800 271.050 411.900 ;
        RECT 247.950 403.950 250.050 406.050 ;
        RECT 244.950 394.950 247.050 397.050 ;
        RECT 253.950 388.950 256.050 391.050 ;
        RECT 247.950 385.950 250.050 388.050 ;
        RECT 238.950 379.950 241.050 382.050 ;
        RECT 241.950 371.100 244.050 373.200 ;
        RECT 242.400 370.050 243.600 371.100 ;
        RECT 248.400 370.050 249.600 385.950 ;
        RECT 254.400 373.200 255.600 388.950 ;
        RECT 256.950 373.950 259.050 376.050 ;
        RECT 253.950 371.100 256.050 373.200 ;
        RECT 241.950 367.950 244.050 370.050 ;
        RECT 244.950 367.950 247.050 370.050 ;
        RECT 247.950 367.950 250.050 370.050 ;
        RECT 250.950 367.950 253.050 370.050 ;
        RECT 245.400 366.000 246.600 367.950 ;
        RECT 244.950 361.950 247.050 366.000 ;
        RECT 251.400 358.050 252.600 367.950 ;
        RECT 253.950 364.950 256.050 367.050 ;
        RECT 238.950 355.950 241.050 358.050 ;
        RECT 250.950 355.950 253.050 358.050 ;
        RECT 239.400 325.050 240.600 355.950 ;
        RECT 254.400 352.050 255.600 364.950 ;
        RECT 257.400 364.050 258.600 373.950 ;
        RECT 256.950 361.950 259.050 364.050 ;
        RECT 260.400 361.050 261.600 406.950 ;
        RECT 275.400 406.050 276.600 416.100 ;
        RECT 287.400 415.050 288.600 417.000 ;
        RECT 277.950 412.950 280.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 412.950 289.050 415.050 ;
        RECT 274.950 403.950 277.050 406.050 ;
        RECT 278.400 400.050 279.600 412.950 ;
        RECT 280.950 406.950 283.050 409.050 ;
        RECT 277.950 397.950 280.050 400.050 ;
        RECT 271.950 390.600 274.050 391.050 ;
        RECT 277.950 390.600 280.050 391.050 ;
        RECT 271.950 389.400 280.050 390.600 ;
        RECT 271.950 388.950 274.050 389.400 ;
        RECT 277.950 388.950 280.050 389.400 ;
        RECT 268.950 387.600 271.050 388.050 ;
        RECT 268.950 386.400 276.600 387.600 ;
        RECT 268.950 385.950 271.050 386.400 ;
        RECT 271.950 382.950 274.050 385.050 ;
        RECT 262.950 379.950 265.050 382.050 ;
        RECT 263.400 373.050 264.600 379.950 ;
        RECT 272.400 379.050 273.600 382.950 ;
        RECT 275.400 382.050 276.600 386.400 ;
        RECT 274.950 379.950 277.050 382.050 ;
        RECT 271.950 376.950 274.050 379.050 ;
        RECT 262.950 370.950 265.050 373.050 ;
        RECT 265.950 372.000 268.050 376.050 ;
        RECT 266.400 370.050 267.600 372.000 ;
        RECT 271.950 371.100 274.050 373.200 ;
        RECT 272.400 370.050 273.600 371.100 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 274.950 367.950 277.050 370.050 ;
        RECT 262.950 364.800 265.050 366.900 ;
        RECT 269.400 366.000 270.600 367.950 ;
        RECT 275.400 366.900 276.600 367.950 ;
        RECT 259.950 358.950 262.050 361.050 ;
        RECT 259.950 355.800 262.050 357.900 ;
        RECT 247.950 349.950 250.050 352.050 ;
        RECT 253.950 349.950 256.050 352.050 ;
        RECT 248.400 346.050 249.600 349.950 ;
        RECT 253.950 346.800 256.050 348.900 ;
        RECT 247.950 343.950 250.050 346.050 ;
        RECT 250.950 343.950 253.050 346.050 ;
        RECT 244.950 339.000 247.050 343.050 ;
        RECT 245.400 337.050 246.600 339.000 ;
        RECT 251.400 337.050 252.600 343.950 ;
        RECT 254.400 340.050 255.600 346.800 ;
        RECT 260.400 346.050 261.600 355.800 ;
        RECT 263.400 346.050 264.600 364.800 ;
        RECT 268.950 361.950 271.050 366.000 ;
        RECT 274.950 364.800 277.050 366.900 ;
        RECT 281.400 361.050 282.600 406.950 ;
        RECT 284.400 406.050 285.600 412.950 ;
        RECT 283.950 403.950 286.050 406.050 ;
        RECT 283.950 397.950 286.050 400.050 ;
        RECT 284.400 373.050 285.600 397.950 ;
        RECT 286.950 388.950 289.050 391.050 ;
        RECT 287.400 373.200 288.600 388.950 ;
        RECT 293.400 382.050 294.600 439.950 ;
        RECT 296.400 418.050 297.600 439.950 ;
        RECT 299.400 421.050 300.600 454.950 ;
        RECT 302.400 451.050 303.600 472.950 ;
        RECT 304.950 451.950 307.050 457.050 ;
        RECT 301.950 448.950 304.050 451.050 ;
        RECT 308.400 448.050 309.600 478.950 ;
        RECT 311.400 460.050 312.600 481.950 ;
        RECT 314.400 466.050 315.600 485.400 ;
        RECT 318.000 484.950 322.050 485.400 ;
        RECT 316.950 478.950 319.050 481.050 ;
        RECT 313.950 463.950 316.050 466.050 ;
        RECT 310.950 457.950 313.050 460.050 ;
        RECT 317.400 451.050 318.600 478.950 ;
        RECT 323.400 475.050 324.600 490.950 ;
        RECT 325.950 487.950 328.050 490.050 ;
        RECT 326.400 478.050 327.600 487.950 ;
        RECT 329.400 487.050 330.600 499.950 ;
        RECT 328.950 484.950 331.050 487.050 ;
        RECT 325.950 475.950 328.050 478.050 ;
        RECT 322.950 472.950 325.050 475.050 ;
        RECT 332.400 469.050 333.600 508.950 ;
        RECT 338.400 505.050 339.600 508.950 ;
        RECT 347.400 508.050 348.600 556.950 ;
        RECT 349.950 553.950 352.050 556.050 ;
        RECT 346.950 505.950 349.050 508.050 ;
        RECT 337.950 502.950 340.050 505.050 ;
        RECT 350.400 502.050 351.600 553.950 ;
        RECT 356.400 547.050 357.600 562.950 ;
        RECT 359.400 562.050 360.600 605.400 ;
        RECT 365.400 604.050 366.600 619.950 ;
        RECT 370.950 613.950 373.050 616.050 ;
        RECT 371.400 610.050 372.600 613.950 ;
        RECT 370.950 606.000 373.050 610.050 ;
        RECT 371.400 604.050 372.600 606.000 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 368.400 574.050 369.600 601.950 ;
        RECT 377.400 577.050 378.600 640.950 ;
        RECT 382.950 640.500 384.000 647.700 ;
        RECT 385.800 644.100 387.900 646.200 ;
        RECT 388.800 645.300 389.700 647.700 ;
        RECT 386.400 641.550 387.600 644.100 ;
        RECT 388.800 643.200 390.900 645.300 ;
        RECT 392.400 641.700 393.300 650.700 ;
        RECT 394.500 646.950 396.600 649.050 ;
        RECT 395.400 644.400 396.600 646.950 ;
        RECT 398.400 643.050 399.600 664.950 ;
        RECT 400.950 658.950 403.050 661.050 ;
        RECT 401.400 652.050 402.600 658.950 ;
        RECT 404.400 655.050 405.600 664.950 ;
        RECT 410.400 664.050 411.600 679.950 ;
        RECT 412.950 676.950 415.050 679.050 ;
        RECT 409.950 661.950 412.050 664.050 ;
        RECT 406.950 658.950 409.050 661.050 ;
        RECT 403.950 652.950 406.050 655.050 ;
        RECT 400.950 649.950 403.050 652.050 ;
        RECT 407.400 649.050 408.600 658.950 ;
        RECT 410.400 658.050 411.600 661.950 ;
        RECT 409.950 655.950 412.050 658.050 ;
        RECT 413.400 654.600 414.600 676.950 ;
        RECT 416.400 661.050 417.600 731.400 ;
        RECT 419.400 724.050 420.600 733.950 ;
        RECT 422.400 730.050 423.600 751.950 ;
        RECT 425.400 745.050 426.600 757.950 ;
        RECT 437.400 757.050 438.600 778.950 ;
        RECT 436.950 754.950 439.050 757.050 ;
        RECT 440.400 756.600 441.600 787.950 ;
        RECT 446.400 778.050 447.600 799.950 ;
        RECT 452.400 787.050 453.600 802.950 ;
        RECT 454.950 799.950 457.050 802.050 ;
        RECT 451.950 784.950 454.050 787.050 ;
        RECT 455.400 780.600 456.600 799.950 ;
        RECT 458.400 784.050 459.600 826.950 ;
        RECT 461.400 820.050 462.600 835.950 ;
        RECT 482.400 834.900 483.600 835.950 ;
        RECT 481.950 832.800 484.050 834.900 ;
        RECT 475.950 823.950 478.050 826.050 ;
        RECT 460.950 817.950 463.050 820.050 ;
        RECT 476.400 811.050 477.600 823.950 ;
        RECT 491.400 817.050 492.600 838.950 ;
        RECT 500.400 838.050 501.600 839.100 ;
        RECT 506.400 838.050 507.600 856.950 ;
        RECT 496.950 835.950 499.050 838.050 ;
        RECT 499.950 835.950 502.050 838.050 ;
        RECT 502.950 835.950 505.050 838.050 ;
        RECT 505.950 835.950 508.050 838.050 ;
        RECT 497.400 834.900 498.600 835.950 ;
        RECT 496.950 832.800 499.050 834.900 ;
        RECT 499.950 826.950 502.050 829.050 ;
        RECT 481.950 814.950 484.050 817.050 ;
        RECT 490.950 814.950 493.050 817.050 ;
        RECT 478.950 811.950 481.050 814.050 ;
        RECT 469.950 807.000 472.050 811.050 ;
        RECT 470.400 805.050 471.600 807.000 ;
        RECT 475.950 805.950 478.050 811.050 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 469.950 802.950 472.050 805.050 ;
        RECT 472.950 802.950 475.050 805.050 ;
        RECT 464.400 793.050 465.600 802.950 ;
        RECT 473.400 801.900 474.600 802.950 ;
        RECT 479.400 802.050 480.600 811.950 ;
        RECT 472.950 799.800 475.050 801.900 ;
        RECT 475.950 799.950 478.050 802.050 ;
        RECT 463.950 790.950 466.050 793.050 ;
        RECT 476.400 787.050 477.600 799.950 ;
        RECT 478.950 796.950 481.050 802.050 ;
        RECT 482.400 793.050 483.600 814.950 ;
        RECT 493.950 807.000 496.050 811.050 ;
        RECT 500.400 808.050 501.600 826.950 ;
        RECT 503.400 823.050 504.600 835.950 ;
        RECT 502.950 820.950 505.050 823.050 ;
        RECT 508.950 820.950 511.050 823.050 ;
        RECT 502.950 817.800 505.050 819.900 ;
        RECT 494.400 805.050 495.600 807.000 ;
        RECT 499.950 805.950 502.050 808.050 ;
        RECT 490.950 802.950 493.050 805.050 ;
        RECT 493.950 802.950 496.050 805.050 ;
        RECT 496.950 802.950 499.050 805.050 ;
        RECT 487.950 799.950 490.050 802.050 ;
        RECT 491.400 801.000 492.600 802.950 ;
        RECT 497.400 801.900 498.600 802.950 ;
        RECT 481.950 790.950 484.050 793.050 ;
        RECT 475.950 784.950 478.050 787.050 ;
        RECT 481.950 784.950 484.050 787.050 ;
        RECT 457.950 781.950 460.050 784.050 ;
        RECT 455.400 779.400 459.600 780.600 ;
        RECT 445.950 775.950 448.050 778.050 ;
        RECT 451.950 775.950 454.050 778.050 ;
        RECT 445.950 772.800 448.050 774.900 ;
        RECT 446.400 763.200 447.600 772.800 ;
        RECT 452.400 763.200 453.600 775.950 ;
        RECT 445.950 761.100 448.050 763.200 ;
        RECT 451.950 761.100 454.050 763.200 ;
        RECT 446.400 760.050 447.600 761.100 ;
        RECT 452.400 760.050 453.600 761.100 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 449.400 756.900 450.600 757.950 ;
        RECT 440.400 755.400 444.600 756.600 ;
        RECT 439.950 745.950 442.050 748.050 ;
        RECT 424.950 742.950 427.050 745.050 ;
        RECT 424.950 733.950 427.050 736.050 ;
        RECT 425.400 730.200 426.600 733.950 ;
        RECT 421.950 727.950 424.050 730.050 ;
        RECT 424.950 728.100 427.050 730.200 ;
        RECT 430.950 728.100 433.050 730.200 ;
        RECT 425.400 727.050 426.600 728.100 ;
        RECT 431.400 727.050 432.600 728.100 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 427.950 724.950 430.050 727.050 ;
        RECT 430.950 724.950 433.050 727.050 ;
        RECT 433.950 724.950 436.050 727.050 ;
        RECT 418.950 721.950 421.050 724.050 ;
        RECT 428.400 723.900 429.600 724.950 ;
        RECT 418.950 718.800 421.050 720.900 ;
        RECT 427.950 718.950 430.050 723.900 ;
        RECT 419.400 685.050 420.600 718.800 ;
        RECT 434.400 712.050 435.600 724.950 ;
        RECT 433.950 709.950 436.050 712.050 ;
        RECT 430.950 694.950 433.050 697.050 ;
        RECT 418.950 682.950 421.050 685.050 ;
        RECT 421.950 683.100 424.050 685.200 ;
        RECT 422.400 682.050 423.600 683.100 ;
        RECT 421.950 679.950 424.050 682.050 ;
        RECT 424.950 679.950 427.050 682.050 ;
        RECT 425.400 678.900 426.600 679.950 ;
        RECT 424.950 676.800 427.050 678.900 ;
        RECT 421.950 673.950 424.050 676.050 ;
        RECT 418.950 664.950 421.050 667.050 ;
        RECT 415.950 658.950 418.050 661.050 ;
        RECT 419.400 658.050 420.600 664.950 ;
        RECT 418.950 655.950 421.050 658.050 ;
        RECT 413.400 654.000 420.600 654.600 ;
        RECT 413.400 653.400 421.050 654.000 ;
        RECT 412.950 650.100 415.050 652.200 ;
        RECT 413.400 649.050 414.600 650.100 ;
        RECT 418.950 649.950 421.050 653.400 ;
        RECT 422.400 651.600 423.600 673.950 ;
        RECT 431.400 670.050 432.600 694.950 ;
        RECT 434.400 685.050 435.600 709.950 ;
        RECT 436.950 703.950 439.050 706.050 ;
        RECT 437.400 688.050 438.600 703.950 ;
        RECT 440.400 697.050 441.600 745.950 ;
        RECT 443.400 745.050 444.600 755.400 ;
        RECT 448.950 754.800 451.050 756.900 ;
        RECT 458.400 756.600 459.600 779.400 ;
        RECT 466.950 772.950 469.050 775.050 ;
        RECT 472.950 772.950 475.050 775.050 ;
        RECT 467.400 760.050 468.600 772.950 ;
        RECT 473.400 760.050 474.600 772.950 ;
        RECT 463.950 757.950 466.050 760.050 ;
        RECT 466.950 757.950 469.050 760.050 ;
        RECT 469.950 757.950 472.050 760.050 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 464.400 756.900 465.600 757.950 ;
        RECT 458.400 755.400 462.600 756.600 ;
        RECT 457.950 751.950 460.050 754.050 ;
        RECT 458.400 745.050 459.600 751.950 ;
        RECT 442.950 742.950 445.050 745.050 ;
        RECT 457.950 742.950 460.050 745.050 ;
        RECT 448.950 733.950 451.050 736.050 ;
        RECT 457.950 733.950 460.050 736.050 ;
        RECT 449.400 727.050 450.600 733.950 ;
        RECT 454.950 728.100 457.050 730.200 ;
        RECT 458.400 730.050 459.600 733.950 ;
        RECT 455.400 727.050 456.600 728.100 ;
        RECT 457.950 727.950 460.050 730.050 ;
        RECT 445.950 724.950 448.050 727.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 451.950 724.950 454.050 727.050 ;
        RECT 454.950 724.950 457.050 727.050 ;
        RECT 446.400 723.000 447.600 724.950 ;
        RECT 445.950 718.950 448.050 723.000 ;
        RECT 439.950 694.950 442.050 697.050 ;
        RECT 439.950 690.600 444.000 691.050 ;
        RECT 439.950 690.000 444.600 690.600 ;
        RECT 439.950 688.950 445.050 690.000 ;
        RECT 436.950 687.600 441.000 688.050 ;
        RECT 436.950 685.950 441.600 687.600 ;
        RECT 442.950 685.950 445.050 688.950 ;
        RECT 433.950 682.950 436.050 685.050 ;
        RECT 440.400 682.050 441.600 685.950 ;
        RECT 446.400 682.050 447.600 718.950 ;
        RECT 452.400 709.050 453.600 724.950 ;
        RECT 454.950 718.950 457.050 721.050 ;
        RECT 451.950 706.950 454.050 709.050 ;
        RECT 455.400 706.050 456.600 718.950 ;
        RECT 454.950 703.950 457.050 706.050 ;
        RECT 451.950 685.950 454.050 688.050 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 439.950 679.950 442.050 682.050 ;
        RECT 442.950 679.950 445.050 682.050 ;
        RECT 445.950 679.950 448.050 682.050 ;
        RECT 433.950 676.950 436.050 679.050 ;
        RECT 437.400 678.900 438.600 679.950 ;
        RECT 443.400 678.900 444.600 679.950 ;
        RECT 452.400 678.900 453.600 685.950 ;
        RECT 430.950 667.950 433.050 670.050 ;
        RECT 427.950 656.400 430.050 658.500 ;
        RECT 422.400 650.400 426.600 651.600 ;
        RECT 425.400 649.050 426.600 650.400 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 415.950 646.950 418.050 649.050 ;
        RECT 424.950 646.950 427.050 649.050 ;
        RECT 403.950 643.950 406.050 646.050 ;
        RECT 382.500 638.400 384.600 640.500 ;
        RECT 392.100 639.600 394.200 641.700 ;
        RECT 397.950 640.950 400.050 643.050 ;
        RECT 404.400 634.050 405.600 643.950 ;
        RECT 410.400 640.050 411.600 646.950 ;
        RECT 409.950 637.950 412.050 640.050 ;
        RECT 397.950 631.950 400.050 634.050 ;
        RECT 403.950 631.950 406.050 634.050 ;
        RECT 385.950 628.950 388.050 631.050 ;
        RECT 379.950 625.950 382.050 628.050 ;
        RECT 380.400 586.050 381.600 625.950 ;
        RECT 386.400 625.050 387.600 628.950 ;
        RECT 385.950 622.950 388.050 625.050 ;
        RECT 394.950 616.950 397.050 619.050 ;
        RECT 391.950 606.000 394.050 610.050 ;
        RECT 395.400 607.050 396.600 616.950 ;
        RECT 398.400 616.050 399.600 631.950 ;
        RECT 406.950 622.950 409.050 625.050 ;
        RECT 397.950 613.950 400.050 616.050 ;
        RECT 400.950 613.950 406.050 616.050 ;
        RECT 400.950 610.800 403.050 612.900 ;
        RECT 397.950 607.950 400.050 610.050 ;
        RECT 392.400 604.050 393.600 606.000 ;
        RECT 394.950 604.950 397.050 607.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 386.400 600.900 387.600 601.950 ;
        RECT 385.950 598.800 388.050 600.900 ;
        RECT 398.400 586.050 399.600 607.950 ;
        RECT 379.950 583.950 382.050 586.050 ;
        RECT 391.950 580.950 394.050 586.050 ;
        RECT 397.950 583.950 400.050 586.050 ;
        RECT 397.950 580.800 400.050 582.900 ;
        RECT 382.950 577.950 385.050 580.050 ;
        RECT 393.000 579.900 396.000 580.050 ;
        RECT 391.950 577.950 397.050 579.900 ;
        RECT 367.950 571.950 370.050 574.050 ;
        RECT 370.950 573.000 373.050 577.050 ;
        RECT 376.950 574.950 379.050 577.050 ;
        RECT 371.400 571.050 372.600 573.000 ;
        RECT 383.400 571.050 384.600 577.950 ;
        RECT 391.950 577.800 394.050 577.950 ;
        RECT 394.950 577.800 397.050 577.950 ;
        RECT 388.950 572.100 391.050 574.200 ;
        RECT 389.400 571.050 390.600 572.100 ;
        RECT 394.950 571.950 397.050 574.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 379.950 568.950 382.050 571.050 ;
        RECT 382.950 568.950 385.050 571.050 ;
        RECT 385.950 568.950 388.050 571.050 ;
        RECT 388.950 568.950 391.050 571.050 ;
        RECT 358.950 559.950 361.050 562.050 ;
        RECT 361.950 550.950 364.050 553.050 ;
        RECT 352.800 544.950 354.900 547.050 ;
        RECT 355.950 544.950 358.050 547.050 ;
        RECT 353.400 529.050 354.600 544.950 ;
        RECT 355.950 535.950 358.050 538.050 ;
        RECT 352.950 526.950 355.050 529.050 ;
        RECT 356.400 526.050 357.600 535.950 ;
        RECT 362.400 529.050 363.600 550.950 ;
        RECT 365.400 550.050 366.600 568.950 ;
        RECT 373.950 565.950 376.050 568.050 ;
        RECT 367.950 562.950 370.050 565.050 ;
        RECT 364.950 547.950 367.050 550.050 ;
        RECT 364.950 538.950 367.050 541.050 ;
        RECT 361.950 526.950 364.050 529.050 ;
        RECT 355.950 523.950 358.050 526.050 ;
        RECT 358.950 523.950 361.050 526.050 ;
        RECT 359.400 522.900 360.600 523.950 ;
        RECT 358.950 520.800 361.050 522.900 ;
        RECT 352.950 517.950 355.050 520.050 ;
        RECT 340.950 499.950 343.050 502.050 ;
        RECT 349.950 499.950 352.050 502.050 ;
        RECT 341.400 493.050 342.600 499.950 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 346.950 490.950 349.050 493.050 ;
        RECT 334.950 487.950 337.050 490.050 ;
        RECT 335.400 481.050 336.600 487.950 ;
        RECT 334.950 478.950 337.050 481.050 ;
        RECT 338.400 475.050 339.600 490.950 ;
        RECT 347.400 481.050 348.600 490.950 ;
        RECT 349.950 484.950 352.050 487.050 ;
        RECT 340.950 478.950 343.050 481.050 ;
        RECT 346.950 478.950 349.050 481.050 ;
        RECT 337.950 472.950 340.050 475.050 ;
        RECT 331.950 466.950 334.050 469.050 ;
        RECT 319.950 463.950 322.050 466.050 ;
        RECT 322.950 463.950 325.050 466.050 ;
        RECT 316.950 448.950 319.050 451.050 ;
        RECT 304.950 445.950 307.050 448.050 ;
        RECT 307.950 445.950 310.050 448.050 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 320.400 447.600 321.600 463.950 ;
        RECT 317.400 446.400 321.600 447.600 ;
        RECT 305.400 444.000 306.600 445.950 ;
        RECT 311.400 444.900 312.600 445.950 ;
        RECT 304.950 439.950 307.050 444.000 ;
        RECT 310.800 442.800 312.900 444.900 ;
        RECT 313.950 442.950 316.050 445.050 ;
        RECT 301.950 430.950 304.050 433.050 ;
        RECT 298.950 418.950 301.050 421.050 ;
        RECT 295.950 415.950 298.050 418.050 ;
        RECT 302.400 415.050 303.600 430.950 ;
        RECT 307.950 427.950 310.050 430.050 ;
        RECT 314.400 429.600 315.600 442.950 ;
        RECT 311.400 428.400 315.600 429.600 ;
        RECT 308.400 424.050 309.600 427.950 ;
        RECT 307.950 421.950 310.050 424.050 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 299.400 411.900 300.600 412.950 ;
        RECT 298.950 409.800 301.050 411.900 ;
        RECT 301.950 406.950 304.050 409.050 ;
        RECT 302.400 403.050 303.600 406.950 ;
        RECT 301.950 400.950 304.050 403.050 ;
        RECT 292.950 379.950 295.050 382.050 ;
        RECT 283.800 370.950 285.900 373.050 ;
        RECT 286.950 371.100 289.050 373.200 ;
        RECT 292.950 372.000 295.050 376.050 ;
        RECT 287.400 370.050 288.600 371.100 ;
        RECT 293.400 370.050 294.600 372.000 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 289.950 367.950 292.050 370.050 ;
        RECT 292.950 367.950 295.050 370.050 ;
        RECT 298.950 367.950 301.050 370.050 ;
        RECT 283.950 364.950 286.050 367.050 ;
        RECT 280.950 358.950 283.050 361.050 ;
        RECT 277.950 355.950 280.050 358.050 ;
        RECT 271.950 346.950 274.050 349.050 ;
        RECT 259.950 343.950 262.050 346.050 ;
        RECT 262.950 343.950 265.050 346.050 ;
        RECT 267.000 345.600 271.050 346.050 ;
        RECT 266.400 343.950 271.050 345.600 ;
        RECT 266.400 340.200 267.600 343.950 ;
        RECT 253.950 337.950 256.050 340.050 ;
        RECT 256.950 338.100 259.050 340.200 ;
        RECT 265.950 338.100 268.050 340.200 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 241.950 331.950 244.050 334.050 ;
        RECT 248.400 333.900 249.600 334.950 ;
        RECT 238.950 322.950 241.050 325.050 ;
        RECT 242.400 322.050 243.600 331.950 ;
        RECT 247.950 331.800 250.050 333.900 ;
        RECT 257.400 328.050 258.600 338.100 ;
        RECT 266.400 337.050 267.600 338.100 ;
        RECT 272.400 337.050 273.600 346.950 ;
        RECT 278.400 343.050 279.600 355.950 ;
        RECT 280.950 349.950 283.050 352.050 ;
        RECT 277.800 340.950 279.900 343.050 ;
        RECT 281.400 340.050 282.600 349.950 ;
        RECT 284.400 340.050 285.600 364.950 ;
        RECT 286.950 361.950 289.050 364.050 ;
        RECT 287.400 352.050 288.600 361.950 ;
        RECT 290.400 361.050 291.600 367.950 ;
        RECT 295.950 364.950 298.050 367.050 ;
        RECT 289.950 358.950 292.050 361.050 ;
        RECT 292.950 355.950 295.050 358.050 ;
        RECT 286.950 349.950 289.050 352.050 ;
        RECT 280.950 337.950 283.050 340.050 ;
        RECT 283.950 337.950 286.050 340.050 ;
        RECT 289.950 339.000 292.050 343.050 ;
        RECT 293.400 340.050 294.600 355.950 ;
        RECT 296.400 355.050 297.600 364.950 ;
        RECT 295.950 352.950 298.050 355.050 ;
        RECT 299.400 342.600 300.600 367.950 ;
        RECT 302.400 367.050 303.600 400.950 ;
        RECT 305.400 394.050 306.600 412.950 ;
        RECT 304.950 391.950 307.050 394.050 ;
        RECT 311.400 391.050 312.600 428.400 ;
        RECT 313.950 424.950 316.050 427.050 ;
        RECT 314.400 418.050 315.600 424.950 ;
        RECT 317.400 418.050 318.600 446.400 ;
        RECT 319.950 442.950 322.050 445.050 ;
        RECT 320.400 424.050 321.600 442.950 ;
        RECT 323.400 433.050 324.600 463.950 ;
        RECT 328.950 460.950 331.050 463.050 ;
        RECT 325.950 454.950 328.050 457.050 ;
        RECT 326.400 451.050 327.600 454.950 ;
        RECT 325.950 448.950 328.050 451.050 ;
        RECT 329.400 448.050 330.600 460.950 ;
        RECT 341.400 460.050 342.600 478.950 ;
        RECT 346.950 475.800 349.050 477.900 ;
        RECT 347.400 466.050 348.600 475.800 ;
        RECT 346.950 463.950 349.050 466.050 ;
        RECT 350.400 462.600 351.600 484.950 ;
        RECT 353.400 478.050 354.600 517.950 ;
        RECT 365.400 508.050 366.600 538.950 ;
        RECT 355.800 505.950 357.900 508.050 ;
        RECT 358.950 505.950 361.050 508.050 ;
        RECT 364.950 505.950 367.050 508.050 ;
        RECT 356.400 499.050 357.600 505.950 ;
        RECT 355.950 496.950 358.050 499.050 ;
        RECT 359.400 496.050 360.600 505.950 ;
        RECT 368.400 505.050 369.600 562.950 ;
        RECT 370.950 541.950 373.050 544.050 ;
        RECT 371.400 534.600 372.600 541.950 ;
        RECT 374.400 541.050 375.600 565.950 ;
        RECT 380.400 556.050 381.600 568.950 ;
        RECT 382.950 562.950 385.050 565.050 ;
        RECT 379.950 553.950 382.050 556.050 ;
        RECT 373.950 538.950 376.050 541.050 ;
        RECT 371.400 533.400 375.600 534.600 ;
        RECT 374.400 526.050 375.600 533.400 ;
        RECT 383.400 529.050 384.600 562.950 ;
        RECT 386.400 562.050 387.600 568.950 ;
        RECT 385.950 559.950 388.050 562.050 ;
        RECT 386.400 532.050 387.600 559.950 ;
        RECT 395.400 549.600 396.600 571.950 ;
        RECT 398.400 565.050 399.600 580.800 ;
        RECT 397.950 562.950 400.050 565.050 ;
        RECT 395.400 548.400 399.600 549.600 ;
        RECT 394.950 544.950 397.050 547.050 ;
        RECT 385.950 529.950 388.050 532.050 ;
        RECT 382.950 528.600 385.050 529.050 ;
        RECT 380.400 527.400 385.050 528.600 ;
        RECT 380.400 526.050 381.600 527.400 ;
        RECT 382.950 526.950 385.050 527.400 ;
        RECT 395.400 528.600 396.600 544.950 ;
        RECT 398.400 541.050 399.600 548.400 ;
        RECT 401.400 544.050 402.600 610.800 ;
        RECT 407.400 604.050 408.600 622.950 ;
        RECT 412.950 605.100 415.050 607.200 ;
        RECT 416.400 607.050 417.600 646.950 ;
        RECT 421.950 643.950 424.050 646.050 ;
        RECT 418.950 640.950 421.050 643.050 ;
        RECT 413.400 604.050 414.600 605.100 ;
        RECT 415.950 604.950 418.050 607.050 ;
        RECT 406.950 601.950 409.050 604.050 ;
        RECT 409.950 601.950 412.050 604.050 ;
        RECT 412.950 601.950 415.050 604.050 ;
        RECT 410.400 600.900 411.600 601.950 ;
        RECT 403.950 598.800 406.050 600.900 ;
        RECT 409.950 598.800 412.050 600.900 ;
        RECT 404.400 580.050 405.600 598.800 ;
        RECT 415.950 595.950 418.050 601.050 ;
        RECT 412.950 580.950 415.050 583.050 ;
        RECT 403.950 577.950 406.050 580.050 ;
        RECT 404.400 574.050 405.600 577.950 ;
        RECT 403.950 571.950 406.050 574.050 ;
        RECT 406.950 573.000 409.050 580.050 ;
        RECT 407.400 571.050 408.600 573.000 ;
        RECT 413.400 571.050 414.600 580.950 ;
        RECT 419.400 580.050 420.600 640.950 ;
        RECT 422.400 610.050 423.600 643.950 ;
        RECT 428.850 641.400 430.050 656.400 ;
        RECT 434.400 654.600 435.600 676.950 ;
        RECT 436.950 676.800 439.050 678.900 ;
        RECT 442.950 676.800 445.050 678.900 ;
        RECT 451.950 676.800 454.050 678.900 ;
        RECT 436.950 670.950 439.050 673.050 ;
        RECT 437.400 658.050 438.600 670.950 ;
        RECT 455.400 667.050 456.600 703.950 ;
        RECT 461.400 700.050 462.600 755.400 ;
        RECT 463.950 754.800 466.050 756.900 ;
        RECT 464.400 723.600 465.600 754.800 ;
        RECT 470.400 739.050 471.600 757.950 ;
        RECT 475.950 754.800 478.050 756.900 ;
        RECT 476.400 742.050 477.600 754.800 ;
        RECT 482.400 754.050 483.600 784.950 ;
        RECT 488.400 783.600 489.600 799.950 ;
        RECT 490.950 796.950 493.050 801.000 ;
        RECT 496.950 796.950 499.050 801.900 ;
        RECT 499.950 784.950 502.050 787.050 ;
        RECT 488.400 782.400 492.600 783.600 ;
        RECT 487.950 778.950 490.050 781.050 ;
        RECT 488.400 760.050 489.600 778.950 ;
        RECT 491.400 772.050 492.600 782.400 ;
        RECT 490.950 769.950 493.050 772.050 ;
        RECT 493.950 761.100 496.050 763.200 ;
        RECT 494.400 760.050 495.600 761.100 ;
        RECT 500.400 760.050 501.600 784.950 ;
        RECT 503.400 784.050 504.600 817.800 ;
        RECT 505.950 808.950 508.050 811.050 ;
        RECT 506.400 802.050 507.600 808.950 ;
        RECT 509.400 808.050 510.600 820.950 ;
        RECT 512.400 811.050 513.600 868.950 ;
        RECT 521.400 868.050 522.600 880.950 ;
        RECT 527.400 879.900 528.600 880.950 ;
        RECT 533.400 880.050 534.600 898.950 ;
        RECT 536.400 898.050 537.600 917.100 ;
        RECT 542.400 916.050 543.600 917.100 ;
        RECT 548.400 916.050 549.600 917.100 ;
        RECT 541.950 913.950 544.050 916.050 ;
        RECT 544.950 913.950 547.050 916.050 ;
        RECT 547.950 913.950 550.050 916.050 ;
        RECT 550.950 913.950 553.050 916.050 ;
        RECT 545.400 907.050 546.600 913.950 ;
        RECT 551.400 912.900 552.600 913.950 ;
        RECT 550.950 910.800 553.050 912.900 ;
        RECT 557.400 907.050 558.600 922.950 ;
        RECT 565.950 917.100 568.050 919.200 ;
        RECT 566.400 916.050 567.600 917.100 ;
        RECT 572.400 916.050 573.600 922.950 ;
        RECT 584.400 919.200 585.600 922.950 ;
        RECT 583.800 917.100 585.900 919.200 ;
        RECT 586.950 917.100 589.050 922.050 ;
        RECT 592.950 917.100 595.050 919.200 ;
        RECT 598.950 917.100 601.050 919.200 ;
        RECT 602.400 919.050 603.600 922.950 ;
        RECT 562.950 913.950 565.050 916.050 ;
        RECT 565.950 913.950 568.050 916.050 ;
        RECT 568.950 913.950 571.050 916.050 ;
        RECT 571.950 913.950 574.050 916.050 ;
        RECT 544.950 904.950 547.050 907.050 ;
        RECT 556.950 904.950 559.050 907.050 ;
        RECT 563.400 898.050 564.600 913.950 ;
        RECT 565.950 901.950 568.050 904.050 ;
        RECT 535.950 895.950 538.050 898.050 ;
        RECT 562.950 895.950 565.050 898.050 ;
        RECT 541.950 885.000 544.050 889.050 ;
        RECT 550.950 886.950 553.050 889.050 ;
        RECT 542.400 883.050 543.600 885.000 ;
        RECT 551.400 883.050 552.600 886.950 ;
        RECT 553.950 883.950 556.050 886.050 ;
        RECT 556.950 885.600 561.000 886.050 ;
        RECT 556.950 883.950 561.600 885.600 ;
        RECT 541.950 880.950 544.050 883.050 ;
        RECT 544.950 880.950 547.050 883.050 ;
        RECT 550.950 880.950 553.050 883.050 ;
        RECT 526.950 877.800 529.050 879.900 ;
        RECT 532.950 877.950 535.050 880.050 ;
        RECT 545.400 879.900 546.600 880.950 ;
        RECT 554.400 879.900 555.600 883.950 ;
        RECT 560.400 883.050 561.600 883.950 ;
        RECT 566.400 883.050 567.600 901.950 ;
        RECT 569.400 901.050 570.600 913.950 ;
        RECT 584.400 913.050 585.600 917.100 ;
        RECT 593.400 916.050 594.600 917.100 ;
        RECT 599.400 916.050 600.600 917.100 ;
        RECT 601.950 916.950 604.050 919.050 ;
        RECT 604.950 917.100 607.050 919.200 ;
        RECT 613.950 917.100 616.050 919.200 ;
        RECT 589.950 913.950 592.050 916.050 ;
        RECT 592.950 913.950 595.050 916.050 ;
        RECT 595.950 913.950 598.050 916.050 ;
        RECT 598.950 913.950 601.050 916.050 ;
        RECT 583.950 910.950 586.050 913.050 ;
        RECT 586.950 909.600 589.050 913.050 ;
        RECT 590.400 912.900 591.600 913.950 ;
        RECT 589.950 910.800 592.050 912.900 ;
        RECT 596.400 912.000 597.600 913.950 ;
        RECT 586.950 909.000 591.600 909.600 ;
        RECT 587.400 908.400 591.600 909.000 ;
        RECT 568.950 898.950 571.050 901.050 ;
        RECT 590.400 883.050 591.600 908.400 ;
        RECT 595.950 907.950 598.050 912.000 ;
        RECT 601.950 907.950 604.050 910.050 ;
        RECT 595.950 889.950 598.050 892.050 ;
        RECT 596.400 883.050 597.600 889.950 ;
        RECT 559.950 880.950 562.050 883.050 ;
        RECT 562.950 880.950 565.050 883.050 ;
        RECT 565.950 880.950 568.050 883.050 ;
        RECT 568.950 880.950 571.050 883.050 ;
        RECT 586.950 880.950 589.050 883.050 ;
        RECT 589.950 880.950 592.050 883.050 ;
        RECT 592.950 880.950 595.050 883.050 ;
        RECT 595.950 880.950 598.050 883.050 ;
        RECT 544.950 877.800 547.050 879.900 ;
        RECT 550.950 877.800 553.050 879.900 ;
        RECT 553.950 877.800 556.050 879.900 ;
        RECT 532.950 871.950 535.050 874.050 ;
        RECT 520.950 865.950 523.050 868.050 ;
        RECT 514.950 847.950 517.050 850.050 ;
        RECT 526.950 847.950 529.050 850.050 ;
        RECT 515.400 832.050 516.600 847.950 ;
        RECT 520.950 839.100 523.050 841.200 ;
        RECT 521.400 838.050 522.600 839.100 ;
        RECT 527.400 838.050 528.600 847.950 ;
        RECT 533.400 841.200 534.600 871.950 ;
        RECT 545.400 867.600 546.600 877.800 ;
        RECT 542.400 866.400 546.600 867.600 ;
        RECT 538.950 862.800 541.050 864.900 ;
        RECT 532.950 839.100 535.050 841.200 ;
        RECT 533.400 838.050 534.600 839.100 ;
        RECT 520.950 835.950 523.050 838.050 ;
        RECT 523.950 835.950 526.050 838.050 ;
        RECT 526.950 835.950 529.050 838.050 ;
        RECT 529.950 835.950 532.050 838.050 ;
        RECT 532.950 835.950 535.050 838.050 ;
        RECT 524.400 834.000 525.600 835.950 ;
        RECT 514.950 829.950 517.050 832.050 ;
        RECT 523.950 829.950 526.050 834.000 ;
        RECT 511.950 808.950 514.050 811.050 ;
        RECT 508.950 805.950 511.050 808.050 ;
        RECT 515.400 805.050 516.600 829.950 ;
        RECT 524.400 826.050 525.600 829.950 ;
        RECT 520.800 823.950 522.900 826.050 ;
        RECT 523.950 823.950 526.050 826.050 ;
        RECT 521.400 805.050 522.600 823.950 ;
        RECT 523.950 820.800 526.050 822.900 ;
        RECT 524.400 811.050 525.600 820.800 ;
        RECT 530.400 820.050 531.600 835.950 ;
        RECT 535.950 832.950 538.050 835.050 ;
        RECT 532.950 829.950 535.050 832.050 ;
        RECT 529.950 817.950 532.050 820.050 ;
        RECT 529.950 811.950 532.050 814.050 ;
        RECT 523.950 808.950 526.050 811.050 ;
        RECT 530.400 808.050 531.600 811.950 ;
        RECT 529.950 805.950 532.050 808.050 ;
        RECT 533.400 805.050 534.600 829.950 ;
        RECT 536.400 823.050 537.600 832.950 ;
        RECT 535.950 820.950 538.050 823.050 ;
        RECT 539.400 820.050 540.600 862.800 ;
        RECT 538.950 817.950 541.050 820.050 ;
        RECT 542.400 813.600 543.600 866.400 ;
        RECT 551.400 850.050 552.600 877.800 ;
        RECT 563.400 876.600 564.600 880.950 ;
        RECT 569.400 879.900 570.600 880.950 ;
        RECT 587.400 879.900 588.600 880.950 ;
        RECT 568.950 877.800 571.050 879.900 ;
        RECT 586.950 877.800 589.050 879.900 ;
        RECT 593.400 877.050 594.600 880.950 ;
        RECT 602.400 877.050 603.600 907.950 ;
        RECT 605.400 892.050 606.600 917.100 ;
        RECT 614.400 916.050 615.600 917.100 ;
        RECT 619.800 916.950 621.900 919.050 ;
        RECT 622.950 917.100 625.050 919.200 ;
        RECT 628.950 917.100 631.050 919.200 ;
        RECT 634.950 917.100 637.050 919.200 ;
        RECT 610.950 913.950 613.050 916.050 ;
        RECT 613.950 913.950 616.050 916.050 ;
        RECT 611.400 913.050 612.600 913.950 ;
        RECT 607.950 911.400 612.600 913.050 ;
        RECT 607.950 910.950 612.000 911.400 ;
        RECT 620.400 910.050 621.600 916.950 ;
        RECT 619.950 907.950 622.050 910.050 ;
        RECT 623.400 904.050 624.600 917.100 ;
        RECT 629.400 916.050 630.600 917.100 ;
        RECT 635.400 916.050 636.600 917.100 ;
        RECT 628.950 913.950 631.050 916.050 ;
        RECT 631.950 913.950 634.050 916.050 ;
        RECT 634.950 913.950 637.050 916.050 ;
        RECT 637.950 913.950 640.050 916.050 ;
        RECT 632.400 907.050 633.600 913.950 ;
        RECT 638.400 912.900 639.600 913.950 ;
        RECT 637.950 910.800 640.050 912.900 ;
        RECT 644.400 912.600 645.600 922.950 ;
        RECT 653.400 919.200 654.600 931.950 ;
        RECT 658.950 922.950 661.050 925.050 ;
        RECT 652.950 917.100 655.050 919.200 ;
        RECT 653.400 916.050 654.600 917.100 ;
        RECT 659.400 916.050 660.600 922.950 ;
        RECT 649.950 913.950 652.050 916.050 ;
        RECT 652.950 913.950 655.050 916.050 ;
        RECT 655.950 913.950 658.050 916.050 ;
        RECT 658.950 913.950 661.050 916.050 ;
        RECT 641.400 911.400 645.600 912.600 ;
        RECT 634.950 907.950 637.050 910.050 ;
        RECT 631.950 904.950 634.050 907.050 ;
        RECT 622.950 901.950 625.050 904.050 ;
        RECT 635.400 901.050 636.600 907.950 ;
        RECT 638.400 903.600 639.600 910.800 ;
        RECT 641.400 907.050 642.600 911.400 ;
        RECT 643.950 907.950 646.050 910.050 ;
        RECT 640.950 904.950 643.050 907.050 ;
        RECT 638.400 902.400 642.600 903.600 ;
        RECT 628.950 898.950 631.050 901.050 ;
        RECT 634.950 898.950 637.050 901.050 ;
        RECT 629.400 895.050 630.600 898.950 ;
        RECT 628.950 892.950 631.050 895.050 ;
        RECT 604.950 889.950 607.050 892.050 ;
        RECT 619.950 889.950 622.050 892.050 ;
        RECT 620.400 886.200 621.600 889.950 ;
        RECT 641.400 889.050 642.600 902.400 ;
        RECT 644.400 889.050 645.600 907.950 ;
        RECT 650.400 904.050 651.600 913.950 ;
        RECT 649.950 901.950 652.050 904.050 ;
        RECT 649.800 898.800 651.900 900.900 ;
        RECT 652.950 898.950 655.050 901.050 ;
        RECT 613.950 884.100 616.050 886.200 ;
        RECT 619.950 884.100 622.050 886.200 ;
        RECT 631.950 884.100 634.050 886.200 ;
        RECT 637.950 885.000 640.050 889.050 ;
        RECT 640.950 886.950 643.050 889.050 ;
        RECT 643.950 886.950 646.050 889.050 ;
        RECT 614.400 883.050 615.600 884.100 ;
        RECT 620.400 883.050 621.600 884.100 ;
        RECT 632.400 883.050 633.600 884.100 ;
        RECT 638.400 883.050 639.600 885.000 ;
        RECT 610.950 880.950 613.050 883.050 ;
        RECT 613.950 880.950 616.050 883.050 ;
        RECT 616.950 880.950 619.050 883.050 ;
        RECT 619.950 880.950 622.050 883.050 ;
        RECT 628.950 880.950 631.050 883.050 ;
        RECT 631.950 880.950 634.050 883.050 ;
        RECT 634.950 880.950 637.050 883.050 ;
        RECT 637.950 880.950 640.050 883.050 ;
        RECT 611.400 879.900 612.600 880.950 ;
        RECT 610.950 877.800 613.050 879.900 ;
        RECT 560.400 875.400 564.600 876.600 ;
        RECT 553.950 856.950 556.050 859.050 ;
        RECT 550.950 847.950 553.050 850.050 ;
        RECT 554.400 841.200 555.600 856.950 ;
        RECT 553.950 839.100 556.050 841.200 ;
        RECT 554.400 838.050 555.600 839.100 ;
        RECT 550.950 835.950 553.050 838.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 544.950 832.950 547.050 835.050 ;
        RECT 551.400 834.900 552.600 835.950 ;
        RECT 545.400 828.600 546.600 832.950 ;
        RECT 550.950 832.800 553.050 834.900 ;
        RECT 547.950 828.600 550.050 829.050 ;
        RECT 545.400 827.400 550.050 828.600 ;
        RECT 547.950 826.950 550.050 827.400 ;
        RECT 544.950 823.800 547.050 825.900 ;
        RECT 545.400 817.050 546.600 823.800 ;
        RECT 544.950 814.950 547.050 817.050 ;
        RECT 542.400 812.400 546.600 813.600 ;
        RECT 538.950 806.100 541.050 808.200 ;
        RECT 545.400 808.050 546.600 812.400 ;
        RECT 539.400 805.050 540.600 806.100 ;
        RECT 544.950 805.950 547.050 808.050 ;
        RECT 511.950 802.950 514.050 805.050 ;
        RECT 514.950 802.950 517.050 805.050 ;
        RECT 517.950 802.950 520.050 805.050 ;
        RECT 520.950 802.950 523.050 805.050 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 532.950 802.950 535.050 805.050 ;
        RECT 535.950 802.950 538.050 805.050 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 541.950 802.950 544.050 805.050 ;
        RECT 505.950 799.950 508.050 802.050 ;
        RECT 508.950 799.950 511.050 802.050 ;
        RECT 512.400 801.900 513.600 802.950 ;
        RECT 505.950 796.800 508.050 798.900 ;
        RECT 502.950 781.950 505.050 784.050 ;
        RECT 487.950 757.950 490.050 760.050 ;
        RECT 490.950 757.950 493.050 760.050 ;
        RECT 493.950 757.950 496.050 760.050 ;
        RECT 496.950 757.950 499.050 760.050 ;
        RECT 499.950 757.950 502.050 760.050 ;
        RECT 491.400 756.900 492.600 757.950 ;
        RECT 490.950 754.800 493.050 756.900 ;
        RECT 497.400 756.000 498.600 757.950 ;
        RECT 481.950 751.950 484.050 754.050 ;
        RECT 487.950 751.950 490.050 754.050 ;
        RECT 496.950 751.950 499.050 756.000 ;
        RECT 502.950 754.800 505.050 756.900 ;
        RECT 481.950 742.950 484.050 745.050 ;
        RECT 475.950 739.950 478.050 742.050 ;
        RECT 469.950 736.950 472.050 739.050 ;
        RECT 472.950 728.100 475.050 730.200 ;
        RECT 473.400 727.050 474.600 728.100 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 475.950 724.950 478.050 727.050 ;
        RECT 464.400 722.400 468.600 723.600 ;
        RECT 470.400 723.000 471.600 724.950 ;
        RECT 476.400 723.000 477.600 724.950 ;
        RECT 460.950 697.950 463.050 700.050 ;
        RECT 463.950 688.950 466.050 691.050 ;
        RECT 464.400 685.050 465.600 688.950 ;
        RECT 463.950 682.950 466.050 685.050 ;
        RECT 467.400 682.050 468.600 722.400 ;
        RECT 469.950 718.950 472.050 723.000 ;
        RECT 475.950 718.950 478.050 723.000 ;
        RECT 478.950 721.800 481.050 723.900 ;
        RECT 479.400 717.600 480.600 721.800 ;
        RECT 482.400 718.050 483.600 742.950 ;
        RECT 484.950 727.950 487.050 730.050 ;
        RECT 476.400 716.400 480.600 717.600 ;
        RECT 472.950 682.950 475.050 685.050 ;
        RECT 460.950 679.950 463.050 682.050 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 461.400 678.900 462.600 679.950 ;
        RECT 460.950 676.800 463.050 678.900 ;
        RECT 469.950 673.950 472.050 676.050 ;
        RECT 439.950 664.950 442.050 667.050 ;
        RECT 454.950 664.950 457.050 667.050 ;
        RECT 436.950 655.950 439.050 658.050 ;
        RECT 434.400 653.400 438.600 654.600 ;
        RECT 433.950 649.950 436.050 652.050 ;
        RECT 427.950 639.300 430.050 641.400 ;
        RECT 428.850 635.700 430.050 639.300 ;
        RECT 427.950 633.600 430.050 635.700 ;
        RECT 430.950 625.950 433.050 628.050 ;
        RECT 424.950 613.050 427.050 616.050 ;
        RECT 424.950 612.000 430.050 613.050 ;
        RECT 425.400 611.400 430.050 612.000 ;
        RECT 426.000 610.950 430.050 611.400 ;
        RECT 421.950 607.950 424.050 610.050 ;
        RECT 427.950 605.100 430.050 607.200 ;
        RECT 431.400 606.600 432.600 625.950 ;
        RECT 434.400 625.050 435.600 649.950 ;
        RECT 433.950 622.950 436.050 625.050 ;
        RECT 431.400 605.400 435.600 606.600 ;
        RECT 428.400 604.050 429.600 605.100 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 425.400 600.900 426.600 601.950 ;
        RECT 424.950 600.600 427.050 600.900 ;
        RECT 422.400 599.400 427.050 600.600 ;
        RECT 418.950 577.950 421.050 580.050 ;
        RECT 418.950 574.800 421.050 576.900 ;
        RECT 406.950 568.950 409.050 571.050 ;
        RECT 409.950 568.950 412.050 571.050 ;
        RECT 412.950 568.950 415.050 571.050 ;
        RECT 403.950 565.950 406.050 568.050 ;
        RECT 400.950 541.950 403.050 544.050 ;
        RECT 397.950 538.950 400.050 541.050 ;
        RECT 395.400 527.400 402.600 528.600 ;
        RECT 395.400 526.050 396.600 527.400 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 379.950 523.950 382.050 526.050 ;
        RECT 385.950 523.950 388.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 370.950 520.950 373.050 523.050 ;
        RECT 377.400 522.000 378.600 523.950 ;
        RECT 367.950 502.950 370.050 505.050 ;
        RECT 355.950 493.800 358.050 495.900 ;
        RECT 358.950 493.950 361.050 496.050 ;
        RECT 364.950 494.100 367.050 496.200 ;
        RECT 371.400 496.050 372.600 520.950 ;
        RECT 376.950 517.950 379.050 522.000 ;
        RECT 386.400 517.050 387.600 523.950 ;
        RECT 388.950 520.950 391.050 523.050 ;
        RECT 385.950 514.950 388.050 517.050 ;
        RECT 376.950 508.950 379.050 511.050 ;
        RECT 373.950 499.950 376.050 505.050 ;
        RECT 352.950 475.950 355.050 478.050 ;
        RECT 356.400 472.050 357.600 493.800 ;
        RECT 365.400 493.050 366.600 494.100 ;
        RECT 370.950 493.950 373.050 496.050 ;
        RECT 361.950 490.950 364.050 493.050 ;
        RECT 364.950 490.950 367.050 493.050 ;
        RECT 367.950 490.950 370.050 493.050 ;
        RECT 358.950 487.950 361.050 490.050 ;
        RECT 362.400 489.000 363.600 490.950 ;
        RECT 359.400 484.050 360.600 487.950 ;
        RECT 361.950 484.950 364.050 489.000 ;
        RECT 358.950 481.950 361.050 484.050 ;
        RECT 364.950 481.950 367.050 484.050 ;
        RECT 355.950 469.950 358.050 472.050 ;
        RECT 361.950 463.950 364.050 466.050 ;
        RECT 347.400 461.400 351.600 462.600 ;
        RECT 340.950 457.950 343.050 460.050 ;
        RECT 343.950 454.950 346.050 457.050 ;
        RECT 334.950 449.100 337.050 451.200 ;
        RECT 335.400 448.050 336.600 449.100 ;
        RECT 344.400 448.050 345.600 454.950 ;
        RECT 347.400 454.050 348.600 461.400 ;
        RECT 358.950 457.950 361.050 460.050 ;
        RECT 346.950 451.950 349.050 454.050 ;
        RECT 349.950 449.100 352.050 451.200 ;
        RECT 350.400 448.050 351.600 449.100 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 331.950 445.950 334.050 448.050 ;
        RECT 334.950 445.950 337.050 448.050 ;
        RECT 343.950 445.950 346.050 448.050 ;
        RECT 346.950 445.950 349.050 448.050 ;
        RECT 349.950 445.950 352.050 448.050 ;
        RECT 352.950 445.950 355.050 448.050 ;
        RECT 325.950 442.950 328.050 445.050 ;
        RECT 326.400 439.050 327.600 442.950 ;
        RECT 328.950 439.950 331.050 442.050 ;
        RECT 325.950 436.950 328.050 439.050 ;
        RECT 322.950 430.950 325.050 433.050 ;
        RECT 325.950 427.950 328.050 430.050 ;
        RECT 319.950 421.950 322.050 424.050 ;
        RECT 326.400 421.050 327.600 427.950 ;
        RECT 329.400 423.600 330.600 439.950 ;
        RECT 332.400 427.050 333.600 445.950 ;
        RECT 340.950 442.950 343.050 445.050 ;
        RECT 334.950 436.950 337.050 442.050 ;
        RECT 334.950 430.950 337.050 433.050 ;
        RECT 331.950 424.950 334.050 427.050 ;
        RECT 329.400 422.400 333.600 423.600 ;
        RECT 325.950 418.950 328.050 421.050 ;
        RECT 313.950 415.950 316.050 418.050 ;
        RECT 316.950 415.950 319.050 418.050 ;
        RECT 319.950 416.100 322.050 418.200 ;
        RECT 320.400 415.050 321.600 416.100 ;
        RECT 326.400 415.050 327.600 418.950 ;
        RECT 313.950 412.800 316.050 414.900 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 325.950 412.950 328.050 415.050 ;
        RECT 310.950 388.950 313.050 391.050 ;
        RECT 304.950 379.950 307.050 382.050 ;
        RECT 301.950 364.950 304.050 367.050 ;
        RECT 301.950 352.950 304.050 355.050 ;
        RECT 302.400 346.050 303.600 352.950 ;
        RECT 301.950 343.950 304.050 346.050 ;
        RECT 301.950 342.600 304.050 342.900 ;
        RECT 299.400 341.400 304.050 342.600 ;
        RECT 301.950 340.800 304.050 341.400 ;
        RECT 290.400 337.050 291.600 339.000 ;
        RECT 292.950 337.950 295.050 340.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 265.950 334.950 268.050 337.050 ;
        RECT 268.950 334.950 271.050 337.050 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 289.950 334.950 292.050 337.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 263.400 334.050 264.600 334.950 ;
        RECT 259.950 332.400 264.600 334.050 ;
        RECT 269.400 333.000 270.600 334.950 ;
        RECT 259.950 331.950 264.000 332.400 ;
        RECT 262.950 328.950 265.050 331.050 ;
        RECT 268.950 328.950 271.050 333.000 ;
        RECT 271.950 328.950 274.050 331.050 ;
        RECT 247.950 325.950 250.050 328.050 ;
        RECT 256.950 325.950 259.050 328.050 ;
        RECT 241.950 319.950 244.050 322.050 ;
        RECT 238.950 310.950 241.050 313.050 ;
        RECT 229.950 307.950 232.050 310.050 ;
        RECT 235.950 307.950 238.050 310.050 ;
        RECT 220.950 298.950 223.050 301.050 ;
        RECT 230.400 295.200 231.600 307.950 ;
        RECT 239.400 307.050 240.600 310.950 ;
        RECT 248.400 310.050 249.600 325.950 ;
        RECT 259.950 322.950 262.050 325.050 ;
        RECT 250.950 319.950 253.050 322.050 ;
        RECT 247.950 307.950 250.050 310.050 ;
        RECT 238.800 304.950 240.900 307.050 ;
        RECT 248.400 304.050 249.600 307.950 ;
        RECT 235.950 301.950 238.050 304.050 ;
        RECT 247.950 301.950 250.050 304.050 ;
        RECT 223.950 292.950 226.050 295.050 ;
        RECT 229.950 293.100 232.050 295.200 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 196.950 280.950 199.050 283.050 ;
        RECT 205.950 280.950 208.050 283.050 ;
        RECT 193.950 259.950 196.050 262.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 178.950 253.950 181.050 256.050 ;
        RECT 185.400 255.900 186.600 256.950 ;
        RECT 175.950 226.950 178.050 229.050 ;
        RECT 163.950 220.950 166.050 223.050 ;
        RECT 172.950 220.950 175.050 223.050 ;
        RECT 164.400 217.050 165.600 220.950 ;
        RECT 163.950 214.950 166.050 217.050 ;
        RECT 169.950 216.000 172.050 220.050 ;
        RECT 179.400 217.200 180.600 253.950 ;
        RECT 184.950 253.800 187.050 255.900 ;
        RECT 191.400 250.050 192.600 256.950 ;
        RECT 190.950 247.950 193.050 250.050 ;
        RECT 197.400 232.050 198.600 280.950 ;
        RECT 208.950 268.950 211.050 271.050 ;
        RECT 199.950 262.950 202.050 265.050 ;
        RECT 200.400 259.050 201.600 262.950 ;
        RECT 209.400 259.050 210.600 268.950 ;
        RECT 215.400 265.050 216.600 289.950 ;
        RECT 224.400 268.050 225.600 292.950 ;
        RECT 230.400 292.050 231.600 293.100 ;
        RECT 236.400 292.050 237.600 301.950 ;
        RECT 251.400 300.600 252.600 319.950 ;
        RECT 256.950 313.950 259.050 316.050 ;
        RECT 257.400 301.050 258.600 313.950 ;
        RECT 248.400 299.400 252.600 300.600 ;
        RECT 241.950 293.100 244.050 295.200 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 229.950 280.950 232.050 283.050 ;
        RECT 217.950 265.950 220.050 268.050 ;
        RECT 223.950 265.950 226.050 268.050 ;
        RECT 214.950 262.950 217.050 265.050 ;
        RECT 199.950 256.950 202.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 208.950 256.950 211.050 259.050 ;
        RECT 214.950 256.950 217.050 259.050 ;
        RECT 206.400 250.050 207.600 256.950 ;
        RECT 205.950 247.950 208.050 250.050 ;
        RECT 211.950 238.950 214.050 241.050 ;
        RECT 196.950 229.950 199.050 232.050 ;
        RECT 184.950 217.950 187.050 223.050 ;
        RECT 199.950 220.950 202.050 223.050 ;
        RECT 205.950 220.950 208.050 223.050 ;
        RECT 178.950 216.600 181.050 217.200 ;
        RECT 170.400 214.050 171.600 216.000 ;
        RECT 176.400 215.400 181.050 216.600 ;
        RECT 176.400 214.050 177.600 215.400 ;
        RECT 178.950 215.100 181.050 215.400 ;
        RECT 185.400 214.050 186.600 217.950 ;
        RECT 190.950 215.100 193.050 217.200 ;
        RECT 191.400 214.050 192.600 215.100 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 184.950 211.950 187.050 214.050 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 163.950 208.950 166.050 211.050 ;
        RECT 160.950 198.600 163.050 199.050 ;
        RECT 158.400 197.400 163.050 198.600 ;
        RECT 154.950 193.950 157.050 196.050 ;
        RECT 154.950 181.950 157.050 184.050 ;
        RECT 151.950 172.950 154.050 175.050 ;
        RECT 148.950 148.950 151.050 151.050 ;
        RECT 155.400 142.050 156.600 181.950 ;
        RECT 158.400 175.050 159.600 197.400 ;
        RECT 160.950 196.950 163.050 197.400 ;
        RECT 164.400 193.050 165.600 208.950 ;
        RECT 167.400 202.050 168.600 211.950 ;
        RECT 173.400 210.000 174.600 211.950 ;
        RECT 188.400 210.000 189.600 211.950 ;
        RECT 172.950 205.950 175.050 210.000 ;
        RECT 187.950 205.950 190.050 210.000 ;
        RECT 166.950 199.950 169.050 202.050 ;
        RECT 187.950 196.950 190.050 199.050 ;
        RECT 163.950 190.950 166.050 193.050 ;
        RECT 169.950 190.950 172.050 193.050 ;
        RECT 178.950 190.950 181.050 193.050 ;
        RECT 163.950 182.100 166.050 184.200 ;
        RECT 164.400 181.050 165.600 182.100 ;
        RECT 170.400 181.050 171.600 190.950 ;
        RECT 163.950 178.950 166.050 181.050 ;
        RECT 166.950 178.950 169.050 181.050 ;
        RECT 169.950 178.950 172.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 160.950 175.950 163.050 178.050 ;
        RECT 157.950 172.950 160.050 175.050 ;
        RECT 157.950 148.950 160.050 151.050 ;
        RECT 151.950 137.100 154.050 142.050 ;
        RECT 154.950 139.950 157.050 142.050 ;
        RECT 152.400 136.050 153.600 137.100 ;
        RECT 158.400 136.050 159.600 148.950 ;
        RECT 161.400 148.050 162.600 175.950 ;
        RECT 167.400 163.050 168.600 178.950 ;
        RECT 173.400 177.000 174.600 178.950 ;
        RECT 172.950 172.950 175.050 177.000 ;
        RECT 179.400 175.050 180.600 190.950 ;
        RECT 188.400 181.050 189.600 196.950 ;
        RECT 194.400 190.050 195.600 211.950 ;
        RECT 200.400 208.050 201.600 220.950 ;
        RECT 199.950 205.950 202.050 208.050 ;
        RECT 202.950 193.950 205.050 196.050 ;
        RECT 193.950 187.950 196.050 190.050 ;
        RECT 199.950 187.950 202.050 190.050 ;
        RECT 193.950 182.100 196.050 184.200 ;
        RECT 194.400 181.050 195.600 182.100 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 185.400 177.000 186.600 178.950 ;
        RECT 178.950 172.950 181.050 175.050 ;
        RECT 184.950 172.950 187.050 177.000 ;
        RECT 191.400 169.050 192.600 178.950 ;
        RECT 196.950 175.950 199.050 178.050 ;
        RECT 190.950 166.950 193.050 169.050 ;
        RECT 191.400 163.050 192.600 166.950 ;
        RECT 166.950 160.950 169.050 163.050 ;
        RECT 190.950 160.950 193.050 163.050 ;
        RECT 178.950 148.950 181.050 151.050 ;
        RECT 160.950 145.950 163.050 148.050 ;
        RECT 161.400 142.050 162.600 145.950 ;
        RECT 179.400 142.050 180.600 148.950 ;
        RECT 184.950 145.950 187.050 148.050 ;
        RECT 160.950 139.950 163.050 142.050 ;
        RECT 163.950 139.950 166.050 142.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 157.950 133.950 160.050 136.050 ;
        RECT 142.950 127.950 145.050 130.050 ;
        RECT 139.950 115.950 142.050 118.050 ;
        RECT 124.800 109.950 126.900 112.050 ;
        RECT 127.950 109.950 130.050 112.050 ;
        RECT 121.950 103.950 124.050 106.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 110.400 99.900 111.600 100.950 ;
        RECT 109.950 97.800 112.050 99.900 ;
        RECT 100.950 94.950 103.050 97.050 ;
        RECT 116.400 94.050 117.600 100.950 ;
        RECT 115.950 91.950 118.050 94.050 ;
        RECT 125.400 88.050 126.600 109.950 ;
        RECT 124.950 85.950 127.050 88.050 ;
        RECT 118.950 70.950 121.050 73.050 ;
        RECT 103.950 59.100 106.050 61.200 ;
        RECT 109.950 59.100 112.050 61.200 ;
        RECT 104.400 58.050 105.600 59.100 ;
        RECT 110.400 58.050 111.600 59.100 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 100.950 52.950 103.050 55.050 ;
        RECT 107.400 54.000 108.600 55.950 ;
        RECT 97.950 49.950 100.050 52.050 ;
        RECT 101.400 49.050 102.600 52.950 ;
        RECT 106.950 49.950 109.050 54.000 ;
        RECT 100.950 46.950 103.050 49.050 ;
        RECT 91.950 43.950 94.050 46.050 ;
        RECT 97.950 40.950 100.050 43.050 ;
        RECT 88.950 31.950 91.050 34.050 ;
        RECT 89.400 21.900 90.600 31.950 ;
        RECT 98.400 25.050 99.600 40.950 ;
        RECT 109.950 37.950 112.050 40.050 ;
        RECT 110.400 30.600 111.600 37.950 ;
        RECT 113.400 34.050 114.600 55.950 ;
        RECT 119.400 55.050 120.600 70.950 ;
        RECT 128.400 70.050 129.600 109.950 ;
        RECT 149.400 106.200 150.600 133.950 ;
        RECT 155.400 132.000 156.600 133.950 ;
        RECT 154.950 127.950 157.050 132.000 ;
        RECT 164.400 121.050 165.600 139.950 ;
        RECT 172.950 138.000 175.050 142.050 ;
        RECT 178.950 138.000 181.050 142.050 ;
        RECT 173.400 136.050 174.600 138.000 ;
        RECT 179.400 136.050 180.600 138.000 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 172.950 133.950 175.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 170.400 132.900 171.600 133.950 ;
        RECT 169.950 130.800 172.050 132.900 ;
        RECT 163.950 118.950 166.050 121.050 ;
        RECT 172.950 118.950 175.050 121.050 ;
        RECT 163.950 109.950 166.050 112.050 ;
        RECT 133.950 104.100 136.050 106.200 ;
        RECT 139.950 104.100 142.050 106.200 ;
        RECT 148.950 104.100 151.050 106.200 ;
        RECT 157.950 104.100 160.050 106.200 ;
        RECT 134.400 103.050 135.600 104.100 ;
        RECT 140.400 103.050 141.600 104.100 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 136.950 100.950 139.050 103.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 130.950 97.950 133.050 100.050 ;
        RECT 137.400 99.900 138.600 100.950 ;
        RECT 131.400 82.050 132.600 97.950 ;
        RECT 136.950 97.800 139.050 99.900 ;
        RECT 137.400 91.050 138.600 97.800 ;
        RECT 136.950 88.950 139.050 91.050 ;
        RECT 143.400 88.050 144.600 100.950 ;
        RECT 149.400 99.600 150.600 104.100 ;
        RECT 158.400 103.050 159.600 104.100 ;
        RECT 164.400 103.050 165.600 109.950 ;
        RECT 169.950 103.950 172.050 106.050 ;
        RECT 154.950 100.950 157.050 103.050 ;
        RECT 157.950 100.950 160.050 103.050 ;
        RECT 160.950 100.950 163.050 103.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 155.400 99.600 156.600 100.950 ;
        RECT 149.400 98.400 156.600 99.600 ;
        RECT 161.400 88.050 162.600 100.950 ;
        RECT 142.950 85.950 145.050 88.050 ;
        RECT 160.950 85.950 163.050 88.050 ;
        RECT 130.950 79.950 133.050 82.050 ;
        RECT 127.950 67.950 130.050 70.050 ;
        RECT 131.400 63.600 132.600 79.950 ;
        RECT 170.400 79.050 171.600 103.950 ;
        RECT 173.400 94.050 174.600 118.950 ;
        RECT 176.400 112.050 177.600 133.950 ;
        RECT 185.400 132.900 186.600 145.950 ;
        RECT 193.950 142.950 196.050 145.050 ;
        RECT 194.400 136.050 195.600 142.950 ;
        RECT 197.400 142.050 198.600 175.950 ;
        RECT 200.400 157.050 201.600 187.950 ;
        RECT 203.400 175.050 204.600 193.950 ;
        RECT 206.400 177.900 207.600 220.950 ;
        RECT 212.400 214.050 213.600 238.950 ;
        RECT 215.400 223.050 216.600 256.950 ;
        RECT 218.400 223.050 219.600 265.950 ;
        RECT 223.950 260.100 226.050 262.200 ;
        RECT 224.400 259.050 225.600 260.100 ;
        RECT 230.400 259.050 231.600 280.950 ;
        RECT 233.400 274.050 234.600 289.950 ;
        RECT 232.950 271.950 235.050 274.050 ;
        RECT 238.950 271.950 241.050 274.050 ;
        RECT 235.950 268.950 238.050 271.050 ;
        RECT 236.400 262.050 237.600 268.950 ;
        RECT 235.950 259.950 238.050 262.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 227.400 247.050 228.600 256.950 ;
        RECT 233.400 255.900 234.600 256.950 ;
        RECT 232.950 253.800 235.050 255.900 ;
        RECT 226.950 244.950 229.050 247.050 ;
        RECT 239.400 238.050 240.600 271.950 ;
        RECT 242.400 268.050 243.600 293.100 ;
        RECT 248.400 292.050 249.600 299.400 ;
        RECT 256.950 298.950 259.050 301.050 ;
        RECT 253.950 293.100 256.050 295.200 ;
        RECT 254.400 292.050 255.600 293.100 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 250.950 289.950 253.050 292.050 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 244.950 286.950 247.050 289.050 ;
        RECT 241.950 265.950 244.050 268.050 ;
        RECT 241.950 262.800 244.050 264.900 ;
        RECT 242.400 250.050 243.600 262.800 ;
        RECT 245.400 262.050 246.600 286.950 ;
        RECT 247.950 271.950 250.050 274.050 ;
        RECT 244.950 259.950 247.050 262.050 ;
        RECT 248.400 259.050 249.600 271.950 ;
        RECT 251.400 271.050 252.600 289.950 ;
        RECT 256.950 286.950 259.050 289.050 ;
        RECT 260.400 288.600 261.600 322.950 ;
        RECT 263.400 295.050 264.600 328.950 ;
        RECT 272.400 297.600 273.600 328.950 ;
        RECT 275.400 316.050 276.600 334.950 ;
        RECT 277.800 331.950 279.900 334.050 ;
        RECT 280.950 331.950 283.050 334.050 ;
        RECT 287.400 333.900 288.600 334.950 ;
        RECT 296.400 334.050 297.600 334.950 ;
        RECT 274.950 313.950 277.050 316.050 ;
        RECT 269.400 296.400 273.600 297.600 ;
        RECT 262.950 292.950 265.050 295.050 ;
        RECT 269.400 292.050 270.600 296.400 ;
        RECT 274.950 294.000 277.050 298.050 ;
        RECT 278.400 295.050 279.600 331.950 ;
        RECT 275.400 292.050 276.600 294.000 ;
        RECT 277.950 292.950 280.050 295.050 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 268.950 289.950 271.050 292.050 ;
        RECT 271.950 289.950 274.050 292.050 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 266.400 288.600 267.600 289.950 ;
        RECT 260.400 287.400 267.600 288.600 ;
        RECT 253.950 280.950 256.050 283.050 ;
        RECT 254.400 274.050 255.600 280.950 ;
        RECT 257.400 280.050 258.600 286.950 ;
        RECT 262.950 283.950 265.050 286.050 ;
        RECT 266.400 285.600 267.600 287.400 ;
        RECT 266.400 284.400 270.600 285.600 ;
        RECT 256.950 277.950 259.050 280.050 ;
        RECT 253.950 271.950 256.050 274.050 ;
        RECT 250.950 268.950 253.050 271.050 ;
        RECT 253.950 261.000 256.050 265.050 ;
        RECT 263.400 262.050 264.600 283.950 ;
        RECT 269.400 280.050 270.600 284.400 ;
        RECT 265.800 277.950 267.900 280.050 ;
        RECT 268.950 277.950 271.050 280.050 ;
        RECT 254.400 259.050 255.600 261.000 ;
        RECT 262.950 259.950 265.050 262.050 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 250.950 256.950 253.050 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 244.950 253.950 247.050 256.050 ;
        RECT 251.400 255.900 252.600 256.950 ;
        RECT 241.950 247.950 244.050 250.050 ;
        RECT 238.950 235.950 241.050 238.050 ;
        RECT 223.950 229.950 226.050 232.050 ;
        RECT 214.950 220.950 217.050 223.050 ;
        RECT 218.400 220.950 223.050 223.050 ;
        RECT 218.400 214.050 219.600 220.950 ;
        RECT 224.400 220.050 225.600 229.950 ;
        RECT 245.400 229.050 246.600 253.950 ;
        RECT 250.950 253.800 253.050 255.900 ;
        RECT 257.400 255.000 258.600 256.950 ;
        RECT 262.950 256.800 265.050 258.900 ;
        RECT 256.950 250.950 259.050 255.000 ;
        RECT 259.950 253.950 262.050 256.050 ;
        RECT 250.950 247.950 253.050 250.050 ;
        RECT 232.950 226.950 235.050 229.050 ;
        RECT 241.800 226.950 243.900 229.050 ;
        RECT 244.950 226.950 247.050 229.050 ;
        RECT 226.950 223.950 229.050 226.050 ;
        RECT 223.950 217.950 226.050 220.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 214.950 211.950 217.050 214.050 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 215.400 210.900 216.600 211.950 ;
        RECT 227.400 210.900 228.600 223.950 ;
        RECT 233.400 214.050 234.600 226.950 ;
        RECT 238.950 223.950 241.050 226.050 ;
        RECT 239.400 214.050 240.600 223.950 ;
        RECT 242.400 220.050 243.600 226.950 ;
        RECT 241.950 217.950 244.050 220.050 ;
        RECT 247.950 217.950 250.050 220.050 ;
        RECT 232.950 211.950 235.050 214.050 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 214.950 208.800 217.050 210.900 ;
        RECT 226.950 208.800 229.050 210.900 ;
        RECT 236.400 210.000 237.600 211.950 ;
        RECT 242.400 210.900 243.600 211.950 ;
        RECT 217.950 205.950 223.050 208.050 ;
        RECT 227.400 190.050 228.600 208.800 ;
        RECT 229.950 205.950 235.050 208.050 ;
        RECT 235.950 205.950 238.050 210.000 ;
        RECT 241.950 208.800 244.050 210.900 ;
        RECT 232.950 193.950 235.050 196.050 ;
        RECT 226.950 187.950 229.050 190.050 ;
        RECT 214.950 182.100 217.050 184.200 ;
        RECT 215.400 181.050 216.600 182.100 ;
        RECT 233.400 181.050 234.600 193.950 ;
        RECT 242.400 189.600 243.600 208.800 ;
        RECT 242.400 188.400 246.600 189.600 ;
        RECT 241.950 184.950 244.050 187.050 ;
        RECT 242.400 181.050 243.600 184.950 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 232.950 178.950 235.050 181.050 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 212.400 177.900 213.600 178.950 ;
        RECT 205.950 175.800 208.050 177.900 ;
        RECT 211.950 175.800 214.050 177.900 ;
        RECT 218.400 177.000 219.600 178.950 ;
        RECT 202.950 172.950 205.050 175.050 ;
        RECT 212.400 166.050 213.600 175.800 ;
        RECT 217.950 172.950 220.050 177.000 ;
        RECT 220.950 175.950 223.050 178.050 ;
        RECT 221.400 169.050 222.600 175.950 ;
        RECT 220.950 166.950 223.050 169.050 ;
        RECT 227.400 166.050 228.600 178.950 ;
        RECT 211.950 163.950 214.050 166.050 ;
        RECT 226.950 163.950 229.050 166.050 ;
        RECT 199.950 154.950 202.050 157.050 ;
        RECT 200.400 145.050 201.600 154.950 ;
        RECT 236.400 148.050 237.600 178.950 ;
        RECT 241.950 160.950 244.050 163.050 ;
        RECT 205.950 147.600 208.050 148.050 ;
        RECT 205.950 146.400 210.600 147.600 ;
        RECT 205.950 145.950 208.050 146.400 ;
        RECT 199.950 142.950 202.050 145.050 ;
        RECT 196.950 139.950 199.050 142.050 ;
        RECT 206.400 139.200 207.600 145.950 ;
        RECT 199.950 137.100 202.050 139.200 ;
        RECT 205.950 137.100 208.050 139.200 ;
        RECT 200.400 136.050 201.600 137.100 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 196.950 133.950 199.050 136.050 ;
        RECT 199.950 133.950 202.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 197.400 132.900 198.600 133.950 ;
        RECT 184.950 130.800 187.050 132.900 ;
        RECT 196.950 130.800 199.050 132.900 ;
        RECT 175.950 109.950 178.050 112.050 ;
        RECT 184.950 109.950 187.050 112.050 ;
        RECT 193.950 109.950 196.050 112.050 ;
        RECT 185.400 106.200 186.600 109.950 ;
        RECT 178.950 104.100 181.050 106.200 ;
        RECT 184.950 104.100 187.050 106.200 ;
        RECT 179.400 103.050 180.600 104.100 ;
        RECT 185.400 103.050 186.600 104.100 ;
        RECT 190.950 103.950 193.050 109.050 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 182.400 99.000 183.600 100.950 ;
        RECT 188.400 99.900 189.600 100.950 ;
        RECT 194.400 99.900 195.600 109.950 ;
        RECT 203.400 106.200 204.600 133.950 ;
        RECT 209.400 127.050 210.600 146.400 ;
        RECT 235.950 145.950 238.050 148.050 ;
        RECT 223.950 138.000 226.050 142.050 ;
        RECT 232.950 139.950 238.050 142.050 ;
        RECT 224.400 136.050 225.600 138.000 ;
        RECT 229.950 137.100 232.050 139.200 ;
        RECT 242.400 139.050 243.600 160.950 ;
        RECT 245.400 154.050 246.600 188.400 ;
        RECT 244.950 151.950 247.050 154.050 ;
        RECT 244.950 142.950 247.050 145.050 ;
        RECT 245.400 139.200 246.600 142.950 ;
        RECT 248.400 142.050 249.600 217.950 ;
        RECT 251.400 211.050 252.600 247.950 ;
        RECT 260.400 244.050 261.600 253.950 ;
        RECT 263.400 247.050 264.600 256.800 ;
        RECT 266.400 250.050 267.600 277.950 ;
        RECT 272.400 274.050 273.600 289.950 ;
        RECT 271.950 271.950 274.050 274.050 ;
        RECT 274.950 261.000 277.050 265.050 ;
        RECT 275.400 259.050 276.600 261.000 ;
        RECT 281.400 259.050 282.600 331.950 ;
        RECT 286.950 331.800 289.050 333.900 ;
        RECT 292.950 331.950 297.600 334.050 ;
        RECT 298.950 331.950 301.050 334.050 ;
        RECT 283.950 325.950 286.050 331.050 ;
        RECT 296.400 325.050 297.600 331.950 ;
        RECT 295.950 322.950 298.050 325.050 ;
        RECT 295.950 319.800 298.050 321.900 ;
        RECT 296.400 313.050 297.600 319.800 ;
        RECT 299.400 316.050 300.600 331.950 ;
        RECT 302.400 316.050 303.600 340.800 ;
        RECT 305.400 325.050 306.600 379.950 ;
        RECT 314.400 376.050 315.600 412.800 ;
        RECT 316.950 409.950 319.050 412.050 ;
        RECT 323.400 411.000 324.600 412.950 ;
        RECT 317.400 387.600 318.600 409.950 ;
        RECT 322.950 406.950 325.050 411.000 ;
        RECT 332.400 409.050 333.600 422.400 ;
        RECT 325.950 406.950 328.050 409.050 ;
        RECT 331.950 406.950 334.050 409.050 ;
        RECT 322.950 397.950 325.050 400.050 ;
        RECT 319.950 387.600 322.050 388.050 ;
        RECT 317.400 386.400 322.050 387.600 ;
        RECT 319.950 385.950 322.050 386.400 ;
        RECT 320.400 382.050 321.600 385.950 ;
        RECT 319.950 379.950 322.050 382.050 ;
        RECT 307.950 375.600 312.000 376.050 ;
        RECT 307.950 373.950 312.600 375.600 ;
        RECT 313.950 373.950 316.050 376.050 ;
        RECT 311.400 370.050 312.600 373.950 ;
        RECT 319.950 372.000 322.050 376.050 ;
        RECT 323.400 373.050 324.600 397.950 ;
        RECT 320.400 370.050 321.600 372.000 ;
        RECT 322.950 370.950 325.050 373.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 314.400 366.900 315.600 367.950 ;
        RECT 313.950 364.800 316.050 366.900 ;
        RECT 307.950 358.950 310.050 361.050 ;
        RECT 308.400 340.050 309.600 358.950 ;
        RECT 314.400 355.050 315.600 364.800 ;
        RECT 313.800 352.950 315.900 355.050 ;
        RECT 316.950 352.950 319.050 355.050 ;
        RECT 317.400 349.050 318.600 352.950 ;
        RECT 316.950 346.950 319.050 349.050 ;
        RECT 326.400 343.050 327.600 406.950 ;
        RECT 331.950 391.950 334.050 394.050 ;
        RECT 328.950 373.950 331.050 376.050 ;
        RECT 329.400 346.050 330.600 373.950 ;
        RECT 332.400 373.050 333.600 391.950 ;
        RECT 335.400 387.600 336.600 430.950 ;
        RECT 337.950 424.950 340.050 427.050 ;
        RECT 338.400 418.050 339.600 424.950 ;
        RECT 341.400 421.050 342.600 442.950 ;
        RECT 347.400 427.050 348.600 445.950 ;
        RECT 353.400 444.000 354.600 445.950 ;
        RECT 349.950 439.950 352.050 442.050 ;
        RECT 352.950 439.950 355.050 444.000 ;
        RECT 355.950 442.950 358.050 445.050 ;
        RECT 350.400 430.050 351.600 439.950 ;
        RECT 356.400 438.600 357.600 442.950 ;
        RECT 359.400 442.050 360.600 457.950 ;
        RECT 358.950 439.950 361.050 442.050 ;
        RECT 353.400 437.400 357.600 438.600 ;
        RECT 349.950 427.950 352.050 430.050 ;
        RECT 346.950 424.950 349.050 427.050 ;
        RECT 343.950 421.950 346.050 424.050 ;
        RECT 340.950 418.950 343.050 421.050 ;
        RECT 337.950 415.950 340.050 418.050 ;
        RECT 344.400 415.050 345.600 421.950 ;
        RECT 353.400 418.050 354.600 437.400 ;
        RECT 362.400 436.050 363.600 463.950 ;
        RECT 365.400 439.050 366.600 481.950 ;
        RECT 368.400 472.050 369.600 490.950 ;
        RECT 370.950 487.950 373.050 490.050 ;
        RECT 367.950 469.950 370.050 472.050 ;
        RECT 371.400 466.050 372.600 487.950 ;
        RECT 374.400 487.050 375.600 499.950 ;
        RECT 373.950 484.950 376.050 487.050 ;
        RECT 377.400 478.050 378.600 508.950 ;
        RECT 379.950 502.950 382.050 505.050 ;
        RECT 382.950 502.950 385.050 508.050 ;
        RECT 376.950 475.950 379.050 478.050 ;
        RECT 370.950 463.950 373.050 466.050 ;
        RECT 370.950 454.950 373.050 457.050 ;
        RECT 371.400 448.050 372.600 454.950 ;
        RECT 380.400 450.600 381.600 502.950 ;
        RECT 389.400 502.050 390.600 520.950 ;
        RECT 392.400 519.600 393.600 523.950 ;
        RECT 401.400 522.600 402.600 527.400 ;
        RECT 398.400 521.400 402.600 522.600 ;
        RECT 392.400 518.400 396.600 519.600 ;
        RECT 395.400 514.050 396.600 518.400 ;
        RECT 394.950 511.950 397.050 514.050 ;
        RECT 382.950 499.800 385.050 501.900 ;
        RECT 388.950 499.950 391.050 502.050 ;
        RECT 383.400 496.050 384.600 499.800 ;
        RECT 382.950 493.950 385.050 496.050 ;
        RECT 388.950 494.100 391.050 496.200 ;
        RECT 395.400 496.050 396.600 511.950 ;
        RECT 389.400 493.050 390.600 494.100 ;
        RECT 394.950 493.950 397.050 496.050 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 388.950 490.950 391.050 493.050 ;
        RECT 391.950 490.950 394.050 493.050 ;
        RECT 386.400 489.900 387.600 490.950 ;
        RECT 385.950 487.800 388.050 489.900 ;
        RECT 392.400 489.000 393.600 490.950 ;
        RECT 384.000 486.750 387.000 487.050 ;
        RECT 382.950 484.950 388.050 486.750 ;
        RECT 391.950 484.950 394.050 489.000 ;
        RECT 394.950 487.950 397.050 490.050 ;
        RECT 382.950 484.650 385.050 484.950 ;
        RECT 385.950 484.650 388.050 484.950 ;
        RECT 388.950 472.950 391.050 475.050 ;
        RECT 385.950 466.950 388.050 469.050 ;
        RECT 386.400 451.050 387.600 466.950 ;
        RECT 380.400 449.400 384.600 450.600 ;
        RECT 370.950 445.950 373.050 448.050 ;
        RECT 376.950 445.950 379.050 448.050 ;
        RECT 377.400 444.900 378.600 445.950 ;
        RECT 376.950 442.800 379.050 444.900 ;
        RECT 367.950 439.950 370.050 442.050 ;
        RECT 364.950 436.950 367.050 439.050 ;
        RECT 361.950 433.950 364.050 436.050 ;
        RECT 358.950 427.950 361.050 430.050 ;
        RECT 352.950 415.950 355.050 418.050 ;
        RECT 359.400 417.600 360.600 427.950 ;
        RECT 368.400 421.050 369.600 439.950 ;
        RECT 370.950 436.950 373.050 439.050 ;
        RECT 367.950 418.950 370.050 421.050 ;
        RECT 361.950 417.600 364.050 418.200 ;
        RECT 359.400 416.400 364.050 417.600 ;
        RECT 361.950 416.100 364.050 416.400 ;
        RECT 362.400 415.050 363.600 416.100 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 355.950 412.950 358.050 415.050 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 337.950 409.950 340.050 412.050 ;
        RECT 338.400 406.050 339.600 409.950 ;
        RECT 337.950 403.950 340.050 406.050 ;
        RECT 341.400 397.050 342.600 412.950 ;
        RECT 347.400 408.600 348.600 412.950 ;
        RECT 349.950 409.950 352.050 412.050 ;
        RECT 344.400 407.400 348.600 408.600 ;
        RECT 340.950 394.950 343.050 397.050 ;
        RECT 335.400 386.400 339.600 387.600 ;
        RECT 334.950 382.950 337.050 385.050 ;
        RECT 331.950 370.950 334.050 373.050 ;
        RECT 335.400 370.050 336.600 382.950 ;
        RECT 338.400 373.050 339.600 386.400 ;
        RECT 344.400 382.050 345.600 407.400 ;
        RECT 346.950 388.950 349.050 391.050 ;
        RECT 343.950 379.950 346.050 382.050 ;
        RECT 337.950 370.950 340.050 373.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 337.950 364.950 340.050 367.050 ;
        RECT 341.400 366.600 342.600 367.950 ;
        RECT 341.400 365.400 345.600 366.600 ;
        RECT 331.950 361.950 334.050 364.050 ;
        RECT 328.950 343.950 331.050 346.050 ;
        RECT 325.950 340.950 328.050 343.050 ;
        RECT 307.950 337.950 310.050 340.050 ;
        RECT 313.950 338.100 316.050 340.200 ;
        RECT 314.400 337.050 315.600 338.100 ;
        RECT 322.800 337.950 324.900 340.050 ;
        RECT 310.950 334.950 313.050 337.050 ;
        RECT 313.950 334.950 316.050 337.050 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 307.950 331.950 310.050 334.050 ;
        RECT 311.400 333.900 312.600 334.950 ;
        RECT 304.950 322.950 307.050 325.050 ;
        RECT 298.800 313.950 300.900 316.050 ;
        RECT 301.950 313.950 304.050 316.050 ;
        RECT 295.950 310.950 298.050 313.050 ;
        RECT 289.950 293.100 292.050 298.050 ;
        RECT 297.000 294.600 301.050 295.050 ;
        RECT 290.400 292.050 291.600 293.100 ;
        RECT 296.400 292.950 301.050 294.600 ;
        RECT 296.400 292.050 297.600 292.950 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 293.400 288.900 294.600 289.950 ;
        RECT 292.950 286.800 295.050 288.900 ;
        RECT 298.950 286.950 301.050 289.050 ;
        RECT 295.950 280.950 298.050 283.050 ;
        RECT 289.950 271.950 292.050 274.050 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 283.950 256.950 286.050 259.050 ;
        RECT 272.400 255.000 273.600 256.950 ;
        RECT 271.950 250.950 274.050 255.000 ;
        RECT 265.950 247.950 268.050 250.050 ;
        RECT 262.950 244.950 265.050 247.050 ;
        RECT 259.950 241.950 262.050 244.050 ;
        RECT 265.800 235.950 267.900 238.050 ;
        RECT 268.950 235.950 271.050 238.050 ;
        RECT 258.000 219.600 262.050 220.050 ;
        RECT 257.400 217.950 262.050 219.600 ;
        RECT 257.400 217.200 258.600 217.950 ;
        RECT 256.950 215.100 259.050 217.200 ;
        RECT 257.400 214.050 258.600 215.100 ;
        RECT 256.950 211.950 259.050 214.050 ;
        RECT 259.950 211.950 262.050 214.050 ;
        RECT 250.950 208.950 253.050 211.050 ;
        RECT 260.400 210.900 261.600 211.950 ;
        RECT 259.950 208.800 262.050 210.900 ;
        RECT 266.400 196.050 267.600 235.950 ;
        RECT 269.400 229.050 270.600 235.950 ;
        RECT 278.400 235.050 279.600 256.950 ;
        RECT 280.950 250.950 283.050 253.050 ;
        RECT 277.950 232.950 280.050 235.050 ;
        RECT 268.950 226.950 271.050 229.050 ;
        RECT 277.950 226.950 280.050 229.050 ;
        RECT 269.400 217.050 270.600 226.950 ;
        RECT 278.400 220.050 279.600 226.950 ;
        RECT 281.400 223.050 282.600 250.950 ;
        RECT 280.950 220.950 283.050 223.050 ;
        RECT 284.400 220.050 285.600 256.950 ;
        RECT 290.400 255.900 291.600 271.950 ;
        RECT 292.950 262.950 295.050 265.050 ;
        RECT 289.950 253.800 292.050 255.900 ;
        RECT 286.950 244.950 289.050 247.050 ;
        RECT 287.400 232.050 288.600 244.950 ;
        RECT 293.400 241.050 294.600 262.950 ;
        RECT 296.400 262.050 297.600 280.950 ;
        RECT 299.400 274.050 300.600 286.950 ;
        RECT 298.950 271.950 301.050 274.050 ;
        RECT 302.400 265.200 303.600 313.950 ;
        RECT 308.400 297.600 309.600 331.950 ;
        RECT 310.950 331.800 313.050 333.900 ;
        RECT 317.400 327.600 318.600 334.950 ;
        RECT 317.400 326.400 321.600 327.600 ;
        RECT 310.950 322.950 313.050 325.050 ;
        RECT 311.400 304.050 312.600 322.950 ;
        RECT 316.950 310.950 319.050 313.050 ;
        RECT 310.950 301.950 313.050 304.050 ;
        RECT 317.400 298.050 318.600 310.950 ;
        RECT 305.400 296.400 309.600 297.600 ;
        RECT 305.400 283.050 306.600 296.400 ;
        RECT 310.950 294.600 313.050 298.050 ;
        RECT 316.950 295.950 319.050 298.050 ;
        RECT 320.400 295.200 321.600 326.400 ;
        RECT 323.400 313.050 324.600 337.950 ;
        RECT 325.950 337.800 328.050 339.900 ;
        RECT 326.400 327.600 327.600 337.800 ;
        RECT 332.400 337.050 333.600 361.950 ;
        RECT 338.400 343.050 339.600 364.950 ;
        RECT 344.400 343.050 345.600 365.400 ;
        RECT 347.400 358.050 348.600 388.950 ;
        RECT 350.400 373.050 351.600 409.950 ;
        RECT 356.400 397.050 357.600 412.950 ;
        RECT 365.400 411.900 366.600 412.950 ;
        RECT 364.950 409.800 367.050 411.900 ;
        RECT 367.950 409.950 370.050 412.050 ;
        RECT 361.950 406.950 364.050 409.050 ;
        RECT 355.950 394.950 358.050 397.050 ;
        RECT 362.400 391.050 363.600 406.950 ;
        RECT 364.950 403.950 367.050 406.050 ;
        RECT 368.400 405.600 369.600 409.950 ;
        RECT 371.400 409.050 372.600 436.950 ;
        RECT 373.950 433.950 376.050 436.050 ;
        RECT 370.950 406.950 373.050 409.050 ;
        RECT 368.400 404.400 372.600 405.600 ;
        RECT 361.950 388.950 364.050 391.050 ;
        RECT 361.950 385.800 364.050 387.900 ;
        RECT 349.950 370.950 352.050 373.050 ;
        RECT 352.950 372.000 355.050 376.050 ;
        RECT 362.400 373.050 363.600 385.800 ;
        RECT 365.400 385.050 366.600 403.950 ;
        RECT 367.950 400.950 370.050 403.050 ;
        RECT 364.950 382.950 367.050 385.050 ;
        RECT 353.400 370.050 354.600 372.000 ;
        RECT 361.950 370.950 364.050 373.050 ;
        RECT 364.950 370.950 367.050 373.050 ;
        RECT 352.950 367.950 355.050 370.050 ;
        RECT 358.950 367.950 361.050 370.050 ;
        RECT 349.950 364.950 352.050 367.050 ;
        RECT 359.400 366.900 360.600 367.950 ;
        RECT 365.400 366.900 366.600 370.950 ;
        RECT 350.400 361.050 351.600 364.950 ;
        RECT 358.950 364.800 361.050 366.900 ;
        RECT 364.950 364.800 367.050 366.900 ;
        RECT 349.950 358.950 352.050 361.050 ;
        RECT 346.950 355.950 349.050 358.050 ;
        RECT 352.950 349.950 355.050 352.050 ;
        RECT 337.950 340.950 340.050 343.050 ;
        RECT 343.950 340.950 346.050 343.050 ;
        RECT 338.400 338.400 345.600 339.600 ;
        RECT 338.400 337.050 339.600 338.400 ;
        RECT 331.950 334.950 334.050 337.050 ;
        RECT 334.950 334.950 337.050 337.050 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 328.950 331.050 331.050 334.050 ;
        RECT 328.800 330.000 331.050 331.050 ;
        RECT 328.800 328.950 330.900 330.000 ;
        RECT 326.400 326.400 330.600 327.600 ;
        RECT 322.950 310.950 325.050 313.050 ;
        RECT 322.950 298.800 325.050 300.900 ;
        RECT 308.400 294.000 313.050 294.600 ;
        RECT 308.400 293.400 312.600 294.000 ;
        RECT 308.400 286.050 309.600 293.400 ;
        RECT 313.950 293.100 316.050 295.200 ;
        RECT 319.950 293.100 322.050 295.200 ;
        RECT 314.400 292.050 315.600 293.100 ;
        RECT 323.400 292.050 324.600 298.800 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 316.950 289.950 319.050 292.050 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 307.950 283.950 310.050 286.050 ;
        RECT 304.950 280.950 307.050 283.050 ;
        RECT 313.950 277.950 316.050 280.050 ;
        RECT 301.950 263.100 304.050 265.200 ;
        RECT 314.400 262.200 315.600 277.950 ;
        RECT 317.400 277.050 318.600 289.950 ;
        RECT 329.400 277.050 330.600 326.400 ;
        RECT 335.400 325.050 336.600 334.950 ;
        RECT 340.950 325.950 343.050 328.050 ;
        RECT 334.950 322.950 337.050 325.050 ;
        RECT 334.950 307.950 337.050 310.050 ;
        RECT 335.400 301.050 336.600 307.950 ;
        RECT 334.950 298.950 337.050 301.050 ;
        RECT 341.400 298.050 342.600 325.950 ;
        RECT 344.400 325.050 345.600 338.400 ;
        RECT 353.400 337.050 354.600 349.950 ;
        RECT 361.800 343.950 363.900 346.050 ;
        RECT 364.950 343.950 367.050 346.050 ;
        RECT 355.950 337.950 358.050 343.050 ;
        RECT 358.950 340.950 361.050 343.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 350.400 331.050 351.600 334.950 ;
        RECT 350.400 330.600 355.050 331.050 ;
        RECT 350.400 329.400 357.600 330.600 ;
        RECT 351.000 328.950 355.050 329.400 ;
        RECT 349.950 325.950 352.050 328.050 ;
        RECT 343.950 322.950 346.050 325.050 ;
        RECT 350.400 304.050 351.600 325.950 ;
        RECT 352.950 322.950 355.050 325.050 ;
        RECT 349.950 301.950 352.050 304.050 ;
        RECT 343.950 298.950 346.050 301.050 ;
        RECT 340.950 295.950 343.050 298.050 ;
        RECT 334.950 293.100 337.050 295.200 ;
        RECT 344.400 294.600 345.600 298.950 ;
        RECT 349.950 295.950 352.050 298.050 ;
        RECT 341.400 293.400 345.600 294.600 ;
        RECT 335.400 292.050 336.600 293.100 ;
        RECT 341.400 292.050 342.600 293.400 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 337.950 289.950 340.050 292.050 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 346.950 289.950 349.050 292.050 ;
        RECT 334.950 283.950 337.050 286.050 ;
        RECT 331.950 277.950 334.050 280.050 ;
        RECT 316.950 274.950 319.050 277.050 ;
        RECT 328.950 274.950 331.050 277.050 ;
        RECT 316.950 265.950 319.050 268.050 ;
        RECT 325.950 265.950 328.050 268.050 ;
        RECT 295.950 259.950 298.050 262.050 ;
        RECT 301.950 259.950 304.050 262.050 ;
        RECT 307.950 260.100 310.050 262.200 ;
        RECT 313.950 260.100 316.050 262.200 ;
        RECT 317.400 262.050 318.600 265.950 ;
        RECT 302.400 259.050 303.600 259.950 ;
        RECT 308.400 259.050 309.600 260.100 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 304.950 256.950 307.050 259.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 299.400 255.900 300.600 256.950 ;
        RECT 298.950 253.800 301.050 255.900 ;
        RECT 305.400 253.050 306.600 256.950 ;
        RECT 305.400 251.400 310.050 253.050 ;
        RECT 306.000 250.950 310.050 251.400 ;
        RECT 310.950 250.950 313.050 256.050 ;
        RECT 314.400 241.050 315.600 260.100 ;
        RECT 316.950 259.950 319.050 262.050 ;
        RECT 319.950 260.100 322.050 262.200 ;
        RECT 320.400 259.050 321.600 260.100 ;
        RECT 326.400 259.050 327.600 265.950 ;
        RECT 332.400 262.050 333.600 277.950 ;
        RECT 331.950 259.950 334.050 262.050 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 322.950 256.950 325.050 259.050 ;
        RECT 325.950 256.950 328.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 316.950 253.950 319.050 256.050 ;
        RECT 323.400 255.900 324.600 256.950 ;
        RECT 329.400 255.900 330.600 256.950 ;
        RECT 292.950 238.950 295.050 241.050 ;
        RECT 313.950 238.950 316.050 241.050 ;
        RECT 286.950 229.950 289.050 232.050 ;
        RECT 289.950 226.950 292.050 229.050 ;
        RECT 317.400 228.600 318.600 253.950 ;
        RECT 322.950 253.800 325.050 255.900 ;
        RECT 328.950 253.800 331.050 255.900 ;
        RECT 319.950 250.950 322.050 253.050 ;
        RECT 320.400 240.600 321.600 250.950 ;
        RECT 323.400 244.050 324.600 253.800 ;
        RECT 322.950 241.950 325.050 244.050 ;
        RECT 320.400 239.400 324.600 240.600 ;
        RECT 323.400 232.050 324.600 239.400 ;
        RECT 322.950 229.950 325.050 232.050 ;
        RECT 319.800 228.600 321.900 229.050 ;
        RECT 317.400 227.400 321.900 228.600 ;
        RECT 319.800 226.950 321.900 227.400 ;
        RECT 271.950 219.600 276.000 220.050 ;
        RECT 271.950 217.950 276.600 219.600 ;
        RECT 277.800 217.950 279.900 220.050 ;
        RECT 268.950 214.950 271.050 217.050 ;
        RECT 275.400 214.050 276.600 217.950 ;
        RECT 280.950 216.000 283.050 219.900 ;
        RECT 283.950 217.950 286.050 220.050 ;
        RECT 281.400 214.050 282.600 216.000 ;
        RECT 286.950 215.100 289.050 217.200 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 280.950 211.950 283.050 214.050 ;
        RECT 272.400 210.900 273.600 211.950 ;
        RECT 271.950 208.800 274.050 210.900 ;
        RECT 278.400 210.000 279.600 211.950 ;
        RECT 277.950 205.950 280.050 210.000 ;
        RECT 287.400 208.050 288.600 215.100 ;
        RECT 290.400 211.050 291.600 226.950 ;
        RECT 307.950 223.950 310.050 226.050 ;
        RECT 295.950 220.950 298.050 223.050 ;
        RECT 296.400 217.050 297.600 220.950 ;
        RECT 295.950 214.950 298.050 217.050 ;
        RECT 301.950 215.100 304.050 217.200 ;
        RECT 302.400 214.050 303.600 215.100 ;
        RECT 308.400 214.050 309.600 223.950 ;
        RECT 320.400 214.050 321.600 226.950 ;
        RECT 322.950 226.800 325.050 228.900 ;
        RECT 323.400 220.050 324.600 226.800 ;
        RECT 322.950 217.950 325.050 220.050 ;
        RECT 325.950 215.100 328.050 217.200 ;
        RECT 329.400 217.050 330.600 253.800 ;
        RECT 335.400 247.050 336.600 283.950 ;
        RECT 338.400 262.050 339.600 289.950 ;
        RECT 347.400 268.050 348.600 289.950 ;
        RECT 350.400 280.050 351.600 295.950 ;
        RECT 349.950 277.950 352.050 280.050 ;
        RECT 346.950 265.950 349.050 268.050 ;
        RECT 337.950 259.950 340.050 262.050 ;
        RECT 343.950 260.100 346.050 262.200 ;
        RECT 344.400 259.050 345.600 260.100 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 337.950 253.950 340.050 256.050 ;
        RECT 334.950 244.950 337.050 247.050 ;
        RECT 338.400 226.050 339.600 253.950 ;
        RECT 341.400 250.050 342.600 256.950 ;
        RECT 347.400 255.900 348.600 256.950 ;
        RECT 346.950 253.800 349.050 255.900 ;
        RECT 340.950 247.950 343.050 250.050 ;
        RECT 343.950 244.950 346.050 247.050 ;
        RECT 344.400 235.050 345.600 244.950 ;
        RECT 346.950 238.950 349.050 241.050 ;
        RECT 343.950 232.950 346.050 235.050 ;
        RECT 331.950 223.950 334.050 226.050 ;
        RECT 337.950 223.950 340.050 226.050 ;
        RECT 326.400 214.050 327.600 215.100 ;
        RECT 328.950 214.950 331.050 217.050 ;
        RECT 298.950 211.950 301.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 307.950 211.950 310.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 289.950 208.950 292.050 211.050 ;
        RECT 295.950 208.950 298.050 211.050 ;
        RECT 286.950 205.950 289.050 208.050 ;
        RECT 271.950 202.950 274.050 205.050 ;
        RECT 272.400 199.050 273.600 202.950 ;
        RECT 296.400 199.050 297.600 208.950 ;
        RECT 299.400 207.600 300.600 211.950 ;
        RECT 305.400 210.900 306.600 211.950 ;
        RECT 304.950 208.800 307.050 210.900 ;
        RECT 313.950 208.800 316.050 210.900 ;
        RECT 299.400 206.400 303.600 207.600 ;
        RECT 298.950 202.950 301.050 205.050 ;
        RECT 271.950 196.950 274.050 199.050 ;
        RECT 295.950 196.950 298.050 199.050 ;
        RECT 265.950 193.950 268.050 196.050 ;
        RECT 277.950 187.950 280.050 190.050 ;
        RECT 253.950 183.000 256.050 187.050 ;
        RECT 278.400 184.200 279.600 187.950 ;
        RECT 296.400 186.600 297.600 196.950 ;
        RECT 293.400 185.400 297.600 186.600 ;
        RECT 254.400 181.050 255.600 183.000 ;
        RECT 259.950 182.100 262.050 184.200 ;
        RECT 260.400 181.050 261.600 182.100 ;
        RECT 268.950 181.950 271.050 184.050 ;
        RECT 277.950 182.100 280.050 184.200 ;
        RECT 253.950 178.950 256.050 181.050 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 259.950 178.950 262.050 181.050 ;
        RECT 262.950 178.950 265.050 181.050 ;
        RECT 253.950 151.950 256.050 154.050 ;
        RECT 247.950 139.950 250.050 142.050 ;
        RECT 230.400 136.050 231.600 137.100 ;
        RECT 235.950 136.800 238.050 138.900 ;
        RECT 241.950 136.950 244.050 139.050 ;
        RECT 244.950 137.100 247.050 139.200 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 208.950 124.950 211.050 127.050 ;
        RECT 202.950 104.100 205.050 106.200 ;
        RECT 208.950 104.100 211.050 106.200 ;
        RECT 221.400 106.050 222.600 133.950 ;
        RECT 227.400 132.900 228.600 133.950 ;
        RECT 236.400 132.900 237.600 136.800 ;
        RECT 245.400 136.050 246.600 137.100 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 248.400 132.900 249.600 133.950 ;
        RECT 254.400 132.900 255.600 151.950 ;
        RECT 257.400 151.050 258.600 178.950 ;
        RECT 256.950 148.950 259.050 151.050 ;
        RECT 257.400 139.200 258.600 148.950 ;
        RECT 263.400 145.050 264.600 178.950 ;
        RECT 269.400 177.900 270.600 181.950 ;
        RECT 278.400 181.050 279.600 182.100 ;
        RECT 286.950 181.950 289.050 184.050 ;
        RECT 274.950 178.950 277.050 181.050 ;
        RECT 277.950 178.950 280.050 181.050 ;
        RECT 275.400 177.900 276.600 178.950 ;
        RECT 268.950 175.800 271.050 177.900 ;
        RECT 274.950 175.800 277.050 177.900 ;
        RECT 262.950 142.950 265.050 145.050 ;
        RECT 256.950 137.100 259.050 139.200 ;
        RECT 262.950 137.100 265.050 139.200 ;
        RECT 263.400 136.050 264.600 137.100 ;
        RECT 269.400 136.050 270.600 175.800 ;
        RECT 259.950 133.950 262.050 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 260.400 132.900 261.600 133.950 ;
        RECT 226.950 130.800 229.050 132.900 ;
        RECT 235.950 130.800 238.050 132.900 ;
        RECT 247.950 130.800 250.050 132.900 ;
        RECT 253.950 130.800 256.050 132.900 ;
        RECT 259.950 127.950 262.050 132.900 ;
        RECT 259.950 121.950 262.050 124.050 ;
        RECT 226.950 118.950 229.050 121.050 ;
        RECT 203.400 103.050 204.600 104.100 ;
        RECT 209.400 103.050 210.600 104.100 ;
        RECT 220.950 103.950 223.050 106.050 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 200.400 100.050 201.600 100.950 ;
        RECT 181.950 94.950 184.050 99.000 ;
        RECT 187.950 97.800 190.050 99.900 ;
        RECT 193.950 97.800 196.050 99.900 ;
        RECT 196.950 98.400 201.600 100.050 ;
        RECT 206.400 99.900 207.600 100.950 ;
        RECT 196.950 97.950 201.000 98.400 ;
        RECT 205.950 97.800 208.050 99.900 ;
        RECT 211.950 97.950 214.050 100.050 ;
        RECT 172.950 91.950 175.050 94.050 ;
        RECT 181.950 79.950 184.050 82.050 ;
        RECT 148.950 76.950 151.050 79.050 ;
        RECT 163.950 76.950 166.050 79.050 ;
        RECT 169.950 76.950 172.050 79.050 ;
        RECT 142.950 73.950 145.050 76.050 ;
        RECT 133.950 67.950 136.050 70.050 ;
        RECT 139.950 67.950 142.050 70.050 ;
        RECT 128.400 62.400 132.600 63.600 ;
        RECT 128.400 58.050 129.600 62.400 ;
        RECT 134.400 58.050 135.600 67.950 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 118.950 52.950 121.050 55.050 ;
        RECT 125.400 54.900 126.600 55.950 ;
        RECT 124.950 52.800 127.050 54.900 ;
        RECT 131.400 54.000 132.600 55.950 ;
        RECT 140.400 54.600 141.600 67.950 ;
        RECT 143.400 55.050 144.600 73.950 ;
        RECT 149.400 58.050 150.600 76.950 ;
        RECT 154.950 73.950 157.050 76.050 ;
        RECT 155.400 58.050 156.600 73.950 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 154.950 55.950 157.050 58.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 130.950 49.950 133.050 54.000 ;
        RECT 137.400 53.400 141.600 54.600 ;
        RECT 121.950 46.950 124.050 49.050 ;
        RECT 112.950 31.950 115.050 34.050 ;
        RECT 122.400 31.050 123.600 46.950 ;
        RECT 137.400 43.050 138.600 53.400 ;
        RECT 142.950 52.950 145.050 55.050 ;
        RECT 152.400 54.900 153.600 55.950 ;
        RECT 151.950 52.800 154.050 54.900 ;
        RECT 139.950 46.950 142.050 52.050 ;
        RECT 136.950 40.950 139.050 43.050 ;
        RECT 124.950 37.950 127.050 40.050 ;
        RECT 133.950 37.950 136.050 40.050 ;
        RECT 110.400 29.400 114.600 30.600 ;
        RECT 104.400 26.400 111.600 27.600 ;
        RECT 104.400 25.050 105.600 26.400 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 97.950 22.950 100.050 25.050 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 103.950 22.950 106.050 25.050 ;
        RECT 95.400 21.900 96.600 22.950 ;
        RECT 88.950 19.800 91.050 21.900 ;
        RECT 94.950 19.800 97.050 21.900 ;
        RECT 101.400 21.000 102.600 22.950 ;
        RECT 85.950 16.950 88.050 19.050 ;
        RECT 100.950 16.950 103.050 21.000 ;
        RECT 110.400 13.050 111.600 26.400 ;
        RECT 109.950 10.950 112.050 13.050 ;
        RECT 46.950 7.950 49.050 10.050 ;
        RECT 113.400 7.050 114.600 29.400 ;
        RECT 121.950 28.950 124.050 31.050 ;
        RECT 118.950 26.100 121.050 28.200 ;
        RECT 119.400 25.050 120.600 26.100 ;
        RECT 125.400 25.050 126.600 37.950 ;
        RECT 130.950 31.950 133.050 34.050 ;
        RECT 131.400 28.050 132.600 31.950 ;
        RECT 130.950 25.950 133.050 28.050 ;
        RECT 118.950 22.950 121.050 25.050 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 122.400 21.900 123.600 22.950 ;
        RECT 128.400 21.900 129.600 22.950 ;
        RECT 121.950 19.800 124.050 21.900 ;
        RECT 127.950 19.800 130.050 21.900 ;
        RECT 134.400 16.050 135.600 37.950 ;
        RECT 137.400 25.050 138.600 40.950 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 140.400 22.050 141.600 46.950 ;
        RECT 158.400 40.050 159.600 55.950 ;
        RECT 148.950 37.950 151.050 40.050 ;
        RECT 157.950 37.950 160.050 40.050 ;
        RECT 149.400 28.200 150.600 37.950 ;
        RECT 164.400 37.050 165.600 76.950 ;
        RECT 175.950 73.950 178.050 76.050 ;
        RECT 176.400 70.050 177.600 73.950 ;
        RECT 175.950 67.950 178.050 70.050 ;
        RECT 166.950 60.600 171.000 61.050 ;
        RECT 166.950 58.950 171.600 60.600 ;
        RECT 170.400 58.050 171.600 58.950 ;
        RECT 176.400 58.050 177.600 67.950 ;
        RECT 182.400 61.050 183.600 79.950 ;
        RECT 205.950 73.950 208.050 76.050 ;
        RECT 190.950 67.950 193.050 70.050 ;
        RECT 181.950 58.950 184.050 61.050 ;
        RECT 191.400 58.050 192.600 67.950 ;
        RECT 196.950 59.100 199.050 61.200 ;
        RECT 197.400 58.050 198.600 59.100 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 166.950 52.950 169.050 55.050 ;
        RECT 173.400 54.900 174.600 55.950 ;
        RECT 179.400 54.900 180.600 55.950 ;
        RECT 188.400 54.900 189.600 55.950 ;
        RECT 167.400 49.050 168.600 52.950 ;
        RECT 172.950 52.800 175.050 54.900 ;
        RECT 178.950 52.800 181.050 54.900 ;
        RECT 187.950 52.800 190.050 54.900 ;
        RECT 166.950 46.950 169.050 49.050 ;
        RECT 190.950 46.950 193.050 49.050 ;
        RECT 184.950 40.950 187.050 43.050 ;
        RECT 163.950 34.950 166.050 37.050 ;
        RECT 175.950 34.950 178.050 37.050 ;
        RECT 164.400 30.600 165.600 34.950 ;
        RECT 161.400 29.400 165.600 30.600 ;
        RECT 148.950 26.100 151.050 28.200 ;
        RECT 149.400 25.050 150.600 26.100 ;
        RECT 161.400 25.050 162.600 29.400 ;
        RECT 166.950 26.100 169.050 28.200 ;
        RECT 167.400 25.050 168.600 26.100 ;
        RECT 172.950 25.950 175.050 28.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 163.950 22.950 166.050 25.050 ;
        RECT 166.950 22.950 169.050 25.050 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 146.400 21.900 147.600 22.950 ;
        RECT 158.400 21.900 159.600 22.950 ;
        RECT 145.950 19.800 148.050 21.900 ;
        RECT 157.950 19.800 160.050 21.900 ;
        RECT 164.400 21.000 165.600 22.950 ;
        RECT 146.400 19.050 147.600 19.800 ;
        RECT 146.400 17.400 151.050 19.050 ;
        RECT 147.000 16.950 151.050 17.400 ;
        RECT 163.950 16.950 166.050 21.000 ;
        RECT 173.400 19.050 174.600 25.950 ;
        RECT 176.400 19.050 177.600 34.950 ;
        RECT 185.400 25.050 186.600 40.950 ;
        RECT 191.400 25.050 192.600 46.950 ;
        RECT 194.400 37.050 195.600 55.950 ;
        RECT 206.400 49.050 207.600 73.950 ;
        RECT 212.400 70.050 213.600 97.950 ;
        RECT 221.400 94.050 222.600 103.950 ;
        RECT 227.400 103.050 228.600 118.950 ;
        RECT 247.950 115.950 250.050 118.050 ;
        RECT 248.400 106.200 249.600 115.950 ;
        RECT 232.950 104.100 235.050 106.200 ;
        RECT 247.950 104.100 250.050 106.200 ;
        RECT 255.000 105.600 259.050 106.050 ;
        RECT 233.400 103.050 234.600 104.100 ;
        RECT 248.400 103.050 249.600 104.100 ;
        RECT 254.400 103.950 259.050 105.600 ;
        RECT 254.400 103.050 255.600 103.950 ;
        RECT 226.950 100.950 229.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 247.950 100.950 250.050 103.050 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 230.400 99.000 231.600 100.950 ;
        RECT 236.400 99.900 237.600 100.950 ;
        RECT 223.950 94.950 226.050 97.050 ;
        RECT 229.950 94.950 232.050 99.000 ;
        RECT 235.950 97.800 238.050 99.900 ;
        RECT 220.950 91.950 223.050 94.050 ;
        RECT 224.400 91.050 225.600 94.950 ;
        RECT 245.400 94.050 246.600 100.950 ;
        RECT 251.400 99.900 252.600 100.950 ;
        RECT 260.400 100.050 261.600 121.950 ;
        RECT 266.400 118.050 267.600 133.950 ;
        RECT 275.400 132.900 276.600 175.800 ;
        RECT 277.950 163.950 280.050 166.050 ;
        RECT 274.950 130.800 277.050 132.900 ;
        RECT 265.950 115.950 268.050 118.050 ;
        RECT 271.950 115.950 274.050 118.050 ;
        RECT 272.400 112.050 273.600 115.950 ;
        RECT 271.950 109.950 274.050 112.050 ;
        RECT 278.400 109.050 279.600 163.950 ;
        RECT 287.400 163.050 288.600 181.950 ;
        RECT 293.400 181.050 294.600 185.400 ;
        RECT 299.400 181.050 300.600 202.950 ;
        RECT 302.400 184.050 303.600 206.400 ;
        RECT 301.950 181.950 304.050 184.050 ;
        RECT 307.950 183.000 310.050 187.050 ;
        RECT 308.400 181.050 309.600 183.000 ;
        RECT 314.400 181.050 315.600 208.800 ;
        RECT 317.400 205.050 318.600 211.950 ;
        RECT 323.400 205.050 324.600 211.950 ;
        RECT 332.400 211.050 333.600 223.950 ;
        RECT 340.950 215.100 343.050 217.200 ;
        RECT 341.400 214.050 342.600 215.100 ;
        RECT 337.950 211.950 340.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 328.950 208.950 331.050 211.050 ;
        RECT 331.950 208.950 334.050 211.050 ;
        RECT 338.400 210.900 339.600 211.950 ;
        RECT 316.950 202.950 319.050 205.050 ;
        RECT 322.950 202.950 325.050 205.050 ;
        RECT 317.400 199.050 318.600 202.950 ;
        RECT 316.950 196.950 319.050 199.050 ;
        RECT 322.950 195.600 325.050 196.050 ;
        RECT 317.400 194.400 325.050 195.600 ;
        RECT 317.400 187.050 318.600 194.400 ;
        RECT 322.950 193.950 325.050 194.400 ;
        RECT 322.950 187.950 325.050 190.050 ;
        RECT 316.950 184.950 319.050 187.050 ;
        RECT 292.950 178.950 295.050 181.050 ;
        RECT 295.950 178.950 298.050 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 313.950 178.950 316.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 286.950 160.950 289.050 163.050 ;
        RECT 287.400 157.050 288.600 160.950 ;
        RECT 286.950 154.950 289.050 157.050 ;
        RECT 283.950 145.950 286.050 148.050 ;
        RECT 284.400 136.050 285.600 145.950 ;
        RECT 289.950 138.000 292.050 142.050 ;
        RECT 296.400 139.050 297.600 178.950 ;
        RECT 304.950 175.950 307.050 178.050 ;
        RECT 311.400 177.000 312.600 178.950 ;
        RECT 317.400 177.900 318.600 178.950 ;
        RECT 323.400 177.900 324.600 187.950 ;
        RECT 329.400 186.600 330.600 208.950 ;
        RECT 337.950 208.800 340.050 210.900 ;
        RECT 331.950 205.800 334.050 207.900 ;
        RECT 332.400 187.050 333.600 205.800 ;
        RECT 347.400 205.050 348.600 238.950 ;
        RECT 349.950 234.600 352.050 235.050 ;
        RECT 353.400 234.600 354.600 322.950 ;
        RECT 356.400 316.050 357.600 329.400 ;
        RECT 355.950 313.950 358.050 316.050 ;
        RECT 359.400 301.050 360.600 340.950 ;
        RECT 362.400 325.050 363.600 343.950 ;
        RECT 365.400 337.050 366.600 343.950 ;
        RECT 368.400 343.050 369.600 400.950 ;
        RECT 371.400 373.050 372.600 404.400 ;
        RECT 374.400 403.050 375.600 433.950 ;
        RECT 379.950 430.950 382.050 433.050 ;
        RECT 376.950 421.950 379.050 424.050 ;
        RECT 377.400 418.050 378.600 421.950 ;
        RECT 380.400 421.050 381.600 430.950 ;
        RECT 383.400 424.050 384.600 449.400 ;
        RECT 385.950 448.950 388.050 451.050 ;
        RECT 389.400 448.050 390.600 472.950 ;
        RECT 395.400 469.050 396.600 487.950 ;
        RECT 394.950 466.950 397.050 469.050 ;
        RECT 394.950 457.950 397.050 460.050 ;
        RECT 395.400 448.050 396.600 457.950 ;
        RECT 398.400 454.050 399.600 521.400 ;
        RECT 400.950 499.950 403.050 502.050 ;
        RECT 401.400 495.600 402.600 499.950 ;
        RECT 404.400 499.050 405.600 565.950 ;
        RECT 410.400 547.050 411.600 568.950 ;
        RECT 419.400 568.050 420.600 574.800 ;
        RECT 422.400 574.050 423.600 599.400 ;
        RECT 424.950 598.800 427.050 599.400 ;
        RECT 430.950 598.950 433.050 601.050 ;
        RECT 431.400 595.050 432.600 598.950 ;
        RECT 430.950 592.950 433.050 595.050 ;
        RECT 434.400 577.050 435.600 605.400 ;
        RECT 437.400 601.050 438.600 653.400 ;
        RECT 440.400 652.050 441.600 664.950 ;
        RECT 457.950 661.950 460.050 664.050 ;
        RECT 448.950 656.400 451.050 658.500 ;
        RECT 439.950 649.950 442.050 652.050 ;
        RECT 442.950 646.950 445.050 649.050 ;
        RECT 443.400 646.050 444.600 646.950 ;
        RECT 443.400 644.400 448.050 646.050 ;
        RECT 444.000 643.950 448.050 644.400 ;
        RECT 449.100 636.600 450.300 656.400 ;
        RECT 458.400 651.600 459.600 661.950 ;
        RECT 463.950 656.400 466.050 658.500 ;
        RECT 458.400 650.400 462.600 651.600 ;
        RECT 461.400 649.050 462.600 650.400 ;
        RECT 451.950 646.950 454.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 452.400 640.050 453.600 646.950 ;
        RECT 464.850 641.400 466.050 656.400 ;
        RECT 451.950 637.950 454.050 640.050 ;
        RECT 463.950 639.300 466.050 641.400 ;
        RECT 448.950 634.500 451.050 636.600 ;
        RECT 464.850 635.700 466.050 639.300 ;
        RECT 463.950 633.600 466.050 635.700 ;
        RECT 442.950 628.950 445.050 631.050 ;
        RECT 470.400 630.600 471.600 673.950 ;
        RECT 467.400 629.400 471.600 630.600 ;
        RECT 443.400 607.050 444.600 628.950 ;
        RECT 451.950 622.950 454.050 625.050 ;
        RECT 439.950 604.950 442.050 607.050 ;
        RECT 442.950 604.950 445.050 607.050 ;
        RECT 436.950 598.950 439.050 601.050 ;
        RECT 440.400 594.600 441.600 604.950 ;
        RECT 452.400 604.050 453.600 622.950 ;
        RECT 460.950 615.300 463.050 617.400 ;
        RECT 461.850 611.700 463.050 615.300 ;
        RECT 460.950 609.600 463.050 611.700 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 457.950 601.950 460.050 604.050 ;
        RECT 442.950 598.950 445.050 601.050 ;
        RECT 446.400 600.900 447.600 601.950 ;
        RECT 437.400 593.400 441.600 594.600 ;
        RECT 437.400 583.050 438.600 593.400 ;
        RECT 439.950 583.950 442.050 586.050 ;
        RECT 436.950 580.950 439.050 583.050 ;
        RECT 433.950 574.950 436.050 577.050 ;
        RECT 421.950 571.950 424.050 574.050 ;
        RECT 427.950 572.100 430.050 574.200 ;
        RECT 437.400 573.600 438.600 580.950 ;
        RECT 434.400 572.400 438.600 573.600 ;
        RECT 428.400 571.050 429.600 572.100 ;
        RECT 434.400 571.050 435.600 572.400 ;
        RECT 424.950 568.950 427.050 571.050 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 433.950 568.950 436.050 571.050 ;
        RECT 418.950 565.950 421.050 568.050 ;
        RECT 425.400 567.900 426.600 568.950 ;
        RECT 424.950 565.800 427.050 567.900 ;
        RECT 418.950 562.800 421.050 564.900 ;
        RECT 427.950 562.950 430.050 565.050 ;
        RECT 419.400 556.050 420.600 562.800 ;
        RECT 418.950 553.950 421.050 556.050 ;
        RECT 409.950 544.950 412.050 547.050 ;
        RECT 406.950 541.950 409.050 544.050 ;
        RECT 407.400 505.050 408.600 541.950 ;
        RECT 419.400 532.050 420.600 553.950 ;
        RECT 428.400 538.050 429.600 562.950 ;
        RECT 431.400 544.050 432.600 568.950 ;
        RECT 440.400 567.900 441.600 583.950 ;
        RECT 443.400 574.050 444.600 598.950 ;
        RECT 445.950 598.800 448.050 600.900 ;
        RECT 458.400 600.600 459.600 601.950 ;
        RECT 455.400 599.400 459.600 600.600 ;
        RECT 455.400 580.050 456.600 599.400 ;
        RECT 461.850 594.600 463.050 609.600 ;
        RECT 460.950 592.500 463.050 594.600 ;
        RECT 467.400 586.050 468.600 629.400 ;
        RECT 473.400 606.600 474.600 682.950 ;
        RECT 476.400 676.050 477.600 716.400 ;
        RECT 481.950 715.950 484.050 718.050 ;
        RECT 485.400 685.050 486.600 727.950 ;
        RECT 488.400 697.050 489.600 751.950 ;
        RECT 493.950 745.950 496.050 748.050 ;
        RECT 494.400 742.050 495.600 745.950 ;
        RECT 493.950 739.950 496.050 742.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 494.400 723.900 495.600 724.950 ;
        RECT 493.950 721.800 496.050 723.900 ;
        RECT 496.950 718.950 499.050 721.050 ;
        RECT 493.950 712.950 496.050 715.050 ;
        RECT 490.950 703.950 493.050 706.050 ;
        RECT 491.400 700.050 492.600 703.950 ;
        RECT 490.950 697.950 493.050 700.050 ;
        RECT 487.950 694.950 490.050 697.050 ;
        RECT 484.950 682.950 487.050 685.050 ;
        RECT 488.400 682.050 489.600 694.950 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 475.950 673.950 478.050 676.050 ;
        RECT 482.400 664.050 483.600 679.950 ;
        RECT 494.400 664.050 495.600 712.950 ;
        RECT 497.400 685.050 498.600 718.950 ;
        RECT 503.400 715.050 504.600 754.800 ;
        RECT 506.400 730.050 507.600 796.800 ;
        RECT 509.400 781.050 510.600 799.950 ;
        RECT 511.950 799.800 514.050 801.900 ;
        RECT 514.950 796.950 517.050 799.050 ;
        RECT 508.950 778.950 511.050 781.050 ;
        RECT 515.400 775.050 516.600 796.950 ;
        RECT 518.400 790.050 519.600 802.950 ;
        RECT 524.400 801.900 525.600 802.950 ;
        RECT 536.400 801.900 537.600 802.950 ;
        RECT 542.400 801.900 543.600 802.950 ;
        RECT 523.950 799.800 526.050 801.900 ;
        RECT 535.950 799.800 538.050 801.900 ;
        RECT 541.950 799.800 544.050 801.900 ;
        RECT 544.950 799.950 547.050 802.050 ;
        RECT 517.950 787.950 520.050 790.050 ;
        RECT 524.400 787.050 525.600 799.800 ;
        RECT 542.400 796.050 543.600 799.800 ;
        RECT 541.950 793.950 544.050 796.050 ;
        RECT 523.950 784.950 526.050 787.050 ;
        RECT 526.950 778.950 529.050 781.050 ;
        RECT 514.950 772.950 517.050 775.050 ;
        RECT 508.950 760.950 511.050 763.050 ;
        RECT 509.400 745.050 510.600 760.950 ;
        RECT 515.400 760.050 516.600 772.950 ;
        RECT 520.950 761.100 523.050 763.200 ;
        RECT 527.400 763.050 528.600 778.950 ;
        RECT 545.400 778.050 546.600 799.950 ;
        RECT 529.950 775.950 532.050 778.050 ;
        RECT 544.950 775.950 547.050 778.050 ;
        RECT 521.400 760.050 522.600 761.100 ;
        RECT 526.950 760.950 529.050 763.050 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 517.950 757.950 520.050 760.050 ;
        RECT 520.950 757.950 523.050 760.050 ;
        RECT 523.950 757.950 526.050 760.050 ;
        RECT 508.950 742.950 511.050 745.050 ;
        RECT 518.400 739.050 519.600 757.950 ;
        RECT 524.400 756.900 525.600 757.950 ;
        RECT 530.400 757.050 531.600 775.950 ;
        RECT 532.950 769.950 535.050 772.050 ;
        RECT 538.950 769.950 541.050 772.050 ;
        RECT 533.400 766.050 534.600 769.950 ;
        RECT 532.950 763.950 535.050 766.050 ;
        RECT 539.400 763.200 540.600 769.950 ;
        RECT 532.950 760.800 535.050 762.900 ;
        RECT 538.950 761.100 541.050 763.200 ;
        RECT 523.950 754.800 526.050 756.900 ;
        RECT 529.950 754.950 532.050 757.050 ;
        RECT 523.950 748.950 526.050 751.050 ;
        RECT 520.950 745.950 523.050 748.050 ;
        RECT 521.400 742.050 522.600 745.950 ;
        RECT 520.950 739.950 523.050 742.050 ;
        RECT 508.950 736.950 511.050 739.050 ;
        RECT 517.950 736.950 520.050 739.050 ;
        RECT 505.950 727.950 508.050 730.050 ;
        RECT 509.400 727.050 510.600 736.950 ;
        RECT 514.950 733.950 517.050 736.050 ;
        RECT 515.400 727.050 516.600 733.950 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 512.400 718.050 513.600 724.950 ;
        RECT 518.400 718.050 519.600 724.950 ;
        RECT 524.400 723.600 525.600 748.950 ;
        RECT 533.400 748.050 534.600 760.800 ;
        RECT 539.400 760.050 540.600 761.100 ;
        RECT 545.400 760.050 546.600 775.950 ;
        RECT 548.400 763.050 549.600 826.950 ;
        RECT 560.400 820.050 561.600 875.400 ;
        RECT 592.950 874.950 595.050 877.050 ;
        RECT 601.950 874.950 604.050 877.050 ;
        RECT 568.950 868.950 571.050 871.050 ;
        RECT 569.400 865.050 570.600 868.950 ;
        RECT 568.950 862.950 571.050 865.050 ;
        RECT 583.950 859.950 586.050 862.050 ;
        RECT 577.950 856.950 580.050 859.050 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 566.400 823.050 567.600 835.950 ;
        RECT 578.400 835.050 579.600 856.950 ;
        RECT 584.400 838.050 585.600 859.950 ;
        RECT 593.400 856.050 594.600 874.950 ;
        RECT 611.400 874.050 612.600 877.800 ;
        RECT 610.950 871.950 613.050 874.050 ;
        RECT 617.400 871.050 618.600 880.950 ;
        RECT 625.800 879.000 627.900 880.050 ;
        RECT 629.400 879.900 630.600 880.950 ;
        RECT 625.800 877.950 628.050 879.000 ;
        RECT 625.950 874.950 628.050 877.950 ;
        RECT 628.950 877.800 631.050 879.900 ;
        RECT 635.400 879.000 636.600 880.950 ;
        RECT 634.950 874.950 637.050 879.000 ;
        RECT 640.950 877.950 643.050 880.050 ;
        RECT 650.400 879.900 651.600 898.800 ;
        RECT 653.400 889.050 654.600 898.950 ;
        RECT 656.400 889.050 657.600 913.950 ;
        RECT 658.950 904.950 661.050 907.050 ;
        RECT 652.950 886.950 655.050 889.050 ;
        RECT 655.950 886.950 658.050 889.050 ;
        RECT 659.400 883.050 660.600 904.950 ;
        RECT 665.400 901.050 666.600 934.950 ;
        RECT 739.950 931.950 742.050 934.050 ;
        RECT 694.500 922.500 696.600 924.600 ;
        RECT 673.950 917.100 676.050 919.200 ;
        RECT 674.400 916.050 675.600 917.100 ;
        RECT 682.950 916.950 685.050 919.050 ;
        RECT 673.950 913.950 676.050 916.050 ;
        RECT 676.950 913.950 679.050 916.050 ;
        RECT 677.400 912.900 678.600 913.950 ;
        RECT 683.400 912.900 684.600 916.950 ;
        RECT 685.950 913.950 688.050 916.050 ;
        RECT 691.950 913.950 694.050 916.050 ;
        RECT 694.950 915.300 696.000 922.500 ;
        RECT 698.400 918.900 699.600 921.450 ;
        RECT 704.100 921.300 706.200 923.400 ;
        RECT 718.950 922.950 721.050 925.050 ;
        RECT 697.800 916.800 699.900 918.900 ;
        RECT 700.800 917.700 702.900 919.800 ;
        RECT 700.800 915.300 701.700 917.700 ;
        RECT 694.950 914.100 701.700 915.300 ;
        RECT 667.950 910.800 670.050 912.900 ;
        RECT 676.950 910.800 679.050 912.900 ;
        RECT 682.950 910.800 685.050 912.900 ;
        RECT 664.950 898.950 667.050 901.050 ;
        RECT 668.400 895.050 669.600 910.800 ;
        RECT 677.400 907.050 678.600 910.800 ;
        RECT 673.800 904.950 675.900 907.050 ;
        RECT 676.950 904.950 679.050 907.050 ;
        RECT 670.950 895.950 673.050 898.050 ;
        RECT 667.950 892.950 670.050 895.050 ;
        RECT 664.950 885.000 667.050 889.050 ;
        RECT 665.400 883.050 666.600 885.000 ;
        RECT 655.950 880.950 658.050 883.050 ;
        RECT 658.950 880.950 661.050 883.050 ;
        RECT 661.950 880.950 664.050 883.050 ;
        RECT 664.950 880.950 667.050 883.050 ;
        RECT 656.400 879.900 657.600 880.950 ;
        RECT 641.400 871.050 642.600 877.950 ;
        RECT 649.950 877.800 652.050 879.900 ;
        RECT 655.950 877.800 658.050 879.900 ;
        RECT 662.400 874.050 663.600 880.950 ;
        RECT 671.400 879.900 672.600 895.950 ;
        RECT 674.400 892.050 675.600 904.950 ;
        RECT 673.950 889.950 676.050 892.050 ;
        RECT 679.950 889.950 682.050 892.050 ;
        RECT 680.400 883.050 681.600 889.950 ;
        RECT 683.400 888.600 684.600 910.800 ;
        RECT 686.400 907.050 687.600 913.950 ;
        RECT 692.400 911.400 693.600 913.950 ;
        RECT 694.950 908.700 695.850 914.100 ;
        RECT 696.750 912.300 698.850 913.200 ;
        RECT 704.400 912.300 705.300 921.300 ;
        RECT 707.400 916.050 708.600 918.600 ;
        RECT 719.400 916.050 720.600 922.950 ;
        RECT 724.950 917.100 727.050 919.200 ;
        RECT 733.950 917.100 736.050 919.200 ;
        RECT 725.400 916.050 726.600 917.100 ;
        RECT 706.500 913.950 708.600 916.050 ;
        RECT 718.950 913.950 721.050 916.050 ;
        RECT 721.950 913.950 724.050 916.050 ;
        RECT 724.950 913.950 727.050 916.050 ;
        RECT 727.950 913.950 730.050 916.050 ;
        RECT 696.750 911.100 705.300 912.300 ;
        RECT 685.950 904.950 688.050 907.050 ;
        RECT 694.500 906.600 696.600 908.700 ;
        RECT 697.800 908.100 699.900 910.200 ;
        RECT 701.700 909.300 703.800 911.100 ;
        RECT 709.950 910.950 712.050 913.050 ;
        RECT 722.400 912.900 723.600 913.950 ;
        RECT 694.950 895.950 697.050 898.050 ;
        RECT 691.950 889.950 694.050 892.050 ;
        RECT 683.400 887.400 687.600 888.600 ;
        RECT 686.400 883.050 687.600 887.400 ;
        RECT 692.400 886.050 693.600 889.950 ;
        RECT 691.950 883.950 694.050 886.050 ;
        RECT 676.950 880.950 679.050 883.050 ;
        RECT 679.950 880.950 682.050 883.050 ;
        RECT 682.950 880.950 685.050 883.050 ;
        RECT 685.950 880.950 688.050 883.050 ;
        RECT 688.950 880.950 691.050 883.050 ;
        RECT 677.400 879.900 678.600 880.950 ;
        RECT 670.950 877.800 673.050 879.900 ;
        RECT 676.950 877.800 679.050 879.900 ;
        RECT 661.950 873.600 664.050 874.050 ;
        RECT 659.400 872.400 664.050 873.600 ;
        RECT 616.950 868.950 619.050 871.050 ;
        RECT 640.950 868.950 643.050 871.050 ;
        RECT 634.950 856.950 637.050 859.050 ;
        RECT 592.950 853.950 595.050 856.050 ;
        RECT 598.950 853.950 601.050 856.050 ;
        RECT 589.950 839.100 592.050 841.200 ;
        RECT 590.400 838.050 591.600 839.100 ;
        RECT 583.950 835.950 586.050 838.050 ;
        RECT 586.950 835.950 589.050 838.050 ;
        RECT 589.950 835.950 592.050 838.050 ;
        RECT 577.800 832.950 579.900 835.050 ;
        RECT 577.950 826.950 580.050 829.050 ;
        RECT 565.950 820.950 568.050 823.050 ;
        RECT 559.950 817.950 562.050 820.050 ;
        RECT 556.950 806.100 559.050 808.200 ;
        RECT 562.950 806.100 565.050 808.200 ;
        RECT 557.400 805.050 558.600 806.100 ;
        RECT 563.400 805.050 564.600 806.100 ;
        RECT 571.800 805.950 573.900 808.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 565.950 802.950 568.050 805.050 ;
        RECT 560.400 790.050 561.600 802.950 ;
        RECT 559.950 787.950 562.050 790.050 ;
        RECT 556.950 784.950 559.050 787.050 ;
        RECT 557.400 775.050 558.600 784.950 ;
        RECT 566.400 784.050 567.600 802.950 ;
        RECT 572.400 796.050 573.600 805.950 ;
        RECT 578.400 805.050 579.600 826.950 ;
        RECT 587.400 823.050 588.600 835.950 ;
        RECT 592.950 832.950 595.050 835.050 ;
        RECT 593.400 825.600 594.600 832.950 ;
        RECT 599.400 829.050 600.600 853.950 ;
        RECT 613.950 839.100 616.050 841.200 ;
        RECT 619.950 839.100 622.050 841.200 ;
        RECT 628.950 839.100 631.050 841.200 ;
        RECT 614.400 838.050 615.600 839.100 ;
        RECT 604.950 835.950 607.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 605.400 829.050 606.600 835.950 ;
        RECT 611.400 829.050 612.600 835.950 ;
        RECT 598.950 826.950 601.050 829.050 ;
        RECT 604.950 826.950 607.050 829.050 ;
        RECT 610.950 826.950 613.050 829.050 ;
        RECT 593.400 824.400 597.600 825.600 ;
        RECT 586.950 820.950 589.050 823.050 ;
        RECT 583.950 817.950 586.050 820.050 ;
        RECT 584.400 805.050 585.600 817.950 ;
        RECT 596.400 817.050 597.600 824.400 ;
        RECT 620.400 822.600 621.600 839.100 ;
        RECT 629.400 838.050 630.600 839.100 ;
        RECT 635.400 838.050 636.600 856.950 ;
        RECT 640.950 839.100 643.050 841.200 ;
        RECT 646.950 839.100 649.050 841.200 ;
        RECT 652.950 839.100 655.050 841.200 ;
        RECT 625.950 835.950 628.050 838.050 ;
        RECT 628.950 835.950 631.050 838.050 ;
        RECT 631.950 835.950 634.050 838.050 ;
        RECT 634.950 835.950 637.050 838.050 ;
        RECT 626.400 834.000 627.600 835.950 ;
        RECT 625.950 829.950 628.050 834.000 ;
        RECT 632.400 823.050 633.600 835.950 ;
        RECT 637.950 829.950 640.050 832.050 ;
        RECT 622.950 822.600 625.050 823.050 ;
        RECT 620.400 821.400 625.050 822.600 ;
        RECT 622.950 820.950 625.050 821.400 ;
        RECT 631.950 820.950 634.050 823.050 ;
        RECT 589.950 814.950 592.050 817.050 ;
        RECT 595.950 814.950 598.050 817.050 ;
        RECT 610.950 814.950 613.050 817.050 ;
        RECT 590.400 808.050 591.600 814.950 ;
        RECT 589.950 807.600 592.050 808.050 ;
        RECT 589.950 806.400 594.600 807.600 ;
        RECT 589.950 805.950 592.050 806.400 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 586.950 802.950 589.050 805.050 ;
        RECT 581.400 798.600 582.600 802.950 ;
        RECT 587.400 801.900 588.600 802.950 ;
        RECT 586.800 799.800 588.900 801.900 ;
        RECT 589.950 799.800 592.050 801.900 ;
        RECT 578.400 797.400 582.600 798.600 ;
        RECT 571.950 793.950 574.050 796.050 ;
        RECT 565.950 781.950 568.050 784.050 ;
        RECT 556.950 772.950 559.050 775.050 ;
        RECT 571.950 774.600 574.050 775.050 ;
        RECT 571.950 773.400 576.600 774.600 ;
        RECT 571.950 772.950 574.050 773.400 ;
        RECT 553.950 766.950 556.050 769.050 ;
        RECT 565.950 766.950 568.050 769.050 ;
        RECT 547.950 760.950 550.050 763.050 ;
        RECT 538.950 757.950 541.050 760.050 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 544.950 757.950 547.050 760.050 ;
        RECT 542.400 756.900 543.600 757.950 ;
        RECT 541.950 754.800 544.050 756.900 ;
        RECT 547.950 754.950 550.050 757.050 ;
        RECT 548.400 748.050 549.600 754.950 ;
        RECT 532.950 745.950 535.050 748.050 ;
        RECT 538.950 745.950 541.050 748.050 ;
        RECT 547.950 745.950 550.050 748.050 ;
        RECT 532.950 728.100 535.050 730.200 ;
        RECT 539.400 730.050 540.600 745.950 ;
        RECT 554.400 733.050 555.600 766.950 ;
        RECT 559.950 761.100 562.050 763.200 ;
        RECT 560.400 760.050 561.600 761.100 ;
        RECT 566.400 760.050 567.600 766.950 ;
        RECT 572.400 760.050 573.600 772.950 ;
        RECT 575.400 769.050 576.600 773.400 ;
        RECT 574.950 766.950 577.050 769.050 ;
        RECT 559.950 757.950 562.050 760.050 ;
        RECT 562.950 757.950 565.050 760.050 ;
        RECT 565.950 757.950 568.050 760.050 ;
        RECT 568.950 757.950 571.050 760.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 556.950 754.950 559.050 757.050 ;
        RECT 557.400 751.050 558.600 754.950 ;
        RECT 563.400 753.600 564.600 757.950 ;
        RECT 563.400 752.400 567.600 753.600 ;
        RECT 556.950 748.950 559.050 751.050 ;
        RECT 562.950 745.950 565.050 748.050 ;
        RECT 553.950 730.950 556.050 733.050 ;
        RECT 533.400 727.050 534.600 728.100 ;
        RECT 538.950 727.950 541.050 730.050 ;
        RECT 541.950 727.950 544.050 730.050 ;
        RECT 547.950 727.950 550.050 730.050 ;
        RECT 556.950 728.100 559.050 730.200 ;
        RECT 563.400 730.050 564.600 745.950 ;
        RECT 566.400 742.050 567.600 752.400 ;
        RECT 569.400 751.050 570.600 757.950 ;
        RECT 578.400 754.050 579.600 797.400 ;
        RECT 587.400 790.050 588.600 799.800 ;
        RECT 586.950 787.950 589.050 790.050 ;
        RECT 590.400 787.050 591.600 799.800 ;
        RECT 580.950 784.950 583.050 787.050 ;
        RECT 589.950 784.950 592.050 787.050 ;
        RECT 581.400 763.050 582.600 784.950 ;
        RECT 593.400 780.600 594.600 806.400 ;
        RECT 601.950 802.950 604.050 805.050 ;
        RECT 602.400 801.900 603.600 802.950 ;
        RECT 601.950 799.800 604.050 801.900 ;
        RECT 611.400 796.050 612.600 814.950 ;
        RECT 613.950 811.950 616.050 814.050 ;
        RECT 598.950 793.950 601.050 796.050 ;
        RECT 610.950 793.950 613.050 796.050 ;
        RECT 595.950 790.950 598.050 793.050 ;
        RECT 596.400 787.050 597.600 790.950 ;
        RECT 595.950 784.950 598.050 787.050 ;
        RECT 590.400 779.400 594.600 780.600 ;
        RECT 583.950 769.950 586.050 772.050 ;
        RECT 580.950 760.950 583.050 763.050 ;
        RECT 584.400 760.050 585.600 769.950 ;
        RECT 590.400 763.050 591.600 779.400 ;
        RECT 592.950 775.950 595.050 778.050 ;
        RECT 593.400 769.050 594.600 775.950 ;
        RECT 592.950 766.950 595.050 769.050 ;
        RECT 589.950 760.950 592.050 763.050 ;
        RECT 596.400 762.600 597.600 784.950 ;
        RECT 593.400 761.400 597.600 762.600 ;
        RECT 593.400 760.050 594.600 761.400 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 586.950 757.950 589.050 760.050 ;
        RECT 592.950 757.950 595.050 760.050 ;
        RECT 587.400 756.000 588.600 757.950 ;
        RECT 577.950 751.950 580.050 754.050 ;
        RECT 583.800 751.950 585.900 754.050 ;
        RECT 586.950 751.950 589.050 756.000 ;
        RECT 595.950 754.950 598.050 757.050 ;
        RECT 568.950 748.950 571.050 751.050 ;
        RECT 571.950 745.950 574.050 748.050 ;
        RECT 572.400 742.050 573.600 745.950 ;
        RECT 565.950 739.950 568.050 742.050 ;
        RECT 571.950 739.950 574.050 742.050 ;
        RECT 568.950 736.950 571.050 739.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 524.400 722.400 528.600 723.600 ;
        RECT 511.950 715.950 514.050 718.050 ;
        RECT 517.950 715.950 520.050 718.050 ;
        RECT 502.950 712.950 505.050 715.050 ;
        RECT 499.950 706.950 502.050 709.050 ;
        RECT 496.950 682.950 499.050 685.050 ;
        RECT 497.400 678.600 498.600 682.950 ;
        RECT 500.400 682.050 501.600 706.950 ;
        RECT 505.800 687.300 507.900 689.400 ;
        RECT 515.400 688.500 517.500 690.600 ;
        RECT 523.950 688.950 526.050 691.050 ;
        RECT 503.400 682.050 504.600 684.600 ;
        RECT 499.950 679.950 502.050 682.050 ;
        RECT 503.400 679.950 505.500 682.050 ;
        RECT 497.400 677.400 501.600 678.600 ;
        RECT 496.950 670.950 499.050 673.050 ;
        RECT 481.950 661.950 484.050 664.050 ;
        RECT 493.950 661.950 496.050 664.050 ;
        RECT 484.950 656.400 487.050 658.500 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 479.400 637.050 480.600 646.950 ;
        RECT 478.950 634.950 481.050 637.050 ;
        RECT 485.100 636.600 486.300 656.400 ;
        RECT 493.950 655.950 496.050 658.050 ;
        RECT 487.950 646.950 490.050 649.050 ;
        RECT 488.400 645.600 489.600 646.950 ;
        RECT 488.400 644.400 492.600 645.600 ;
        RECT 491.400 640.050 492.600 644.400 ;
        RECT 490.950 637.950 493.050 640.050 ;
        RECT 484.950 634.500 487.050 636.600 ;
        RECT 487.950 628.950 490.050 631.050 ;
        RECT 488.400 619.050 489.600 628.950 ;
        RECT 487.950 616.950 490.050 619.050 ;
        RECT 481.950 614.400 484.050 616.500 ;
        RECT 470.400 605.400 474.600 606.600 ;
        RECT 475.950 605.400 478.050 607.500 ;
        RECT 466.950 583.950 469.050 586.050 ;
        RECT 470.400 580.050 471.600 605.400 ;
        RECT 476.400 604.050 477.600 605.400 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 472.950 598.950 475.050 601.050 ;
        RECT 454.950 577.950 457.050 580.050 ;
        RECT 460.950 577.950 463.050 580.050 ;
        RECT 469.950 577.950 472.050 580.050 ;
        RECT 442.950 571.950 445.050 574.050 ;
        RECT 448.950 573.000 451.050 577.050 ;
        RECT 457.950 574.950 460.050 577.050 ;
        RECT 449.400 571.050 450.600 573.000 ;
        RECT 445.950 568.950 448.050 571.050 ;
        RECT 448.950 568.950 451.050 571.050 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 446.400 567.900 447.600 568.950 ;
        RECT 452.400 567.900 453.600 568.950 ;
        RECT 439.950 565.800 442.050 567.900 ;
        RECT 445.950 565.800 448.050 567.900 ;
        RECT 451.950 565.800 454.050 567.900 ;
        RECT 458.400 565.050 459.600 574.950 ;
        RECT 433.950 562.950 436.050 565.050 ;
        RECT 457.950 562.950 460.050 565.050 ;
        RECT 434.400 553.050 435.600 562.950 ;
        RECT 448.950 553.950 451.050 556.050 ;
        RECT 433.950 550.950 436.050 553.050 ;
        RECT 436.950 547.950 439.050 550.050 ;
        RECT 430.950 541.950 433.050 544.050 ;
        RECT 427.950 535.950 430.050 538.050 ;
        RECT 412.950 528.000 415.050 532.050 ;
        RECT 418.950 529.950 421.050 532.050 ;
        RECT 413.400 526.050 414.600 528.000 ;
        RECT 419.400 526.050 420.600 529.950 ;
        RECT 427.950 526.950 430.050 532.050 ;
        RECT 430.950 528.000 433.050 532.050 ;
        RECT 431.400 526.050 432.600 528.000 ;
        RECT 437.400 526.050 438.600 547.950 ;
        RECT 449.400 529.200 450.600 553.950 ;
        RECT 454.950 550.950 457.050 553.050 ;
        RECT 451.950 535.950 454.050 538.050 ;
        RECT 442.950 527.100 445.050 529.200 ;
        RECT 448.950 527.100 451.050 529.200 ;
        RECT 443.400 526.050 444.600 527.100 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 433.950 523.950 436.050 526.050 ;
        RECT 436.950 523.950 439.050 526.050 ;
        RECT 439.950 523.950 442.050 526.050 ;
        RECT 442.950 523.950 445.050 526.050 ;
        RECT 416.400 514.050 417.600 523.950 ;
        RECT 421.950 514.950 424.050 517.050 ;
        RECT 415.950 511.950 418.050 514.050 ;
        RECT 409.950 505.950 412.050 508.050 ;
        RECT 406.950 502.950 409.050 505.050 ;
        RECT 403.950 496.950 406.050 499.050 ;
        RECT 410.400 496.050 411.600 505.950 ;
        RECT 415.950 502.950 418.050 505.050 ;
        RECT 412.950 496.950 415.050 499.050 ;
        RECT 401.400 494.400 405.600 495.600 ;
        RECT 404.400 493.050 405.600 494.400 ;
        RECT 409.950 493.950 412.050 496.050 ;
        RECT 403.950 490.950 406.050 493.050 ;
        RECT 406.950 490.950 409.050 493.050 ;
        RECT 400.950 487.950 403.050 490.050 ;
        RECT 401.400 469.050 402.600 487.950 ;
        RECT 407.400 484.050 408.600 490.950 ;
        RECT 409.950 487.950 412.050 490.050 ;
        RECT 406.950 481.950 409.050 484.050 ;
        RECT 403.950 478.950 406.050 481.050 ;
        RECT 400.950 466.950 403.050 469.050 ;
        RECT 397.950 451.950 400.050 454.050 ;
        RECT 401.400 450.600 402.600 466.950 ;
        RECT 404.400 457.050 405.600 478.950 ;
        RECT 403.950 454.950 406.050 457.050 ;
        RECT 406.950 451.950 409.050 454.050 ;
        RECT 401.400 449.400 405.600 450.600 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 391.950 445.950 394.050 448.050 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 392.400 444.000 393.600 445.950 ;
        RECT 388.950 439.950 391.050 442.050 ;
        RECT 391.950 439.950 394.050 444.000 ;
        RECT 382.950 421.950 385.050 424.050 ;
        RECT 376.950 415.950 379.050 418.050 ;
        RECT 379.950 417.000 382.050 421.050 ;
        RECT 380.400 415.050 381.600 417.000 ;
        RECT 389.400 415.050 390.600 439.950 ;
        RECT 398.400 430.050 399.600 445.950 ;
        RECT 404.400 445.050 405.600 449.400 ;
        RECT 403.950 442.950 406.050 445.050 ;
        RECT 407.400 439.050 408.600 451.950 ;
        RECT 410.400 451.050 411.600 487.950 ;
        RECT 413.400 466.050 414.600 496.950 ;
        RECT 416.400 487.050 417.600 502.950 ;
        RECT 422.400 499.050 423.600 514.950 ;
        RECT 425.400 505.050 426.600 523.950 ;
        RECT 434.400 522.900 435.600 523.950 ;
        RECT 433.950 520.800 436.050 522.900 ;
        RECT 440.400 511.050 441.600 523.950 ;
        RECT 445.950 517.950 448.050 520.050 ;
        RECT 439.950 508.950 442.050 511.050 ;
        RECT 433.950 505.950 436.050 508.050 ;
        RECT 424.950 502.950 427.050 505.050 ;
        RECT 421.950 496.950 424.050 499.050 ;
        RECT 424.950 494.100 427.050 496.200 ;
        RECT 425.400 493.050 426.600 494.100 ;
        RECT 430.950 493.950 433.050 499.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 427.950 490.950 430.050 493.050 ;
        RECT 422.400 489.900 423.600 490.950 ;
        RECT 428.400 489.900 429.600 490.950 ;
        RECT 421.950 487.800 424.050 489.900 ;
        RECT 415.950 484.950 418.050 487.050 ;
        RECT 427.950 484.950 430.050 489.900 ;
        RECT 434.400 487.050 435.600 505.950 ;
        RECT 446.400 502.050 447.600 517.950 ;
        RECT 449.400 517.050 450.600 527.100 ;
        RECT 448.950 514.950 451.050 517.050 ;
        RECT 452.400 508.050 453.600 535.950 ;
        RECT 451.950 505.950 454.050 508.050 ;
        RECT 455.400 505.050 456.600 550.950 ;
        RECT 457.950 544.950 460.050 547.050 ;
        RECT 458.400 528.600 459.600 544.950 ;
        RECT 461.400 535.050 462.600 577.950 ;
        RECT 463.950 571.950 466.050 574.050 ;
        RECT 464.400 565.050 465.600 571.950 ;
        RECT 473.400 571.050 474.600 598.950 ;
        RECT 482.100 594.600 483.300 614.400 ;
        RECT 484.950 605.400 487.050 607.500 ;
        RECT 485.400 604.050 486.600 605.400 ;
        RECT 484.950 601.950 487.050 604.050 ;
        RECT 491.400 603.600 492.600 637.950 ;
        RECT 494.400 613.050 495.600 655.950 ;
        RECT 497.400 616.050 498.600 670.950 ;
        RECT 500.400 658.050 501.600 677.400 ;
        RECT 506.700 678.300 507.600 687.300 ;
        RECT 509.100 683.700 511.200 685.800 ;
        RECT 512.400 684.900 513.600 687.450 ;
        RECT 510.300 681.300 511.200 683.700 ;
        RECT 512.100 682.800 514.200 684.900 ;
        RECT 516.000 681.300 517.050 688.500 ;
        RECT 524.400 682.050 525.600 688.950 ;
        RECT 527.400 685.050 528.600 722.400 ;
        RECT 536.400 712.050 537.600 724.950 ;
        RECT 538.950 721.950 541.050 724.050 ;
        RECT 535.950 709.950 538.050 712.050 ;
        RECT 532.950 700.950 535.050 703.050 ;
        RECT 533.400 697.050 534.600 700.950 ;
        RECT 536.400 697.050 537.600 709.950 ;
        RECT 532.800 694.950 534.900 697.050 ;
        RECT 535.950 694.950 538.050 697.050 ;
        RECT 526.950 682.950 529.050 685.050 ;
        RECT 539.400 682.050 540.600 721.950 ;
        RECT 542.400 718.050 543.600 727.950 ;
        RECT 548.400 718.050 549.600 727.950 ;
        RECT 557.400 727.050 558.600 728.100 ;
        RECT 562.950 727.950 565.050 730.050 ;
        RECT 569.400 727.050 570.600 736.950 ;
        RECT 574.950 728.100 577.050 730.200 ;
        RECT 575.400 727.050 576.600 728.100 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 568.950 724.950 571.050 727.050 ;
        RECT 571.950 724.950 574.050 727.050 ;
        RECT 574.950 724.950 577.050 727.050 ;
        RECT 577.950 724.950 580.050 727.050 ;
        RECT 541.950 715.950 544.050 718.050 ;
        RECT 547.950 715.950 550.050 718.050 ;
        RECT 554.400 706.050 555.600 724.950 ;
        RECT 572.400 723.900 573.600 724.950 ;
        RECT 571.950 721.800 574.050 723.900 ;
        RECT 568.950 718.950 571.050 721.050 ;
        RECT 565.950 706.950 568.050 709.050 ;
        RECT 541.950 703.950 544.050 706.050 ;
        RECT 553.950 703.950 556.050 706.050 ;
        RECT 542.400 685.050 543.600 703.950 ;
        RECT 547.950 700.950 550.050 703.050 ;
        RECT 541.950 682.950 544.050 685.050 ;
        RECT 510.300 680.100 517.050 681.300 ;
        RECT 513.150 678.300 515.250 679.200 ;
        RECT 506.700 677.100 515.250 678.300 ;
        RECT 508.200 675.300 510.300 677.100 ;
        RECT 512.100 674.100 514.200 676.200 ;
        RECT 516.150 674.700 517.050 680.100 ;
        RECT 517.950 679.950 520.050 682.050 ;
        RECT 523.950 679.950 526.050 682.050 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 538.950 679.950 541.050 682.050 ;
        RECT 518.400 677.400 519.600 679.950 ;
        RECT 512.400 661.050 513.600 674.100 ;
        RECT 515.400 672.600 517.500 674.700 ;
        RECT 523.950 673.950 526.050 676.050 ;
        RECT 511.950 658.950 514.050 661.050 ;
        RECT 499.950 655.950 502.050 658.050 ;
        RECT 517.950 655.950 520.050 658.050 ;
        RECT 505.950 650.100 508.050 652.200 ;
        RECT 511.950 650.100 514.050 652.200 ;
        RECT 506.400 649.050 507.600 650.100 ;
        RECT 512.400 649.050 513.600 650.100 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 508.950 646.950 511.050 649.050 ;
        RECT 511.950 646.950 514.050 649.050 ;
        RECT 496.950 613.950 499.050 616.050 ;
        RECT 493.950 610.950 496.050 613.050 ;
        RECT 499.950 610.950 502.050 613.050 ;
        RECT 500.400 604.050 501.600 610.950 ;
        RECT 503.400 610.050 504.600 646.950 ;
        RECT 502.950 607.950 505.050 610.050 ;
        RECT 505.950 606.600 508.050 607.200 ;
        RECT 509.400 606.600 510.600 646.950 ;
        RECT 518.400 637.050 519.600 655.950 ;
        RECT 524.400 652.200 525.600 673.950 ;
        RECT 533.400 673.050 534.600 679.950 ;
        RECT 532.950 670.950 535.050 673.050 ;
        RECT 541.950 670.950 544.050 673.050 ;
        RECT 535.950 664.950 538.050 667.050 ;
        RECT 529.950 655.950 532.050 658.050 ;
        RECT 523.950 650.100 526.050 652.200 ;
        RECT 524.400 649.050 525.600 650.100 ;
        RECT 530.400 649.050 531.600 655.950 ;
        RECT 536.400 652.050 537.600 664.950 ;
        RECT 538.950 658.950 541.050 661.050 ;
        RECT 535.950 649.950 538.050 652.050 ;
        RECT 523.950 646.950 526.050 649.050 ;
        RECT 526.950 646.950 529.050 649.050 ;
        RECT 529.950 646.950 532.050 649.050 ;
        RECT 532.950 646.950 535.050 649.050 ;
        RECT 517.950 634.950 520.050 637.050 ;
        RECT 527.400 619.050 528.600 646.950 ;
        RECT 533.400 645.900 534.600 646.950 ;
        RECT 532.950 643.800 535.050 645.900 ;
        RECT 535.950 640.950 538.050 643.050 ;
        RECT 536.400 631.050 537.600 640.950 ;
        RECT 535.950 628.950 538.050 631.050 ;
        RECT 539.400 622.050 540.600 658.950 ;
        RECT 542.400 640.050 543.600 670.950 ;
        RECT 548.400 651.600 549.600 700.950 ;
        RECT 553.950 700.800 556.050 702.900 ;
        RECT 554.400 682.050 555.600 700.800 ;
        RECT 559.950 683.100 562.050 685.200 ;
        RECT 560.400 682.050 561.600 683.100 ;
        RECT 553.950 679.950 556.050 682.050 ;
        RECT 556.950 679.950 559.050 682.050 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 557.400 667.050 558.600 679.950 ;
        RECT 566.400 679.050 567.600 706.950 ;
        RECT 565.950 676.950 568.050 679.050 ;
        RECT 556.950 664.950 559.050 667.050 ;
        RECT 556.950 658.950 559.050 661.050 ;
        RECT 557.400 654.600 558.600 658.950 ;
        RECT 562.950 656.400 565.050 658.500 ;
        RECT 557.400 653.400 561.600 654.600 ;
        RECT 560.400 652.500 561.600 653.400 ;
        RECT 545.400 650.400 549.600 651.600 ;
        RECT 541.950 637.950 544.050 640.050 ;
        RECT 545.400 628.050 546.600 650.400 ;
        RECT 553.950 650.100 556.050 652.200 ;
        RECT 559.950 650.400 562.050 652.500 ;
        RECT 554.400 649.050 555.600 650.100 ;
        RECT 560.400 649.050 561.600 650.400 ;
        RECT 550.950 646.950 553.050 649.050 ;
        RECT 553.950 646.950 556.050 649.050 ;
        RECT 559.950 646.950 562.050 649.050 ;
        RECT 551.400 640.050 552.600 646.950 ;
        RECT 556.950 643.950 559.050 646.050 ;
        RECT 550.800 637.950 552.900 640.050 ;
        RECT 553.950 637.950 556.050 640.050 ;
        RECT 544.950 625.950 547.050 628.050 ;
        RECT 538.950 619.950 541.050 622.050 ;
        RECT 547.950 619.950 550.050 622.050 ;
        RECT 517.950 615.300 520.050 617.400 ;
        RECT 526.950 616.950 529.050 619.050 ;
        RECT 518.850 611.700 520.050 615.300 ;
        RECT 523.950 613.950 526.050 616.050 ;
        RECT 538.950 614.400 541.050 616.500 ;
        RECT 517.950 609.600 520.050 611.700 ;
        RECT 505.950 605.400 510.600 606.600 ;
        RECT 505.950 605.100 508.050 605.400 ;
        RECT 506.400 604.050 507.600 605.100 ;
        RECT 493.950 603.600 496.050 604.050 ;
        RECT 491.400 602.400 496.050 603.600 ;
        RECT 493.950 601.950 496.050 602.400 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 502.950 601.950 505.050 604.050 ;
        RECT 505.950 601.950 508.050 604.050 ;
        RECT 514.950 601.950 517.050 604.050 ;
        RECT 494.400 595.050 495.600 601.950 ;
        RECT 503.400 600.900 504.600 601.950 ;
        RECT 502.950 598.800 505.050 600.900 ;
        RECT 508.950 598.950 511.050 601.050 ;
        RECT 515.400 600.600 516.600 601.950 ;
        RECT 481.950 592.500 484.050 594.600 ;
        RECT 493.950 592.950 496.050 595.050 ;
        RECT 509.400 589.050 510.600 598.950 ;
        RECT 514.950 598.500 517.050 600.600 ;
        RECT 511.950 592.950 514.050 595.050 ;
        RECT 518.850 594.600 520.050 609.600 ;
        RECT 524.400 600.600 525.600 613.950 ;
        RECT 526.950 604.950 529.050 607.050 ;
        RECT 532.950 605.400 535.050 607.500 ;
        RECT 523.950 598.500 526.050 600.600 ;
        RECT 493.950 586.950 496.050 589.050 ;
        RECT 508.950 586.950 511.050 589.050 ;
        RECT 478.950 583.950 481.050 586.050 ;
        RECT 479.400 580.050 480.600 583.950 ;
        RECT 481.950 580.950 484.050 583.050 ;
        RECT 478.950 577.950 481.050 580.050 ;
        RECT 479.400 571.050 480.600 577.950 ;
        RECT 482.400 574.050 483.600 580.950 ;
        RECT 487.950 578.400 490.050 580.500 ;
        RECT 481.950 573.600 486.000 574.050 ;
        RECT 481.950 571.950 486.600 573.600 ;
        RECT 485.400 571.050 486.600 571.950 ;
        RECT 469.950 568.950 472.050 571.050 ;
        RECT 472.950 568.950 475.050 571.050 ;
        RECT 475.950 568.950 478.050 571.050 ;
        RECT 478.950 568.950 481.050 571.050 ;
        RECT 484.950 568.950 487.050 571.050 ;
        RECT 470.400 567.000 471.600 568.950 ;
        RECT 476.400 567.900 477.600 568.950 ;
        RECT 463.950 562.950 466.050 565.050 ;
        RECT 469.950 562.950 472.050 567.000 ;
        RECT 475.950 565.800 478.050 567.900 ;
        RECT 476.400 562.050 477.600 565.800 ;
        RECT 481.950 562.950 484.050 565.050 ;
        RECT 488.850 563.400 490.050 578.400 ;
        RECT 475.950 559.950 478.050 562.050 ;
        RECT 478.950 553.950 481.050 556.050 ;
        RECT 475.950 544.950 478.050 547.050 ;
        RECT 476.400 541.050 477.600 544.950 ;
        RECT 479.400 541.050 480.600 553.950 ;
        RECT 475.800 538.950 477.900 541.050 ;
        RECT 478.950 538.950 481.050 541.050 ;
        RECT 482.400 535.050 483.600 562.950 ;
        RECT 487.950 561.300 490.050 563.400 ;
        RECT 488.850 557.700 490.050 561.300 ;
        RECT 494.400 561.600 495.600 586.950 ;
        RECT 512.400 586.050 513.600 592.950 ;
        RECT 517.950 592.500 520.050 594.600 ;
        RECT 524.400 592.050 525.600 598.500 ;
        RECT 523.950 589.950 526.050 592.050 ;
        RECT 527.400 589.050 528.600 604.950 ;
        RECT 533.400 604.050 534.600 605.400 ;
        RECT 532.950 601.950 535.050 604.050 ;
        RECT 539.100 594.600 540.300 614.400 ;
        RECT 541.950 605.400 544.050 607.500 ;
        RECT 542.400 604.050 543.600 605.400 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 544.950 598.950 547.050 601.050 ;
        RECT 545.400 595.050 546.600 598.950 ;
        RECT 538.950 592.500 541.050 594.600 ;
        RECT 544.950 592.950 547.050 595.050 ;
        RECT 514.950 586.950 517.050 589.050 ;
        RECT 526.950 586.950 529.050 589.050 ;
        RECT 511.950 583.950 514.050 586.050 ;
        RECT 508.950 578.400 511.050 580.500 ;
        RECT 496.950 574.950 499.050 577.050 ;
        RECT 497.400 568.050 498.600 574.950 ;
        RECT 502.950 568.950 505.050 571.050 ;
        RECT 496.950 565.950 499.050 568.050 ;
        RECT 503.400 567.600 504.600 568.950 ;
        RECT 502.800 565.500 504.900 567.600 ;
        RECT 505.950 565.950 508.050 568.050 ;
        RECT 496.950 561.600 499.050 562.050 ;
        RECT 506.400 561.600 507.600 565.950 ;
        RECT 494.400 560.400 499.050 561.600 ;
        RECT 496.950 559.950 499.050 560.400 ;
        RECT 503.400 560.400 507.600 561.600 ;
        RECT 487.950 555.600 490.050 557.700 ;
        RECT 497.400 550.050 498.600 559.950 ;
        RECT 503.400 553.050 504.600 560.400 ;
        RECT 509.100 558.600 510.300 578.400 ;
        RECT 515.400 574.050 516.600 586.950 ;
        RECT 517.950 583.950 520.050 586.050 ;
        RECT 541.950 583.950 544.050 586.050 ;
        RECT 514.950 571.950 517.050 574.050 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 512.400 567.600 513.600 568.950 ;
        RECT 518.400 567.600 519.600 583.950 ;
        RECT 520.950 580.950 523.050 583.050 ;
        RECT 511.950 565.500 514.050 567.600 ;
        RECT 517.950 565.500 520.050 567.600 ;
        RECT 521.400 565.050 522.600 580.950 ;
        RECT 523.950 576.600 526.050 577.050 ;
        RECT 523.950 575.400 534.600 576.600 ;
        RECT 523.950 574.950 526.050 575.400 ;
        RECT 526.950 572.100 529.050 574.200 ;
        RECT 527.400 571.050 528.600 572.100 ;
        RECT 533.400 571.050 534.600 575.400 ;
        RECT 526.950 568.950 529.050 571.050 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 520.950 562.950 523.050 565.050 ;
        RECT 508.950 556.500 511.050 558.600 ;
        RECT 502.950 550.950 505.050 553.050 ;
        RECT 490.950 547.950 493.050 550.050 ;
        RECT 496.950 547.950 499.050 550.050 ;
        RECT 487.950 544.950 490.050 547.050 ;
        RECT 484.950 538.950 487.050 541.050 ;
        RECT 460.950 532.950 463.050 535.050 ;
        RECT 472.950 532.950 475.050 535.050 ;
        RECT 481.950 532.950 484.050 535.050 ;
        RECT 458.400 527.400 462.600 528.600 ;
        RECT 461.400 526.050 462.600 527.400 ;
        RECT 466.950 527.100 469.050 529.200 ;
        RECT 473.400 529.050 474.600 532.950 ;
        RECT 467.400 526.050 468.600 527.100 ;
        RECT 472.950 526.950 475.050 529.050 ;
        RECT 478.950 527.100 481.050 529.200 ;
        RECT 479.400 526.050 480.600 527.100 ;
        RECT 485.400 526.050 486.600 538.950 ;
        RECT 488.400 529.050 489.600 544.950 ;
        RECT 487.950 526.950 490.050 529.050 ;
        RECT 460.950 523.950 463.050 526.050 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 469.950 523.950 472.050 526.050 ;
        RECT 478.950 523.950 481.050 526.050 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 454.950 502.950 457.050 505.050 ;
        RECT 436.950 499.950 439.050 502.050 ;
        RECT 445.950 499.950 448.050 502.050 ;
        RECT 460.950 499.950 463.050 502.050 ;
        RECT 433.950 484.950 436.050 487.050 ;
        RECT 416.400 475.050 417.600 484.950 ;
        RECT 430.950 481.950 433.050 484.050 ;
        RECT 427.950 478.950 430.050 481.050 ;
        RECT 415.950 472.950 418.050 475.050 ;
        RECT 421.950 472.950 424.050 475.050 ;
        RECT 412.950 463.950 415.050 466.050 ;
        RECT 413.400 454.050 414.600 463.950 ;
        RECT 422.400 454.200 423.600 472.950 ;
        RECT 424.950 466.950 427.050 469.050 ;
        RECT 425.400 463.050 426.600 466.950 ;
        RECT 424.950 460.950 427.050 463.050 ;
        RECT 412.950 451.950 415.050 454.050 ;
        RECT 421.950 452.100 424.050 454.200 ;
        RECT 409.950 448.950 412.050 451.050 ;
        RECT 415.950 449.100 418.050 451.200 ;
        RECT 416.400 448.050 417.600 449.100 ;
        RECT 421.950 448.950 424.050 451.050 ;
        RECT 422.400 448.050 423.600 448.950 ;
        RECT 412.950 445.950 415.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 413.400 441.600 414.600 445.950 ;
        RECT 413.400 440.400 417.600 441.600 ;
        RECT 406.950 436.950 409.050 439.050 ;
        RECT 397.950 427.950 400.050 430.050 ;
        RECT 409.950 424.950 412.050 427.050 ;
        RECT 410.400 421.050 411.600 424.950 ;
        RECT 391.950 415.950 394.050 418.050 ;
        RECT 403.950 416.100 406.050 418.200 ;
        RECT 409.950 417.000 412.050 421.050 ;
        RECT 379.950 412.950 382.050 415.050 ;
        RECT 382.950 412.950 385.050 415.050 ;
        RECT 388.950 412.950 391.050 415.050 ;
        RECT 376.950 406.950 379.050 409.050 ;
        RECT 373.950 400.950 376.050 403.050 ;
        RECT 377.400 382.050 378.600 406.950 ;
        RECT 379.950 403.950 382.050 409.050 ;
        RECT 383.400 403.050 384.600 412.950 ;
        RECT 385.950 409.950 388.050 412.050 ;
        RECT 382.950 400.950 385.050 403.050 ;
        RECT 386.400 400.050 387.600 409.950 ;
        RECT 392.400 409.050 393.600 415.950 ;
        RECT 404.400 415.050 405.600 416.100 ;
        RECT 410.400 415.050 411.600 417.000 ;
        RECT 394.950 412.950 397.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 391.950 406.950 394.050 409.050 ;
        RECT 395.400 405.600 396.600 412.950 ;
        RECT 401.400 411.900 402.600 412.950 ;
        RECT 407.400 411.900 408.600 412.950 ;
        RECT 400.950 409.800 403.050 411.900 ;
        RECT 406.950 409.800 409.050 411.900 ;
        RECT 392.400 404.400 396.600 405.600 ;
        RECT 397.950 405.600 400.050 409.050 ;
        RECT 412.950 408.600 415.050 412.050 ;
        RECT 416.400 411.900 417.600 440.400 ;
        RECT 419.400 439.050 420.600 445.950 ;
        RECT 424.950 442.950 427.050 445.050 ;
        RECT 418.950 436.950 421.050 439.050 ;
        RECT 418.950 433.800 421.050 435.900 ;
        RECT 419.400 418.050 420.600 433.800 ;
        RECT 425.400 418.200 426.600 442.950 ;
        RECT 428.400 436.050 429.600 478.950 ;
        RECT 431.400 469.050 432.600 481.950 ;
        RECT 433.950 475.950 436.050 478.050 ;
        RECT 430.950 466.950 433.050 469.050 ;
        RECT 434.400 457.050 435.600 475.950 ;
        RECT 437.400 460.050 438.600 499.950 ;
        RECT 454.950 496.950 457.050 499.050 ;
        RECT 445.950 494.100 448.050 496.200 ;
        RECT 446.400 493.050 447.600 494.100 ;
        RECT 442.950 490.950 445.050 493.050 ;
        RECT 445.950 490.950 448.050 493.050 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 439.950 487.950 442.050 490.050 ;
        RECT 443.400 489.900 444.600 490.950 ;
        RECT 440.400 484.050 441.600 487.950 ;
        RECT 442.950 487.800 445.050 489.900 ;
        RECT 439.950 481.950 442.050 484.050 ;
        RECT 439.950 472.950 442.050 475.050 ;
        RECT 436.950 457.950 439.050 460.050 ;
        RECT 433.950 454.950 436.050 457.050 ;
        RECT 433.950 450.000 436.050 453.900 ;
        RECT 434.400 448.050 435.600 450.000 ;
        RECT 440.400 448.050 441.600 472.950 ;
        RECT 449.400 463.050 450.600 490.950 ;
        RECT 451.950 481.950 454.050 484.050 ;
        RECT 448.950 460.950 451.050 463.050 ;
        RECT 445.950 450.000 448.050 454.050 ;
        RECT 449.400 451.050 450.600 460.950 ;
        RECT 446.400 448.050 447.600 450.000 ;
        RECT 448.950 448.950 451.050 451.050 ;
        RECT 433.950 445.950 436.050 448.050 ;
        RECT 436.950 445.950 439.050 448.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 430.950 442.950 433.050 445.050 ;
        RECT 437.400 444.900 438.600 445.950 ;
        RECT 427.950 433.950 430.050 436.050 ;
        RECT 431.400 430.050 432.600 442.950 ;
        RECT 436.950 442.800 439.050 444.900 ;
        RECT 443.400 433.050 444.600 445.950 ;
        RECT 452.400 439.050 453.600 481.950 ;
        RECT 455.400 481.050 456.600 496.950 ;
        RECT 461.400 493.050 462.600 499.950 ;
        RECT 464.400 499.050 465.600 523.950 ;
        RECT 470.400 514.050 471.600 523.950 ;
        RECT 472.800 520.950 474.900 523.050 ;
        RECT 475.950 520.950 478.050 523.050 ;
        RECT 473.400 517.050 474.600 520.950 ;
        RECT 472.950 514.950 475.050 517.050 ;
        RECT 469.950 511.950 472.050 514.050 ;
        RECT 466.950 508.950 469.050 511.050 ;
        RECT 463.950 496.950 466.050 499.050 ;
        RECT 467.400 493.050 468.600 508.950 ;
        RECT 470.400 502.050 471.600 511.950 ;
        RECT 469.950 499.950 472.050 502.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 466.950 490.950 469.050 493.050 ;
        RECT 469.950 490.950 472.050 493.050 ;
        RECT 464.400 484.050 465.600 490.950 ;
        RECT 470.400 489.900 471.600 490.950 ;
        RECT 469.950 487.800 472.050 489.900 ;
        RECT 463.950 481.950 466.050 484.050 ;
        RECT 454.950 478.950 457.050 481.050 ;
        RECT 469.950 475.950 472.050 478.050 ;
        RECT 454.950 471.600 457.050 472.050 ;
        RECT 460.950 471.600 463.050 472.050 ;
        RECT 454.950 470.400 463.050 471.600 ;
        RECT 454.950 469.950 457.050 470.400 ;
        RECT 460.950 469.950 463.050 470.400 ;
        RECT 457.950 466.950 460.050 469.050 ;
        RECT 454.950 457.950 457.050 460.050 ;
        RECT 455.400 445.050 456.600 457.950 ;
        RECT 458.400 451.050 459.600 466.950 ;
        RECT 470.400 466.050 471.600 475.950 ;
        RECT 476.400 466.050 477.600 520.950 ;
        RECT 478.950 517.950 481.050 520.050 ;
        RECT 479.400 511.050 480.600 517.950 ;
        RECT 482.400 517.050 483.600 523.950 ;
        RECT 487.950 520.950 490.050 523.050 ;
        RECT 481.950 514.950 484.050 517.050 ;
        RECT 488.400 514.050 489.600 520.950 ;
        RECT 491.400 520.050 492.600 547.950 ;
        RECT 530.400 544.050 531.600 568.950 ;
        RECT 536.400 562.050 537.600 568.950 ;
        RECT 535.950 559.950 538.050 562.050 ;
        RECT 542.400 544.050 543.600 583.950 ;
        RECT 548.400 577.050 549.600 619.950 ;
        RECT 550.950 616.950 553.050 619.050 ;
        RECT 551.400 586.050 552.600 616.950 ;
        RECT 554.400 607.050 555.600 637.950 ;
        RECT 557.400 625.050 558.600 643.950 ;
        RECT 563.850 641.400 565.050 656.400 ;
        RECT 562.950 639.300 565.050 641.400 ;
        RECT 563.850 635.700 565.050 639.300 ;
        RECT 562.950 633.600 565.050 635.700 ;
        RECT 569.400 625.050 570.600 718.950 ;
        RECT 578.400 718.050 579.600 724.950 ;
        RECT 580.950 721.950 583.050 724.050 ;
        RECT 577.950 715.950 580.050 718.050 ;
        RECT 571.950 691.950 574.050 694.050 ;
        RECT 572.400 685.200 573.600 691.950 ;
        RECT 581.400 691.050 582.600 721.950 ;
        RECT 580.950 688.950 583.050 691.050 ;
        RECT 584.400 687.600 585.600 751.950 ;
        RECT 589.950 736.950 592.050 739.050 ;
        RECT 586.950 733.950 589.050 736.050 ;
        RECT 587.400 703.050 588.600 733.950 ;
        RECT 590.400 709.050 591.600 736.950 ;
        RECT 596.400 733.050 597.600 754.950 ;
        RECT 599.400 739.050 600.600 793.950 ;
        RECT 604.950 781.950 607.050 784.050 ;
        RECT 605.400 778.050 606.600 781.950 ;
        RECT 604.950 775.950 607.050 778.050 ;
        RECT 601.950 772.950 604.050 775.050 ;
        RECT 602.400 769.050 603.600 772.950 ;
        RECT 601.950 766.950 604.050 769.050 ;
        RECT 605.400 760.050 606.600 775.950 ;
        RECT 607.800 768.000 609.900 769.050 ;
        RECT 607.800 766.950 610.050 768.000 ;
        RECT 610.950 766.950 613.050 769.050 ;
        RECT 607.950 763.950 610.050 766.950 ;
        RECT 611.400 760.050 612.600 766.950 ;
        RECT 614.400 766.050 615.600 811.950 ;
        RECT 623.400 805.050 624.600 820.950 ;
        RECT 628.950 806.100 631.050 808.200 ;
        RECT 629.400 805.050 630.600 806.100 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 620.400 801.900 621.600 802.950 ;
        RECT 626.400 801.900 627.600 802.950 ;
        RECT 619.950 799.800 622.050 801.900 ;
        RECT 625.950 799.800 628.050 801.900 ;
        RECT 632.400 796.050 633.600 802.950 ;
        RECT 638.400 802.050 639.600 829.950 ;
        RECT 641.400 802.050 642.600 839.100 ;
        RECT 647.400 838.050 648.600 839.100 ;
        RECT 653.400 838.050 654.600 839.100 ;
        RECT 646.950 835.950 649.050 838.050 ;
        RECT 649.950 835.950 652.050 838.050 ;
        RECT 652.950 835.950 655.050 838.050 ;
        RECT 650.400 834.900 651.600 835.950 ;
        RECT 649.950 832.800 652.050 834.900 ;
        RECT 655.950 826.950 658.050 829.050 ;
        RECT 651.000 807.600 655.050 808.050 ;
        RECT 650.400 805.950 655.050 807.600 ;
        RECT 650.400 805.050 651.600 805.950 ;
        RECT 646.950 802.950 649.050 805.050 ;
        RECT 649.950 802.950 652.050 805.050 ;
        RECT 634.950 799.950 637.050 802.050 ;
        RECT 637.950 799.950 640.050 802.050 ;
        RECT 640.950 801.600 643.050 802.050 ;
        RECT 647.400 801.900 648.600 802.950 ;
        RECT 656.400 802.050 657.600 826.950 ;
        RECT 659.400 817.050 660.600 872.400 ;
        RECT 661.950 871.950 664.050 872.400 ;
        RECT 683.400 853.050 684.600 880.950 ;
        RECT 689.400 879.900 690.600 880.950 ;
        RECT 695.400 879.900 696.600 895.950 ;
        RECT 688.950 877.800 691.050 879.900 ;
        RECT 694.950 877.800 697.050 879.900 ;
        RECT 688.950 853.950 691.050 856.050 ;
        RECT 661.950 850.950 664.050 853.050 ;
        RECT 682.950 850.950 685.050 853.050 ;
        RECT 658.950 814.950 661.050 817.050 ;
        RECT 662.400 814.050 663.600 850.950 ;
        RECT 676.950 844.950 679.050 847.050 ;
        RECT 664.950 839.100 667.050 841.200 ;
        RECT 670.950 839.100 673.050 841.200 ;
        RECT 665.400 829.050 666.600 839.100 ;
        RECT 671.400 838.050 672.600 839.100 ;
        RECT 677.400 838.050 678.600 844.950 ;
        RECT 689.400 838.050 690.600 853.950 ;
        RECT 694.950 839.100 697.050 841.200 ;
        RECT 698.400 840.600 699.600 908.100 ;
        RECT 700.950 904.950 703.050 907.050 ;
        RECT 701.400 886.050 702.600 904.950 ;
        RECT 710.400 898.050 711.600 910.950 ;
        RECT 721.950 910.800 724.050 912.900 ;
        RECT 728.400 901.050 729.600 913.950 ;
        RECT 734.400 901.050 735.600 917.100 ;
        RECT 740.400 907.050 741.600 931.950 ;
        RECT 841.950 925.950 844.050 928.050 ;
        RECT 745.950 922.950 748.050 925.050 ;
        RECT 790.950 922.950 793.050 925.050 ;
        RECT 746.400 916.050 747.600 922.950 ;
        RECT 751.950 918.000 754.050 922.050 ;
        RECT 781.950 919.950 784.050 922.050 ;
        RECT 752.400 916.050 753.600 918.000 ;
        RECT 769.950 917.100 772.050 919.200 ;
        RECT 770.400 916.050 771.600 917.100 ;
        RECT 745.950 913.950 748.050 916.050 ;
        RECT 748.950 913.950 751.050 916.050 ;
        RECT 751.950 913.950 754.050 916.050 ;
        RECT 754.950 913.950 757.050 916.050 ;
        RECT 766.950 913.950 769.050 916.050 ;
        RECT 769.950 913.950 772.050 916.050 ;
        RECT 772.950 913.950 775.050 916.050 ;
        RECT 739.950 904.950 742.050 907.050 ;
        RECT 718.950 898.950 721.050 901.050 ;
        RECT 727.950 898.950 730.050 901.050 ;
        RECT 733.950 898.950 736.050 901.050 ;
        RECT 709.950 897.600 712.050 898.050 ;
        RECT 709.950 896.400 714.600 897.600 ;
        RECT 709.950 895.950 712.050 896.400 ;
        RECT 706.950 892.950 709.050 895.050 ;
        RECT 700.950 883.950 703.050 886.050 ;
        RECT 707.400 883.050 708.600 892.950 ;
        RECT 713.400 886.050 714.600 896.400 ;
        RECT 715.950 892.950 718.050 895.050 ;
        RECT 712.950 883.950 715.050 886.050 ;
        RECT 703.950 880.950 706.050 883.050 ;
        RECT 706.950 880.950 709.050 883.050 ;
        RECT 709.950 880.950 712.050 883.050 ;
        RECT 704.400 879.900 705.600 880.950 ;
        RECT 710.400 879.900 711.600 880.950 ;
        RECT 716.400 879.900 717.600 892.950 ;
        RECT 719.400 886.050 720.600 898.950 ;
        RECT 749.400 898.050 750.600 913.950 ;
        RECT 755.400 912.900 756.600 913.950 ;
        RECT 767.400 912.900 768.600 913.950 ;
        RECT 754.950 910.800 757.050 912.900 ;
        RECT 766.950 910.800 769.050 912.900 ;
        RECT 767.400 907.050 768.600 910.800 ;
        RECT 766.950 904.950 769.050 907.050 ;
        RECT 773.400 904.050 774.600 913.950 ;
        RECT 782.400 913.050 783.600 919.950 ;
        RECT 791.400 916.050 792.600 922.950 ;
        RECT 808.950 917.100 811.050 919.200 ;
        RECT 814.950 918.000 817.050 922.050 ;
        RECT 820.950 921.600 823.050 922.050 ;
        RECT 826.950 921.600 829.050 922.050 ;
        RECT 820.950 920.400 829.050 921.600 ;
        RECT 820.950 919.950 823.050 920.400 ;
        RECT 826.950 919.950 829.050 920.400 ;
        RECT 809.400 916.050 810.600 917.100 ;
        RECT 815.400 916.050 816.600 918.000 ;
        RECT 823.950 917.100 826.050 919.200 ;
        RECT 832.950 918.000 835.050 922.050 ;
        RECT 824.400 916.050 825.600 917.100 ;
        RECT 833.400 916.050 834.600 918.000 ;
        RECT 838.950 916.950 841.050 925.050 ;
        RECT 787.950 913.950 790.050 916.050 ;
        RECT 790.950 913.950 793.050 916.050 ;
        RECT 808.950 913.950 811.050 916.050 ;
        RECT 811.950 913.950 814.050 916.050 ;
        RECT 814.950 913.950 817.050 916.050 ;
        RECT 823.950 913.950 826.050 916.050 ;
        RECT 826.950 913.950 829.050 916.050 ;
        RECT 832.950 913.950 835.050 916.050 ;
        RECT 835.950 913.950 838.050 916.050 ;
        RECT 775.950 907.950 778.050 913.050 ;
        RECT 781.950 910.950 784.050 913.050 ;
        RECT 788.400 912.000 789.600 913.950 ;
        RECT 787.950 907.950 790.050 912.000 ;
        RECT 793.950 910.950 796.050 913.050 ;
        RECT 805.950 910.950 808.050 913.050 ;
        RECT 781.950 904.950 784.050 907.050 ;
        RECT 772.950 901.950 775.050 904.050 ;
        RECT 782.400 901.050 783.600 904.950 ;
        RECT 781.950 898.950 784.050 901.050 ;
        RECT 748.950 895.950 751.050 898.050 ;
        RECT 766.950 892.950 769.050 895.050 ;
        RECT 724.950 889.950 727.050 892.050 ;
        RECT 736.950 889.950 739.050 892.050 ;
        RECT 718.950 883.950 721.050 886.050 ;
        RECT 725.400 883.050 726.600 889.950 ;
        RECT 730.950 884.100 733.050 886.200 ;
        RECT 731.400 883.050 732.600 884.100 ;
        RECT 721.950 880.950 724.050 883.050 ;
        RECT 724.950 880.950 727.050 883.050 ;
        RECT 727.950 880.950 730.050 883.050 ;
        RECT 730.950 880.950 733.050 883.050 ;
        RECT 722.400 879.900 723.600 880.950 ;
        RECT 728.400 879.900 729.600 880.950 ;
        RECT 703.950 877.800 706.050 879.900 ;
        RECT 709.950 877.800 712.050 879.900 ;
        RECT 715.950 877.800 718.050 879.900 ;
        RECT 721.950 877.800 724.050 879.900 ;
        RECT 727.950 877.800 730.050 879.900 ;
        RECT 721.950 871.950 724.050 874.050 ;
        RECT 722.400 862.050 723.600 871.950 ;
        RECT 721.950 859.950 724.050 862.050 ;
        RECT 709.950 856.950 712.050 859.050 ;
        RECT 703.950 844.950 706.050 847.050 ;
        RECT 698.400 839.400 702.600 840.600 ;
        RECT 695.400 838.050 696.600 839.100 ;
        RECT 670.950 835.950 673.050 838.050 ;
        RECT 673.950 835.950 676.050 838.050 ;
        RECT 676.950 835.950 679.050 838.050 ;
        RECT 688.950 835.950 691.050 838.050 ;
        RECT 691.950 835.950 694.050 838.050 ;
        RECT 694.950 835.950 697.050 838.050 ;
        RECT 674.400 834.900 675.600 835.950 ;
        RECT 673.950 832.800 676.050 834.900 ;
        RECT 692.400 834.000 693.600 835.950 ;
        RECT 691.950 829.950 694.050 834.000 ;
        RECT 697.950 832.950 700.050 835.050 ;
        RECT 664.950 826.950 667.050 829.050 ;
        RECT 688.950 826.950 691.050 829.050 ;
        RECT 694.950 826.950 697.050 829.050 ;
        RECT 661.950 811.950 664.050 814.050 ;
        RECT 689.400 808.200 690.600 826.950 ;
        RECT 695.400 823.050 696.600 826.950 ;
        RECT 694.950 820.950 697.050 823.050 ;
        RECT 698.400 819.600 699.600 832.950 ;
        RECT 701.400 823.050 702.600 839.400 ;
        RECT 704.400 826.050 705.600 844.950 ;
        RECT 710.400 838.050 711.600 856.950 ;
        RECT 727.950 853.950 730.050 856.050 ;
        RECT 721.950 850.950 724.050 853.050 ;
        RECT 715.950 839.100 718.050 841.200 ;
        RECT 722.400 841.050 723.600 850.950 ;
        RECT 724.950 844.950 727.050 847.050 ;
        RECT 716.400 838.050 717.600 839.100 ;
        RECT 721.950 838.950 724.050 841.050 ;
        RECT 709.950 835.950 712.050 838.050 ;
        RECT 712.950 835.950 715.050 838.050 ;
        RECT 715.950 835.950 718.050 838.050 ;
        RECT 718.950 835.950 721.050 838.050 ;
        RECT 703.950 823.950 706.050 826.050 ;
        RECT 700.950 820.950 703.050 823.050 ;
        RECT 698.400 818.400 702.600 819.600 ;
        RECT 691.950 811.950 694.050 814.050 ;
        RECT 664.950 806.100 667.050 808.200 ;
        RECT 665.400 805.050 666.600 806.100 ;
        RECT 673.950 805.950 676.050 808.050 ;
        RECT 682.950 806.100 685.050 808.200 ;
        RECT 688.950 806.100 691.050 808.200 ;
        RECT 664.950 802.950 667.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 640.950 801.000 645.600 801.600 ;
        RECT 640.950 800.400 646.050 801.000 ;
        RECT 640.950 799.950 643.050 800.400 ;
        RECT 631.950 793.950 634.050 796.050 ;
        RECT 632.400 786.600 633.600 793.950 ;
        RECT 635.400 790.050 636.600 799.950 ;
        RECT 643.950 796.950 646.050 800.400 ;
        RECT 646.950 799.800 649.050 801.900 ;
        RECT 652.950 799.950 655.050 802.050 ;
        RECT 655.950 799.950 658.050 802.050 ;
        RECT 653.400 796.050 654.600 799.950 ;
        RECT 668.400 796.050 669.600 802.950 ;
        RECT 674.400 801.900 675.600 805.950 ;
        RECT 683.400 805.050 684.600 806.100 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 682.950 802.950 685.050 805.050 ;
        RECT 685.950 802.950 688.050 805.050 ;
        RECT 680.400 801.900 681.600 802.950 ;
        RECT 673.950 799.800 676.050 801.900 ;
        RECT 679.950 799.800 682.050 801.900 ;
        RECT 652.950 793.950 655.050 796.050 ;
        RECT 667.950 793.950 670.050 796.050 ;
        RECT 634.950 787.950 637.050 790.050 ;
        RECT 632.400 785.400 636.600 786.600 ;
        RECT 622.950 781.950 625.050 784.050 ;
        RECT 623.400 778.050 624.600 781.950 ;
        RECT 625.950 778.950 628.050 781.050 ;
        RECT 622.950 775.950 625.050 778.050 ;
        RECT 619.950 772.950 622.050 775.050 ;
        RECT 620.400 766.050 621.600 772.950 ;
        RECT 613.950 763.950 616.050 766.050 ;
        RECT 619.950 763.950 622.050 766.050 ;
        RECT 616.950 761.100 619.050 763.200 ;
        RECT 617.400 760.050 618.600 761.100 ;
        RECT 604.950 757.950 607.050 760.050 ;
        RECT 607.950 757.950 610.050 760.050 ;
        RECT 610.950 757.950 613.050 760.050 ;
        RECT 613.950 757.950 616.050 760.050 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 601.950 754.950 604.050 757.050 ;
        RECT 602.400 748.050 603.600 754.950 ;
        RECT 601.950 745.950 604.050 748.050 ;
        RECT 608.400 739.050 609.600 757.950 ;
        RECT 610.950 751.950 613.050 754.050 ;
        RECT 598.950 736.950 601.050 739.050 ;
        RECT 607.950 736.950 610.050 739.050 ;
        RECT 595.950 730.950 598.050 733.050 ;
        RECT 598.950 728.100 601.050 730.200 ;
        RECT 604.950 729.000 607.050 733.050 ;
        RECT 611.400 730.200 612.600 751.950 ;
        RECT 614.400 748.050 615.600 757.950 ;
        RECT 619.950 754.950 622.050 757.050 ;
        RECT 616.950 748.950 619.050 751.050 ;
        RECT 613.950 745.950 616.050 748.050 ;
        RECT 617.400 739.050 618.600 748.950 ;
        RECT 620.400 742.050 621.600 754.950 ;
        RECT 619.950 739.950 622.050 742.050 ;
        RECT 616.950 736.950 619.050 739.050 ;
        RECT 626.400 736.050 627.600 778.950 ;
        RECT 628.950 777.600 633.000 778.050 ;
        RECT 628.950 775.950 633.600 777.600 ;
        RECT 628.950 772.800 631.050 774.900 ;
        RECT 629.400 763.050 630.600 772.800 ;
        RECT 628.950 760.950 631.050 763.050 ;
        RECT 632.400 760.050 633.600 775.950 ;
        RECT 635.400 766.050 636.600 785.400 ;
        RECT 649.950 784.950 652.050 787.050 ;
        RECT 650.400 781.050 651.600 784.950 ;
        RECT 643.950 778.950 646.050 781.050 ;
        RECT 649.950 778.950 652.050 781.050 ;
        RECT 637.950 775.950 640.050 778.050 ;
        RECT 634.950 763.950 637.050 766.050 ;
        RECT 638.400 760.050 639.600 775.950 ;
        RECT 644.400 760.050 645.600 778.950 ;
        RECT 653.400 762.600 654.600 793.950 ;
        RECT 670.950 787.950 673.050 790.050 ;
        RECT 655.950 781.950 658.050 784.050 ;
        RECT 667.950 781.950 670.050 784.050 ;
        RECT 650.400 761.400 654.600 762.600 ;
        RECT 631.950 757.950 634.050 760.050 ;
        RECT 634.950 757.950 637.050 760.050 ;
        RECT 637.950 757.950 640.050 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 643.950 757.950 646.050 760.050 ;
        RECT 628.950 754.950 631.050 757.050 ;
        RECT 635.400 756.900 636.600 757.950 ;
        RECT 629.400 745.050 630.600 754.950 ;
        RECT 634.950 754.800 637.050 756.900 ;
        RECT 631.950 748.950 634.050 751.050 ;
        RECT 628.950 742.950 631.050 745.050 ;
        RECT 628.950 736.950 631.050 739.050 ;
        RECT 625.950 733.950 628.050 736.050 ;
        RECT 629.400 733.050 630.600 736.950 ;
        RECT 628.950 730.950 631.050 733.050 ;
        RECT 599.400 727.050 600.600 728.100 ;
        RECT 605.400 727.050 606.600 729.000 ;
        RECT 610.950 728.100 613.050 730.200 ;
        RECT 619.950 728.100 622.050 730.200 ;
        RECT 627.000 729.900 630.000 730.050 ;
        RECT 627.000 729.600 631.050 729.900 ;
        RECT 595.950 724.950 598.050 727.050 ;
        RECT 598.950 724.950 601.050 727.050 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 604.950 724.950 607.050 727.050 ;
        RECT 596.400 723.900 597.600 724.950 ;
        RECT 602.400 723.900 603.600 724.950 ;
        RECT 611.400 724.050 612.600 728.100 ;
        RECT 620.400 727.050 621.600 728.100 ;
        RECT 626.400 727.950 631.050 729.600 ;
        RECT 626.400 727.050 627.600 727.950 ;
        RECT 628.950 727.800 631.050 727.950 ;
        RECT 632.400 727.050 633.600 748.950 ;
        RECT 641.400 748.050 642.600 757.950 ;
        RECT 646.950 754.950 649.050 757.050 ;
        RECT 640.950 745.950 643.050 748.050 ;
        RECT 647.400 745.050 648.600 754.950 ;
        RECT 634.950 742.950 637.050 745.050 ;
        RECT 646.950 742.950 649.050 745.050 ;
        RECT 616.950 724.950 619.050 727.050 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 622.950 724.950 625.050 727.050 ;
        RECT 625.950 724.950 628.050 727.050 ;
        RECT 631.950 724.950 634.050 727.050 ;
        RECT 595.950 721.800 598.050 723.900 ;
        RECT 601.950 721.800 604.050 723.900 ;
        RECT 610.950 721.950 613.050 724.050 ;
        RECT 617.400 723.000 618.600 724.950 ;
        RECT 623.400 723.900 624.600 724.950 ;
        RECT 592.950 712.950 595.050 715.050 ;
        RECT 589.950 706.950 592.050 709.050 ;
        RECT 593.400 705.600 594.600 712.950 ;
        RECT 590.400 704.400 594.600 705.600 ;
        RECT 586.950 700.950 589.050 703.050 ;
        RECT 581.400 686.400 585.600 687.600 ;
        RECT 571.950 683.100 574.050 685.200 ;
        RECT 556.950 622.950 559.050 625.050 ;
        RECT 568.950 622.950 571.050 625.050 ;
        RECT 553.950 604.950 556.050 607.050 ;
        RECT 557.400 604.050 558.600 622.950 ;
        RECT 572.400 619.050 573.600 683.100 ;
        RECT 581.400 682.050 582.600 686.400 ;
        RECT 577.950 679.950 580.050 682.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 574.950 676.950 577.050 679.050 ;
        RECT 575.400 652.050 576.600 676.950 ;
        RECT 578.400 673.050 579.600 679.950 ;
        RECT 577.950 670.950 580.050 673.050 ;
        RECT 590.400 670.050 591.600 704.400 ;
        RECT 598.950 703.950 601.050 706.050 ;
        RECT 599.400 700.050 600.600 703.950 ;
        RECT 598.950 697.950 601.050 700.050 ;
        RECT 602.400 685.200 603.600 721.800 ;
        RECT 616.950 718.950 619.050 723.000 ;
        RECT 622.950 721.800 625.050 723.900 ;
        RECT 628.950 721.950 631.050 724.050 ;
        RECT 625.950 718.950 628.050 721.050 ;
        RECT 610.950 715.950 613.050 718.050 ;
        RECT 607.950 706.950 610.050 709.050 ;
        RECT 601.950 683.100 604.050 685.200 ;
        RECT 602.400 682.050 603.600 683.100 ;
        RECT 595.950 679.950 598.050 682.050 ;
        RECT 601.950 679.950 604.050 682.050 ;
        RECT 596.400 678.600 597.600 679.950 ;
        RECT 593.400 677.400 597.600 678.600 ;
        RECT 589.950 667.950 592.050 670.050 ;
        RECT 593.400 661.050 594.600 677.400 ;
        RECT 598.950 673.950 601.050 676.050 ;
        RECT 595.950 661.950 598.050 664.050 ;
        RECT 592.950 658.950 595.050 661.050 ;
        RECT 583.950 656.400 586.050 658.500 ;
        RECT 574.950 649.950 577.050 652.050 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 578.400 646.050 579.600 646.950 ;
        RECT 574.950 643.950 577.050 646.050 ;
        RECT 578.400 644.400 583.050 646.050 ;
        RECT 579.000 643.950 583.050 644.400 ;
        RECT 571.950 616.950 574.050 619.050 ;
        RECT 575.400 615.600 576.600 643.950 ;
        RECT 584.100 636.600 585.300 656.400 ;
        RECT 592.950 652.950 595.050 655.050 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 587.400 640.050 588.600 646.950 ;
        RECT 586.950 637.950 589.050 640.050 ;
        RECT 583.950 634.500 586.050 636.600 ;
        RECT 572.400 614.400 576.600 615.600 ;
        RECT 562.950 610.950 565.050 613.050 ;
        RECT 563.400 604.050 564.600 610.950 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 560.400 600.900 561.600 601.950 ;
        RECT 559.950 598.800 562.050 600.900 ;
        RECT 550.950 583.950 553.050 586.050 ;
        RECT 547.950 574.950 550.050 577.050 ;
        RECT 559.950 574.950 562.050 577.050 ;
        RECT 550.950 572.100 553.050 574.200 ;
        RECT 551.400 571.050 552.600 572.100 ;
        RECT 547.950 568.950 550.050 571.050 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 553.950 568.950 556.050 571.050 ;
        RECT 548.400 567.000 549.600 568.950 ;
        RECT 547.950 562.950 550.050 567.000 ;
        RECT 499.950 541.950 502.050 544.050 ;
        RECT 529.950 541.950 532.050 544.050 ;
        RECT 541.950 541.950 544.050 544.050 ;
        RECT 500.400 529.200 501.600 541.950 ;
        RECT 548.400 541.050 549.600 562.950 ;
        RECT 554.400 556.050 555.600 568.950 ;
        RECT 553.950 553.950 556.050 556.050 ;
        RECT 547.950 538.950 550.050 541.050 ;
        RECT 535.950 532.950 538.050 535.050 ;
        RECT 499.950 527.100 502.050 529.200 ;
        RECT 514.950 527.100 517.050 529.200 ;
        RECT 523.950 527.100 526.050 529.200 ;
        RECT 529.950 527.100 532.050 529.200 ;
        RECT 500.400 526.050 501.600 527.100 ;
        RECT 496.950 523.950 499.050 526.050 ;
        RECT 499.950 523.950 502.050 526.050 ;
        RECT 502.950 523.950 505.050 526.050 ;
        RECT 493.950 520.950 496.050 523.050 ;
        RECT 497.400 522.000 498.600 523.950 ;
        RECT 490.950 517.950 493.050 520.050 ;
        RECT 487.950 511.950 490.050 514.050 ;
        RECT 478.950 508.950 481.050 511.050 ;
        RECT 494.400 508.050 495.600 520.950 ;
        RECT 496.950 517.950 499.050 522.000 ;
        RECT 487.950 505.950 490.050 508.050 ;
        RECT 493.950 505.950 496.050 508.050 ;
        RECT 481.950 499.950 484.050 502.050 ;
        RECT 478.950 496.950 481.050 499.050 ;
        RECT 469.950 463.950 472.050 466.050 ;
        RECT 475.950 463.950 478.050 466.050 ;
        RECT 479.400 457.050 480.600 496.950 ;
        RECT 482.400 489.900 483.600 499.950 ;
        RECT 488.400 493.050 489.600 505.950 ;
        RECT 493.950 494.100 496.050 496.200 ;
        RECT 494.400 493.050 495.600 494.100 ;
        RECT 487.950 490.950 490.050 493.050 ;
        RECT 490.950 490.950 493.050 493.050 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 491.400 489.900 492.600 490.950 ;
        RECT 481.950 487.800 484.050 489.900 ;
        RECT 490.950 487.800 493.050 489.900 ;
        RECT 484.950 484.950 487.050 487.050 ;
        RECT 493.950 484.950 496.050 487.050 ;
        RECT 485.400 460.050 486.600 484.950 ;
        RECT 490.950 478.950 493.050 481.050 ;
        RECT 487.950 475.950 490.050 478.050 ;
        RECT 488.400 469.050 489.600 475.950 ;
        RECT 487.950 466.950 490.050 469.050 ;
        RECT 484.950 457.950 487.050 460.050 ;
        RECT 475.800 454.950 477.900 457.050 ;
        RECT 478.950 454.950 481.050 457.050 ;
        RECT 457.950 448.950 460.050 451.050 ;
        RECT 463.950 449.100 466.050 454.050 ;
        RECT 472.950 449.100 475.050 451.200 ;
        RECT 476.400 451.050 477.600 454.950 ;
        RECT 464.400 448.050 465.600 449.100 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 463.950 445.950 466.050 448.050 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 454.950 444.600 457.050 445.050 ;
        RECT 461.400 444.900 462.600 445.950 ;
        RECT 454.950 443.400 459.600 444.600 ;
        RECT 454.950 442.950 457.050 443.400 ;
        RECT 454.950 439.800 457.050 441.900 ;
        RECT 451.950 436.950 454.050 439.050 ;
        RECT 442.950 430.950 445.050 433.050 ;
        RECT 430.950 427.950 433.050 430.050 ;
        RECT 433.950 421.950 436.050 424.050 ;
        RECT 445.950 421.950 448.050 424.050 ;
        RECT 418.950 415.950 421.050 418.050 ;
        RECT 424.950 416.100 427.050 418.200 ;
        RECT 425.400 415.050 426.600 416.100 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 415.950 409.800 418.050 411.900 ;
        RECT 410.400 408.000 415.050 408.600 ;
        RECT 410.400 407.400 414.600 408.000 ;
        RECT 397.950 405.000 402.600 405.600 ;
        RECT 398.400 404.400 402.600 405.000 ;
        RECT 385.950 397.950 388.050 400.050 ;
        RECT 388.950 394.950 391.050 397.050 ;
        RECT 382.950 391.950 385.050 394.050 ;
        RECT 376.950 379.950 379.050 382.050 ;
        RECT 376.950 376.800 379.050 378.900 ;
        RECT 370.950 370.950 373.050 373.050 ;
        RECT 377.400 370.050 378.600 376.800 ;
        RECT 383.400 370.050 384.600 391.950 ;
        RECT 373.950 367.950 376.050 370.050 ;
        RECT 376.950 367.950 379.050 370.050 ;
        RECT 379.950 367.950 382.050 370.050 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 370.950 364.950 373.050 367.050 ;
        RECT 371.400 349.050 372.600 364.950 ;
        RECT 374.400 358.050 375.600 367.950 ;
        RECT 380.400 366.900 381.600 367.950 ;
        RECT 379.950 364.800 382.050 366.900 ;
        RECT 373.950 355.950 376.050 358.050 ;
        RECT 389.400 355.050 390.600 394.950 ;
        RECT 392.400 373.200 393.600 404.400 ;
        RECT 394.950 400.950 397.050 403.050 ;
        RECT 395.400 376.050 396.600 400.950 ;
        RECT 401.400 396.600 402.600 404.400 ;
        RECT 410.400 402.600 411.600 407.400 ;
        RECT 412.950 403.950 415.050 406.050 ;
        RECT 407.400 401.400 411.600 402.600 ;
        RECT 407.400 400.050 408.600 401.400 ;
        RECT 403.950 398.400 408.600 400.050 ;
        RECT 403.950 397.950 408.000 398.400 ;
        RECT 406.950 396.600 409.050 397.050 ;
        RECT 401.400 395.400 409.050 396.600 ;
        RECT 406.950 394.950 409.050 395.400 ;
        RECT 403.950 391.950 406.050 394.050 ;
        RECT 404.400 388.050 405.600 391.950 ;
        RECT 413.400 390.600 414.600 403.950 ;
        RECT 410.400 389.400 414.600 390.600 ;
        RECT 403.950 385.950 406.050 388.050 ;
        RECT 400.950 382.950 403.050 385.050 ;
        RECT 401.400 376.050 402.600 382.950 ;
        RECT 406.950 376.950 409.050 379.050 ;
        RECT 394.950 373.950 397.050 376.050 ;
        RECT 401.400 374.400 406.050 376.050 ;
        RECT 402.000 373.950 406.050 374.400 ;
        RECT 391.950 371.100 394.050 373.200 ;
        RECT 395.400 370.050 396.600 373.950 ;
        RECT 400.950 371.100 403.050 373.200 ;
        RECT 407.400 373.050 408.600 376.950 ;
        RECT 401.400 370.050 402.600 371.100 ;
        RECT 406.950 370.950 409.050 373.050 ;
        RECT 394.950 367.950 397.050 370.050 ;
        RECT 397.950 367.950 400.050 370.050 ;
        RECT 400.950 367.950 403.050 370.050 ;
        RECT 403.950 367.950 406.050 370.050 ;
        RECT 398.400 355.050 399.600 367.950 ;
        RECT 404.400 367.050 405.600 367.950 ;
        RECT 404.400 364.950 409.050 367.050 ;
        RECT 373.950 352.800 376.050 354.900 ;
        RECT 388.950 352.950 391.050 355.050 ;
        RECT 397.950 352.950 400.050 355.050 ;
        RECT 370.950 346.950 373.050 349.050 ;
        RECT 367.950 340.950 370.050 343.050 ;
        RECT 374.400 337.050 375.600 352.800 ;
        RECT 400.950 349.950 403.050 352.050 ;
        RECT 388.950 346.950 391.050 349.050 ;
        RECT 364.950 334.950 367.050 337.050 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 379.950 334.950 382.050 337.050 ;
        RECT 364.950 331.800 367.050 333.900 ;
        RECT 361.950 322.950 364.050 325.050 ;
        RECT 365.400 322.050 366.600 331.800 ;
        RECT 364.950 319.950 367.050 322.050 ;
        RECT 371.400 319.050 372.600 334.950 ;
        RECT 361.950 316.950 364.050 319.050 ;
        RECT 370.950 316.950 373.050 319.050 ;
        RECT 358.950 298.950 361.050 301.050 ;
        RECT 362.400 292.050 363.600 316.950 ;
        RECT 380.400 313.050 381.600 334.950 ;
        RECT 382.950 328.950 385.050 331.050 ;
        RECT 383.400 316.050 384.600 328.950 ;
        RECT 382.950 313.950 385.050 316.050 ;
        RECT 379.950 312.600 382.050 313.050 ;
        RECT 379.950 311.400 384.600 312.600 ;
        RECT 379.950 310.950 382.050 311.400 ;
        RECT 367.950 301.950 370.050 304.050 ;
        RECT 364.950 295.950 367.050 301.050 ;
        RECT 368.400 292.050 369.600 301.950 ;
        RECT 370.950 298.950 373.050 301.050 ;
        RECT 376.950 298.950 382.050 301.050 ;
        RECT 371.400 295.050 372.600 298.950 ;
        RECT 370.800 292.950 372.900 295.050 ;
        RECT 376.950 294.600 379.050 297.900 ;
        RECT 383.400 297.600 384.600 311.400 ;
        RECT 389.400 298.050 390.600 346.950 ;
        RECT 401.400 337.050 402.600 349.950 ;
        RECT 404.400 340.050 405.600 364.950 ;
        RECT 406.950 358.950 409.050 363.900 ;
        RECT 406.950 343.950 409.050 346.050 ;
        RECT 403.950 337.950 406.050 340.050 ;
        RECT 407.400 337.050 408.600 343.950 ;
        RECT 400.950 334.950 403.050 337.050 ;
        RECT 406.950 334.950 409.050 337.050 ;
        RECT 406.950 331.800 409.050 333.900 ;
        RECT 394.950 325.950 397.050 328.050 ;
        RECT 407.400 327.600 408.600 331.800 ;
        RECT 410.400 331.050 411.600 389.400 ;
        RECT 412.950 373.950 415.050 376.050 ;
        RECT 413.400 366.750 414.600 373.950 ;
        RECT 416.400 373.050 417.600 409.800 ;
        RECT 422.400 406.050 423.600 412.950 ;
        RECT 428.400 411.900 429.600 412.950 ;
        RECT 434.400 412.050 435.600 421.950 ;
        RECT 436.950 415.950 439.050 418.050 ;
        RECT 427.950 409.800 430.050 411.900 ;
        RECT 433.950 409.950 436.050 412.050 ;
        RECT 421.950 403.950 424.050 406.050 ;
        RECT 418.950 397.950 421.050 400.050 ;
        RECT 419.400 388.050 420.600 397.950 ;
        RECT 428.400 391.050 429.600 409.800 ;
        RECT 437.400 408.600 438.600 415.950 ;
        RECT 446.400 415.050 447.600 421.950 ;
        RECT 451.950 416.100 454.050 418.200 ;
        RECT 455.400 418.050 456.600 439.800 ;
        RECT 452.400 415.050 453.600 416.100 ;
        RECT 454.950 415.950 457.050 418.050 ;
        RECT 442.950 412.950 445.050 415.050 ;
        RECT 445.950 412.950 448.050 415.050 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 434.400 407.400 438.600 408.600 ;
        RECT 434.400 400.050 435.600 407.400 ;
        RECT 443.400 406.050 444.600 412.950 ;
        RECT 449.400 411.900 450.600 412.950 ;
        RECT 448.950 409.800 451.050 411.900 ;
        RECT 454.950 409.950 457.050 412.050 ;
        RECT 436.950 403.950 439.050 406.050 ;
        RECT 442.950 403.950 445.050 406.050 ;
        RECT 433.950 397.950 436.050 400.050 ;
        RECT 427.950 388.950 430.050 391.050 ;
        RECT 418.950 385.950 421.050 388.050 ;
        RECT 427.950 382.950 430.050 385.050 ;
        RECT 424.950 376.950 427.050 379.050 ;
        RECT 415.950 370.950 418.050 373.050 ;
        RECT 425.400 369.900 426.600 376.950 ;
        RECT 428.400 376.050 429.600 382.950 ;
        RECT 427.950 373.950 430.050 376.050 ;
        RECT 437.400 373.050 438.600 403.950 ;
        RECT 443.400 400.050 444.600 403.950 ;
        RECT 445.950 400.950 448.050 403.050 ;
        RECT 442.950 397.950 445.050 400.050 ;
        RECT 439.950 385.950 442.050 388.050 ;
        RECT 433.950 370.950 436.050 373.050 ;
        RECT 436.950 370.950 439.050 373.050 ;
        RECT 434.400 369.900 435.600 370.950 ;
        RECT 440.400 370.050 441.600 385.950 ;
        RECT 446.400 375.600 447.600 400.950 ;
        RECT 455.400 376.050 456.600 409.950 ;
        RECT 458.400 388.050 459.600 443.400 ;
        RECT 460.950 442.800 463.050 444.900 ;
        RECT 467.400 439.050 468.600 445.950 ;
        RECT 473.400 442.050 474.600 449.100 ;
        RECT 475.950 448.950 478.050 451.050 ;
        RECT 478.950 449.100 481.050 451.200 ;
        RECT 484.950 449.100 487.050 451.200 ;
        RECT 491.400 451.050 492.600 478.950 ;
        RECT 479.400 448.050 480.600 449.100 ;
        RECT 485.400 448.050 486.600 449.100 ;
        RECT 490.950 448.950 493.050 451.050 ;
        RECT 478.950 445.950 481.050 448.050 ;
        RECT 481.950 445.950 484.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 475.950 442.950 478.050 445.050 ;
        RECT 482.400 444.900 483.600 445.950 ;
        RECT 488.400 444.900 489.600 445.950 ;
        RECT 494.400 445.050 495.600 484.950 ;
        RECT 497.400 475.050 498.600 490.950 ;
        RECT 496.950 472.950 499.050 475.050 ;
        RECT 503.400 454.050 504.600 523.950 ;
        RECT 508.950 520.950 511.050 523.050 ;
        RECT 515.400 522.600 516.600 527.100 ;
        RECT 524.400 526.050 525.600 527.100 ;
        RECT 530.400 526.050 531.600 527.100 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 523.950 523.950 526.050 526.050 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 529.950 523.950 532.050 526.050 ;
        RECT 521.400 522.900 522.600 523.950 ;
        RECT 515.400 521.400 519.600 522.600 ;
        RECT 509.400 502.050 510.600 520.950 ;
        RECT 514.950 511.950 517.050 514.050 ;
        RECT 508.950 499.950 511.050 502.050 ;
        RECT 515.400 499.050 516.600 511.950 ;
        RECT 514.950 496.950 517.050 499.050 ;
        RECT 511.950 494.100 514.050 496.200 ;
        RECT 512.400 493.050 513.600 494.100 ;
        RECT 518.400 493.050 519.600 521.400 ;
        RECT 520.950 520.800 523.050 522.900 ;
        RECT 520.950 508.950 523.050 511.050 ;
        RECT 521.400 496.050 522.600 508.950 ;
        RECT 523.950 496.950 526.050 499.050 ;
        RECT 520.950 493.950 523.050 496.050 ;
        RECT 508.950 490.950 511.050 493.050 ;
        RECT 511.950 490.950 514.050 493.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 509.400 475.050 510.600 490.950 ;
        RECT 515.400 489.900 516.600 490.950 ;
        RECT 524.400 489.900 525.600 496.950 ;
        RECT 514.950 487.800 517.050 489.900 ;
        RECT 523.950 487.800 526.050 489.900 ;
        RECT 527.400 484.050 528.600 523.950 ;
        RECT 536.400 522.900 537.600 532.950 ;
        RECT 560.400 532.050 561.600 574.950 ;
        RECT 572.400 574.050 573.600 614.400 ;
        RECT 586.950 610.950 589.050 613.050 ;
        RECT 574.950 605.100 577.050 607.200 ;
        RECT 580.950 605.100 583.050 607.200 ;
        RECT 575.400 601.050 576.600 605.100 ;
        RECT 581.400 604.050 582.600 605.100 ;
        RECT 587.400 604.050 588.600 610.950 ;
        RECT 593.400 607.050 594.600 652.950 ;
        RECT 596.400 640.050 597.600 661.950 ;
        RECT 599.400 645.900 600.600 673.950 ;
        RECT 608.400 664.050 609.600 706.950 ;
        RECT 607.950 661.950 610.050 664.050 ;
        RECT 611.400 655.050 612.600 715.950 ;
        RECT 622.950 691.950 625.050 694.050 ;
        RECT 616.950 683.100 619.050 685.200 ;
        RECT 617.400 682.050 618.600 683.100 ;
        RECT 623.400 682.050 624.600 691.950 ;
        RECT 626.400 685.050 627.600 718.950 ;
        RECT 629.400 709.050 630.600 721.950 ;
        RECT 628.950 706.950 631.050 709.050 ;
        RECT 632.400 706.050 633.600 724.950 ;
        RECT 635.400 712.050 636.600 742.950 ;
        RECT 643.950 739.950 646.050 742.050 ;
        RECT 644.400 727.050 645.600 739.950 ;
        RECT 650.400 730.050 651.600 761.400 ;
        RECT 656.400 760.050 657.600 781.950 ;
        RECT 661.950 762.000 664.050 766.050 ;
        RECT 662.400 760.050 663.600 762.000 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 652.950 754.950 655.050 757.050 ;
        RECT 649.950 727.950 652.050 730.050 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 646.950 724.950 649.050 727.050 ;
        RECT 641.400 712.050 642.600 724.950 ;
        RECT 647.400 723.900 648.600 724.950 ;
        RECT 646.950 721.800 649.050 723.900 ;
        RECT 649.950 721.950 652.050 724.050 ;
        RECT 650.400 718.050 651.600 721.950 ;
        RECT 649.950 715.950 652.050 718.050 ;
        RECT 634.950 709.950 637.050 712.050 ;
        RECT 640.950 709.950 643.050 712.050 ;
        RECT 631.950 703.950 634.050 706.050 ;
        RECT 641.400 694.050 642.600 709.950 ;
        RECT 653.400 706.050 654.600 754.950 ;
        RECT 655.950 745.950 658.050 748.050 ;
        RECT 656.400 715.050 657.600 745.950 ;
        RECT 659.400 736.050 660.600 757.950 ;
        RECT 664.950 751.950 667.050 754.050 ;
        RECT 658.950 733.950 661.050 736.050 ;
        RECT 665.400 730.200 666.600 751.950 ;
        RECT 668.400 748.050 669.600 781.950 ;
        RECT 667.950 745.950 670.050 748.050 ;
        RECT 671.400 733.050 672.600 787.950 ;
        RECT 673.950 784.950 676.050 787.050 ;
        RECT 674.400 763.050 675.600 784.950 ;
        RECT 676.950 778.950 679.050 781.050 ;
        RECT 677.400 763.200 678.600 778.950 ;
        RECT 682.950 775.950 685.050 778.050 ;
        RECT 683.400 769.050 684.600 775.950 ;
        RECT 686.400 775.050 687.600 802.950 ;
        RECT 685.950 772.950 688.050 775.050 ;
        RECT 682.950 766.950 685.050 769.050 ;
        RECT 673.800 760.950 675.900 763.050 ;
        RECT 676.950 761.100 679.050 763.200 ;
        RECT 685.950 761.100 688.050 766.050 ;
        RECT 677.400 760.050 678.600 761.100 ;
        RECT 686.400 760.050 687.600 761.100 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 682.950 757.950 685.050 760.050 ;
        RECT 685.950 757.950 688.050 760.050 ;
        RECT 673.950 754.950 676.050 757.050 ;
        RECT 679.950 754.950 682.050 757.050 ;
        RECT 670.950 730.950 673.050 733.050 ;
        RECT 664.950 728.100 667.050 730.200 ;
        RECT 674.400 730.050 675.600 754.950 ;
        RECT 676.950 730.950 679.050 733.050 ;
        RECT 665.400 727.050 666.600 728.100 ;
        RECT 673.950 727.950 676.050 730.050 ;
        RECT 661.950 724.950 664.050 727.050 ;
        RECT 664.950 724.950 667.050 727.050 ;
        RECT 670.950 724.950 673.050 727.050 ;
        RECT 662.400 723.900 663.600 724.950 ;
        RECT 671.400 724.050 672.600 724.950 ;
        RECT 661.950 721.800 664.050 723.900 ;
        RECT 667.950 721.950 670.050 724.050 ;
        RECT 671.400 722.400 676.050 724.050 ;
        RECT 672.000 721.950 676.050 722.400 ;
        RECT 668.400 718.050 669.600 721.950 ;
        RECT 667.950 715.950 670.050 718.050 ;
        RECT 677.400 715.050 678.600 730.950 ;
        RECT 680.400 730.050 681.600 754.950 ;
        RECT 683.400 745.050 684.600 757.950 ;
        RECT 682.950 742.950 685.050 745.050 ;
        RECT 683.400 736.050 684.600 742.950 ;
        RECT 692.400 742.050 693.600 811.950 ;
        RECT 701.400 805.050 702.600 818.400 ;
        RECT 713.400 816.600 714.600 835.950 ;
        RECT 719.400 826.050 720.600 835.950 ;
        RECT 721.950 832.950 724.050 835.050 ;
        RECT 715.800 823.950 717.900 826.050 ;
        RECT 718.950 823.950 721.050 826.050 ;
        RECT 716.400 820.050 717.600 823.950 ;
        RECT 715.950 817.950 718.050 820.050 ;
        RECT 722.400 816.600 723.600 832.950 ;
        RECT 725.400 829.050 726.600 844.950 ;
        RECT 724.950 826.950 727.050 829.050 ;
        RECT 728.400 826.050 729.600 853.950 ;
        RECT 737.400 844.200 738.600 889.950 ;
        RECT 742.950 886.950 745.050 889.050 ;
        RECT 739.950 883.950 742.050 886.050 ;
        RECT 740.400 853.050 741.600 883.950 ;
        RECT 743.400 879.600 744.600 886.950 ;
        RECT 767.400 886.050 768.600 892.950 ;
        RECT 766.950 883.950 769.050 886.050 ;
        RECT 772.950 884.100 775.050 886.200 ;
        RECT 782.400 886.050 783.600 898.950 ;
        RECT 787.950 889.950 790.050 892.050 ;
        RECT 773.400 883.050 774.600 884.100 ;
        RECT 781.950 883.950 784.050 886.050 ;
        RECT 788.400 883.050 789.600 889.950 ;
        RECT 794.400 886.050 795.600 910.950 ;
        RECT 806.400 901.050 807.600 910.950 ;
        RECT 812.400 907.050 813.600 913.950 ;
        RECT 820.950 910.950 823.050 913.050 ;
        RECT 827.400 912.900 828.600 913.950 ;
        RECT 836.400 912.900 837.600 913.950 ;
        RECT 811.950 904.950 814.050 907.050 ;
        RECT 821.400 904.050 822.600 910.950 ;
        RECT 826.950 910.800 829.050 912.900 ;
        RECT 835.950 910.800 838.050 912.900 ;
        RECT 820.950 901.950 823.050 904.050 ;
        RECT 805.950 898.950 808.050 901.050 ;
        RECT 811.950 898.950 814.050 901.050 ;
        RECT 793.950 883.950 796.050 886.050 ;
        RECT 796.950 884.100 799.050 886.200 ;
        RECT 805.950 884.100 808.050 886.200 ;
        RECT 748.950 880.950 751.050 883.050 ;
        RECT 769.950 880.950 772.050 883.050 ;
        RECT 772.950 880.950 775.050 883.050 ;
        RECT 775.950 880.950 778.050 883.050 ;
        RECT 784.950 880.950 787.050 883.050 ;
        RECT 787.950 880.950 790.050 883.050 ;
        RECT 790.950 880.950 793.050 883.050 ;
        RECT 749.400 879.600 750.600 880.950 ;
        RECT 770.400 879.900 771.600 880.950 ;
        RECT 743.400 878.400 750.600 879.600 ;
        RECT 769.950 877.800 772.050 879.900 ;
        RECT 776.400 879.600 777.600 880.950 ;
        RECT 785.400 879.900 786.600 880.950 ;
        RECT 791.400 879.900 792.600 880.950 ;
        RECT 776.400 878.400 780.600 879.600 ;
        RECT 779.400 874.050 780.600 878.400 ;
        RECT 784.950 877.800 787.050 879.900 ;
        RECT 790.950 877.800 793.050 879.900 ;
        RECT 793.950 877.950 796.050 880.050 ;
        RECT 794.400 874.050 795.600 877.950 ;
        RECT 778.950 871.950 781.050 874.050 ;
        RECT 793.950 871.950 796.050 874.050 ;
        RECT 772.950 865.950 775.050 868.050 ;
        RECT 763.950 862.950 766.050 865.050 ;
        RECT 742.950 859.950 745.050 862.050 ;
        RECT 739.950 850.950 742.050 853.050 ;
        RECT 730.950 841.950 733.050 844.050 ;
        RECT 736.950 842.100 739.050 844.200 ;
        RECT 727.950 823.950 730.050 826.050 ;
        RECT 731.400 820.050 732.600 841.950 ;
        RECT 736.950 838.950 739.050 841.050 ;
        RECT 737.400 838.050 738.600 838.950 ;
        RECT 743.400 838.050 744.600 859.950 ;
        RECT 757.950 840.000 760.050 844.050 ;
        RECT 758.400 838.050 759.600 840.000 ;
        RECT 764.400 838.050 765.600 862.950 ;
        RECT 773.400 862.050 774.600 865.950 ;
        RECT 779.400 865.050 780.600 871.950 ;
        RECT 778.950 862.950 781.050 865.050 ;
        RECT 772.950 859.950 775.050 862.050 ;
        RECT 784.950 856.950 787.050 859.050 ;
        RECT 769.950 853.950 772.050 856.050 ;
        RECT 770.400 838.050 771.600 853.950 ;
        RECT 772.950 847.950 775.050 850.050 ;
        RECT 773.400 841.050 774.600 847.950 ;
        RECT 785.400 844.050 786.600 856.950 ;
        RECT 797.400 856.050 798.600 884.100 ;
        RECT 806.400 883.050 807.600 884.100 ;
        RECT 812.400 883.050 813.600 898.950 ;
        RECT 829.950 892.950 832.050 895.050 ;
        RECT 823.950 889.950 826.050 892.050 ;
        RECT 820.950 884.100 823.050 886.200 ;
        RECT 805.950 880.950 808.050 883.050 ;
        RECT 808.950 880.950 811.050 883.050 ;
        RECT 811.950 880.950 814.050 883.050 ;
        RECT 814.950 880.950 817.050 883.050 ;
        RECT 809.400 879.900 810.600 880.950 ;
        RECT 808.950 877.800 811.050 879.900 ;
        RECT 815.400 879.000 816.600 880.950 ;
        RECT 814.950 874.950 817.050 879.000 ;
        RECT 821.400 874.050 822.600 884.100 ;
        RECT 820.950 871.950 823.050 874.050 ;
        RECT 817.950 865.950 820.050 868.050 ;
        RECT 818.400 856.050 819.600 865.950 ;
        RECT 821.400 859.050 822.600 871.950 ;
        RECT 820.950 856.950 823.050 859.050 ;
        RECT 787.950 853.950 790.050 856.050 ;
        RECT 796.950 853.950 799.050 856.050 ;
        RECT 817.950 853.950 820.050 856.050 ;
        RECT 784.950 841.950 787.050 844.050 ;
        RECT 772.950 838.950 775.050 841.050 ;
        RECT 788.400 838.050 789.600 853.950 ;
        RECT 790.950 847.950 793.050 850.050 ;
        RECT 791.400 841.050 792.600 847.950 ;
        RECT 790.950 838.950 793.050 841.050 ;
        RECT 797.400 838.050 798.600 853.950 ;
        RECT 808.500 844.500 810.600 846.600 ;
        RECT 736.950 835.950 739.050 838.050 ;
        RECT 739.950 835.950 742.050 838.050 ;
        RECT 742.950 835.950 745.050 838.050 ;
        RECT 745.950 835.950 748.050 838.050 ;
        RECT 757.950 835.950 760.050 838.050 ;
        RECT 760.950 835.950 763.050 838.050 ;
        RECT 763.950 835.950 766.050 838.050 ;
        RECT 766.950 835.950 769.050 838.050 ;
        RECT 769.950 835.950 772.050 838.050 ;
        RECT 784.950 835.950 787.050 838.050 ;
        RECT 787.950 835.950 790.050 838.050 ;
        RECT 796.950 835.950 799.050 838.050 ;
        RECT 805.950 835.950 808.050 838.050 ;
        RECT 808.950 837.300 810.000 844.500 ;
        RECT 812.400 840.900 813.600 843.450 ;
        RECT 818.100 843.300 820.200 845.400 ;
        RECT 811.800 838.800 813.900 840.900 ;
        RECT 814.800 839.700 816.900 841.800 ;
        RECT 814.800 837.300 815.700 839.700 ;
        RECT 808.950 836.100 815.700 837.300 ;
        RECT 733.950 832.950 736.050 835.050 ;
        RECT 740.400 834.900 741.600 835.950 ;
        RECT 727.800 817.950 729.900 820.050 ;
        RECT 730.950 817.950 733.050 820.050 ;
        RECT 713.400 815.400 723.600 816.600 ;
        RECT 728.400 814.050 729.600 817.950 ;
        RECT 712.950 811.950 715.050 814.050 ;
        RECT 724.800 811.950 726.900 814.050 ;
        RECT 727.950 811.950 730.050 814.050 ;
        RECT 697.950 802.950 700.050 805.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 698.400 801.900 699.600 802.950 ;
        RECT 697.950 799.800 700.050 801.900 ;
        RECT 704.400 801.000 705.600 802.950 ;
        RECT 703.950 796.950 706.050 801.000 ;
        RECT 713.400 799.050 714.600 811.950 ;
        RECT 718.950 806.100 721.050 808.200 ;
        RECT 719.400 805.050 720.600 806.100 ;
        RECT 725.400 805.050 726.600 811.950 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 721.950 802.950 724.050 805.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 706.950 796.950 709.050 799.050 ;
        RECT 712.950 796.950 715.050 799.050 ;
        RECT 715.950 796.950 721.050 799.050 ;
        RECT 694.950 772.950 697.050 775.050 ;
        RECT 695.400 754.050 696.600 772.950 ;
        RECT 707.400 765.600 708.600 796.950 ;
        RECT 715.950 775.950 718.050 778.050 ;
        RECT 707.400 764.400 711.600 765.600 ;
        RECT 703.950 761.100 706.050 763.200 ;
        RECT 710.400 763.050 711.600 764.400 ;
        RECT 704.400 760.050 705.600 761.100 ;
        RECT 710.400 760.950 715.050 763.050 ;
        RECT 710.400 760.050 711.600 760.950 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 694.950 751.950 697.050 754.050 ;
        RECT 701.400 748.050 702.600 757.950 ;
        RECT 707.400 756.900 708.600 757.950 ;
        RECT 706.950 754.800 709.050 756.900 ;
        RECT 716.400 754.050 717.600 775.950 ;
        RECT 722.400 766.050 723.600 802.950 ;
        RECT 734.400 790.050 735.600 832.950 ;
        RECT 739.950 832.800 742.050 834.900 ;
        RECT 736.950 820.950 739.050 823.050 ;
        RECT 733.950 787.950 736.050 790.050 ;
        RECT 737.400 781.050 738.600 820.950 ;
        RECT 746.400 819.600 747.600 835.950 ;
        RECT 761.400 834.900 762.600 835.950 ;
        RECT 767.400 834.900 768.600 835.950 ;
        RECT 760.950 832.800 763.050 834.900 ;
        RECT 766.950 832.800 769.050 834.900 ;
        RECT 781.950 834.600 784.050 834.900 ;
        RECT 785.400 834.600 786.600 835.950 ;
        RECT 781.950 833.400 786.600 834.600 ;
        RECT 806.400 833.400 807.600 835.950 ;
        RECT 781.950 832.800 784.050 833.400 ;
        RECT 754.950 826.950 757.050 829.050 ;
        RECT 746.400 818.400 750.600 819.600 ;
        RECT 749.400 808.050 750.600 818.400 ;
        RECT 751.950 810.600 754.050 814.050 ;
        RECT 755.400 810.600 756.600 826.950 ;
        RECT 778.950 826.800 781.050 828.900 ;
        RECT 779.400 823.050 780.600 826.800 ;
        RECT 778.950 820.950 781.050 823.050 ;
        RECT 760.950 817.950 763.050 820.050 ;
        RECT 751.950 810.000 756.600 810.600 ;
        RECT 752.400 809.400 756.600 810.000 ;
        RECT 748.950 805.950 751.050 808.050 ;
        RECT 752.400 805.050 753.600 809.400 ;
        RECT 745.950 802.950 748.050 805.050 ;
        RECT 751.950 802.950 754.050 805.050 ;
        RECT 746.400 801.000 747.600 802.950 ;
        RECT 745.950 796.950 748.050 801.000 ;
        RECT 748.950 799.950 751.050 802.050 ;
        RECT 736.950 778.950 739.050 781.050 ;
        RECT 749.400 775.050 750.600 799.950 ;
        RECT 761.400 793.050 762.600 817.950 ;
        RECT 782.400 808.050 783.600 832.800 ;
        RECT 808.950 830.700 809.850 836.100 ;
        RECT 810.750 834.300 812.850 835.200 ;
        RECT 818.400 834.300 819.300 843.300 ;
        RECT 821.400 838.050 822.600 840.600 ;
        RECT 824.400 838.050 825.600 889.950 ;
        RECT 830.400 886.200 831.600 892.950 ;
        RECT 829.950 884.100 832.050 886.200 ;
        RECT 835.950 884.100 838.050 886.200 ;
        RECT 830.400 883.050 831.600 884.100 ;
        RECT 836.400 883.050 837.600 884.100 ;
        RECT 829.950 880.950 832.050 883.050 ;
        RECT 832.950 880.950 835.050 883.050 ;
        RECT 835.950 880.950 838.050 883.050 ;
        RECT 833.400 879.900 834.600 880.950 ;
        RECT 832.950 877.800 835.050 879.900 ;
        RECT 826.950 874.950 829.050 877.050 ;
        RECT 827.400 865.050 828.600 874.950 ;
        RECT 826.950 862.950 829.050 865.050 ;
        RECT 829.950 853.950 832.050 856.050 ;
        RECT 842.400 855.600 843.600 925.950 ;
        RECT 848.400 907.050 849.600 934.950 ;
        RECT 874.950 925.950 877.050 928.050 ;
        RECT 853.950 918.000 856.050 922.050 ;
        RECT 854.400 916.050 855.600 918.000 ;
        RECT 859.950 917.100 862.050 919.200 ;
        RECT 860.400 916.050 861.600 917.100 ;
        RECT 875.400 916.050 876.600 925.950 ;
        RECT 853.950 913.950 856.050 916.050 ;
        RECT 856.950 913.950 859.050 916.050 ;
        RECT 859.950 913.950 862.050 916.050 ;
        RECT 862.950 913.950 865.050 916.050 ;
        RECT 868.950 913.950 871.050 916.050 ;
        RECT 874.950 913.950 877.050 916.050 ;
        RECT 877.950 913.950 880.050 916.050 ;
        RECT 895.950 913.950 898.050 916.050 ;
        RECT 857.400 912.900 858.600 913.950 ;
        RECT 856.950 910.800 859.050 912.900 ;
        RECT 863.400 912.000 864.600 913.950 ;
        RECT 862.950 907.950 865.050 912.000 ;
        RECT 847.950 904.950 850.050 907.050 ;
        RECT 859.950 904.950 862.050 907.050 ;
        RECT 860.400 898.050 861.600 904.950 ;
        RECT 869.400 901.050 870.600 913.950 ;
        RECT 862.950 898.950 865.050 901.050 ;
        RECT 868.950 898.950 871.050 901.050 ;
        RECT 859.950 895.950 862.050 898.050 ;
        RECT 847.950 892.950 850.050 895.050 ;
        RECT 848.400 883.050 849.600 892.950 ;
        RECT 853.950 889.950 856.050 892.050 ;
        RECT 854.400 883.050 855.600 889.950 ;
        RECT 847.950 880.950 850.050 883.050 ;
        RECT 850.950 880.950 853.050 883.050 ;
        RECT 853.950 880.950 856.050 883.050 ;
        RECT 856.950 880.950 859.050 883.050 ;
        RECT 851.400 879.900 852.600 880.950 ;
        RECT 857.400 879.900 858.600 880.950 ;
        RECT 850.950 877.800 853.050 879.900 ;
        RECT 856.950 877.800 859.050 879.900 ;
        RECT 851.400 871.050 852.600 877.800 ;
        RECT 850.950 868.950 853.050 871.050 ;
        RECT 842.400 854.400 846.600 855.600 ;
        RECT 826.950 838.950 829.050 841.050 ;
        RECT 820.500 835.950 822.600 838.050 ;
        RECT 823.950 835.950 826.050 838.050 ;
        RECT 810.750 833.100 819.300 834.300 ;
        RECT 808.500 828.600 810.600 830.700 ;
        RECT 811.800 830.100 813.900 832.200 ;
        RECT 815.700 831.300 817.800 833.100 ;
        RECT 823.950 832.800 826.050 834.900 ;
        RECT 812.400 828.000 813.600 830.100 ;
        RECT 796.950 823.950 799.050 826.050 ;
        RECT 811.950 823.950 814.050 828.000 ;
        RECT 814.950 826.950 817.050 829.050 ;
        RECT 781.950 805.950 784.050 808.050 ;
        RECT 790.950 807.000 793.050 811.050 ;
        RECT 791.400 805.050 792.600 807.000 ;
        RECT 766.950 802.950 769.050 805.050 ;
        RECT 787.950 802.950 790.050 805.050 ;
        RECT 790.950 802.950 793.050 805.050 ;
        RECT 760.950 790.950 763.050 793.050 ;
        RECT 757.950 781.950 760.050 784.050 ;
        RECT 739.950 772.950 742.050 775.050 ;
        RECT 748.950 772.950 751.050 775.050 ;
        RECT 724.950 766.950 727.050 769.050 ;
        RECT 721.950 763.950 724.050 766.050 ;
        RECT 725.400 760.050 726.600 766.950 ;
        RECT 736.950 763.950 739.050 766.050 ;
        RECT 730.950 761.100 733.050 763.200 ;
        RECT 731.400 760.050 732.600 761.100 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 724.950 757.950 727.050 760.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 718.950 754.950 721.050 757.050 ;
        RECT 722.400 756.900 723.600 757.950 ;
        RECT 709.950 750.600 712.050 754.050 ;
        RECT 715.950 751.950 718.050 754.050 ;
        RECT 707.400 750.000 712.050 750.600 ;
        RECT 707.400 749.400 711.600 750.000 ;
        RECT 700.950 745.950 703.050 748.050 ;
        RECT 707.400 747.600 708.600 749.400 ;
        RECT 704.400 746.400 708.600 747.600 ;
        RECT 691.950 739.950 694.050 742.050 ;
        RECT 694.950 736.950 697.050 739.050 ;
        RECT 682.950 733.950 685.050 736.050 ;
        RECT 695.400 733.050 696.600 736.950 ;
        RECT 697.950 733.950 700.050 736.050 ;
        RECT 694.950 730.950 697.050 733.050 ;
        RECT 679.950 727.950 682.050 730.050 ;
        RECT 682.950 728.100 685.050 730.200 ;
        RECT 688.950 728.100 691.050 730.200 ;
        RECT 683.400 727.050 684.600 728.100 ;
        RECT 689.400 727.050 690.600 728.100 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 685.950 724.950 688.050 727.050 ;
        RECT 688.950 724.950 691.050 727.050 ;
        RECT 691.950 724.950 694.050 727.050 ;
        RECT 679.950 721.950 682.050 724.050 ;
        RECT 680.400 715.050 681.600 721.950 ;
        RECT 682.950 718.950 685.050 721.050 ;
        RECT 655.950 712.950 658.050 715.050 ;
        RECT 661.950 712.950 664.050 715.050 ;
        RECT 670.950 712.950 673.050 715.050 ;
        RECT 676.950 712.950 679.050 715.050 ;
        RECT 679.950 712.950 682.050 715.050 ;
        RECT 652.950 703.950 655.050 706.050 ;
        RECT 649.950 700.950 652.050 703.050 ;
        RECT 650.400 697.050 651.600 700.950 ;
        RECT 649.950 694.950 652.050 697.050 ;
        RECT 640.950 691.950 643.050 694.050 ;
        RECT 625.950 682.950 628.050 685.050 ;
        RECT 637.950 683.100 640.050 685.200 ;
        RECT 643.950 683.100 646.050 685.200 ;
        RECT 647.400 683.400 654.600 684.600 ;
        RECT 638.400 682.050 639.600 683.100 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 619.950 679.950 622.050 682.050 ;
        RECT 622.950 679.950 625.050 682.050 ;
        RECT 637.950 679.950 640.050 682.050 ;
        RECT 620.400 678.000 621.600 679.950 ;
        RECT 619.950 676.050 622.050 678.000 ;
        RECT 619.800 675.000 622.050 676.050 ;
        RECT 619.800 673.950 621.900 675.000 ;
        RECT 622.950 673.950 625.050 676.050 ;
        RECT 610.950 652.950 613.050 655.050 ;
        RECT 607.950 650.100 610.050 652.200 ;
        RECT 613.950 650.100 616.050 652.200 ;
        RECT 608.400 649.050 609.600 650.100 ;
        RECT 614.400 649.050 615.600 650.100 ;
        RECT 623.400 649.050 624.600 673.950 ;
        RECT 644.400 673.050 645.600 683.100 ;
        RECT 647.400 673.050 648.600 683.400 ;
        RECT 653.400 682.050 654.600 683.400 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 631.950 670.950 634.050 673.050 ;
        RECT 643.800 670.950 645.900 673.050 ;
        RECT 646.950 670.950 649.050 673.050 ;
        RECT 604.950 646.950 607.050 649.050 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 610.950 646.950 613.050 649.050 ;
        RECT 613.950 646.950 616.050 649.050 ;
        RECT 622.950 646.950 625.050 649.050 ;
        RECT 625.950 646.950 628.050 649.050 ;
        RECT 605.400 645.900 606.600 646.950 ;
        RECT 598.950 643.800 601.050 645.900 ;
        RECT 604.950 643.800 607.050 645.900 ;
        RECT 595.950 637.950 598.050 640.050 ;
        RECT 601.950 622.950 604.050 625.050 ;
        RECT 602.400 613.050 603.600 622.950 ;
        RECT 611.400 619.050 612.600 646.950 ;
        RECT 619.950 643.950 622.050 646.050 ;
        RECT 613.950 637.950 616.050 640.050 ;
        RECT 610.950 616.950 613.050 619.050 ;
        RECT 595.950 610.950 598.050 613.050 ;
        RECT 601.950 610.950 604.050 613.050 ;
        RECT 592.950 604.950 595.050 607.050 ;
        RECT 580.950 601.950 583.050 604.050 ;
        RECT 583.950 601.950 586.050 604.050 ;
        RECT 586.950 601.950 589.050 604.050 ;
        RECT 589.950 601.950 592.050 604.050 ;
        RECT 574.950 598.950 577.050 601.050 ;
        RECT 577.950 595.950 580.050 598.050 ;
        RECT 574.950 589.950 577.050 592.050 ;
        RECT 562.800 571.950 564.900 574.050 ;
        RECT 571.950 571.950 574.050 574.050 ;
        RECT 563.400 562.050 564.600 571.950 ;
        RECT 575.400 571.050 576.600 589.950 ;
        RECT 578.400 574.050 579.600 595.950 ;
        RECT 584.400 589.050 585.600 601.950 ;
        RECT 590.400 589.050 591.600 601.950 ;
        RECT 583.950 586.950 586.050 589.050 ;
        RECT 589.950 586.950 592.050 589.050 ;
        RECT 580.950 577.950 583.050 580.050 ;
        RECT 577.950 571.950 580.050 574.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 569.400 567.900 570.600 568.950 ;
        RECT 568.950 565.800 571.050 567.900 ;
        RECT 577.950 565.950 580.050 568.050 ;
        RECT 569.400 564.600 570.600 565.800 ;
        RECT 566.400 563.400 570.600 564.600 ;
        RECT 562.950 559.950 565.050 562.050 ;
        RECT 553.950 529.950 556.050 532.050 ;
        RECT 559.950 529.950 562.050 532.050 ;
        RECT 544.950 527.100 547.050 529.200 ;
        RECT 545.400 526.050 546.600 527.100 ;
        RECT 544.950 523.950 547.050 526.050 ;
        RECT 547.950 523.950 550.050 526.050 ;
        RECT 548.400 522.900 549.600 523.950 ;
        RECT 554.400 522.900 555.600 529.950 ;
        RECT 562.950 527.100 565.050 529.200 ;
        RECT 566.400 529.050 567.600 563.400 ;
        RECT 578.400 558.600 579.600 565.950 ;
        RECT 575.400 557.400 579.600 558.600 ;
        RECT 563.400 526.050 564.600 527.100 ;
        RECT 565.950 526.950 568.050 529.050 ;
        RECT 568.950 526.950 571.050 529.050 ;
        RECT 571.950 526.950 574.050 529.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 535.950 520.800 538.050 522.900 ;
        RECT 547.950 520.800 550.050 522.900 ;
        RECT 553.950 520.800 556.050 522.900 ;
        RECT 536.400 517.050 537.600 520.800 ;
        RECT 560.400 517.050 561.600 523.950 ;
        RECT 565.950 520.950 568.050 523.050 ;
        RECT 535.950 514.950 538.050 517.050 ;
        RECT 559.950 514.950 562.050 517.050 ;
        RECT 532.950 495.000 535.050 499.050 ;
        RECT 541.950 496.950 544.050 499.050 ;
        RECT 533.400 493.050 534.600 495.000 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 536.400 489.900 537.600 490.950 ;
        RECT 542.400 490.050 543.600 496.950 ;
        RECT 553.950 495.000 556.050 499.050 ;
        RECT 559.950 495.000 562.050 499.050 ;
        RECT 554.400 493.050 555.600 495.000 ;
        RECT 560.400 493.050 561.600 495.000 ;
        RECT 550.950 490.950 553.050 493.050 ;
        RECT 553.950 490.950 556.050 493.050 ;
        RECT 556.950 490.950 559.050 493.050 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 535.950 487.800 538.050 489.900 ;
        RECT 541.950 487.950 544.050 490.050 ;
        RECT 551.400 489.900 552.600 490.950 ;
        RECT 550.950 487.800 553.050 489.900 ;
        RECT 547.950 484.950 550.050 487.050 ;
        RECT 526.950 481.950 529.050 484.050 ;
        RECT 508.950 472.950 511.050 475.050 ;
        RECT 538.950 463.950 541.050 466.050 ;
        RECT 529.950 457.950 532.050 460.050 ;
        RECT 517.950 454.950 520.050 457.050 ;
        RECT 496.950 451.950 499.050 454.050 ;
        RECT 502.950 451.950 505.050 454.050 ;
        RECT 472.950 439.950 475.050 442.050 ;
        RECT 460.950 436.950 463.050 439.050 ;
        RECT 466.950 436.950 469.050 439.050 ;
        RECT 457.950 385.950 460.050 388.050 ;
        RECT 461.400 379.050 462.600 436.950 ;
        RECT 476.400 436.050 477.600 442.950 ;
        RECT 481.950 442.800 484.050 444.900 ;
        RECT 487.950 442.800 490.050 444.900 ;
        RECT 490.950 442.950 493.050 445.050 ;
        RECT 493.950 442.950 496.050 445.050 ;
        RECT 484.950 439.950 487.050 442.050 ;
        RECT 475.950 433.950 478.050 436.050 ;
        RECT 475.950 423.000 478.050 427.050 ;
        RECT 472.500 420.300 474.600 422.400 ;
        RECT 476.400 420.900 477.600 423.000 ;
        RECT 470.400 415.050 471.600 417.600 ;
        RECT 463.950 412.950 466.050 415.050 ;
        RECT 469.950 412.950 472.050 415.050 ;
        RECT 472.950 414.900 473.850 420.300 ;
        RECT 475.800 418.800 477.900 420.900 ;
        RECT 479.700 417.900 481.800 419.700 ;
        RECT 474.750 416.700 483.300 417.900 ;
        RECT 474.750 415.800 476.850 416.700 ;
        RECT 472.950 413.700 479.700 414.900 ;
        RECT 464.400 400.050 465.600 412.950 ;
        RECT 472.950 406.500 474.000 413.700 ;
        RECT 475.800 410.100 477.900 412.200 ;
        RECT 478.800 411.300 479.700 413.700 ;
        RECT 476.400 407.550 477.600 410.100 ;
        RECT 478.800 409.200 480.900 411.300 ;
        RECT 482.400 407.700 483.300 416.700 ;
        RECT 485.400 415.050 486.600 439.950 ;
        RECT 484.500 412.950 486.600 415.050 ;
        RECT 487.950 412.950 490.050 415.050 ;
        RECT 484.950 409.800 487.050 412.950 ;
        RECT 472.500 404.400 474.600 406.500 ;
        RECT 482.100 405.600 484.200 407.700 ;
        RECT 488.400 402.600 489.600 412.950 ;
        RECT 491.400 403.050 492.600 442.950 ;
        RECT 493.950 433.950 496.050 436.050 ;
        RECT 494.400 418.050 495.600 433.950 ;
        RECT 497.400 421.050 498.600 451.950 ;
        RECT 505.950 449.100 508.050 451.200 ;
        RECT 506.400 448.050 507.600 449.100 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 503.400 430.050 504.600 445.950 ;
        RECT 509.400 430.050 510.600 445.950 ;
        RECT 518.400 444.900 519.600 454.950 ;
        RECT 523.950 449.100 526.050 451.200 ;
        RECT 524.400 448.050 525.600 449.100 ;
        RECT 530.400 448.050 531.600 457.950 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 529.950 445.950 532.050 448.050 ;
        RECT 532.950 445.950 535.050 448.050 ;
        RECT 527.400 444.900 528.600 445.950 ;
        RECT 517.950 442.800 520.050 444.900 ;
        RECT 526.950 442.800 529.050 444.900 ;
        RECT 502.950 427.950 505.050 430.050 ;
        RECT 508.950 427.950 511.050 430.050 ;
        RECT 517.950 427.950 520.050 430.050 ;
        RECT 496.950 418.950 499.050 421.050 ;
        RECT 493.950 415.950 496.050 418.050 ;
        RECT 502.950 416.100 505.050 418.200 ;
        RECT 509.400 418.050 510.600 427.950 ;
        RECT 511.950 418.950 514.050 421.050 ;
        RECT 503.400 415.050 504.600 416.100 ;
        RECT 508.950 415.950 511.050 418.050 ;
        RECT 496.950 412.950 499.050 415.050 ;
        RECT 502.950 412.950 505.050 415.050 ;
        RECT 505.950 412.950 508.050 415.050 ;
        RECT 493.950 409.950 496.050 412.050 ;
        RECT 485.400 401.400 489.600 402.600 ;
        RECT 463.950 397.950 466.050 400.050 ;
        RECT 466.950 388.950 469.050 391.050 ;
        RECT 460.950 378.600 463.050 379.050 ;
        RECT 460.950 377.400 465.600 378.600 ;
        RECT 460.950 376.950 463.050 377.400 ;
        RECT 443.400 374.400 447.600 375.600 ;
        RECT 454.950 375.600 457.050 376.050 ;
        RECT 454.950 374.400 459.600 375.600 ;
        RECT 418.950 367.800 421.050 369.900 ;
        RECT 424.950 367.800 427.050 369.900 ;
        RECT 427.950 367.800 430.050 369.900 ;
        RECT 433.950 367.800 436.050 369.900 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 419.400 366.750 420.600 367.800 ;
        RECT 412.950 364.650 415.050 366.750 ;
        RECT 418.800 364.650 420.900 366.750 ;
        RECT 421.950 361.950 424.050 367.050 ;
        RECT 428.400 358.050 429.600 367.800 ;
        RECT 436.950 361.950 439.050 367.050 ;
        RECT 427.950 355.950 430.050 358.050 ;
        RECT 424.950 352.950 427.050 355.050 ;
        RECT 425.400 349.050 426.600 352.950 ;
        RECT 424.950 346.950 427.050 349.050 ;
        RECT 421.950 343.950 424.050 346.050 ;
        RECT 422.400 337.050 423.600 343.950 ;
        RECT 440.400 340.200 441.600 367.950 ;
        RECT 433.950 338.100 436.050 340.200 ;
        RECT 439.950 338.100 442.050 340.200 ;
        RECT 434.400 337.050 435.600 338.100 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 421.950 334.950 424.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 436.950 334.950 439.050 337.050 ;
        RECT 416.400 334.050 417.600 334.950 ;
        RECT 412.950 332.400 417.600 334.050 ;
        RECT 437.400 333.900 438.600 334.950 ;
        RECT 412.950 331.950 417.000 332.400 ;
        RECT 436.950 331.800 439.050 333.900 ;
        RECT 409.950 328.950 412.050 331.050 ;
        RECT 415.950 328.950 418.050 331.050 ;
        RECT 407.400 326.400 411.600 327.600 ;
        RECT 391.950 322.950 394.050 325.050 ;
        RECT 374.400 293.400 379.050 294.600 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 361.950 289.950 364.050 292.050 ;
        RECT 364.950 289.950 367.050 292.050 ;
        RECT 367.950 289.950 370.050 292.050 ;
        RECT 359.400 288.000 360.600 289.950 ;
        RECT 365.400 288.900 366.600 289.950 ;
        RECT 374.400 288.900 375.600 293.400 ;
        RECT 376.950 293.100 379.050 293.400 ;
        RECT 380.400 296.400 384.600 297.600 ;
        RECT 380.400 292.050 381.600 296.400 ;
        RECT 388.950 295.950 391.050 298.050 ;
        RECT 385.950 293.100 388.050 295.200 ;
        RECT 386.400 292.050 387.600 293.100 ;
        RECT 379.950 289.950 382.050 292.050 ;
        RECT 382.950 289.950 385.050 292.050 ;
        RECT 385.950 289.950 388.050 292.050 ;
        RECT 358.950 283.950 361.050 288.000 ;
        RECT 364.950 286.800 367.050 288.900 ;
        RECT 373.950 286.800 376.050 288.900 ;
        RECT 383.400 280.050 384.600 289.950 ;
        RECT 367.950 277.950 370.050 280.050 ;
        RECT 382.950 277.950 385.050 280.050 ;
        RECT 355.950 274.950 358.050 277.050 ;
        RECT 356.400 255.900 357.600 274.950 ;
        RECT 358.800 271.950 360.900 274.050 ;
        RECT 361.950 271.950 364.050 274.050 ;
        RECT 359.400 265.050 360.600 271.950 ;
        RECT 362.400 268.050 363.600 271.950 ;
        RECT 361.950 265.950 364.050 268.050 ;
        RECT 358.950 262.950 361.050 265.050 ;
        RECT 362.400 259.050 363.600 265.950 ;
        RECT 368.400 259.050 369.600 277.950 ;
        RECT 373.950 268.950 376.050 271.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 364.950 256.950 367.050 259.050 ;
        RECT 367.950 256.950 370.050 259.050 ;
        RECT 355.950 253.800 358.050 255.900 ;
        RECT 365.400 252.600 366.600 256.950 ;
        RECT 370.950 253.950 373.050 256.050 ;
        RECT 365.400 251.400 369.600 252.600 ;
        RECT 349.950 233.400 354.600 234.600 ;
        RECT 349.950 232.950 352.050 233.400 ;
        RECT 340.950 202.950 343.050 205.050 ;
        RECT 346.950 202.950 349.050 205.050 ;
        RECT 326.400 186.000 330.600 186.600 ;
        RECT 325.950 185.400 330.600 186.000 ;
        RECT 325.950 184.050 328.050 185.400 ;
        RECT 331.800 184.950 333.900 187.050 ;
        RECT 325.800 183.000 328.050 184.050 ;
        RECT 325.800 181.950 327.900 183.000 ;
        RECT 328.950 182.100 331.050 184.200 ;
        RECT 334.950 183.000 337.050 187.050 ;
        RECT 341.400 184.050 342.600 202.950 ;
        RECT 347.400 196.050 348.600 202.950 ;
        RECT 346.950 193.950 349.050 196.050 ;
        RECT 350.400 189.600 351.600 232.950 ;
        RECT 361.950 229.950 364.050 232.050 ;
        RECT 355.950 215.100 358.050 217.200 ;
        RECT 356.400 214.050 357.600 215.100 ;
        RECT 362.400 214.050 363.600 229.950 ;
        RECT 364.950 226.950 367.050 229.050 ;
        RECT 365.400 223.050 366.600 226.950 ;
        RECT 364.950 220.950 367.050 223.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 347.400 188.400 351.600 189.600 ;
        RECT 329.400 181.050 330.600 182.100 ;
        RECT 335.400 181.050 336.600 183.000 ;
        RECT 340.950 181.950 343.050 184.050 ;
        RECT 343.950 181.950 346.050 184.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 334.950 178.950 337.050 181.050 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 332.400 177.900 333.600 178.950 ;
        RECT 338.400 177.900 339.600 178.950 ;
        RECT 344.400 177.900 345.600 181.950 ;
        RECT 305.400 163.050 306.600 175.950 ;
        RECT 310.950 172.950 313.050 177.000 ;
        RECT 316.950 175.800 319.050 177.900 ;
        RECT 322.950 175.800 325.050 177.900 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 337.950 175.800 340.050 177.900 ;
        RECT 343.950 175.800 346.050 177.900 ;
        RECT 304.950 160.950 307.050 163.050 ;
        RECT 298.950 142.950 301.050 145.050 ;
        RECT 290.400 136.050 291.600 138.000 ;
        RECT 295.950 136.950 298.050 139.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 292.950 133.950 295.050 136.050 ;
        RECT 287.400 132.900 288.600 133.950 ;
        RECT 293.400 132.900 294.600 133.950 ;
        RECT 299.400 132.900 300.600 142.950 ;
        RECT 305.400 139.200 306.600 160.950 ;
        RECT 313.950 154.950 316.050 157.050 ;
        RECT 310.950 148.950 313.050 151.050 ;
        RECT 301.950 136.950 304.050 139.050 ;
        RECT 304.950 137.100 307.050 139.200 ;
        RECT 286.950 130.800 289.050 132.900 ;
        RECT 292.950 130.800 295.050 132.900 ;
        RECT 298.950 130.800 301.050 132.900 ;
        RECT 292.950 121.950 295.050 124.050 ;
        RECT 293.400 118.050 294.600 121.950 ;
        RECT 289.800 117.000 291.900 118.050 ;
        RECT 289.800 115.950 292.050 117.000 ;
        RECT 292.950 115.950 295.050 118.050 ;
        RECT 286.950 112.950 289.050 115.050 ;
        RECT 289.950 114.600 292.050 115.950 ;
        RECT 289.950 114.000 294.600 114.600 ;
        RECT 290.400 113.400 294.600 114.000 ;
        RECT 262.950 103.950 265.050 106.050 ;
        RECT 268.950 104.100 271.050 106.200 ;
        RECT 274.950 105.000 277.050 109.050 ;
        RECT 277.950 106.950 280.050 109.050 ;
        RECT 283.950 106.950 286.050 109.050 ;
        RECT 250.950 94.950 253.050 99.900 ;
        RECT 259.950 97.950 262.050 100.050 ;
        RECT 263.400 97.050 264.600 103.950 ;
        RECT 269.400 103.050 270.600 104.100 ;
        RECT 275.400 103.050 276.600 105.000 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 274.950 100.950 277.050 103.050 ;
        RECT 277.950 100.950 280.050 103.050 ;
        RECT 262.950 94.950 265.050 97.050 ;
        RECT 265.950 94.950 268.050 100.050 ;
        RECT 244.950 91.950 247.050 94.050 ;
        RECT 223.950 88.950 226.050 91.050 ;
        RECT 247.950 85.950 250.050 88.050 ;
        RECT 241.950 82.950 244.050 85.050 ;
        RECT 211.950 67.950 214.050 70.050 ;
        RECT 215.100 64.200 217.200 66.300 ;
        RECT 224.100 64.500 226.200 66.600 ;
        RECT 235.950 64.950 238.050 67.050 ;
        RECT 208.950 61.950 211.050 64.050 ;
        RECT 209.400 52.050 210.600 61.950 ;
        RECT 212.400 58.050 213.600 60.450 ;
        RECT 211.950 57.900 214.050 58.050 ;
        RECT 211.950 55.950 214.500 57.900 ;
        RECT 212.400 55.800 214.500 55.950 ;
        RECT 208.950 49.950 211.050 52.050 ;
        RECT 215.400 51.600 216.300 64.200 ;
        RECT 221.400 61.200 222.600 63.450 ;
        RECT 220.950 60.900 223.050 61.200 ;
        RECT 220.950 59.100 223.500 60.900 ;
        RECT 221.400 58.800 223.500 59.100 ;
        RECT 217.200 57.900 219.300 58.200 ;
        RECT 225.150 57.900 226.050 64.500 ;
        RECT 217.200 57.000 226.050 57.900 ;
        RECT 217.200 56.100 219.300 57.000 ;
        RECT 222.150 55.200 224.250 56.100 ;
        RECT 217.200 54.000 224.250 55.200 ;
        RECT 217.200 53.100 219.300 54.000 ;
        RECT 214.650 49.500 216.750 51.600 ;
        RECT 221.400 50.100 223.500 52.200 ;
        RECT 225.150 51.900 226.050 57.000 ;
        RECT 226.950 55.800 229.050 57.900 ;
        RECT 227.400 53.400 228.600 55.800 ;
        RECT 205.950 46.950 208.050 49.050 ;
        RECT 221.400 40.050 222.600 50.100 ;
        RECT 224.700 49.800 226.800 51.900 ;
        RECT 223.950 43.950 226.050 46.050 ;
        RECT 220.950 37.950 223.050 40.050 ;
        RECT 193.950 34.950 196.050 37.050 ;
        RECT 199.950 26.100 202.050 28.200 ;
        RECT 208.950 26.100 211.050 28.200 ;
        RECT 214.950 26.100 217.050 28.200 ;
        RECT 181.950 22.950 184.050 25.050 ;
        RECT 184.950 22.950 187.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 190.950 22.950 193.050 25.050 ;
        RECT 182.400 21.900 183.600 22.950 ;
        RECT 181.950 19.800 184.050 21.900 ;
        RECT 188.400 21.000 189.600 22.950 ;
        RECT 172.800 16.950 174.900 19.050 ;
        RECT 175.950 16.950 178.050 19.050 ;
        RECT 187.950 16.950 190.050 21.000 ;
        RECT 190.950 16.950 193.050 19.050 ;
        RECT 133.950 13.950 136.050 16.050 ;
        RECT 181.950 12.600 184.050 16.050 ;
        RECT 186.000 15.900 189.000 16.050 ;
        RECT 184.950 13.950 190.050 15.900 ;
        RECT 184.950 13.800 187.050 13.950 ;
        RECT 187.950 13.800 190.050 13.950 ;
        RECT 191.400 12.600 192.600 16.950 ;
        RECT 181.950 12.000 192.600 12.600 ;
        RECT 182.400 11.400 192.600 12.000 ;
        RECT 200.400 7.050 201.600 26.100 ;
        RECT 209.400 25.050 210.600 26.100 ;
        RECT 215.400 25.050 216.600 26.100 ;
        RECT 220.950 25.950 223.050 28.050 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 206.400 21.000 207.600 22.950 ;
        RECT 212.400 21.900 213.600 22.950 ;
        RECT 221.400 21.900 222.600 25.950 ;
        RECT 205.950 16.950 208.050 21.000 ;
        RECT 211.950 19.800 214.050 21.900 ;
        RECT 220.950 19.800 223.050 21.900 ;
        RECT 224.400 13.050 225.600 43.950 ;
        RECT 229.950 40.950 232.050 43.050 ;
        RECT 226.950 34.950 229.050 37.050 ;
        RECT 227.400 21.900 228.600 34.950 ;
        RECT 230.400 28.050 231.600 40.950 ;
        RECT 229.950 25.950 232.050 28.050 ;
        RECT 236.400 25.050 237.600 64.950 ;
        RECT 242.400 61.050 243.600 82.950 ;
        RECT 248.400 61.200 249.600 85.950 ;
        RECT 272.400 82.050 273.600 100.950 ;
        RECT 278.400 99.900 279.600 100.950 ;
        RECT 277.950 97.800 280.050 99.900 ;
        RECT 271.950 79.950 274.050 82.050 ;
        RECT 253.950 73.950 256.050 76.050 ;
        RECT 238.950 58.950 243.600 61.050 ;
        RECT 247.950 59.100 250.050 61.200 ;
        RECT 242.400 58.050 243.600 58.950 ;
        RECT 248.400 58.050 249.600 59.100 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 241.950 34.950 244.050 37.050 ;
        RECT 242.400 28.050 243.600 34.950 ;
        RECT 245.400 34.050 246.600 55.950 ;
        RECT 254.400 52.050 255.600 73.950 ;
        RECT 278.400 73.050 279.600 97.800 ;
        RECT 284.400 88.050 285.600 106.950 ;
        RECT 287.400 106.050 288.600 112.950 ;
        RECT 286.950 103.950 289.050 106.050 ;
        RECT 293.400 103.050 294.600 113.400 ;
        RECT 298.950 109.950 301.050 112.050 ;
        RECT 299.400 103.050 300.600 109.950 ;
        RECT 302.400 105.600 303.600 136.950 ;
        RECT 311.400 136.050 312.600 148.950 ;
        RECT 314.400 141.600 315.600 154.950 ;
        RECT 328.950 148.950 331.050 151.050 ;
        RECT 322.950 145.950 325.050 148.050 ;
        RECT 316.950 142.950 322.050 145.050 ;
        RECT 314.400 140.400 318.600 141.600 ;
        RECT 317.400 136.050 318.600 140.400 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 310.950 133.950 313.050 136.050 ;
        RECT 313.950 133.950 316.050 136.050 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 308.400 132.000 309.600 133.950 ;
        RECT 314.400 132.900 315.600 133.950 ;
        RECT 323.400 132.900 324.600 145.950 ;
        RECT 325.950 142.950 328.050 148.050 ;
        RECT 307.950 127.950 310.050 132.000 ;
        RECT 313.950 130.800 316.050 132.900 ;
        RECT 322.950 130.800 325.050 132.900 ;
        RECT 310.950 118.950 313.050 121.050 ;
        RECT 322.950 118.950 325.050 121.050 ;
        RECT 311.400 106.050 312.600 118.950 ;
        RECT 302.400 104.400 306.600 105.600 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 292.950 100.950 295.050 103.050 ;
        RECT 295.950 100.950 298.050 103.050 ;
        RECT 298.950 100.950 301.050 103.050 ;
        RECT 290.400 99.900 291.600 100.950 ;
        RECT 289.950 97.800 292.050 99.900 ;
        RECT 296.400 91.050 297.600 100.950 ;
        RECT 301.950 97.950 304.050 100.050 ;
        RECT 295.950 88.950 298.050 91.050 ;
        RECT 283.950 85.950 286.050 88.050 ;
        RECT 302.400 82.050 303.600 97.950 ;
        RECT 305.400 85.050 306.600 104.400 ;
        RECT 307.950 103.950 310.050 106.050 ;
        RECT 310.950 103.950 313.050 106.050 ;
        RECT 316.950 104.100 319.050 106.200 ;
        RECT 304.950 82.950 307.050 85.050 ;
        RECT 301.950 79.950 304.050 82.050 ;
        RECT 304.950 76.950 307.050 79.050 ;
        RECT 277.950 70.950 280.050 73.050 ;
        RECT 256.950 67.950 259.050 70.050 ;
        RECT 271.950 67.950 274.050 70.050 ;
        RECT 253.950 49.950 256.050 52.050 ;
        RECT 250.950 43.950 253.050 46.050 ;
        RECT 251.400 37.050 252.600 43.950 ;
        RECT 257.400 43.050 258.600 67.950 ;
        RECT 259.950 59.100 262.050 61.200 ;
        RECT 265.950 59.100 268.050 61.200 ;
        RECT 260.400 52.050 261.600 59.100 ;
        RECT 266.400 58.050 267.600 59.100 ;
        RECT 272.400 58.050 273.600 67.950 ;
        RECT 295.950 64.950 298.050 67.050 ;
        RECT 277.950 59.100 280.050 61.200 ;
        RECT 289.950 59.100 292.050 61.200 ;
        RECT 278.400 58.050 279.600 59.100 ;
        RECT 290.400 58.050 291.600 59.100 ;
        RECT 296.400 58.050 297.600 64.950 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 295.950 55.950 298.050 58.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 269.400 54.000 270.600 55.950 ;
        RECT 275.400 54.900 276.600 55.950 ;
        RECT 293.400 54.900 294.600 55.950 ;
        RECT 259.950 49.950 262.050 52.050 ;
        RECT 268.950 49.950 271.050 54.000 ;
        RECT 274.950 52.800 277.050 54.900 ;
        RECT 292.950 49.950 295.050 54.900 ;
        RECT 299.400 49.050 300.600 55.950 ;
        RECT 305.400 52.050 306.600 76.950 ;
        RECT 308.400 61.200 309.600 103.950 ;
        RECT 317.400 103.050 318.600 104.100 ;
        RECT 323.400 103.050 324.600 118.950 ;
        RECT 329.400 118.050 330.600 148.950 ;
        RECT 334.950 137.100 337.050 139.200 ;
        RECT 344.400 139.050 345.600 175.800 ;
        RECT 347.400 175.050 348.600 188.400 ;
        RECT 359.400 187.050 360.600 211.950 ;
        RECT 361.950 205.950 364.050 208.050 ;
        RECT 349.950 184.950 352.050 187.050 ;
        RECT 358.950 184.950 361.050 187.050 ;
        RECT 346.950 172.950 349.050 175.050 ;
        RECT 350.400 166.050 351.600 184.950 ;
        RECT 355.950 182.100 358.050 184.200 ;
        RECT 356.400 181.050 357.600 182.100 ;
        RECT 362.400 181.050 363.600 205.950 ;
        RECT 368.400 186.600 369.600 251.400 ;
        RECT 371.400 220.050 372.600 253.950 ;
        RECT 374.400 250.050 375.600 268.950 ;
        RECT 382.950 260.100 385.050 262.200 ;
        RECT 383.400 259.050 384.600 260.100 ;
        RECT 379.950 256.950 382.050 259.050 ;
        RECT 382.950 256.950 385.050 259.050 ;
        RECT 385.950 256.950 388.050 259.050 ;
        RECT 380.400 255.900 381.600 256.950 ;
        RECT 379.950 253.800 382.050 255.900 ;
        RECT 373.950 247.950 376.050 250.050 ;
        RECT 374.400 220.050 375.600 247.950 ;
        RECT 386.400 247.050 387.600 256.950 ;
        RECT 392.400 255.900 393.600 322.950 ;
        RECT 395.400 271.050 396.600 325.950 ;
        RECT 400.950 313.950 403.050 316.050 ;
        RECT 401.400 295.200 402.600 313.950 ;
        RECT 406.950 301.950 409.050 304.050 ;
        RECT 400.950 293.100 403.050 295.200 ;
        RECT 401.400 292.050 402.600 293.100 ;
        RECT 407.400 292.050 408.600 301.950 ;
        RECT 410.400 295.050 411.600 326.400 ;
        RECT 412.950 310.950 415.050 313.050 ;
        RECT 409.950 292.950 412.050 295.050 ;
        RECT 413.400 292.050 414.600 310.950 ;
        RECT 400.950 289.950 403.050 292.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 406.950 289.950 409.050 292.050 ;
        RECT 412.950 289.950 415.050 292.050 ;
        RECT 397.950 286.950 400.050 289.050 ;
        RECT 394.950 268.950 397.050 271.050 ;
        RECT 394.950 262.950 397.050 265.050 ;
        RECT 395.400 256.050 396.600 262.950 ;
        RECT 398.400 262.050 399.600 286.950 ;
        RECT 404.400 271.050 405.600 289.950 ;
        RECT 416.400 288.600 417.600 328.950 ;
        RECT 443.400 322.050 444.600 374.400 ;
        RECT 454.950 373.950 457.050 374.400 ;
        RECT 445.950 370.950 448.050 373.050 ;
        RECT 451.950 371.100 454.050 373.200 ;
        RECT 446.400 361.050 447.600 370.950 ;
        RECT 452.400 370.050 453.600 371.100 ;
        RECT 458.400 370.050 459.600 374.400 ;
        RECT 464.400 373.050 465.600 377.400 ;
        RECT 463.950 370.950 466.050 373.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 457.950 367.950 460.050 370.050 ;
        RECT 460.950 367.950 463.050 370.050 ;
        RECT 448.950 364.950 451.050 367.050 ;
        RECT 455.400 366.000 456.600 367.950 ;
        RECT 461.400 366.900 462.600 367.950 ;
        RECT 445.950 358.950 448.050 361.050 ;
        RECT 445.950 352.950 448.050 355.050 ;
        RECT 446.400 325.050 447.600 352.950 ;
        RECT 449.400 349.050 450.600 364.950 ;
        RECT 454.950 361.950 457.050 366.000 ;
        RECT 460.950 364.800 463.050 366.900 ;
        RECT 460.950 361.650 463.050 363.750 ;
        RECT 448.950 346.950 451.050 349.050 ;
        RECT 454.950 346.950 457.050 349.050 ;
        RECT 448.950 338.100 451.050 340.200 ;
        RECT 449.400 334.050 450.600 338.100 ;
        RECT 455.400 337.050 456.600 346.950 ;
        RECT 461.400 340.200 462.600 361.650 ;
        RECT 467.400 355.050 468.600 388.950 ;
        RECT 475.950 371.100 478.050 373.200 ;
        RECT 476.400 370.050 477.600 371.100 ;
        RECT 472.950 367.950 475.050 370.050 ;
        RECT 475.950 367.950 478.050 370.050 ;
        RECT 473.400 367.050 474.600 367.950 ;
        RECT 469.950 365.400 474.600 367.050 ;
        RECT 469.950 364.950 474.000 365.400 ;
        RECT 469.950 355.950 472.050 358.050 ;
        RECT 466.950 352.950 469.050 355.050 ;
        RECT 460.950 338.100 463.050 340.200 ;
        RECT 461.400 337.050 462.600 338.100 ;
        RECT 470.400 337.050 471.600 355.950 ;
        RECT 475.950 338.100 478.050 340.200 ;
        RECT 476.400 337.050 477.600 338.100 ;
        RECT 454.950 334.950 457.050 337.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 460.950 334.950 463.050 337.050 ;
        RECT 469.950 334.950 472.050 337.050 ;
        RECT 472.950 334.950 475.050 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 448.950 331.950 451.050 334.050 ;
        RECT 458.400 333.000 459.600 334.950 ;
        RECT 473.400 333.000 474.600 334.950 ;
        RECT 457.950 328.950 460.050 333.000 ;
        RECT 472.950 328.950 475.050 333.000 ;
        RECT 485.400 328.050 486.600 401.400 ;
        RECT 490.950 400.950 493.050 403.050 ;
        RECT 491.400 382.050 492.600 400.950 ;
        RECT 494.400 391.050 495.600 409.950 ;
        RECT 497.400 409.050 498.600 412.950 ;
        RECT 499.950 409.950 502.050 412.050 ;
        RECT 496.950 406.950 499.050 409.050 ;
        RECT 497.400 397.050 498.600 406.950 ;
        RECT 496.950 394.950 499.050 397.050 ;
        RECT 493.950 388.950 496.050 391.050 ;
        RECT 500.400 385.050 501.600 409.950 ;
        RECT 506.400 397.050 507.600 412.950 ;
        RECT 505.950 394.950 508.050 397.050 ;
        RECT 505.950 388.950 508.050 391.050 ;
        RECT 499.950 382.950 502.050 385.050 ;
        RECT 490.950 379.950 493.050 382.050 ;
        RECT 502.950 379.950 505.050 382.050 ;
        RECT 493.950 372.000 496.050 376.050 ;
        RECT 503.400 373.050 504.600 379.950 ;
        RECT 494.400 370.050 495.600 372.000 ;
        RECT 502.950 370.950 505.050 373.050 ;
        RECT 490.950 367.950 493.050 370.050 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 491.400 366.900 492.600 367.950 ;
        RECT 490.950 364.800 493.050 366.900 ;
        RECT 497.400 366.000 498.600 367.950 ;
        RECT 496.950 361.950 499.050 366.000 ;
        RECT 506.400 349.050 507.600 388.950 ;
        RECT 512.400 382.050 513.600 418.950 ;
        RECT 518.400 415.050 519.600 427.950 ;
        RECT 523.950 416.100 526.050 418.200 ;
        RECT 524.400 415.050 525.600 416.100 ;
        RECT 517.950 412.950 520.050 415.050 ;
        RECT 520.950 412.950 523.050 415.050 ;
        RECT 523.950 412.950 526.050 415.050 ;
        RECT 521.400 411.000 522.600 412.950 ;
        RECT 520.950 406.950 523.050 411.000 ;
        RECT 511.950 379.950 514.050 382.050 ;
        RECT 533.400 376.050 534.600 445.950 ;
        RECT 539.400 444.900 540.600 463.950 ;
        RECT 548.400 448.050 549.600 484.950 ;
        RECT 557.400 469.050 558.600 490.950 ;
        RECT 566.400 489.900 567.600 520.950 ;
        RECT 569.400 502.050 570.600 526.950 ;
        RECT 568.950 499.950 571.050 502.050 ;
        RECT 572.400 495.600 573.600 526.950 ;
        RECT 575.400 514.050 576.600 557.400 ;
        RECT 581.400 532.050 582.600 577.950 ;
        RECT 589.950 572.100 592.050 574.200 ;
        RECT 596.400 574.050 597.600 610.950 ;
        RECT 602.400 604.050 603.600 610.950 ;
        RECT 607.950 606.000 610.050 610.050 ;
        RECT 608.400 604.050 609.600 606.000 ;
        RECT 610.950 604.950 613.050 610.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 604.950 601.950 607.050 604.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 605.400 600.900 606.600 601.950 ;
        RECT 604.950 598.800 607.050 600.900 ;
        RECT 614.400 598.050 615.600 637.950 ;
        RECT 620.400 631.050 621.600 643.950 ;
        RECT 619.950 628.950 622.050 631.050 ;
        RECT 616.950 610.950 619.050 613.050 ;
        RECT 598.950 595.950 601.050 598.050 ;
        RECT 613.950 595.950 616.050 598.050 ;
        RECT 590.400 571.050 591.600 572.100 ;
        RECT 595.950 571.950 598.050 574.050 ;
        RECT 599.400 571.050 600.600 595.950 ;
        RECT 610.950 577.950 613.050 580.050 ;
        RECT 601.950 572.400 604.050 574.500 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 598.950 568.950 601.050 571.050 ;
        RECT 583.950 565.950 586.050 568.050 ;
        RECT 584.400 553.050 585.600 565.950 ;
        RECT 583.950 550.950 586.050 553.050 ;
        RECT 587.400 549.600 588.600 568.950 ;
        RECT 593.400 567.900 594.600 568.950 ;
        RECT 592.950 565.800 595.050 567.900 ;
        RECT 598.950 565.800 601.050 567.900 ;
        RECT 602.400 567.600 603.600 572.400 ;
        RECT 611.400 571.050 612.600 577.950 ;
        RECT 617.400 577.050 618.600 610.950 ;
        RECT 620.400 607.050 621.600 628.950 ;
        RECT 626.400 619.050 627.600 646.950 ;
        RECT 628.950 643.950 631.050 646.050 ;
        RECT 629.400 628.050 630.600 643.950 ;
        RECT 628.950 625.950 631.050 628.050 ;
        RECT 625.950 616.950 628.050 619.050 ;
        RECT 632.400 610.050 633.600 670.950 ;
        RECT 634.950 661.950 637.050 664.050 ;
        RECT 635.400 625.050 636.600 661.950 ;
        RECT 643.950 655.950 646.050 658.050 ;
        RECT 640.650 653.400 642.750 655.500 ;
        RECT 638.400 647.100 640.500 649.200 ;
        RECT 638.400 637.050 639.600 647.100 ;
        RECT 641.400 640.800 642.300 653.400 ;
        RECT 644.400 651.900 645.600 655.950 ;
        RECT 647.400 654.900 648.600 657.450 ;
        RECT 647.400 652.800 649.500 654.900 ;
        RECT 650.700 653.100 652.800 655.200 ;
        RECT 643.200 651.000 645.600 651.900 ;
        RECT 643.200 649.800 650.250 651.000 ;
        RECT 648.150 648.900 650.250 649.800 ;
        RECT 643.200 648.000 645.300 648.900 ;
        RECT 651.150 648.000 652.050 653.100 ;
        RECT 658.950 652.950 661.050 655.050 ;
        RECT 653.400 649.200 654.600 651.600 ;
        RECT 643.200 647.100 652.050 648.000 ;
        RECT 652.950 647.100 655.050 649.200 ;
        RECT 643.200 646.800 645.300 647.100 ;
        RECT 647.400 644.100 649.500 646.200 ;
        RECT 641.100 638.700 643.200 640.800 ;
        RECT 637.950 634.950 640.050 637.050 ;
        RECT 634.950 622.950 637.050 625.050 ;
        RECT 647.400 619.050 648.600 644.100 ;
        RECT 651.150 640.500 652.050 647.100 ;
        RECT 650.100 638.400 652.200 640.500 ;
        RECT 634.950 616.950 637.050 619.050 ;
        RECT 646.950 616.950 649.050 619.050 ;
        RECT 619.950 604.950 622.050 607.050 ;
        RECT 622.950 606.000 625.050 610.050 ;
        RECT 628.800 609.000 630.900 610.050 ;
        RECT 628.800 607.950 631.050 609.000 ;
        RECT 631.950 607.950 634.050 610.050 ;
        RECT 623.400 604.050 624.600 606.000 ;
        RECT 628.950 605.100 631.050 607.950 ;
        RECT 635.400 607.050 636.600 616.950 ;
        RECT 652.950 613.950 655.050 616.050 ;
        RECT 645.000 609.600 649.050 610.050 ;
        RECT 644.400 607.950 649.050 609.600 ;
        RECT 629.400 604.050 630.600 605.100 ;
        RECT 634.950 604.950 637.050 607.050 ;
        RECT 637.950 605.100 640.050 607.200 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 625.950 601.950 628.050 604.050 ;
        RECT 628.950 601.950 631.050 604.050 ;
        RECT 631.950 601.950 634.050 604.050 ;
        RECT 619.950 598.950 622.050 601.050 ;
        RECT 616.950 574.950 619.050 577.050 ;
        RECT 620.400 573.600 621.600 598.950 ;
        RECT 626.400 586.050 627.600 601.950 ;
        RECT 632.400 600.900 633.600 601.950 ;
        RECT 631.950 598.800 634.050 600.900 ;
        RECT 638.400 600.600 639.600 605.100 ;
        RECT 644.400 604.050 645.600 607.950 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 646.950 601.950 649.050 604.050 ;
        RECT 647.400 600.900 648.600 601.950 ;
        RECT 653.400 600.900 654.600 613.950 ;
        RECT 655.950 610.950 658.050 613.050 ;
        RECT 635.400 599.400 639.600 600.600 ;
        RECT 632.400 589.050 633.600 598.800 ;
        RECT 631.950 586.950 634.050 589.050 ;
        RECT 625.950 583.950 628.050 586.050 ;
        RECT 631.950 583.800 634.050 585.900 ;
        RECT 625.950 578.400 628.050 580.500 ;
        RECT 617.400 572.400 621.600 573.600 ;
        RECT 622.950 572.400 625.050 574.500 ;
        RECT 617.400 571.050 618.600 572.400 ;
        RECT 623.400 571.050 624.600 572.400 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 616.950 568.950 619.050 571.050 ;
        RECT 622.950 568.950 625.050 571.050 ;
        RECT 602.400 566.400 606.600 567.600 ;
        RECT 593.400 564.600 594.600 565.800 ;
        RECT 584.400 548.400 588.600 549.600 ;
        RECT 590.400 563.400 594.600 564.600 ;
        RECT 584.400 547.050 585.600 548.400 ;
        RECT 583.950 544.950 586.050 547.050 ;
        RECT 580.950 529.950 583.050 532.050 ;
        RECT 584.400 528.600 585.600 544.950 ;
        RECT 590.400 529.050 591.600 563.400 ;
        RECT 599.400 555.600 600.600 565.800 ;
        RECT 601.950 555.600 604.050 556.050 ;
        RECT 599.400 554.400 604.050 555.600 ;
        RECT 601.950 553.950 604.050 554.400 ;
        RECT 595.950 537.300 598.050 539.400 ;
        RECT 596.850 533.700 598.050 537.300 ;
        RECT 595.950 531.600 598.050 533.700 ;
        RECT 581.400 527.400 585.600 528.600 ;
        RECT 581.400 526.050 582.600 527.400 ;
        RECT 589.950 526.950 592.050 529.050 ;
        RECT 580.950 523.950 583.050 526.050 ;
        RECT 586.950 523.950 589.050 526.050 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 574.950 511.950 577.050 514.050 ;
        RECT 587.400 511.050 588.600 523.950 ;
        RECT 593.400 522.600 594.600 523.950 ;
        RECT 592.950 520.500 595.050 522.600 ;
        RECT 596.850 516.600 598.050 531.600 ;
        RECT 602.400 526.050 603.600 553.950 ;
        RECT 601.950 523.950 604.050 526.050 ;
        RECT 605.400 520.050 606.600 566.400 ;
        RECT 608.400 553.050 609.600 568.950 ;
        RECT 614.400 559.050 615.600 568.950 ;
        RECT 626.850 563.400 628.050 578.400 ;
        RECT 632.400 568.050 633.600 583.800 ;
        RECT 631.950 565.950 634.050 568.050 ;
        RECT 625.950 561.300 628.050 563.400 ;
        RECT 631.950 562.800 634.050 564.900 ;
        RECT 613.950 556.950 616.050 559.050 ;
        RECT 626.850 557.700 628.050 561.300 ;
        RECT 625.950 555.600 628.050 557.700 ;
        RECT 607.950 550.950 610.050 553.050 ;
        RECT 622.950 547.950 625.050 550.050 ;
        RECT 616.950 536.400 619.050 538.500 ;
        RECT 610.950 528.000 613.050 532.050 ;
        RECT 611.400 526.050 612.600 528.000 ;
        RECT 610.950 523.950 613.050 526.050 ;
        RECT 604.950 517.950 607.050 520.050 ;
        RECT 610.950 517.950 613.050 520.050 ;
        RECT 595.950 514.500 598.050 516.600 ;
        RECT 607.950 511.950 610.050 514.050 ;
        RECT 586.950 508.950 589.050 511.050 ;
        RECT 598.950 502.950 601.050 505.050 ;
        RECT 580.950 499.950 583.050 502.050 ;
        RECT 569.400 494.400 573.600 495.600 ;
        RECT 565.950 487.800 568.050 489.900 ;
        RECT 556.950 466.950 559.050 469.050 ;
        RECT 569.400 466.050 570.600 494.400 ;
        RECT 574.950 494.100 577.050 496.200 ;
        RECT 575.400 493.050 576.600 494.100 ;
        RECT 581.400 493.050 582.600 499.950 ;
        RECT 589.950 496.950 592.050 499.050 ;
        RECT 574.950 490.950 577.050 493.050 ;
        RECT 577.950 490.950 580.050 493.050 ;
        RECT 580.950 490.950 583.050 493.050 ;
        RECT 583.950 490.950 586.050 493.050 ;
        RECT 578.400 489.900 579.600 490.950 ;
        RECT 584.400 489.900 585.600 490.950 ;
        RECT 590.400 489.900 591.600 496.950 ;
        RECT 599.400 493.050 600.600 502.950 ;
        RECT 604.950 494.100 607.050 496.200 ;
        RECT 608.400 496.050 609.600 511.950 ;
        RECT 605.400 493.050 606.600 494.100 ;
        RECT 607.950 493.950 610.050 496.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 598.950 490.950 601.050 493.050 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 604.950 490.950 607.050 493.050 ;
        RECT 577.950 484.950 580.050 489.900 ;
        RECT 583.950 487.800 586.050 489.900 ;
        RECT 589.950 487.800 592.050 489.900 ;
        RECT 596.400 489.000 597.600 490.950 ;
        RECT 602.400 489.900 603.600 490.950 ;
        RECT 574.950 483.600 577.050 484.050 ;
        RECT 580.950 483.600 583.050 487.050 ;
        RECT 595.950 484.950 598.050 489.000 ;
        RECT 601.950 487.800 604.050 489.900 ;
        RECT 607.950 487.950 610.050 490.050 ;
        RECT 574.950 483.000 583.050 483.600 ;
        RECT 574.950 482.400 582.600 483.000 ;
        RECT 574.950 481.950 577.050 482.400 ;
        RECT 598.950 481.950 601.050 487.050 ;
        RECT 574.950 475.950 577.050 478.050 ;
        RECT 575.400 472.050 576.600 475.950 ;
        RECT 574.950 469.950 577.050 472.050 ;
        RECT 568.950 463.950 571.050 466.050 ;
        RECT 565.950 459.300 568.050 461.400 ;
        RECT 571.950 460.950 574.050 463.050 ;
        RECT 566.850 455.700 568.050 459.300 ;
        RECT 565.950 453.600 568.050 455.700 ;
        RECT 553.950 449.100 556.050 451.200 ;
        RECT 554.400 448.050 555.600 449.100 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 553.950 445.950 556.050 448.050 ;
        RECT 562.950 445.950 565.050 448.050 ;
        RECT 545.400 444.900 546.600 445.950 ;
        RECT 538.950 442.800 541.050 444.900 ;
        RECT 544.950 442.800 547.050 444.900 ;
        RECT 535.950 439.950 538.050 442.050 ;
        RECT 536.400 391.050 537.600 439.950 ;
        RECT 551.400 430.050 552.600 445.950 ;
        RECT 563.400 444.600 564.600 445.950 ;
        RECT 560.400 443.400 565.050 444.600 ;
        RECT 560.400 436.050 561.600 443.400 ;
        RECT 562.950 442.500 565.050 443.400 ;
        RECT 566.850 438.600 568.050 453.600 ;
        RECT 572.400 451.200 573.600 460.950 ;
        RECT 571.950 449.100 574.050 451.200 ;
        RECT 565.950 436.500 568.050 438.600 ;
        RECT 559.950 433.950 562.050 436.050 ;
        RECT 572.400 433.050 573.600 449.100 ;
        RECT 575.400 444.600 576.600 469.950 ;
        RECT 608.400 469.050 609.600 487.950 ;
        RECT 611.400 478.050 612.600 517.950 ;
        RECT 617.100 516.600 618.300 536.400 ;
        RECT 623.400 528.600 624.600 547.950 ;
        RECT 625.950 535.950 628.050 538.050 ;
        RECT 620.400 527.400 624.600 528.600 ;
        RECT 620.400 526.050 621.600 527.400 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 616.950 514.500 619.050 516.600 ;
        RECT 626.400 499.050 627.600 535.950 ;
        RECT 632.400 508.050 633.600 562.800 ;
        RECT 635.400 559.050 636.600 599.400 ;
        RECT 646.950 598.800 649.050 600.900 ;
        RECT 652.950 598.800 655.050 600.900 ;
        RECT 637.950 595.950 640.050 598.050 ;
        RECT 638.400 574.050 639.600 595.950 ;
        RECT 646.950 578.400 649.050 580.500 ;
        RECT 637.950 571.950 640.050 574.050 ;
        RECT 640.950 568.950 643.050 571.050 ;
        RECT 641.400 567.600 642.600 568.950 ;
        RECT 640.950 565.500 643.050 567.600 ;
        RECT 634.950 556.950 637.050 559.050 ;
        RECT 647.100 558.600 648.300 578.400 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 650.400 567.600 651.600 568.950 ;
        RECT 650.400 566.400 654.600 567.600 ;
        RECT 635.400 529.050 636.600 556.950 ;
        RECT 646.950 556.500 649.050 558.600 ;
        RECT 653.400 550.050 654.600 566.400 ;
        RECT 652.950 547.950 655.050 550.050 ;
        RECT 649.950 544.950 652.050 547.050 ;
        RECT 637.950 541.950 640.050 544.050 ;
        RECT 634.950 526.950 637.050 529.050 ;
        RECT 638.400 526.050 639.600 541.950 ;
        RECT 637.950 523.950 640.050 526.050 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 631.950 505.950 634.050 508.050 ;
        RECT 613.950 496.950 616.050 499.050 ;
        RECT 625.950 496.950 628.050 499.050 ;
        RECT 610.950 475.950 613.050 478.050 ;
        RECT 607.950 466.950 610.050 469.050 ;
        RECT 601.950 463.950 604.050 466.050 ;
        RECT 586.950 458.400 589.050 460.500 ;
        RECT 580.950 454.950 583.050 457.050 ;
        RECT 581.400 448.050 582.600 454.950 ;
        RECT 580.950 445.950 583.050 448.050 ;
        RECT 575.400 443.400 579.600 444.600 ;
        RECT 565.950 430.950 568.050 433.050 ;
        RECT 571.950 430.950 574.050 433.050 ;
        RECT 550.950 427.950 553.050 430.050 ;
        RECT 559.950 427.950 562.050 430.050 ;
        RECT 541.950 416.100 544.050 418.200 ;
        RECT 547.950 416.100 550.050 418.200 ;
        RECT 542.400 415.050 543.600 416.100 ;
        RECT 548.400 415.050 549.600 416.100 ;
        RECT 556.950 415.950 559.050 418.050 ;
        RECT 541.950 412.950 544.050 415.050 ;
        RECT 544.950 412.950 547.050 415.050 ;
        RECT 547.950 412.950 550.050 415.050 ;
        RECT 550.950 412.950 553.050 415.050 ;
        RECT 541.950 400.950 544.050 403.050 ;
        RECT 535.950 388.950 538.050 391.050 ;
        RECT 523.950 373.950 526.050 376.050 ;
        RECT 532.950 373.950 535.050 376.050 ;
        RECT 517.950 371.100 520.050 373.200 ;
        RECT 518.400 370.050 519.600 371.100 ;
        RECT 511.950 367.950 514.050 370.050 ;
        RECT 517.950 367.950 520.050 370.050 ;
        RECT 512.400 367.050 513.600 367.950 ;
        RECT 508.950 365.400 513.600 367.050 ;
        RECT 508.950 364.950 513.000 365.400 ;
        RECT 520.950 364.950 523.050 367.050 ;
        RECT 505.950 346.950 508.050 349.050 ;
        RECT 511.950 340.950 514.050 343.050 ;
        RECT 490.950 337.950 493.050 340.050 ;
        RECT 502.950 338.100 505.050 340.200 ;
        RECT 508.950 338.100 511.050 340.200 ;
        RECT 491.400 331.050 492.600 337.950 ;
        RECT 503.400 337.050 504.600 338.100 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 490.950 328.950 493.050 331.050 ;
        RECT 475.950 325.950 478.050 328.050 ;
        RECT 484.950 325.950 487.050 328.050 ;
        RECT 445.950 322.950 448.050 325.050 ;
        RECT 442.950 319.950 445.050 322.050 ;
        RECT 418.950 294.600 423.000 295.050 ;
        RECT 418.950 292.950 423.600 294.600 ;
        RECT 427.950 294.000 430.050 298.050 ;
        RECT 422.400 292.050 423.600 292.950 ;
        RECT 428.400 292.050 429.600 294.000 ;
        RECT 436.950 293.100 439.050 295.200 ;
        RECT 442.950 293.100 445.050 295.200 ;
        RECT 451.950 293.100 454.050 295.200 ;
        RECT 460.950 293.100 463.050 295.200 ;
        RECT 467.400 293.400 474.600 294.600 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 424.950 289.950 427.050 292.050 ;
        RECT 427.950 289.950 430.050 292.050 ;
        RECT 430.950 289.950 433.050 292.050 ;
        RECT 413.400 287.400 417.600 288.600 ;
        RECT 406.950 274.950 409.050 277.050 ;
        RECT 403.950 268.950 406.050 271.050 ;
        RECT 407.400 268.050 408.600 274.950 ;
        RECT 413.400 274.050 414.600 287.400 ;
        RECT 418.950 286.950 421.050 289.050 ;
        RECT 415.950 283.950 418.050 286.050 ;
        RECT 412.950 271.950 415.050 274.050 ;
        RECT 406.950 265.950 409.050 268.050 ;
        RECT 397.950 259.950 400.050 262.050 ;
        RECT 403.950 260.100 406.050 262.200 ;
        RECT 404.400 259.050 405.600 260.100 ;
        RECT 400.950 256.950 403.050 259.050 ;
        RECT 403.950 256.950 406.050 259.050 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 391.800 253.800 393.900 255.900 ;
        RECT 394.950 253.950 397.050 256.050 ;
        RECT 401.400 255.900 402.600 256.950 ;
        RECT 410.400 255.900 411.600 256.950 ;
        RECT 400.950 253.800 403.050 255.900 ;
        RECT 409.950 253.800 412.050 255.900 ;
        RECT 392.400 247.050 393.600 253.800 ;
        RECT 416.400 253.050 417.600 283.950 ;
        RECT 419.400 271.050 420.600 286.950 ;
        RECT 425.400 280.050 426.600 289.950 ;
        RECT 431.400 288.000 432.600 289.950 ;
        RECT 430.950 283.950 433.050 288.000 ;
        RECT 437.400 286.050 438.600 293.100 ;
        RECT 443.400 292.050 444.600 293.100 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 445.950 289.950 448.050 292.050 ;
        RECT 446.400 288.900 447.600 289.950 ;
        RECT 445.950 286.800 448.050 288.900 ;
        RECT 436.950 283.950 439.050 286.050 ;
        RECT 445.800 285.000 447.900 285.750 ;
        RECT 445.800 283.650 448.050 285.000 ;
        RECT 448.950 283.950 451.050 286.050 ;
        RECT 445.950 280.950 448.050 283.650 ;
        RECT 424.950 277.950 427.050 280.050 ;
        RECT 436.950 274.950 439.050 277.050 ;
        RECT 418.950 268.950 421.050 271.050 ;
        RECT 427.950 265.950 430.050 268.050 ;
        RECT 428.400 259.050 429.600 265.950 ;
        RECT 421.950 256.950 424.050 259.050 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 430.950 256.950 433.050 259.050 ;
        RECT 422.400 255.900 423.600 256.950 ;
        RECT 421.950 253.800 424.050 255.900 ;
        RECT 409.950 250.650 412.050 252.750 ;
        RECT 415.950 250.950 418.050 253.050 ;
        RECT 400.950 247.950 403.050 250.050 ;
        RECT 385.950 244.950 388.050 247.050 ;
        RECT 391.950 244.950 394.050 247.050 ;
        RECT 370.800 217.950 372.900 220.050 ;
        RECT 373.950 217.950 376.050 220.050 ;
        RECT 370.950 214.800 373.050 216.900 ;
        RECT 376.950 215.100 379.050 217.200 ;
        RECT 385.950 216.000 388.050 220.050 ;
        RECT 394.950 216.000 397.050 220.050 ;
        RECT 401.400 217.200 402.600 247.950 ;
        RECT 371.400 190.050 372.600 214.800 ;
        RECT 377.400 214.050 378.600 215.100 ;
        RECT 386.400 214.050 387.600 216.000 ;
        RECT 395.400 214.050 396.600 216.000 ;
        RECT 400.950 215.100 403.050 217.200 ;
        RECT 401.400 214.050 402.600 215.100 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 379.950 211.950 382.050 214.050 ;
        RECT 385.950 211.950 388.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 400.950 211.950 403.050 214.050 ;
        RECT 380.400 210.900 381.600 211.950 ;
        RECT 379.950 208.800 382.050 210.900 ;
        RECT 376.950 202.950 379.050 205.050 ;
        RECT 391.950 202.950 394.050 205.050 ;
        RECT 370.950 187.950 373.050 190.050 ;
        RECT 377.400 187.050 378.600 202.950 ;
        RECT 368.400 185.400 372.600 186.600 ;
        RECT 355.950 178.950 358.050 181.050 ;
        RECT 358.950 178.950 361.050 181.050 ;
        RECT 361.950 178.950 364.050 181.050 ;
        RECT 364.950 178.950 367.050 181.050 ;
        RECT 352.950 175.950 355.050 178.050 ;
        RECT 359.400 177.900 360.600 178.950 ;
        RECT 365.400 177.900 366.600 178.950 ;
        RECT 349.950 163.950 352.050 166.050 ;
        RECT 349.950 160.800 352.050 162.900 ;
        RECT 343.950 138.600 346.050 139.050 ;
        RECT 341.400 137.400 346.050 138.600 ;
        RECT 335.400 136.050 336.600 137.100 ;
        RECT 341.400 136.050 342.600 137.400 ;
        RECT 343.950 136.950 346.050 137.400 ;
        RECT 350.400 136.050 351.600 160.800 ;
        RECT 353.400 157.050 354.600 175.950 ;
        RECT 358.950 175.800 361.050 177.900 ;
        RECT 364.950 175.800 367.050 177.900 ;
        RECT 371.400 177.600 372.600 185.400 ;
        RECT 376.950 183.000 379.050 187.050 ;
        RECT 377.400 181.050 378.600 183.000 ;
        RECT 382.950 182.100 385.050 184.200 ;
        RECT 383.400 181.050 384.600 182.100 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 382.950 178.950 385.050 181.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 368.400 176.400 372.600 177.600 ;
        RECT 380.400 177.000 381.600 178.950 ;
        RECT 386.400 177.000 387.600 178.950 ;
        RECT 392.400 177.600 393.600 202.950 ;
        RECT 398.400 196.050 399.600 211.950 ;
        RECT 410.400 205.050 411.600 250.650 ;
        RECT 422.400 247.050 423.600 253.800 ;
        RECT 421.950 244.950 424.050 247.050 ;
        RECT 431.400 232.050 432.600 256.950 ;
        RECT 433.950 253.800 436.050 255.900 ;
        RECT 430.950 229.950 433.050 232.050 ;
        RECT 412.950 215.100 415.050 217.200 ;
        RECT 418.950 215.100 421.050 217.200 ;
        RECT 424.950 216.000 427.050 220.050 ;
        RECT 413.400 208.050 414.600 215.100 ;
        RECT 419.400 214.050 420.600 215.100 ;
        RECT 425.400 214.050 426.600 216.000 ;
        RECT 418.950 211.950 421.050 214.050 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 424.950 211.950 427.050 214.050 ;
        RECT 427.950 211.950 430.050 214.050 ;
        RECT 412.950 205.950 415.050 208.050 ;
        RECT 418.950 205.950 421.050 208.050 ;
        RECT 409.950 202.950 412.050 205.050 ;
        RECT 411.000 201.600 415.050 202.050 ;
        RECT 410.400 199.950 415.050 201.600 ;
        RECT 400.950 196.950 403.050 199.050 ;
        RECT 397.950 193.950 400.050 196.050 ;
        RECT 394.950 181.950 397.050 184.050 ;
        RECT 352.950 154.950 355.050 157.050 ;
        RECT 368.400 154.050 369.600 176.400 ;
        RECT 379.950 172.950 382.050 177.000 ;
        RECT 385.950 172.950 388.050 177.000 ;
        RECT 389.400 176.400 393.600 177.600 ;
        RECT 376.950 157.950 379.050 160.050 ;
        RECT 367.950 151.950 370.050 154.050 ;
        RECT 367.950 142.950 370.050 145.050 ;
        RECT 358.950 137.100 361.050 139.200 ;
        RECT 359.400 136.050 360.600 137.100 ;
        RECT 364.950 136.950 367.050 139.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 349.950 133.950 352.050 136.050 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 338.400 124.050 339.600 133.950 ;
        RECT 356.400 132.900 357.600 133.950 ;
        RECT 355.950 130.800 358.050 132.900 ;
        RECT 337.950 121.950 340.050 124.050 ;
        RECT 328.950 115.950 331.050 118.050 ;
        RECT 338.400 112.050 339.600 121.950 ;
        RECT 358.950 118.950 361.050 121.050 ;
        RECT 355.950 112.950 358.050 115.050 ;
        RECT 328.950 109.950 331.050 112.050 ;
        RECT 337.950 109.950 340.050 112.050 ;
        RECT 343.950 109.950 346.050 112.050 ;
        RECT 352.950 109.950 355.050 112.050 ;
        RECT 313.950 100.950 316.050 103.050 ;
        RECT 316.950 100.950 319.050 103.050 ;
        RECT 319.950 100.950 322.050 103.050 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 314.400 99.000 315.600 100.950 ;
        RECT 313.950 94.950 316.050 99.000 ;
        RECT 320.400 91.050 321.600 100.950 ;
        RECT 325.950 97.950 328.050 100.050 ;
        RECT 319.950 88.950 322.050 91.050 ;
        RECT 307.950 59.100 310.050 61.200 ;
        RECT 316.950 60.000 319.050 64.050 ;
        RECT 326.400 60.600 327.600 97.950 ;
        RECT 329.400 97.050 330.600 109.950 ;
        RECT 331.950 106.950 334.050 109.050 ;
        RECT 332.400 99.900 333.600 106.950 ;
        RECT 334.950 105.600 339.000 106.050 ;
        RECT 334.950 103.950 339.600 105.600 ;
        RECT 338.400 103.050 339.600 103.950 ;
        RECT 344.400 103.050 345.600 109.950 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 340.950 100.950 343.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 341.400 99.900 342.600 100.950 ;
        RECT 347.400 99.900 348.600 100.950 ;
        RECT 331.950 97.800 334.050 99.900 ;
        RECT 340.950 97.800 343.050 99.900 ;
        RECT 346.950 97.800 349.050 99.900 ;
        RECT 328.950 94.950 331.050 97.050 ;
        RECT 340.950 82.950 343.050 85.050 ;
        RECT 341.400 64.050 342.600 82.950 ;
        RECT 353.400 82.050 354.600 109.950 ;
        RECT 356.400 106.050 357.600 112.950 ;
        RECT 355.950 103.950 358.050 106.050 ;
        RECT 359.400 103.050 360.600 118.950 ;
        RECT 365.400 117.600 366.600 136.950 ;
        RECT 368.400 133.050 369.600 142.950 ;
        RECT 377.400 136.050 378.600 157.950 ;
        RECT 382.950 145.950 385.050 148.050 ;
        RECT 379.950 139.950 382.050 145.050 ;
        RECT 383.400 139.200 384.600 145.950 ;
        RECT 382.950 137.100 385.050 139.200 ;
        RECT 383.400 136.050 384.600 137.100 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 382.950 133.950 385.050 136.050 ;
        RECT 367.950 130.950 370.050 133.050 ;
        RECT 370.950 121.950 373.050 124.050 ;
        RECT 362.400 116.400 366.600 117.600 ;
        RECT 362.400 109.050 363.600 116.400 ;
        RECT 364.950 109.950 367.050 112.050 ;
        RECT 361.950 106.950 364.050 109.050 ;
        RECT 365.400 103.050 366.600 109.950 ;
        RECT 371.400 106.050 372.600 121.950 ;
        RECT 370.950 103.950 373.050 106.050 ;
        RECT 358.950 100.950 361.050 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 362.400 94.050 363.600 100.950 ;
        RECT 368.400 99.900 369.600 100.950 ;
        RECT 367.950 97.800 370.050 99.900 ;
        RECT 374.400 94.050 375.600 133.950 ;
        RECT 380.400 132.900 381.600 133.950 ;
        RECT 379.950 130.800 382.050 132.900 ;
        RECT 389.400 130.050 390.600 176.400 ;
        RECT 395.400 160.050 396.600 181.950 ;
        RECT 401.400 181.050 402.600 196.950 ;
        RECT 406.950 183.000 409.050 187.050 ;
        RECT 410.400 184.050 411.600 199.950 ;
        RECT 419.400 196.050 420.600 205.950 ;
        RECT 422.400 202.050 423.600 211.950 ;
        RECT 428.400 202.050 429.600 211.950 ;
        RECT 430.950 208.950 433.050 211.050 ;
        RECT 421.950 199.950 424.050 202.050 ;
        RECT 427.950 199.950 430.050 202.050 ;
        RECT 412.950 193.950 415.050 196.050 ;
        RECT 418.950 193.950 421.050 196.050 ;
        RECT 407.400 181.050 408.600 183.000 ;
        RECT 409.950 181.950 412.050 184.050 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 394.950 157.950 397.050 160.050 ;
        RECT 400.950 157.950 403.050 160.050 ;
        RECT 394.950 138.000 397.050 142.050 ;
        RECT 395.400 136.050 396.600 138.000 ;
        RECT 401.400 136.050 402.600 157.950 ;
        RECT 404.400 148.050 405.600 178.950 ;
        RECT 413.400 175.050 414.600 193.950 ;
        RECT 415.950 190.950 418.050 193.050 ;
        RECT 412.950 172.950 415.050 175.050 ;
        RECT 403.950 145.950 406.050 148.050 ;
        RECT 394.950 133.950 397.050 136.050 ;
        RECT 397.950 133.950 400.050 136.050 ;
        RECT 400.950 133.950 403.050 136.050 ;
        RECT 403.950 133.950 406.050 136.050 ;
        RECT 398.400 132.900 399.600 133.950 ;
        RECT 397.950 130.800 400.050 132.900 ;
        RECT 388.950 127.950 391.050 130.050 ;
        RECT 394.950 127.950 397.050 130.050 ;
        RECT 382.950 112.950 385.050 115.050 ;
        RECT 383.400 103.050 384.600 112.950 ;
        RECT 388.950 104.100 391.050 106.200 ;
        RECT 389.400 103.050 390.600 104.100 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 380.400 99.900 381.600 100.950 ;
        RECT 379.950 97.800 382.050 99.900 ;
        RECT 361.950 91.950 364.050 94.050 ;
        RECT 373.950 91.950 376.050 94.050 ;
        RECT 386.400 82.050 387.600 100.950 ;
        RECT 352.950 79.950 355.050 82.050 ;
        RECT 385.950 79.950 388.050 82.050 ;
        RECT 353.400 73.050 354.600 79.950 ;
        RECT 352.950 70.950 355.050 73.050 ;
        RECT 355.950 64.950 358.050 67.050 ;
        RECT 367.950 64.950 370.050 67.050 ;
        RECT 391.950 64.950 394.050 67.050 ;
        RECT 317.400 58.050 318.600 60.000 ;
        RECT 323.400 59.400 330.600 60.600 ;
        RECT 323.400 58.050 324.600 59.400 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 319.950 55.950 322.050 58.050 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 314.400 54.900 315.600 55.950 ;
        RECT 320.400 54.900 321.600 55.950 ;
        RECT 329.400 54.900 330.600 59.400 ;
        RECT 331.950 58.950 334.050 64.050 ;
        RECT 334.950 59.100 337.050 61.200 ;
        RECT 340.950 60.000 343.050 64.050 ;
        RECT 335.400 58.050 336.600 59.100 ;
        RECT 341.400 58.050 342.600 60.000 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 343.950 55.950 346.050 58.050 ;
        RECT 338.400 54.900 339.600 55.950 ;
        RECT 344.400 54.900 345.600 55.950 ;
        RECT 356.400 55.050 357.600 64.950 ;
        RECT 361.950 59.100 364.050 61.200 ;
        RECT 362.400 58.050 363.600 59.100 ;
        RECT 368.400 58.050 369.600 64.950 ;
        RECT 385.950 59.100 388.050 61.200 ;
        RECT 386.400 58.050 387.600 59.100 ;
        RECT 361.950 55.950 364.050 58.050 ;
        RECT 364.950 55.950 367.050 58.050 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 382.950 55.950 385.050 58.050 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 313.950 52.800 316.050 54.900 ;
        RECT 319.950 52.800 322.050 54.900 ;
        RECT 325.800 54.000 327.900 54.900 ;
        RECT 325.800 52.800 328.050 54.000 ;
        RECT 328.950 52.800 331.050 54.900 ;
        RECT 337.950 52.800 340.050 54.900 ;
        RECT 343.950 52.800 346.050 54.900 ;
        RECT 355.950 52.950 358.050 55.050 ;
        RECT 304.950 49.950 307.050 52.050 ;
        RECT 325.950 49.950 328.050 52.800 ;
        RECT 299.400 47.400 304.050 49.050 ;
        RECT 300.000 46.950 304.050 47.400 ;
        RECT 307.950 46.950 313.050 49.050 ;
        RECT 259.950 43.950 262.050 46.050 ;
        RECT 262.950 43.950 268.050 46.050 ;
        RECT 256.950 40.950 259.050 43.050 ;
        RECT 250.950 34.950 253.050 37.050 ;
        RECT 244.950 31.950 247.050 34.050 ;
        RECT 253.950 31.950 256.050 34.050 ;
        RECT 247.950 28.950 250.050 31.050 ;
        RECT 241.950 25.950 244.050 28.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 233.400 21.900 234.600 22.950 ;
        RECT 226.950 19.800 229.050 21.900 ;
        RECT 232.950 19.800 235.050 21.900 ;
        RECT 239.400 16.050 240.600 22.950 ;
        RECT 248.400 16.050 249.600 28.950 ;
        RECT 254.400 25.050 255.600 31.950 ;
        RECT 260.400 28.200 261.600 43.950 ;
        RECT 298.950 40.950 301.050 43.050 ;
        RECT 299.400 34.050 300.600 40.950 ;
        RECT 301.950 37.950 304.050 40.050 ;
        RECT 316.950 37.950 319.050 40.050 ;
        RECT 268.950 31.950 271.050 34.050 ;
        RECT 298.950 31.950 301.050 34.050 ;
        RECT 259.950 26.100 262.050 28.200 ;
        RECT 260.400 25.050 261.600 26.100 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 257.400 21.900 258.600 22.950 ;
        RECT 256.950 19.800 259.050 21.900 ;
        RECT 263.400 21.000 264.600 22.950 ;
        RECT 238.950 13.950 241.050 16.050 ;
        RECT 247.950 13.950 250.050 16.050 ;
        RECT 223.950 10.950 226.050 13.050 ;
        RECT 257.400 10.050 258.600 19.800 ;
        RECT 262.950 16.950 265.050 21.000 ;
        RECT 269.400 13.050 270.600 31.950 ;
        RECT 292.950 28.950 295.050 31.050 ;
        RECT 277.950 26.100 280.050 28.200 ;
        RECT 283.950 26.100 286.050 28.200 ;
        RECT 278.400 25.050 279.600 26.100 ;
        RECT 284.400 25.050 285.600 26.100 ;
        RECT 289.950 25.950 292.050 28.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 283.950 22.950 286.050 25.050 ;
        RECT 275.400 21.900 276.600 22.950 ;
        RECT 281.400 21.900 282.600 22.950 ;
        RECT 274.950 19.800 277.050 21.900 ;
        RECT 280.950 16.950 283.050 21.900 ;
        RECT 290.400 16.050 291.600 25.950 ;
        RECT 293.400 21.900 294.600 28.950 ;
        RECT 302.400 25.050 303.600 37.950 ;
        RECT 313.950 31.950 316.050 34.050 ;
        RECT 307.950 26.100 310.050 28.200 ;
        RECT 308.400 25.050 309.600 26.100 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 304.950 22.950 307.050 25.050 ;
        RECT 307.950 22.950 310.050 25.050 ;
        RECT 299.400 21.900 300.600 22.950 ;
        RECT 305.400 21.900 306.600 22.950 ;
        RECT 314.400 22.050 315.600 31.950 ;
        RECT 292.950 19.800 295.050 21.900 ;
        RECT 298.950 19.800 301.050 21.900 ;
        RECT 304.950 19.800 307.050 21.900 ;
        RECT 310.950 16.950 313.050 21.900 ;
        RECT 313.950 19.950 316.050 22.050 ;
        RECT 317.400 21.900 318.600 37.950 ;
        RECT 365.400 37.050 366.600 55.950 ;
        RECT 371.400 54.900 372.600 55.950 ;
        RECT 383.400 54.900 384.600 55.950 ;
        RECT 392.400 55.050 393.600 64.950 ;
        RECT 370.950 52.800 373.050 54.900 ;
        RECT 382.950 52.800 385.050 54.900 ;
        RECT 391.950 52.950 394.050 55.050 ;
        RECT 388.950 40.950 391.050 43.050 ;
        RECT 382.950 37.950 385.050 40.050 ;
        RECT 337.950 34.950 340.050 37.050 ;
        RECT 364.950 34.950 367.050 37.050 ;
        RECT 331.950 31.950 334.050 34.050 ;
        RECT 325.950 27.000 328.050 31.050 ;
        RECT 326.400 25.050 327.600 27.000 ;
        RECT 332.400 25.050 333.600 31.950 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 325.950 22.950 328.050 25.050 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 331.950 22.950 334.050 25.050 ;
        RECT 316.950 19.800 319.050 21.900 ;
        RECT 319.950 19.950 322.050 22.050 ;
        RECT 323.400 21.900 324.600 22.950 ;
        RECT 329.400 21.900 330.600 22.950 ;
        RECT 338.400 21.900 339.600 34.950 ;
        RECT 361.950 33.600 364.050 34.050 ;
        RECT 367.950 33.600 370.050 34.050 ;
        RECT 361.950 32.400 370.050 33.600 ;
        RECT 361.950 31.950 364.050 32.400 ;
        RECT 367.950 31.950 370.050 32.400 ;
        RECT 343.950 26.100 346.050 28.200 ;
        RECT 352.950 26.100 355.050 28.200 ;
        RECT 364.950 27.000 367.050 31.050 ;
        RECT 344.400 25.050 345.600 26.100 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 347.400 21.900 348.600 22.950 ;
        RECT 289.950 13.950 292.050 16.050 ;
        RECT 268.950 10.950 271.050 13.050 ;
        RECT 256.950 7.950 259.050 10.050 ;
        RECT 320.400 7.050 321.600 19.950 ;
        RECT 322.950 19.800 325.050 21.900 ;
        RECT 328.950 16.950 331.050 21.900 ;
        RECT 337.950 19.800 340.050 21.900 ;
        RECT 346.950 19.800 349.050 21.900 ;
        RECT 353.400 16.050 354.600 26.100 ;
        RECT 365.400 25.050 366.600 27.000 ;
        RECT 370.950 26.100 373.050 28.200 ;
        RECT 379.950 26.100 382.050 28.200 ;
        RECT 383.400 28.050 384.600 37.950 ;
        RECT 371.400 25.050 372.600 26.100 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 367.950 22.950 370.050 25.050 ;
        RECT 370.950 22.950 373.050 25.050 ;
        RECT 373.950 22.950 376.050 25.050 ;
        RECT 361.950 16.950 364.050 19.050 ;
        RECT 352.950 13.950 355.050 16.050 ;
        RECT 362.400 10.050 363.600 16.950 ;
        RECT 368.400 16.050 369.600 22.950 ;
        RECT 374.400 22.050 375.600 22.950 ;
        RECT 374.400 20.400 379.050 22.050 ;
        RECT 375.000 19.950 379.050 20.400 ;
        RECT 380.400 19.050 381.600 26.100 ;
        RECT 382.950 25.950 385.050 28.050 ;
        RECT 389.400 25.050 390.600 40.950 ;
        RECT 395.400 31.050 396.600 127.950 ;
        RECT 397.950 118.950 400.050 121.050 ;
        RECT 398.400 85.050 399.600 118.950 ;
        RECT 404.400 115.050 405.600 133.950 ;
        RECT 413.400 132.900 414.600 172.950 ;
        RECT 416.400 138.600 417.600 190.950 ;
        RECT 427.950 189.600 430.050 190.050 ;
        RECT 431.400 189.600 432.600 208.950 ;
        RECT 434.400 208.050 435.600 253.800 ;
        RECT 437.400 241.050 438.600 274.950 ;
        RECT 449.400 268.050 450.600 283.950 ;
        RECT 452.400 277.050 453.600 293.100 ;
        RECT 461.400 292.050 462.600 293.100 ;
        RECT 467.400 292.050 468.600 293.400 ;
        RECT 457.950 289.950 460.050 292.050 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 463.950 289.950 466.050 292.050 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 458.400 286.050 459.600 289.950 ;
        RECT 454.950 284.400 459.600 286.050 ;
        RECT 454.950 283.950 459.000 284.400 ;
        RECT 454.950 277.950 457.050 280.050 ;
        RECT 451.950 274.950 454.050 277.050 ;
        RECT 448.950 265.950 451.050 268.050 ;
        RECT 439.950 259.950 442.050 262.050 ;
        RECT 440.400 247.050 441.600 259.950 ;
        RECT 449.400 259.050 450.600 265.950 ;
        RECT 445.950 256.950 448.050 259.050 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 439.950 244.950 442.050 247.050 ;
        RECT 436.950 238.950 439.050 241.050 ;
        RECT 446.400 235.050 447.600 256.950 ;
        RECT 445.950 232.950 448.050 235.050 ;
        RECT 436.950 216.600 441.000 217.050 ;
        RECT 436.950 214.950 441.600 216.600 ;
        RECT 445.950 216.000 448.050 220.050 ;
        RECT 455.400 217.050 456.600 277.950 ;
        RECT 460.950 268.950 463.050 271.050 ;
        RECT 461.400 259.050 462.600 268.950 ;
        RECT 464.400 265.050 465.600 289.950 ;
        RECT 473.400 289.050 474.600 293.400 ;
        RECT 472.950 286.950 475.050 289.050 ;
        RECT 466.950 280.950 469.050 283.050 ;
        RECT 472.950 280.950 475.050 283.050 ;
        RECT 467.400 268.050 468.600 280.950 ;
        RECT 466.950 265.950 469.050 268.050 ;
        RECT 463.950 262.950 466.050 265.050 ;
        RECT 467.400 259.050 468.600 265.950 ;
        RECT 460.950 256.950 463.050 259.050 ;
        RECT 463.950 256.950 466.050 259.050 ;
        RECT 466.950 256.950 469.050 259.050 ;
        RECT 464.400 255.900 465.600 256.950 ;
        RECT 463.950 253.800 466.050 255.900 ;
        RECT 473.400 250.050 474.600 280.950 ;
        RECT 472.950 247.950 475.050 250.050 ;
        RECT 460.950 241.950 463.050 244.050 ;
        RECT 461.400 220.050 462.600 241.950 ;
        RECT 440.400 214.050 441.600 214.950 ;
        RECT 446.400 214.050 447.600 216.000 ;
        RECT 454.950 214.950 457.050 217.050 ;
        RECT 460.950 216.000 463.050 220.050 ;
        RECT 461.400 214.050 462.600 216.000 ;
        RECT 466.950 215.100 469.050 217.200 ;
        RECT 472.800 215.100 474.900 217.200 ;
        RECT 476.400 217.050 477.600 325.950 ;
        RECT 487.950 322.950 490.050 325.050 ;
        RECT 481.950 301.950 484.050 304.050 ;
        RECT 482.400 292.050 483.600 301.950 ;
        RECT 488.400 295.200 489.600 322.950 ;
        RECT 509.400 310.050 510.600 338.100 ;
        RECT 508.950 307.950 511.050 310.050 ;
        RECT 512.400 301.050 513.600 340.950 ;
        RECT 521.400 340.050 522.600 364.950 ;
        RECT 524.400 343.050 525.600 373.950 ;
        RECT 535.950 371.100 538.050 373.200 ;
        RECT 536.400 370.050 537.600 371.100 ;
        RECT 542.400 370.050 543.600 400.950 ;
        RECT 545.400 397.050 546.600 412.950 ;
        RECT 544.950 394.950 547.050 397.050 ;
        RECT 547.950 373.950 550.050 376.050 ;
        RECT 526.950 367.950 529.050 370.050 ;
        RECT 532.950 367.950 535.050 370.050 ;
        RECT 535.950 367.950 538.050 370.050 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 527.400 364.050 528.600 367.950 ;
        RECT 526.950 361.950 529.050 364.050 ;
        RECT 533.400 361.050 534.600 367.950 ;
        RECT 532.950 358.950 535.050 361.050 ;
        RECT 526.950 346.950 529.050 349.050 ;
        RECT 523.950 340.950 526.050 343.050 ;
        RECT 520.950 337.950 523.050 340.050 ;
        RECT 527.400 339.600 528.600 346.950 ;
        RECT 529.950 343.950 532.050 346.050 ;
        RECT 524.400 338.400 528.600 339.600 ;
        RECT 524.400 337.050 525.600 338.400 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 518.400 313.050 519.600 334.950 ;
        RECT 526.950 331.950 529.050 334.050 ;
        RECT 517.950 310.950 520.050 313.050 ;
        RECT 518.400 303.600 519.600 310.950 ;
        RECT 518.400 302.400 522.600 303.600 ;
        RECT 502.800 298.950 504.900 301.050 ;
        RECT 505.950 298.950 508.050 301.050 ;
        RECT 511.950 298.950 514.050 301.050 ;
        RECT 517.950 298.950 520.050 301.050 ;
        RECT 503.400 295.200 504.600 298.950 ;
        RECT 487.950 293.100 490.050 295.200 ;
        RECT 493.950 293.100 496.050 295.200 ;
        RECT 502.950 293.100 505.050 295.200 ;
        RECT 488.400 292.050 489.600 293.100 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 487.950 289.950 490.050 292.050 ;
        RECT 485.400 288.900 486.600 289.950 ;
        RECT 478.950 286.800 481.050 288.900 ;
        RECT 484.950 286.800 487.050 288.900 ;
        RECT 479.400 220.050 480.600 286.800 ;
        RECT 494.400 286.050 495.600 293.100 ;
        RECT 506.400 292.050 507.600 298.950 ;
        RECT 511.950 293.100 514.050 295.200 ;
        RECT 512.400 292.050 513.600 293.100 ;
        RECT 505.950 289.950 508.050 292.050 ;
        RECT 508.950 289.950 511.050 292.050 ;
        RECT 511.950 289.950 514.050 292.050 ;
        RECT 493.950 283.950 496.050 286.050 ;
        RECT 494.400 280.050 495.600 283.950 ;
        RECT 493.950 277.950 496.050 280.050 ;
        RECT 509.400 274.050 510.600 289.950 ;
        RECT 508.950 271.950 511.050 274.050 ;
        RECT 499.950 268.950 502.050 271.050 ;
        RECT 487.950 265.950 490.050 268.050 ;
        RECT 488.400 262.200 489.600 265.950 ;
        RECT 487.950 260.100 490.050 262.200 ;
        RECT 488.400 259.050 489.600 260.100 ;
        RECT 484.950 256.950 487.050 259.050 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 493.950 256.950 496.050 259.050 ;
        RECT 485.400 244.050 486.600 256.950 ;
        RECT 494.400 255.900 495.600 256.950 ;
        RECT 500.400 256.050 501.600 268.950 ;
        RECT 508.950 260.100 511.050 262.200 ;
        RECT 518.400 262.050 519.600 298.950 ;
        RECT 509.400 259.050 510.600 260.100 ;
        RECT 517.950 259.950 520.050 262.050 ;
        RECT 505.950 256.950 508.050 259.050 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 514.950 256.950 517.050 259.050 ;
        RECT 493.950 253.800 496.050 255.900 ;
        RECT 499.950 253.950 502.050 256.050 ;
        RECT 506.400 255.900 507.600 256.950 ;
        RECT 505.950 253.800 508.050 255.900 ;
        RECT 511.950 253.950 514.050 256.050 ;
        RECT 499.950 250.800 502.050 252.900 ;
        RECT 484.950 241.950 487.050 244.050 ;
        RECT 487.950 238.950 490.050 241.050 ;
        RECT 488.400 226.050 489.600 238.950 ;
        RECT 490.950 226.950 493.050 229.050 ;
        RECT 487.950 223.950 490.050 226.050 ;
        RECT 467.400 214.050 468.600 215.100 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 442.950 211.950 445.050 214.050 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 448.950 211.950 451.050 214.050 ;
        RECT 457.950 211.950 460.050 214.050 ;
        RECT 460.950 211.950 463.050 214.050 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 436.950 208.950 439.050 211.050 ;
        RECT 443.400 210.900 444.600 211.950 ;
        RECT 449.400 210.900 450.600 211.950 ;
        RECT 458.400 210.900 459.600 211.950 ;
        RECT 433.950 205.950 436.050 208.050 ;
        RECT 427.950 188.400 432.600 189.600 ;
        RECT 427.950 187.950 430.050 188.400 ;
        RECT 421.950 182.100 424.050 184.200 ;
        RECT 422.400 181.050 423.600 182.100 ;
        RECT 428.400 181.050 429.600 187.950 ;
        RECT 437.400 184.200 438.600 208.950 ;
        RECT 442.950 208.800 445.050 210.900 ;
        RECT 448.950 210.600 451.050 210.900 ;
        RECT 448.950 209.400 453.600 210.600 ;
        RECT 448.950 205.950 451.050 209.400 ;
        RECT 442.950 199.950 445.050 202.050 ;
        RECT 436.950 182.100 439.050 184.200 ;
        RECT 421.950 178.950 424.050 181.050 ;
        RECT 424.950 178.950 427.050 181.050 ;
        RECT 427.950 178.950 430.050 181.050 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 418.950 175.950 421.050 178.050 ;
        RECT 425.400 177.000 426.600 178.950 ;
        RECT 431.400 177.900 432.600 178.950 ;
        RECT 437.400 177.900 438.600 182.100 ;
        RECT 443.400 181.050 444.600 199.950 ;
        RECT 442.950 178.950 445.050 181.050 ;
        RECT 445.950 178.950 448.050 181.050 ;
        RECT 446.400 177.900 447.600 178.950 ;
        RECT 419.400 154.050 420.600 175.950 ;
        RECT 424.950 172.950 427.050 177.000 ;
        RECT 430.950 175.800 433.050 177.900 ;
        RECT 436.950 175.800 439.050 177.900 ;
        RECT 445.950 175.800 448.050 177.900 ;
        RECT 452.400 175.050 453.600 209.400 ;
        RECT 457.950 208.800 460.050 210.900 ;
        RECT 464.400 205.050 465.600 211.950 ;
        RECT 463.950 202.950 466.050 205.050 ;
        RECT 469.950 202.950 472.050 205.050 ;
        RECT 463.950 193.950 466.050 196.050 ;
        RECT 454.950 187.950 457.050 190.050 ;
        RECT 455.400 184.050 456.600 187.950 ;
        RECT 464.400 187.050 465.600 193.950 ;
        RECT 463.950 184.950 466.050 187.050 ;
        RECT 454.950 181.950 457.050 184.050 ;
        RECT 460.950 182.100 463.050 184.200 ;
        RECT 466.950 182.100 469.050 184.200 ;
        RECT 470.400 183.600 471.600 202.950 ;
        RECT 473.400 202.050 474.600 215.100 ;
        RECT 475.950 214.950 478.050 217.050 ;
        RECT 478.950 216.000 481.050 220.050 ;
        RECT 479.400 214.050 480.600 216.000 ;
        RECT 487.950 215.100 490.050 217.200 ;
        RECT 491.400 217.050 492.600 226.950 ;
        RECT 493.950 217.950 496.050 220.050 ;
        RECT 488.400 214.050 489.600 215.100 ;
        RECT 490.950 214.950 493.050 217.050 ;
        RECT 478.950 211.950 481.050 214.050 ;
        RECT 484.950 211.950 487.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 475.950 208.950 478.050 211.050 ;
        RECT 481.800 208.950 483.900 211.050 ;
        RECT 485.400 210.900 486.600 211.950 ;
        RECT 494.400 211.050 495.600 217.950 ;
        RECT 496.800 215.100 498.900 217.200 ;
        RECT 500.400 217.050 501.600 250.800 ;
        RECT 512.400 235.050 513.600 253.950 ;
        RECT 515.400 246.600 516.600 256.950 ;
        RECT 521.400 255.900 522.600 302.400 ;
        RECT 527.400 301.050 528.600 331.950 ;
        RECT 530.400 331.050 531.600 343.950 ;
        RECT 539.400 343.050 540.600 367.950 ;
        RECT 548.400 352.050 549.600 373.950 ;
        RECT 551.400 367.050 552.600 412.950 ;
        RECT 557.400 372.600 558.600 415.950 ;
        RECT 560.400 376.200 561.600 427.950 ;
        RECT 562.950 421.950 565.050 424.050 ;
        RECT 563.400 403.050 564.600 421.950 ;
        RECT 566.400 418.050 567.600 430.950 ;
        RECT 565.950 415.950 568.050 418.050 ;
        RECT 571.950 416.100 574.050 418.200 ;
        RECT 572.400 415.050 573.600 416.100 ;
        RECT 568.950 412.950 571.050 415.050 ;
        RECT 571.950 412.950 574.050 415.050 ;
        RECT 569.400 411.900 570.600 412.950 ;
        RECT 568.950 409.800 571.050 411.900 ;
        RECT 574.950 409.800 577.050 411.900 ;
        RECT 562.950 400.950 565.050 403.050 ;
        RECT 562.950 388.950 565.050 391.050 ;
        RECT 563.400 382.050 564.600 388.950 ;
        RECT 565.950 382.950 568.050 385.050 ;
        RECT 562.950 379.950 565.050 382.050 ;
        RECT 559.950 374.100 562.050 376.200 ;
        RECT 554.400 371.400 558.600 372.600 ;
        RECT 550.950 364.950 553.050 367.050 ;
        RECT 541.950 349.950 544.050 352.050 ;
        RECT 547.950 349.950 550.050 352.050 ;
        RECT 554.400 351.600 555.600 371.400 ;
        RECT 559.950 370.950 562.050 373.050 ;
        RECT 560.400 370.050 561.600 370.950 ;
        RECT 566.400 370.050 567.600 382.950 ;
        RECT 575.400 373.050 576.600 409.800 ;
        RECT 578.400 406.050 579.600 443.400 ;
        RECT 587.100 438.600 588.300 458.400 ;
        RECT 598.950 457.950 601.050 460.050 ;
        RECT 589.950 449.400 592.050 451.500 ;
        RECT 595.950 449.400 598.050 451.500 ;
        RECT 590.400 448.050 591.600 449.400 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 586.950 436.500 589.050 438.600 ;
        RECT 589.950 421.950 592.050 424.050 ;
        RECT 580.950 416.100 583.050 418.200 ;
        RECT 581.400 412.050 582.600 416.100 ;
        RECT 590.400 415.050 591.600 421.950 ;
        RECT 596.400 421.050 597.600 449.400 ;
        RECT 599.400 445.050 600.600 457.950 ;
        RECT 602.400 451.050 603.600 463.950 ;
        RECT 601.950 448.950 604.050 451.050 ;
        RECT 604.950 449.100 607.050 451.200 ;
        RECT 610.950 449.100 613.050 451.200 ;
        RECT 614.400 451.050 615.600 496.950 ;
        RECT 644.400 496.200 645.600 523.950 ;
        RECT 650.400 522.600 651.600 544.950 ;
        RECT 656.400 538.050 657.600 610.950 ;
        RECT 659.400 607.050 660.600 652.950 ;
        RECT 662.400 613.050 663.600 712.950 ;
        RECT 671.400 691.050 672.600 712.950 ;
        RECT 673.800 706.950 675.900 709.050 ;
        RECT 674.400 700.050 675.600 706.950 ;
        RECT 673.950 697.950 676.050 700.050 ;
        RECT 667.800 688.950 669.900 691.050 ;
        RECT 670.950 688.950 673.050 691.050 ;
        RECT 668.400 685.200 669.600 688.950 ;
        RECT 667.950 683.100 670.050 685.200 ;
        RECT 668.400 682.050 669.600 683.100 ;
        RECT 674.400 682.050 675.600 697.950 ;
        RECT 680.400 694.050 681.600 712.950 ;
        RECT 679.950 691.950 682.050 694.050 ;
        RECT 667.950 679.950 670.050 682.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 673.950 679.950 676.050 682.050 ;
        RECT 676.950 679.950 679.050 682.050 ;
        RECT 671.400 664.050 672.600 679.950 ;
        RECT 677.400 678.600 678.600 679.950 ;
        RECT 677.400 677.400 681.600 678.600 ;
        RECT 673.950 667.950 676.050 670.050 ;
        RECT 670.950 661.950 673.050 664.050 ;
        RECT 667.950 658.950 670.050 661.050 ;
        RECT 668.400 652.050 669.600 658.950 ;
        RECT 664.950 649.950 669.600 652.050 ;
        RECT 668.400 649.050 669.600 649.950 ;
        RECT 674.400 649.050 675.600 667.950 ;
        RECT 676.950 664.950 679.050 667.050 ;
        RECT 677.400 658.050 678.600 664.950 ;
        RECT 680.400 658.050 681.600 677.400 ;
        RECT 676.800 655.950 678.900 658.050 ;
        RECT 679.950 655.950 682.050 658.050 ;
        RECT 683.400 655.050 684.600 718.950 ;
        RECT 686.400 718.050 687.600 724.950 ;
        RECT 685.950 715.950 688.050 718.050 ;
        RECT 692.400 703.050 693.600 724.950 ;
        RECT 698.400 715.050 699.600 733.950 ;
        RECT 704.400 733.050 705.600 746.400 ;
        RECT 709.950 745.950 712.050 748.050 ;
        RECT 706.950 742.950 709.050 745.050 ;
        RECT 707.400 733.050 708.600 742.950 ;
        RECT 710.400 742.050 711.600 745.950 ;
        RECT 716.400 742.050 717.600 751.950 ;
        RECT 709.950 739.950 712.050 742.050 ;
        RECT 715.950 739.950 718.050 742.050 ;
        RECT 703.950 730.950 706.050 733.050 ;
        RECT 707.400 731.400 712.050 733.050 ;
        RECT 708.000 730.950 712.050 731.400 ;
        RECT 706.950 728.100 709.050 730.200 ;
        RECT 712.950 728.100 715.050 730.200 ;
        RECT 719.400 730.050 720.600 754.950 ;
        RECT 721.950 754.800 724.050 756.900 ;
        RECT 728.400 751.050 729.600 757.950 ;
        RECT 727.950 748.950 730.050 751.050 ;
        RECT 724.950 745.950 727.050 748.050 ;
        RECT 707.400 727.050 708.600 728.100 ;
        RECT 713.400 727.050 714.600 728.100 ;
        RECT 719.400 727.950 724.050 730.050 ;
        RECT 719.400 727.050 720.600 727.950 ;
        RECT 700.950 724.800 703.050 726.900 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 709.950 724.950 712.050 727.050 ;
        RECT 712.950 724.950 715.050 727.050 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 718.950 724.950 721.050 727.050 ;
        RECT 701.400 718.050 702.600 724.800 ;
        RECT 710.400 720.600 711.600 724.950 ;
        RECT 716.400 723.900 717.600 724.950 ;
        RECT 715.950 721.800 718.050 723.900 ;
        RECT 721.950 721.950 724.050 724.050 ;
        RECT 707.400 719.400 711.600 720.600 ;
        RECT 700.950 715.950 703.050 718.050 ;
        RECT 697.950 712.950 700.050 715.050 ;
        RECT 703.950 706.950 706.050 709.050 ;
        RECT 691.950 700.950 694.050 703.050 ;
        RECT 691.950 697.800 694.050 699.900 ;
        RECT 685.950 688.950 688.050 691.050 ;
        RECT 686.400 685.050 687.600 688.950 ;
        RECT 685.950 682.950 688.050 685.050 ;
        RECT 692.400 682.050 693.600 697.800 ;
        RECT 694.950 691.950 697.050 694.050 ;
        RECT 697.950 691.950 700.050 697.050 ;
        RECT 695.400 688.050 696.600 691.950 ;
        RECT 694.950 685.950 697.050 688.050 ;
        RECT 699.000 684.600 703.050 685.050 ;
        RECT 698.400 682.950 703.050 684.600 ;
        RECT 698.400 682.050 699.600 682.950 ;
        RECT 688.950 679.950 691.050 682.050 ;
        RECT 691.950 679.950 694.050 682.050 ;
        RECT 694.950 679.950 697.050 682.050 ;
        RECT 697.950 679.950 700.050 682.050 ;
        RECT 689.400 679.050 690.600 679.950 ;
        RECT 685.950 677.400 690.600 679.050 ;
        RECT 685.950 676.950 690.000 677.400 ;
        RECT 688.950 673.950 691.050 676.050 ;
        RECT 685.950 670.950 688.050 673.050 ;
        RECT 682.950 652.950 685.050 655.050 ;
        RECT 682.950 649.800 685.050 651.900 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 670.950 646.950 673.050 649.050 ;
        RECT 673.950 646.950 676.050 649.050 ;
        RECT 676.950 646.950 679.050 649.050 ;
        RECT 671.400 637.050 672.600 646.950 ;
        RECT 677.400 645.000 678.600 646.950 ;
        RECT 683.400 646.050 684.600 649.800 ;
        RECT 686.400 646.050 687.600 670.950 ;
        RECT 689.400 667.050 690.600 673.950 ;
        RECT 691.950 670.950 694.050 673.050 ;
        RECT 688.950 664.950 691.050 667.050 ;
        RECT 692.400 664.050 693.600 670.950 ;
        RECT 695.400 667.050 696.600 679.950 ;
        RECT 700.950 676.950 703.050 679.050 ;
        RECT 704.400 678.900 705.600 706.950 ;
        RECT 707.400 706.050 708.600 719.400 ;
        RECT 706.800 703.950 708.900 706.050 ;
        RECT 709.950 703.950 712.050 706.050 ;
        RECT 710.400 694.050 711.600 703.950 ;
        RECT 722.400 703.050 723.600 721.950 ;
        RECT 721.950 700.950 724.050 703.050 ;
        RECT 709.950 691.950 712.050 694.050 ;
        RECT 725.400 693.600 726.600 745.950 ;
        RECT 727.950 729.600 730.050 733.050 ;
        RECT 737.400 730.050 738.600 763.950 ;
        RECT 740.400 736.050 741.600 772.950 ;
        RECT 748.950 757.950 751.050 760.050 ;
        RECT 749.400 756.900 750.600 757.950 ;
        RECT 748.950 754.800 751.050 756.900 ;
        RECT 754.950 754.950 757.050 757.050 ;
        RECT 742.950 745.950 745.050 748.050 ;
        RECT 739.950 733.950 742.050 736.050 ;
        RECT 727.950 729.000 732.600 729.600 ;
        RECT 728.400 728.400 732.600 729.000 ;
        RECT 731.400 727.050 732.600 728.400 ;
        RECT 736.950 727.950 739.050 730.050 ;
        RECT 739.950 727.950 742.050 730.050 ;
        RECT 730.950 724.950 733.050 727.050 ;
        RECT 733.950 724.950 736.050 727.050 ;
        RECT 734.400 723.900 735.600 724.950 ;
        RECT 733.950 721.800 736.050 723.900 ;
        RECT 730.950 715.950 733.050 718.050 ;
        RECT 731.400 703.050 732.600 715.950 ;
        RECT 734.400 715.050 735.600 721.800 ;
        RECT 733.950 712.950 736.050 715.050 ;
        RECT 730.950 700.950 733.050 703.050 ;
        RECT 722.400 693.000 726.600 693.600 ;
        RECT 721.950 692.400 726.600 693.000 ;
        RECT 709.950 688.800 712.050 690.900 ;
        RECT 706.950 685.950 709.050 688.050 ;
        RECT 697.950 673.950 700.050 676.050 ;
        RECT 694.950 664.950 697.050 667.050 ;
        RECT 691.950 661.950 694.050 664.050 ;
        RECT 688.950 652.950 691.050 658.050 ;
        RECT 692.400 651.600 693.600 661.950 ;
        RECT 695.400 661.050 696.600 664.950 ;
        RECT 698.400 664.050 699.600 673.950 ;
        RECT 701.400 673.050 702.600 676.950 ;
        RECT 703.950 676.800 706.050 678.900 ;
        RECT 700.950 670.950 703.050 673.050 ;
        RECT 697.950 661.950 700.050 664.050 ;
        RECT 694.950 658.950 697.050 661.050 ;
        RECT 704.400 655.050 705.600 676.800 ;
        RECT 689.400 650.400 693.600 651.600 ;
        RECT 676.950 640.950 679.050 645.000 ;
        RECT 682.800 643.950 684.900 646.050 ;
        RECT 685.950 643.950 688.050 646.050 ;
        RECT 689.400 643.050 690.600 650.400 ;
        RECT 694.950 650.100 697.050 652.200 ;
        RECT 700.950 650.100 703.050 655.050 ;
        RECT 703.950 652.950 706.050 655.050 ;
        RECT 707.400 652.050 708.600 685.950 ;
        RECT 710.400 682.050 711.600 688.800 ;
        RECT 715.800 687.300 717.900 689.400 ;
        RECT 721.950 688.950 724.050 692.400 ;
        RECT 725.400 688.500 727.500 690.600 ;
        RECT 713.400 682.050 714.600 684.600 ;
        RECT 709.950 679.950 712.050 682.050 ;
        RECT 713.400 679.950 715.500 682.050 ;
        RECT 710.400 664.050 711.600 679.950 ;
        RECT 716.700 678.300 717.600 687.300 ;
        RECT 719.100 683.700 721.200 685.800 ;
        RECT 722.400 684.900 723.600 687.450 ;
        RECT 720.300 681.300 721.200 683.700 ;
        RECT 722.100 682.800 724.200 684.900 ;
        RECT 726.000 681.300 727.050 688.500 ;
        RECT 733.950 685.950 736.050 688.050 ;
        RECT 720.300 680.100 727.050 681.300 ;
        RECT 723.150 678.300 725.250 679.200 ;
        RECT 716.700 677.100 725.250 678.300 ;
        RECT 718.200 675.300 720.300 677.100 ;
        RECT 722.100 674.100 724.200 676.200 ;
        RECT 726.150 674.700 727.050 680.100 ;
        RECT 727.950 679.950 730.050 682.050 ;
        RECT 728.400 677.400 729.600 679.950 ;
        RECT 715.950 670.950 718.050 673.050 ;
        RECT 722.400 672.600 723.600 674.100 ;
        RECT 725.400 672.600 727.500 674.700 ;
        RECT 719.400 671.400 723.600 672.600 ;
        RECT 712.950 667.950 715.050 670.050 ;
        RECT 709.950 661.950 712.050 664.050 ;
        RECT 709.950 658.800 712.050 660.900 ;
        RECT 695.400 649.050 696.600 650.100 ;
        RECT 701.400 649.050 702.600 650.100 ;
        RECT 706.950 649.950 709.050 652.050 ;
        RECT 694.950 646.950 697.050 649.050 ;
        RECT 697.950 646.950 700.050 649.050 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 703.950 646.950 706.050 649.050 ;
        RECT 691.950 643.950 694.050 646.050 ;
        RECT 698.400 645.000 699.600 646.950 ;
        RECT 704.400 645.900 705.600 646.950 ;
        RECT 688.950 640.950 691.050 643.050 ;
        RECT 670.950 634.950 673.050 637.050 ;
        RECT 676.950 631.950 679.050 634.050 ;
        RECT 667.950 616.950 670.050 619.050 ;
        RECT 661.950 610.950 664.050 613.050 ;
        RECT 658.950 604.950 661.050 607.050 ;
        RECT 661.950 606.000 664.050 609.900 ;
        RECT 662.400 604.050 663.600 606.000 ;
        RECT 668.400 604.050 669.600 616.950 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 658.950 598.950 661.050 601.050 ;
        RECT 659.400 565.050 660.600 598.950 ;
        RECT 661.950 589.950 664.050 592.050 ;
        RECT 662.400 574.200 663.600 589.950 ;
        RECT 665.400 586.050 666.600 601.950 ;
        RECT 671.400 600.600 672.600 601.950 ;
        RECT 677.400 600.600 678.600 631.950 ;
        RECT 682.950 616.950 685.050 619.050 ;
        RECT 683.400 604.050 684.600 616.950 ;
        RECT 688.950 605.100 691.050 607.200 ;
        RECT 692.400 607.050 693.600 643.950 ;
        RECT 694.950 640.950 697.050 643.050 ;
        RECT 697.950 640.950 700.050 645.000 ;
        RECT 703.950 643.800 706.050 645.900 ;
        RECT 700.950 640.950 703.050 643.050 ;
        RECT 695.400 622.050 696.600 640.950 ;
        RECT 694.950 619.950 697.050 622.050 ;
        RECT 694.950 616.800 697.050 618.900 ;
        RECT 689.400 604.050 690.600 605.100 ;
        RECT 691.950 604.950 694.050 607.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 686.400 600.900 687.600 601.950 ;
        RECT 671.400 600.000 675.600 600.600 ;
        RECT 671.400 599.400 676.050 600.000 ;
        RECT 677.400 599.400 681.600 600.600 ;
        RECT 673.950 595.950 676.050 599.400 ;
        RECT 664.950 583.950 667.050 586.050 ;
        RECT 661.950 572.100 664.050 574.200 ;
        RECT 673.950 572.100 676.050 574.200 ;
        RECT 658.950 562.950 661.050 565.050 ;
        RECT 662.400 559.050 663.600 572.100 ;
        RECT 674.400 571.050 675.600 572.100 ;
        RECT 667.950 568.950 670.050 571.050 ;
        RECT 673.950 568.950 676.050 571.050 ;
        RECT 668.400 567.000 669.600 568.950 ;
        RECT 680.400 567.600 681.600 599.400 ;
        RECT 685.950 598.800 688.050 600.900 ;
        RECT 691.950 598.950 694.050 601.050 ;
        RECT 682.950 597.600 685.050 598.050 ;
        RECT 682.950 597.000 690.600 597.600 ;
        RECT 682.950 596.400 691.050 597.000 ;
        RECT 682.950 595.950 685.050 596.400 ;
        RECT 682.950 592.800 685.050 594.900 ;
        RECT 688.950 592.950 691.050 596.400 ;
        RECT 683.400 574.050 684.600 592.800 ;
        RECT 692.400 583.050 693.600 598.950 ;
        RECT 695.400 598.050 696.600 616.800 ;
        RECT 698.400 616.050 699.600 640.950 ;
        RECT 701.400 619.050 702.600 640.950 ;
        RECT 710.400 625.050 711.600 658.800 ;
        RECT 713.400 643.050 714.600 667.950 ;
        RECT 716.400 661.050 717.600 670.950 ;
        RECT 715.950 658.950 718.050 661.050 ;
        RECT 719.400 657.600 720.600 671.400 ;
        RECT 721.950 667.950 724.050 670.050 ;
        RECT 722.400 658.050 723.600 667.950 ;
        RECT 716.400 657.000 720.600 657.600 ;
        RECT 715.950 656.400 720.600 657.000 ;
        RECT 715.950 652.950 718.050 656.400 ;
        RECT 721.950 655.950 724.050 658.050 ;
        RECT 734.400 652.200 735.600 685.950 ;
        RECT 740.400 682.050 741.600 727.950 ;
        RECT 743.400 688.050 744.600 745.950 ;
        RECT 748.950 739.950 751.050 742.050 ;
        RECT 749.400 730.200 750.600 739.950 ;
        RECT 755.400 739.050 756.600 754.950 ;
        RECT 758.400 754.050 759.600 781.950 ;
        RECT 760.950 778.950 763.050 781.050 ;
        RECT 757.950 751.950 760.050 754.050 ;
        RECT 754.950 736.950 757.050 739.050 ;
        RECT 748.950 728.100 751.050 730.200 ;
        RECT 754.950 728.100 757.050 730.200 ;
        RECT 761.400 730.050 762.600 778.950 ;
        RECT 767.400 775.050 768.600 802.950 ;
        RECT 788.400 801.900 789.600 802.950 ;
        RECT 787.950 799.800 790.050 801.900 ;
        RECT 781.950 790.950 784.050 793.050 ;
        RECT 769.950 784.950 772.050 787.050 ;
        RECT 766.950 772.950 769.050 775.050 ;
        RECT 766.950 765.600 769.050 766.050 ;
        RECT 770.400 765.600 771.600 784.950 ;
        RECT 766.950 764.400 771.600 765.600 ;
        RECT 766.950 763.950 769.050 764.400 ;
        RECT 767.400 760.050 768.600 763.950 ;
        RECT 772.950 762.000 775.050 766.050 ;
        RECT 773.400 760.050 774.600 762.000 ;
        RECT 778.950 760.950 781.050 766.050 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 769.950 757.950 772.050 760.050 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 775.950 757.950 778.050 760.050 ;
        RECT 770.400 745.050 771.600 757.950 ;
        RECT 776.400 756.900 777.600 757.950 ;
        RECT 775.950 754.800 778.050 756.900 ;
        RECT 772.950 751.950 775.050 754.050 ;
        RECT 769.950 742.950 772.050 745.050 ;
        RECT 766.950 736.950 769.050 739.050 ;
        RECT 749.400 727.050 750.600 728.100 ;
        RECT 755.400 727.050 756.600 728.100 ;
        RECT 760.950 727.950 763.050 730.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 754.950 724.950 757.050 727.050 ;
        RECT 757.950 724.950 760.050 727.050 ;
        RECT 745.950 721.950 748.050 724.050 ;
        RECT 746.400 691.050 747.600 721.950 ;
        RECT 748.950 718.950 751.050 721.050 ;
        RECT 745.950 688.950 748.050 691.050 ;
        RECT 742.950 685.950 745.050 688.050 ;
        RECT 749.400 687.600 750.600 718.950 ;
        RECT 752.400 709.050 753.600 724.950 ;
        RECT 758.400 723.000 759.600 724.950 ;
        RECT 757.950 718.950 760.050 723.000 ;
        RECT 760.950 721.950 763.050 724.050 ;
        RECT 767.400 723.900 768.600 736.950 ;
        RECT 773.400 730.050 774.600 751.950 ;
        RECT 776.400 733.050 777.600 754.800 ;
        RECT 782.400 748.050 783.600 790.950 ;
        RECT 797.400 784.050 798.600 823.950 ;
        RECT 802.950 811.950 805.050 814.050 ;
        RECT 803.400 808.050 804.600 811.950 ;
        RECT 802.950 805.950 805.050 808.050 ;
        RECT 808.950 807.000 811.050 811.050 ;
        RECT 815.400 808.200 816.600 826.950 ;
        RECT 824.400 825.600 825.600 832.800 ;
        RECT 827.400 832.050 828.600 838.950 ;
        RECT 826.950 829.950 829.050 832.050 ;
        RECT 824.400 824.400 828.600 825.600 ;
        RECT 823.950 817.950 826.050 820.050 ;
        RECT 809.400 805.050 810.600 807.000 ;
        RECT 814.950 806.100 817.050 808.200 ;
        RECT 815.400 805.050 816.600 806.100 ;
        RECT 824.400 805.050 825.600 817.950 ;
        RECT 827.400 810.600 828.600 824.400 ;
        RECT 830.400 814.050 831.600 853.950 ;
        RECT 841.950 850.950 844.050 853.050 ;
        RECT 835.950 839.100 838.050 841.200 ;
        RECT 842.400 841.050 843.600 850.950 ;
        RECT 836.400 838.050 837.600 839.100 ;
        RECT 841.950 838.950 844.050 841.050 ;
        RECT 835.950 835.950 838.050 838.050 ;
        RECT 838.950 835.950 841.050 838.050 ;
        RECT 839.400 834.900 840.600 835.950 ;
        RECT 838.950 832.800 841.050 834.900 ;
        RECT 835.950 829.950 838.050 832.050 ;
        RECT 829.950 811.950 832.050 814.050 ;
        RECT 827.400 809.400 831.600 810.600 ;
        RECT 830.400 805.050 831.600 809.400 ;
        RECT 836.400 808.050 837.600 829.950 ;
        RECT 845.400 816.600 846.600 854.400 ;
        RECT 851.400 841.050 852.600 868.950 ;
        RECT 857.400 865.050 858.600 877.800 ;
        RECT 856.950 862.950 859.050 865.050 ;
        RECT 863.400 856.050 864.600 898.950 ;
        RECT 868.950 895.800 871.050 897.900 ;
        RECT 869.400 883.050 870.600 895.800 ;
        RECT 878.400 895.050 879.600 913.950 ;
        RECT 892.950 907.950 895.050 910.050 ;
        RECT 889.950 895.950 892.050 898.050 ;
        RECT 877.950 892.950 880.050 895.050 ;
        RECT 890.400 892.050 891.600 895.950 ;
        RECT 889.950 889.950 892.050 892.050 ;
        RECT 893.400 886.200 894.600 907.950 ;
        RECT 896.400 901.050 897.600 913.950 ;
        RECT 895.950 898.950 898.050 901.050 ;
        RECT 896.400 888.600 897.600 898.950 ;
        RECT 916.950 892.950 919.050 895.050 ;
        RECT 904.950 889.950 907.050 892.050 ;
        RECT 896.400 887.400 900.600 888.600 ;
        RECT 874.950 884.100 877.050 886.200 ;
        RECT 892.950 884.100 895.050 886.200 ;
        RECT 875.400 883.050 876.600 884.100 ;
        RECT 893.400 883.050 894.600 884.100 ;
        RECT 899.400 883.050 900.600 887.400 ;
        RECT 868.950 880.950 871.050 883.050 ;
        RECT 871.950 880.950 874.050 883.050 ;
        RECT 874.950 880.950 877.050 883.050 ;
        RECT 877.950 880.950 880.050 883.050 ;
        RECT 892.950 880.950 895.050 883.050 ;
        RECT 895.950 880.950 898.050 883.050 ;
        RECT 898.950 880.950 901.050 883.050 ;
        RECT 872.400 871.050 873.600 880.950 ;
        RECT 878.400 874.050 879.600 880.950 ;
        RECT 880.950 877.950 883.050 880.050 ;
        RECT 896.400 879.900 897.600 880.950 ;
        RECT 905.400 880.050 906.600 889.950 ;
        RECT 877.950 871.950 880.050 874.050 ;
        RECT 871.950 868.950 874.050 871.050 ;
        RECT 862.950 853.950 865.050 856.050 ;
        RECT 877.950 853.950 880.050 856.050 ;
        RECT 856.950 850.950 859.050 853.050 ;
        RECT 850.950 838.950 853.050 841.050 ;
        RECT 857.400 838.050 858.600 850.950 ;
        RECT 874.950 844.950 877.050 847.050 ;
        RECT 875.400 841.200 876.600 844.950 ;
        RECT 878.400 843.600 879.600 853.950 ;
        RECT 881.400 847.050 882.600 877.950 ;
        RECT 895.950 877.800 898.050 879.900 ;
        RECT 904.950 877.950 907.050 880.050 ;
        RECT 913.950 877.950 916.050 880.050 ;
        RECT 889.950 850.950 892.050 853.050 ;
        RECT 880.950 844.950 883.050 847.050 ;
        RECT 878.400 842.400 882.600 843.600 ;
        RECT 862.950 839.100 865.050 841.200 ;
        RECT 874.950 839.100 877.050 841.200 ;
        RECT 863.400 838.050 864.600 839.100 ;
        RECT 875.400 838.050 876.600 839.100 ;
        RECT 881.400 838.050 882.600 842.400 ;
        RECT 853.950 835.950 856.050 838.050 ;
        RECT 856.950 835.950 859.050 838.050 ;
        RECT 859.950 835.950 862.050 838.050 ;
        RECT 862.950 835.950 865.050 838.050 ;
        RECT 871.950 835.950 874.050 838.050 ;
        RECT 874.950 835.950 877.050 838.050 ;
        RECT 877.950 835.950 880.050 838.050 ;
        RECT 880.950 835.950 883.050 838.050 ;
        RECT 854.400 835.050 855.600 835.950 ;
        RECT 850.950 833.400 855.600 835.050 ;
        RECT 860.400 834.000 861.600 835.950 ;
        RECT 868.950 834.600 871.050 835.050 ;
        RECT 872.400 834.600 873.600 835.950 ;
        RECT 878.400 834.900 879.600 835.950 ;
        RECT 890.400 835.050 891.600 850.950 ;
        RECT 898.950 844.950 901.050 847.050 ;
        RECT 899.400 838.050 900.600 844.950 ;
        RECT 898.950 835.950 901.050 838.050 ;
        RECT 850.950 832.950 855.000 833.400 ;
        RECT 859.950 829.950 862.050 834.000 ;
        RECT 868.950 833.400 873.600 834.600 ;
        RECT 868.950 832.950 871.050 833.400 ;
        RECT 842.400 815.400 846.600 816.600 ;
        RECT 835.950 805.950 838.050 808.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 823.950 802.950 826.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 829.950 802.950 832.050 805.050 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 812.400 801.900 813.600 802.950 ;
        RECT 827.400 801.900 828.600 802.950 ;
        RECT 833.400 801.900 834.600 802.950 ;
        RECT 811.950 799.800 814.050 801.900 ;
        RECT 826.950 799.800 829.050 801.900 ;
        RECT 832.950 799.800 835.050 801.900 ;
        RECT 835.950 799.950 838.050 802.050 ;
        RECT 812.400 793.050 813.600 799.800 ;
        RECT 823.950 793.950 826.050 796.050 ;
        RECT 811.950 790.950 814.050 793.050 ;
        RECT 812.400 787.050 813.600 790.950 ;
        RECT 811.950 784.950 814.050 787.050 ;
        RECT 796.950 781.950 799.050 784.050 ;
        RECT 787.950 778.950 790.050 781.050 ;
        RECT 788.400 763.200 789.600 778.950 ;
        RECT 808.950 775.950 811.050 778.050 ;
        RECT 787.950 761.100 790.050 763.200 ;
        RECT 793.950 761.100 796.050 763.200 ;
        RECT 802.800 761.100 804.900 763.200 ;
        RECT 805.950 761.100 808.050 763.200 ;
        RECT 809.400 763.050 810.600 775.950 ;
        RECT 820.950 766.950 823.050 769.050 ;
        RECT 788.400 760.050 789.600 761.100 ;
        RECT 794.400 760.050 795.600 761.100 ;
        RECT 787.950 757.950 790.050 760.050 ;
        RECT 790.950 757.950 793.050 760.050 ;
        RECT 793.950 757.950 796.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 787.950 753.600 790.050 754.050 ;
        RECT 791.400 753.600 792.600 757.950 ;
        RECT 787.950 752.400 792.600 753.600 ;
        RECT 787.950 751.950 790.050 752.400 ;
        RECT 781.950 745.950 784.050 748.050 ;
        RECT 775.950 730.950 778.050 733.050 ;
        RECT 769.950 727.950 772.050 730.050 ;
        RECT 772.950 727.950 775.050 730.050 ;
        RECT 778.950 728.100 781.050 730.200 ;
        RECT 784.950 729.000 787.050 733.050 ;
        RECT 788.400 730.050 789.600 751.950 ;
        RECT 797.400 751.050 798.600 757.950 ;
        RECT 799.950 754.950 802.050 757.050 ;
        RECT 796.950 748.950 799.050 751.050 ;
        RECT 800.400 748.050 801.600 754.950 ;
        RECT 799.950 745.950 802.050 748.050 ;
        RECT 803.400 745.050 804.600 761.100 ;
        RECT 806.400 748.050 807.600 761.100 ;
        RECT 808.950 760.950 811.050 763.050 ;
        RECT 811.950 761.100 814.050 763.200 ;
        RECT 812.400 760.050 813.600 761.100 ;
        RECT 811.950 757.950 814.050 760.050 ;
        RECT 811.950 748.950 814.050 751.050 ;
        RECT 805.950 745.950 808.050 748.050 ;
        RECT 802.950 742.950 805.050 745.050 ;
        RECT 805.950 739.950 808.050 742.050 ;
        RECT 790.950 730.950 793.050 733.050 ;
        RECT 799.950 730.950 802.050 736.050 ;
        RECT 751.950 706.950 754.050 709.050 ;
        RECT 761.400 699.600 762.600 721.950 ;
        RECT 766.950 718.950 769.050 723.900 ;
        RECT 770.400 718.050 771.600 727.950 ;
        RECT 779.400 727.050 780.600 728.100 ;
        RECT 785.400 727.050 786.600 729.000 ;
        RECT 787.950 727.950 790.050 730.050 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 778.950 724.950 781.050 727.050 ;
        RECT 781.950 724.950 784.050 727.050 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 772.950 721.950 775.050 724.050 ;
        RECT 776.400 723.900 777.600 724.950 ;
        RECT 769.950 715.950 772.050 718.050 ;
        RECT 758.400 698.400 762.600 699.600 ;
        RECT 758.400 688.050 759.600 698.400 ;
        RECT 773.400 697.050 774.600 721.950 ;
        RECT 775.950 721.800 778.050 723.900 ;
        RECT 782.400 712.050 783.600 724.950 ;
        RECT 787.950 721.950 790.050 724.050 ;
        RECT 791.400 723.900 792.600 730.950 ;
        RECT 800.400 727.050 801.600 730.950 ;
        RECT 806.400 727.050 807.600 739.950 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 802.950 724.950 805.050 727.050 ;
        RECT 805.950 724.950 808.050 727.050 ;
        RECT 797.400 723.900 798.600 724.950 ;
        RECT 784.950 718.950 787.050 721.050 ;
        RECT 775.950 709.950 778.050 712.050 ;
        RECT 781.950 709.950 784.050 712.050 ;
        RECT 776.400 700.050 777.600 709.950 ;
        RECT 781.950 703.950 784.050 706.050 ;
        RECT 775.950 697.950 778.050 700.050 ;
        RECT 782.400 697.050 783.600 703.950 ;
        RECT 760.950 694.950 763.050 697.050 ;
        RECT 772.950 694.950 775.050 697.050 ;
        RECT 781.950 694.950 784.050 697.050 ;
        RECT 746.400 686.400 750.600 687.600 ;
        RECT 746.400 682.050 747.600 686.400 ;
        RECT 757.950 685.950 760.050 688.050 ;
        RECT 761.400 685.050 762.600 694.950 ;
        RECT 757.950 682.800 760.050 684.900 ;
        RECT 760.950 682.950 763.050 685.050 ;
        RECT 766.950 683.100 769.050 688.050 ;
        RECT 772.950 683.100 775.050 685.200 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 754.950 679.950 757.050 682.050 ;
        RECT 736.950 676.950 739.050 679.050 ;
        RECT 743.400 678.900 744.600 679.950 ;
        RECT 737.400 667.050 738.600 676.950 ;
        RECT 742.950 676.800 745.050 678.900 ;
        RECT 749.400 678.000 750.600 679.950 ;
        RECT 748.950 673.950 751.050 678.000 ;
        RECT 751.950 676.950 754.050 679.050 ;
        RECT 736.950 664.950 739.050 667.050 ;
        RECT 748.950 652.950 751.050 655.050 ;
        RECT 718.950 650.100 721.050 652.200 ;
        RECT 724.950 650.100 727.050 652.200 ;
        RECT 733.950 650.100 736.050 652.200 ;
        RECT 719.400 649.050 720.600 650.100 ;
        RECT 725.400 649.050 726.600 650.100 ;
        RECT 745.950 649.950 748.050 652.050 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 724.950 646.950 727.050 649.050 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 739.950 646.950 742.050 649.050 ;
        RECT 715.950 643.950 718.050 646.050 ;
        RECT 722.400 645.900 723.600 646.950 ;
        RECT 712.950 640.950 715.050 643.050 ;
        RECT 709.950 622.950 712.050 625.050 ;
        RECT 700.950 616.950 703.050 619.050 ;
        RECT 697.950 613.950 700.050 616.050 ;
        RECT 703.950 605.100 706.050 607.200 ;
        RECT 704.400 604.050 705.600 605.100 ;
        RECT 712.950 604.950 715.050 607.050 ;
        RECT 700.950 601.950 703.050 604.050 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 701.400 600.600 702.600 601.950 ;
        RECT 707.400 600.900 708.600 601.950 ;
        RECT 713.400 600.900 714.600 604.950 ;
        RECT 698.400 599.400 702.600 600.600 ;
        RECT 694.950 595.950 697.050 598.050 ;
        RECT 694.950 592.800 697.050 594.900 ;
        RECT 691.950 580.950 694.050 583.050 ;
        RECT 682.950 571.950 685.050 574.050 ;
        RECT 685.950 568.950 688.050 571.050 ;
        RECT 686.400 567.900 687.600 568.950 ;
        RECT 667.950 562.950 670.050 567.000 ;
        RECT 677.400 566.400 681.600 567.600 ;
        RECT 673.950 559.950 676.050 562.050 ;
        RECT 661.950 556.950 664.050 559.050 ;
        RECT 667.950 556.950 670.050 559.050 ;
        RECT 655.950 535.950 658.050 538.050 ;
        RECT 655.950 527.100 658.050 529.200 ;
        RECT 656.400 526.050 657.600 527.100 ;
        RECT 655.950 523.950 658.050 526.050 ;
        RECT 661.950 523.950 664.050 526.050 ;
        RECT 650.400 521.400 654.600 522.600 ;
        RECT 622.950 494.100 625.050 496.200 ;
        RECT 628.950 494.100 631.050 496.200 ;
        RECT 623.400 493.050 624.600 494.100 ;
        RECT 629.400 493.050 630.600 494.100 ;
        RECT 634.800 493.950 636.900 496.050 ;
        RECT 637.950 494.100 640.050 496.200 ;
        RECT 643.950 494.100 646.050 496.200 ;
        RECT 653.400 496.050 654.600 521.400 ;
        RECT 658.950 520.950 661.050 523.050 ;
        RECT 662.400 522.000 663.600 523.950 ;
        RECT 655.950 496.950 658.050 499.050 ;
        RECT 619.950 490.950 622.050 493.050 ;
        RECT 622.950 490.950 625.050 493.050 ;
        RECT 625.950 490.950 628.050 493.050 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 616.950 487.800 619.050 489.900 ;
        RECT 617.400 484.050 618.600 487.800 ;
        RECT 616.950 481.950 619.050 484.050 ;
        RECT 616.950 472.950 619.050 475.050 ;
        RECT 605.400 448.050 606.600 449.100 ;
        RECT 611.400 448.050 612.600 449.100 ;
        RECT 613.950 448.950 616.050 451.050 ;
        RECT 604.950 445.950 607.050 448.050 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 598.950 442.950 601.050 445.050 ;
        RECT 601.950 442.950 604.050 445.050 ;
        RECT 608.400 444.900 609.600 445.950 ;
        RECT 598.950 433.950 601.050 436.050 ;
        RECT 595.950 418.950 598.050 421.050 ;
        RECT 599.400 417.600 600.600 433.950 ;
        RECT 596.400 416.400 600.600 417.600 ;
        RECT 596.400 415.050 597.600 416.400 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 580.950 409.950 583.050 412.050 ;
        RECT 587.400 411.900 588.600 412.950 ;
        RECT 586.950 409.800 589.050 411.900 ;
        RECT 577.950 403.950 580.050 406.050 ;
        RECT 589.950 403.950 592.050 406.050 ;
        RECT 577.950 397.950 580.050 400.050 ;
        RECT 574.950 370.950 577.050 373.050 ;
        RECT 559.950 367.950 562.050 370.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 565.950 367.950 568.050 370.050 ;
        RECT 568.950 367.950 571.050 370.050 ;
        RECT 563.400 366.900 564.600 367.950 ;
        RECT 569.400 366.900 570.600 367.950 ;
        RECT 562.950 364.800 565.050 366.900 ;
        RECT 568.950 364.800 571.050 366.900 ;
        RECT 575.400 352.050 576.600 370.950 ;
        RECT 554.400 350.400 558.600 351.600 ;
        RECT 532.950 340.950 535.050 343.050 ;
        RECT 538.950 340.950 541.050 343.050 ;
        RECT 529.950 328.950 532.050 331.050 ;
        RECT 533.400 307.050 534.600 340.950 ;
        RECT 542.400 340.200 543.600 349.950 ;
        RECT 550.950 344.400 553.050 346.500 ;
        RECT 541.950 338.100 544.050 340.200 ;
        RECT 547.950 338.400 550.050 340.500 ;
        RECT 542.400 337.050 543.600 338.100 ;
        RECT 548.400 337.050 549.600 338.400 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 539.400 328.050 540.600 334.950 ;
        RECT 551.850 329.400 553.050 344.400 ;
        RECT 538.950 325.950 541.050 328.050 ;
        RECT 550.950 327.300 553.050 329.400 ;
        RECT 551.850 323.700 553.050 327.300 ;
        RECT 557.400 325.050 558.600 350.400 ;
        RECT 559.950 349.950 562.050 352.050 ;
        RECT 574.950 349.950 577.050 352.050 ;
        RECT 550.950 321.600 553.050 323.700 ;
        RECT 556.950 322.950 559.050 325.050 ;
        RECT 538.950 310.950 541.050 313.050 ;
        RECT 532.950 304.950 535.050 307.050 ;
        RECT 526.950 298.950 529.050 301.050 ;
        RECT 527.400 292.050 528.600 298.950 ;
        RECT 532.950 294.000 535.050 298.050 ;
        RECT 533.400 292.050 534.600 294.000 ;
        RECT 539.400 292.050 540.600 310.950 ;
        RECT 547.950 304.950 550.050 307.050 ;
        RECT 544.950 295.950 547.050 298.050 ;
        RECT 526.950 289.950 529.050 292.050 ;
        RECT 529.950 289.950 532.050 292.050 ;
        RECT 532.950 289.950 535.050 292.050 ;
        RECT 535.950 289.950 538.050 292.050 ;
        RECT 538.950 289.950 541.050 292.050 ;
        RECT 530.400 288.900 531.600 289.950 ;
        RECT 529.950 286.800 532.050 288.900 ;
        RECT 530.400 283.050 531.600 286.800 ;
        RECT 529.950 280.950 532.050 283.050 ;
        RECT 536.400 280.050 537.600 289.950 ;
        RECT 545.400 288.900 546.600 295.950 ;
        RECT 544.950 286.800 547.050 288.900 ;
        RECT 535.950 279.600 538.050 280.050 ;
        RECT 535.950 278.400 540.600 279.600 ;
        RECT 535.950 277.950 538.050 278.400 ;
        RECT 523.950 260.100 526.050 265.050 ;
        RECT 529.950 260.100 532.050 262.200 ;
        RECT 530.400 259.050 531.600 260.100 ;
        RECT 535.950 259.950 538.050 265.050 ;
        RECT 526.950 256.950 529.050 259.050 ;
        RECT 529.950 256.950 532.050 259.050 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 520.950 253.800 523.050 255.900 ;
        RECT 523.950 253.950 526.050 256.050 ;
        RECT 527.400 255.900 528.600 256.950 ;
        RECT 515.400 245.400 519.600 246.600 ;
        RECT 511.950 232.950 514.050 235.050 ;
        RECT 514.950 226.950 517.050 232.050 ;
        RECT 472.950 199.950 475.050 202.050 ;
        RECT 470.400 182.400 474.600 183.600 ;
        RECT 461.400 181.050 462.600 182.100 ;
        RECT 467.400 181.050 468.600 182.100 ;
        RECT 457.950 178.950 460.050 181.050 ;
        RECT 460.950 178.950 463.050 181.050 ;
        RECT 463.950 178.950 466.050 181.050 ;
        RECT 466.950 178.950 469.050 181.050 ;
        RECT 458.400 178.050 459.600 178.950 ;
        RECT 454.950 176.400 459.600 178.050 ;
        RECT 464.400 177.900 465.600 178.950 ;
        RECT 454.950 175.950 459.000 176.400 ;
        RECT 463.950 175.800 466.050 177.900 ;
        RECT 469.950 175.950 472.050 178.050 ;
        RECT 451.950 172.950 454.050 175.050 ;
        RECT 433.950 154.950 436.050 157.050 ;
        RECT 418.950 151.950 421.050 154.050 ;
        RECT 424.950 145.950 427.050 148.050 ;
        RECT 416.400 137.400 420.600 138.600 ;
        RECT 419.400 136.050 420.600 137.400 ;
        RECT 425.400 136.050 426.600 145.950 ;
        RECT 434.400 145.050 435.600 154.950 ;
        RECT 470.400 151.050 471.600 175.950 ;
        RECT 473.400 157.050 474.600 182.400 ;
        RECT 472.950 154.950 475.050 157.050 ;
        RECT 472.950 151.800 475.050 153.900 ;
        RECT 469.950 148.950 472.050 151.050 ;
        RECT 457.950 145.950 460.050 148.050 ;
        RECT 433.950 142.950 436.050 145.050 ;
        RECT 448.950 142.950 451.050 145.050 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 421.950 133.950 424.050 136.050 ;
        RECT 424.950 133.950 427.050 136.050 ;
        RECT 412.950 130.800 415.050 132.900 ;
        RECT 403.950 112.950 406.050 115.050 ;
        RECT 403.950 108.600 406.050 111.900 ;
        RECT 406.950 108.600 409.050 109.050 ;
        RECT 403.950 108.000 409.050 108.600 ;
        RECT 404.400 107.400 409.050 108.000 ;
        RECT 406.950 106.950 409.050 107.400 ;
        RECT 407.400 103.050 408.600 106.950 ;
        RECT 413.400 104.400 420.600 105.600 ;
        RECT 413.400 103.050 414.600 104.400 ;
        RECT 403.950 100.950 406.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 404.400 99.900 405.600 100.950 ;
        RECT 403.950 97.800 406.050 99.900 ;
        RECT 410.400 88.050 411.600 100.950 ;
        RECT 409.950 85.950 412.050 88.050 ;
        RECT 397.950 82.950 400.050 85.050 ;
        RECT 397.950 76.950 400.050 79.050 ;
        RECT 398.400 55.050 399.600 76.950 ;
        RECT 412.950 67.950 415.050 70.050 ;
        RECT 406.950 60.000 409.050 64.050 ;
        RECT 413.400 61.200 414.600 67.950 ;
        RECT 419.400 64.050 420.600 104.400 ;
        RECT 422.400 100.050 423.600 133.950 ;
        RECT 434.400 103.050 435.600 142.950 ;
        RECT 442.950 137.100 445.050 139.200 ;
        RECT 443.400 136.050 444.600 137.100 ;
        RECT 449.400 136.050 450.600 142.950 ;
        RECT 439.950 133.950 442.050 136.050 ;
        RECT 442.950 133.950 445.050 136.050 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 440.400 132.900 441.600 133.950 ;
        RECT 439.950 130.800 442.050 132.900 ;
        RECT 446.400 124.050 447.600 133.950 ;
        RECT 458.400 132.900 459.600 145.950 ;
        RECT 466.950 142.950 469.050 145.050 ;
        RECT 467.400 139.200 468.600 142.950 ;
        RECT 466.950 137.100 469.050 139.200 ;
        RECT 467.400 136.050 468.600 137.100 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 464.400 132.900 465.600 133.950 ;
        RECT 457.950 130.800 460.050 132.900 ;
        RECT 463.950 130.800 466.050 132.900 ;
        RECT 469.950 124.950 472.050 127.050 ;
        RECT 445.950 121.950 448.050 124.050 ;
        RECT 470.400 121.050 471.600 124.950 ;
        RECT 469.950 118.950 472.050 121.050 ;
        RECT 451.950 109.950 454.050 112.050 ;
        RECT 442.950 103.950 445.050 106.050 ;
        RECT 445.950 103.950 448.050 109.050 ;
        RECT 448.950 106.950 451.050 109.050 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 421.950 97.950 424.050 100.050 ;
        RECT 428.400 99.900 429.600 100.950 ;
        RECT 427.950 97.800 430.050 99.900 ;
        RECT 428.400 67.050 429.600 97.800 ;
        RECT 437.400 94.050 438.600 100.950 ;
        RECT 436.950 91.950 439.050 94.050 ;
        RECT 443.400 88.050 444.600 103.950 ;
        RECT 449.400 99.900 450.600 106.950 ;
        RECT 452.400 106.050 453.600 109.950 ;
        RECT 451.950 103.950 454.050 106.050 ;
        RECT 457.950 105.000 460.050 109.050 ;
        RECT 458.400 103.050 459.600 105.000 ;
        RECT 463.950 104.100 466.050 106.200 ;
        RECT 464.400 103.050 465.600 104.100 ;
        RECT 473.400 103.050 474.600 151.800 ;
        RECT 476.400 132.900 477.600 208.950 ;
        RECT 478.950 199.950 481.050 202.050 ;
        RECT 479.400 184.050 480.600 199.950 ;
        RECT 482.400 187.050 483.600 208.950 ;
        RECT 484.950 208.800 487.050 210.900 ;
        RECT 490.800 210.000 492.900 210.900 ;
        RECT 490.800 208.800 493.050 210.000 ;
        RECT 493.950 208.950 496.050 211.050 ;
        RECT 490.950 205.950 493.050 208.800 ;
        RECT 497.400 205.050 498.600 215.100 ;
        RECT 499.950 214.950 502.050 217.050 ;
        RECT 505.950 215.100 508.050 217.200 ;
        RECT 506.400 214.050 507.600 215.100 ;
        RECT 511.950 214.950 514.050 220.050 ;
        RECT 502.950 211.950 505.050 214.050 ;
        RECT 505.950 211.950 508.050 214.050 ;
        RECT 508.950 211.950 511.050 214.050 ;
        RECT 503.400 210.900 504.600 211.950 ;
        RECT 509.400 210.900 510.600 211.950 ;
        RECT 515.400 211.050 516.600 226.950 ;
        RECT 502.950 208.800 505.050 210.900 ;
        RECT 508.950 208.800 511.050 210.900 ;
        RECT 511.950 208.950 514.050 211.050 ;
        RECT 514.950 208.950 517.050 211.050 ;
        RECT 496.950 202.950 499.050 205.050 ;
        RECT 499.950 190.950 502.050 193.050 ;
        RECT 484.950 187.950 487.050 190.050 ;
        RECT 481.950 184.950 484.050 187.050 ;
        RECT 478.950 181.950 481.050 184.050 ;
        RECT 485.400 181.050 486.600 187.950 ;
        RECT 491.400 182.400 498.600 183.600 ;
        RECT 491.400 181.050 492.600 182.400 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 484.950 178.950 487.050 181.050 ;
        RECT 487.950 178.950 490.050 181.050 ;
        RECT 490.950 178.950 493.050 181.050 ;
        RECT 482.400 177.900 483.600 178.950 ;
        RECT 488.400 177.900 489.600 178.950 ;
        RECT 481.950 175.800 484.050 177.900 ;
        RECT 487.950 175.800 490.050 177.900 ;
        RECT 478.950 172.950 481.050 175.050 ;
        RECT 479.400 154.050 480.600 172.950 ;
        RECT 478.950 151.950 481.050 154.050 ;
        RECT 487.950 138.000 490.050 142.050 ;
        RECT 497.400 139.200 498.600 182.400 ;
        RECT 500.400 181.050 501.600 190.950 ;
        RECT 512.400 187.050 513.600 208.950 ;
        RECT 514.950 205.800 517.050 207.900 ;
        RECT 511.950 184.950 514.050 187.050 ;
        RECT 502.950 181.950 505.050 184.050 ;
        RECT 508.950 182.100 511.050 184.200 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 503.400 142.050 504.600 181.950 ;
        RECT 509.400 181.050 510.600 182.100 ;
        RECT 515.400 181.050 516.600 205.800 ;
        RECT 518.400 193.050 519.600 245.400 ;
        RECT 524.400 232.050 525.600 253.950 ;
        RECT 526.950 253.800 529.050 255.900 ;
        RECT 533.400 247.050 534.600 256.950 ;
        RECT 539.400 255.900 540.600 278.400 ;
        RECT 548.400 271.050 549.600 304.950 ;
        RECT 553.950 293.100 556.050 295.200 ;
        RECT 560.400 294.600 561.600 349.950 ;
        RECT 571.950 344.400 574.050 346.500 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 566.400 322.050 567.600 334.950 ;
        RECT 572.100 324.600 573.300 344.400 ;
        RECT 578.400 340.050 579.600 397.950 ;
        RECT 590.400 381.600 591.600 403.950 ;
        RECT 593.400 385.050 594.600 412.950 ;
        RECT 598.950 409.950 601.050 412.050 ;
        RECT 599.400 400.050 600.600 409.950 ;
        RECT 598.950 397.950 601.050 400.050 ;
        RECT 592.950 382.950 595.050 385.050 ;
        RECT 602.400 382.050 603.600 442.950 ;
        RECT 607.950 442.800 610.050 444.900 ;
        RECT 613.950 442.950 616.050 445.050 ;
        RECT 614.400 433.050 615.600 442.950 ;
        RECT 617.400 436.050 618.600 472.950 ;
        RECT 620.400 463.050 621.600 490.950 ;
        RECT 626.400 489.900 627.600 490.950 ;
        RECT 625.950 487.800 628.050 489.900 ;
        RECT 622.950 481.950 625.050 484.050 ;
        RECT 619.950 460.950 622.050 463.050 ;
        RECT 619.950 454.950 622.050 457.050 ;
        RECT 620.400 448.050 621.600 454.950 ;
        RECT 619.950 445.950 622.050 448.050 ;
        RECT 623.400 442.050 624.600 481.950 ;
        RECT 631.950 475.950 634.050 478.050 ;
        RECT 632.400 466.050 633.600 475.950 ;
        RECT 631.950 463.950 634.050 466.050 ;
        RECT 625.950 457.950 628.050 460.050 ;
        RECT 626.400 450.600 627.600 457.950 ;
        RECT 635.400 457.050 636.600 493.950 ;
        RECT 638.400 490.050 639.600 494.100 ;
        RECT 644.400 493.050 645.600 494.100 ;
        RECT 652.950 493.950 655.050 496.050 ;
        RECT 643.950 490.950 646.050 493.050 ;
        RECT 649.950 490.950 652.050 493.050 ;
        RECT 637.950 487.950 640.050 490.050 ;
        RECT 646.950 487.950 649.050 490.050 ;
        RECT 650.400 489.000 651.600 490.950 ;
        RECT 647.400 463.050 648.600 487.950 ;
        RECT 649.950 484.950 652.050 489.000 ;
        RECT 652.950 487.950 655.050 490.050 ;
        RECT 653.400 472.050 654.600 487.950 ;
        RECT 656.400 484.050 657.600 496.950 ;
        RECT 659.400 487.050 660.600 520.950 ;
        RECT 661.950 517.950 664.050 522.000 ;
        RECT 664.950 520.950 667.050 523.050 ;
        RECT 662.400 511.050 663.600 517.950 ;
        RECT 665.400 517.050 666.600 520.950 ;
        RECT 664.950 514.950 667.050 517.050 ;
        RECT 661.950 508.950 664.050 511.050 ;
        RECT 661.950 499.950 664.050 502.050 ;
        RECT 662.400 490.050 663.600 499.950 ;
        RECT 668.400 499.050 669.600 556.950 ;
        RECT 674.400 547.050 675.600 559.950 ;
        RECT 673.950 544.950 676.050 547.050 ;
        RECT 677.400 541.050 678.600 566.400 ;
        RECT 685.950 565.800 688.050 567.900 ;
        RECT 695.400 559.050 696.600 592.800 ;
        RECT 698.400 592.050 699.600 599.400 ;
        RECT 706.950 598.800 709.050 600.900 ;
        RECT 712.950 598.800 715.050 600.900 ;
        RECT 700.950 595.950 703.050 598.050 ;
        RECT 697.950 589.950 700.050 592.050 ;
        RECT 698.400 562.050 699.600 589.950 ;
        RECT 697.950 559.950 700.050 562.050 ;
        RECT 682.950 556.950 685.050 559.050 ;
        RECT 694.950 556.950 697.050 559.050 ;
        RECT 679.950 544.950 682.050 547.050 ;
        RECT 676.950 538.950 679.050 541.050 ;
        RECT 680.400 535.050 681.600 544.950 ;
        RECT 670.950 532.950 673.050 535.050 ;
        RECT 679.950 532.950 682.050 535.050 ;
        RECT 671.400 529.050 672.600 532.950 ;
        RECT 670.950 526.950 673.050 529.050 ;
        RECT 673.950 527.100 676.050 529.200 ;
        RECT 674.400 526.050 675.600 527.100 ;
        RECT 680.400 526.050 681.600 532.950 ;
        RECT 683.400 529.050 684.600 556.950 ;
        RECT 697.950 553.950 700.050 556.050 ;
        RECT 688.950 537.300 691.050 539.400 ;
        RECT 694.950 538.950 697.050 541.050 ;
        RECT 689.850 533.700 691.050 537.300 ;
        RECT 688.950 531.600 691.050 533.700 ;
        RECT 682.950 526.950 685.050 529.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 670.950 520.950 673.050 523.050 ;
        RECT 671.400 502.050 672.600 520.950 ;
        RECT 677.400 511.050 678.600 523.950 ;
        RECT 686.400 522.600 687.600 523.950 ;
        RECT 683.400 521.400 687.600 522.600 ;
        RECT 679.950 517.950 682.050 520.050 ;
        RECT 676.950 508.950 679.050 511.050 ;
        RECT 670.950 499.950 673.050 502.050 ;
        RECT 667.950 496.950 670.050 499.050 ;
        RECT 670.950 494.100 673.050 496.200 ;
        RECT 671.400 493.050 672.600 494.100 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 673.950 490.950 676.050 493.050 ;
        RECT 661.950 487.950 664.050 490.050 ;
        RECT 668.400 489.000 669.600 490.950 ;
        RECT 658.950 486.900 663.000 487.050 ;
        RECT 658.950 484.950 664.050 486.900 ;
        RECT 664.950 484.950 667.050 487.050 ;
        RECT 667.950 484.950 670.050 489.000 ;
        RECT 661.950 484.800 664.050 484.950 ;
        RECT 655.950 481.950 658.050 484.050 ;
        RECT 658.950 481.800 661.050 483.900 ;
        RECT 652.950 469.950 655.050 472.050 ;
        RECT 646.950 460.950 649.050 463.050 ;
        RECT 659.400 460.050 660.600 481.800 ;
        RECT 661.950 466.950 664.050 469.050 ;
        RECT 643.950 457.950 646.050 460.050 ;
        RECT 658.950 457.950 661.050 460.050 ;
        RECT 634.950 454.950 637.050 457.050 ;
        RECT 640.950 454.950 643.050 457.050 ;
        RECT 626.400 449.400 630.600 450.600 ;
        RECT 629.400 448.050 630.600 449.400 ;
        RECT 634.950 449.100 637.050 451.200 ;
        RECT 641.400 451.050 642.600 454.950 ;
        RECT 635.400 448.050 636.600 449.100 ;
        RECT 640.950 448.950 643.050 451.050 ;
        RECT 628.950 445.950 631.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 634.950 445.950 637.050 448.050 ;
        RECT 637.950 445.950 640.050 448.050 ;
        RECT 625.950 442.950 628.050 445.050 ;
        RECT 632.400 444.900 633.600 445.950 ;
        RECT 622.950 439.950 625.050 442.050 ;
        RECT 616.950 433.950 619.050 436.050 ;
        RECT 613.950 430.950 616.050 433.050 ;
        RECT 604.950 424.950 607.050 427.050 ;
        RECT 605.400 406.050 606.600 424.950 ;
        RECT 614.400 418.050 615.600 430.950 ;
        RECT 626.400 430.050 627.600 442.950 ;
        RECT 631.950 442.800 634.050 444.900 ;
        RECT 638.400 444.000 639.600 445.950 ;
        RECT 637.950 439.950 640.050 444.000 ;
        RECT 640.950 442.950 643.050 445.050 ;
        RECT 641.400 433.050 642.600 442.950 ;
        RECT 644.400 439.050 645.600 457.950 ;
        RECT 662.400 454.050 663.600 466.950 ;
        RECT 661.950 451.950 664.050 454.050 ;
        RECT 652.950 449.100 655.050 451.200 ;
        RECT 658.950 449.100 661.050 451.200 ;
        RECT 665.400 451.050 666.600 484.950 ;
        RECT 674.400 469.050 675.600 490.950 ;
        RECT 676.950 469.950 679.050 472.050 ;
        RECT 673.950 466.950 676.050 469.050 ;
        RECT 670.950 459.300 673.050 461.400 ;
        RECT 671.850 455.700 673.050 459.300 ;
        RECT 670.950 453.600 673.050 455.700 ;
        RECT 653.400 448.050 654.600 449.100 ;
        RECT 659.400 448.050 660.600 449.100 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 652.950 445.950 655.050 448.050 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 646.950 442.950 649.050 445.050 ;
        RECT 643.950 436.950 646.050 439.050 ;
        RECT 640.950 430.950 643.050 433.050 ;
        RECT 625.950 427.950 628.050 430.050 ;
        RECT 637.950 427.950 640.050 430.050 ;
        RECT 638.400 424.050 639.600 427.950 ;
        RECT 637.950 421.950 640.050 424.050 ;
        RECT 613.950 415.950 616.050 418.050 ;
        RECT 616.950 417.000 619.050 421.050 ;
        RECT 617.400 415.050 618.600 417.000 ;
        RECT 622.950 415.950 625.050 418.050 ;
        RECT 628.950 416.100 631.050 418.200 ;
        RECT 634.950 416.100 637.050 418.200 ;
        RECT 641.400 418.050 642.600 430.950 ;
        RECT 647.400 426.600 648.600 442.950 ;
        RECT 650.400 439.050 651.600 445.950 ;
        RECT 656.400 439.050 657.600 445.950 ;
        RECT 661.950 441.600 664.050 445.050 ;
        RECT 668.400 444.600 669.600 445.950 ;
        RECT 659.400 441.000 664.050 441.600 ;
        RECT 665.400 443.400 670.050 444.600 ;
        RECT 659.400 440.400 663.600 441.000 ;
        RECT 649.950 436.950 652.050 439.050 ;
        RECT 655.950 436.950 658.050 439.050 ;
        RECT 649.950 430.950 652.050 433.050 ;
        RECT 644.400 425.400 648.600 426.600 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 616.950 412.950 619.050 415.050 ;
        RECT 611.400 411.900 612.600 412.950 ;
        RECT 610.950 409.800 613.050 411.900 ;
        RECT 604.950 403.950 607.050 406.050 ;
        RECT 610.950 385.950 613.050 388.050 ;
        RECT 590.400 380.400 594.600 381.600 ;
        RECT 583.950 371.100 586.050 373.200 ;
        RECT 584.400 370.050 585.600 371.100 ;
        RECT 583.950 367.950 586.050 370.050 ;
        RECT 586.950 367.950 589.050 370.050 ;
        RECT 587.400 361.050 588.600 367.950 ;
        RECT 586.950 358.950 589.050 361.050 ;
        RECT 593.400 358.050 594.600 380.400 ;
        RECT 601.950 379.950 604.050 382.050 ;
        RECT 602.400 375.600 603.600 379.950 ;
        RECT 599.400 374.400 603.600 375.600 ;
        RECT 599.400 370.050 600.600 374.400 ;
        RECT 604.950 372.000 607.050 376.050 ;
        RECT 611.400 373.050 612.600 385.950 ;
        RECT 613.950 379.950 616.050 382.050 ;
        RECT 605.400 370.050 606.600 372.000 ;
        RECT 610.950 370.950 613.050 373.050 ;
        RECT 598.950 367.950 601.050 370.050 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 604.950 367.950 607.050 370.050 ;
        RECT 607.950 367.950 610.050 370.050 ;
        RECT 602.400 366.900 603.600 367.950 ;
        RECT 601.950 364.800 604.050 366.900 ;
        RECT 608.400 366.000 609.600 367.950 ;
        RECT 607.950 361.950 610.050 366.000 ;
        RECT 610.950 364.800 613.050 366.900 ;
        RECT 592.950 355.950 595.050 358.050 ;
        RECT 601.950 355.950 604.050 358.050 ;
        RECT 580.950 343.950 583.050 346.050 ;
        RECT 581.400 340.050 582.600 343.950 ;
        RECT 577.950 337.950 580.050 340.050 ;
        RECT 580.950 337.950 583.050 340.050 ;
        RECT 589.950 339.000 592.050 343.050 ;
        RECT 590.400 337.050 591.600 339.000 ;
        RECT 595.950 338.100 598.050 340.200 ;
        RECT 602.400 340.050 603.600 355.950 ;
        RECT 607.950 349.950 610.050 352.050 ;
        RECT 596.400 337.050 597.600 338.100 ;
        RECT 601.950 337.950 604.050 340.050 ;
        RECT 604.950 338.100 607.050 340.200 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 575.400 333.600 576.600 334.950 ;
        RECT 580.950 334.800 583.050 336.900 ;
        RECT 586.950 334.950 589.050 337.050 ;
        RECT 589.950 334.950 592.050 337.050 ;
        RECT 592.950 334.950 595.050 337.050 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 574.950 331.500 577.050 333.600 ;
        RECT 581.400 325.050 582.600 334.800 ;
        RECT 583.950 331.950 586.050 334.050 ;
        RECT 571.950 322.500 574.050 324.600 ;
        RECT 580.950 322.950 583.050 325.050 ;
        RECT 565.950 319.950 568.050 322.050 ;
        RECT 577.950 321.600 580.050 322.050 ;
        RECT 584.400 321.600 585.600 331.950 ;
        RECT 587.400 328.050 588.600 334.950 ;
        RECT 593.400 333.900 594.600 334.950 ;
        RECT 599.400 333.900 600.600 334.950 ;
        RECT 592.950 331.800 595.050 333.900 ;
        RECT 598.950 331.800 601.050 333.900 ;
        RECT 601.950 331.950 604.050 334.050 ;
        RECT 589.950 328.950 592.050 331.050 ;
        RECT 586.950 325.950 589.050 328.050 ;
        RECT 590.400 325.050 591.600 328.950 ;
        RECT 602.400 328.050 603.600 331.950 ;
        RECT 592.950 325.950 595.050 328.050 ;
        RECT 601.950 325.950 604.050 328.050 ;
        RECT 589.950 322.950 592.050 325.050 ;
        RECT 577.950 320.400 585.600 321.600 ;
        RECT 577.950 319.950 580.050 320.400 ;
        RECT 586.950 316.950 589.050 319.050 ;
        RECT 587.400 298.050 588.600 316.950 ;
        RECT 586.950 295.950 589.050 298.050 ;
        RECT 560.400 293.400 564.600 294.600 ;
        RECT 554.400 292.050 555.600 293.100 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 556.950 289.950 559.050 292.050 ;
        RECT 557.400 288.900 558.600 289.950 ;
        RECT 556.950 286.800 559.050 288.900 ;
        RECT 557.400 277.050 558.600 286.800 ;
        RECT 556.950 274.950 559.050 277.050 ;
        RECT 547.950 268.950 550.050 271.050 ;
        RECT 541.950 265.950 544.050 268.050 ;
        RECT 538.950 253.800 541.050 255.900 ;
        RECT 542.400 255.600 543.600 265.950 ;
        RECT 547.950 264.600 552.000 265.050 ;
        RECT 547.950 262.950 552.600 264.600 ;
        RECT 551.400 259.050 552.600 262.950 ;
        RECT 547.950 256.950 550.050 259.050 ;
        RECT 550.950 256.950 553.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 548.400 255.600 549.600 256.950 ;
        RECT 542.400 254.400 549.600 255.600 ;
        RECT 557.400 255.600 558.600 256.950 ;
        RECT 557.400 254.400 561.600 255.600 ;
        RECT 532.950 244.950 535.050 247.050 ;
        RECT 541.950 232.950 544.050 235.050 ;
        RECT 523.950 229.950 526.050 232.050 ;
        RECT 526.950 223.950 529.050 226.050 ;
        RECT 520.950 215.100 523.050 217.200 ;
        RECT 521.400 205.050 522.600 215.100 ;
        RECT 527.400 214.050 528.600 223.950 ;
        RECT 532.950 215.100 535.050 217.200 ;
        RECT 533.400 214.050 534.600 215.100 ;
        RECT 526.950 211.950 529.050 214.050 ;
        RECT 529.950 211.950 532.050 214.050 ;
        RECT 532.950 211.950 535.050 214.050 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 523.950 205.950 526.050 211.050 ;
        RECT 520.950 202.950 523.050 205.050 ;
        RECT 517.950 190.950 520.050 193.050 ;
        RECT 521.400 184.050 522.600 202.950 ;
        RECT 530.400 196.050 531.600 211.950 ;
        RECT 536.400 205.050 537.600 211.950 ;
        RECT 542.400 211.050 543.600 232.950 ;
        RECT 545.400 223.050 546.600 254.400 ;
        RECT 547.950 238.950 550.050 241.050 ;
        RECT 544.950 220.950 547.050 223.050 ;
        RECT 548.400 214.050 549.600 238.950 ;
        RECT 560.400 226.050 561.600 254.400 ;
        RECT 559.950 223.950 562.050 226.050 ;
        RECT 553.950 215.100 556.050 217.200 ;
        RECT 554.400 214.050 555.600 215.100 ;
        RECT 547.950 211.950 550.050 214.050 ;
        RECT 550.950 211.950 553.050 214.050 ;
        RECT 553.950 211.950 556.050 214.050 ;
        RECT 541.950 208.950 544.050 211.050 ;
        RECT 551.400 205.050 552.600 211.950 ;
        RECT 556.950 208.950 559.050 211.050 ;
        RECT 535.950 202.950 538.050 205.050 ;
        RECT 544.950 202.950 547.050 205.050 ;
        RECT 550.950 202.950 553.050 205.050 ;
        RECT 529.950 193.950 532.050 196.050 ;
        RECT 541.950 193.950 544.050 196.050 ;
        RECT 535.950 187.950 538.050 190.050 ;
        RECT 523.950 184.950 526.050 187.050 ;
        RECT 520.950 181.950 523.050 184.050 ;
        RECT 508.950 178.950 511.050 181.050 ;
        RECT 511.950 178.950 514.050 181.050 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 517.950 178.950 520.050 181.050 ;
        RECT 512.400 177.900 513.600 178.950 ;
        RECT 511.950 175.800 514.050 177.900 ;
        RECT 518.400 172.050 519.600 178.950 ;
        RECT 524.400 177.900 525.600 184.950 ;
        RECT 529.950 183.000 532.050 187.050 ;
        RECT 530.400 181.050 531.600 183.000 ;
        RECT 536.400 181.050 537.600 187.950 ;
        RECT 542.400 184.050 543.600 193.950 ;
        RECT 541.950 181.950 544.050 184.050 ;
        RECT 529.950 178.950 532.050 181.050 ;
        RECT 532.950 178.950 535.050 181.050 ;
        RECT 535.950 178.950 538.050 181.050 ;
        RECT 538.950 178.950 541.050 181.050 ;
        RECT 533.400 177.900 534.600 178.950 ;
        RECT 539.400 177.900 540.600 178.950 ;
        RECT 545.400 177.900 546.600 202.950 ;
        RECT 551.400 181.050 552.600 202.950 ;
        RECT 557.400 184.050 558.600 208.950 ;
        RECT 556.950 181.950 559.050 184.050 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 523.950 175.800 526.050 177.900 ;
        RECT 532.950 175.800 535.050 177.900 ;
        RECT 538.950 175.800 541.050 177.900 ;
        RECT 544.950 175.800 547.050 177.900 ;
        RECT 547.950 175.950 550.050 178.050 ;
        RECT 554.400 177.900 555.600 178.950 ;
        RECT 517.950 169.950 520.050 172.050 ;
        RECT 538.950 154.950 541.050 157.050 ;
        RECT 532.950 148.950 535.050 151.050 ;
        RECT 502.950 139.950 505.050 142.050 ;
        RECT 496.950 138.600 499.050 139.200 ;
        RECT 488.400 136.050 489.600 138.000 ;
        RECT 494.400 137.400 499.050 138.600 ;
        RECT 494.400 136.050 495.600 137.400 ;
        RECT 496.950 137.100 499.050 137.400 ;
        RECT 503.400 136.050 504.600 139.950 ;
        RECT 508.950 137.100 511.050 139.200 ;
        RECT 509.400 136.050 510.600 137.100 ;
        RECT 533.400 136.050 534.600 148.950 ;
        RECT 539.400 136.050 540.600 154.950 ;
        RECT 548.400 142.050 549.600 175.950 ;
        RECT 553.950 175.800 556.050 177.900 ;
        RECT 554.400 172.050 555.600 175.800 ;
        RECT 560.400 175.050 561.600 223.950 ;
        RECT 559.950 172.950 562.050 175.050 ;
        RECT 553.950 169.950 556.050 172.050 ;
        RECT 563.400 159.600 564.600 293.400 ;
        RECT 568.950 293.100 571.050 295.200 ;
        RECT 574.950 293.100 577.050 295.200 ;
        RECT 583.950 293.100 586.050 295.200 ;
        RECT 569.400 292.050 570.600 293.100 ;
        RECT 575.400 292.050 576.600 293.100 ;
        RECT 568.950 289.950 571.050 292.050 ;
        RECT 571.950 289.950 574.050 292.050 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 577.950 289.950 580.050 292.050 ;
        RECT 565.950 280.950 568.050 283.050 ;
        RECT 566.400 217.200 567.600 280.950 ;
        RECT 572.400 280.050 573.600 289.950 ;
        RECT 571.950 277.950 574.050 280.050 ;
        RECT 568.950 268.950 571.050 271.050 ;
        RECT 569.400 262.050 570.600 268.950 ;
        RECT 578.400 268.050 579.600 289.950 ;
        RECT 584.400 283.050 585.600 293.100 ;
        RECT 583.950 280.950 586.050 283.050 ;
        RECT 577.950 265.950 580.050 268.050 ;
        RECT 587.400 264.600 588.600 295.950 ;
        RECT 593.400 295.200 594.600 325.950 ;
        RECT 598.950 310.950 601.050 313.050 ;
        RECT 592.950 293.100 595.050 295.200 ;
        RECT 593.400 292.050 594.600 293.100 ;
        RECT 599.400 292.050 600.600 310.950 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 595.950 289.950 598.050 292.050 ;
        RECT 598.950 289.950 601.050 292.050 ;
        RECT 596.400 283.050 597.600 289.950 ;
        RECT 605.400 289.050 606.600 338.100 ;
        RECT 604.950 286.950 607.050 289.050 ;
        RECT 595.950 280.950 598.050 283.050 ;
        RECT 608.400 280.050 609.600 349.950 ;
        RECT 611.400 340.050 612.600 364.800 ;
        RECT 614.400 343.050 615.600 379.950 ;
        RECT 623.400 376.050 624.600 415.950 ;
        RECT 629.400 415.050 630.600 416.100 ;
        RECT 635.400 415.050 636.600 416.100 ;
        RECT 640.950 415.950 643.050 418.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 632.400 406.050 633.600 412.950 ;
        RECT 631.950 403.950 634.050 406.050 ;
        RECT 638.400 403.050 639.600 412.950 ;
        RECT 640.950 409.950 643.050 412.050 ;
        RECT 637.950 400.950 640.050 403.050 ;
        RECT 625.950 391.950 628.050 394.050 ;
        RECT 616.950 373.950 619.050 376.050 ;
        RECT 622.950 373.950 625.050 376.050 ;
        RECT 617.400 367.050 618.600 373.950 ;
        RECT 626.400 370.050 627.600 391.950 ;
        RECT 641.400 373.200 642.600 409.950 ;
        RECT 631.950 371.100 634.050 373.200 ;
        RECT 640.950 371.100 643.050 373.200 ;
        RECT 632.400 370.050 633.600 371.100 ;
        RECT 622.950 367.950 625.050 370.050 ;
        RECT 625.950 367.950 628.050 370.050 ;
        RECT 628.950 367.950 631.050 370.050 ;
        RECT 631.950 367.950 634.050 370.050 ;
        RECT 616.950 364.950 619.050 367.050 ;
        RECT 623.400 366.000 624.600 367.950 ;
        RECT 622.950 361.950 625.050 366.000 ;
        RECT 629.400 355.050 630.600 367.950 ;
        RECT 628.950 352.950 631.050 355.050 ;
        RECT 644.400 352.050 645.600 425.400 ;
        RECT 646.950 421.950 649.050 424.050 ;
        RECT 647.400 382.050 648.600 421.950 ;
        RECT 650.400 388.050 651.600 430.950 ;
        RECT 659.400 415.050 660.600 440.400 ;
        RECT 665.400 433.050 666.600 443.400 ;
        RECT 667.950 442.500 670.050 443.400 ;
        RECT 671.850 438.600 673.050 453.600 ;
        RECT 670.950 436.500 673.050 438.600 ;
        RECT 664.950 430.950 667.050 433.050 ;
        RECT 677.400 424.050 678.600 469.950 ;
        RECT 680.400 436.050 681.600 517.950 ;
        RECT 683.400 499.050 684.600 521.400 ;
        RECT 689.850 516.600 691.050 531.600 ;
        RECT 695.400 520.050 696.600 538.950 ;
        RECT 698.400 522.600 699.600 553.950 ;
        RECT 701.400 529.050 702.600 595.950 ;
        RECT 716.400 547.050 717.600 643.950 ;
        RECT 721.950 643.800 724.050 645.900 ;
        RECT 728.400 640.050 729.600 646.950 ;
        RECT 740.400 645.900 741.600 646.950 ;
        RECT 739.950 643.800 742.050 645.900 ;
        RECT 742.950 643.950 745.050 646.050 ;
        RECT 743.400 640.050 744.600 643.950 ;
        RECT 727.950 637.950 730.050 640.050 ;
        RECT 733.950 637.950 736.050 640.050 ;
        RECT 742.950 637.950 745.050 640.050 ;
        RECT 718.950 631.950 721.050 634.050 ;
        RECT 724.950 631.950 727.050 634.050 ;
        RECT 719.400 628.050 720.600 631.950 ;
        RECT 718.950 625.950 721.050 628.050 ;
        RECT 718.950 622.800 721.050 624.900 ;
        RECT 719.400 592.050 720.600 622.800 ;
        RECT 725.400 607.200 726.600 631.950 ;
        RECT 724.950 605.100 727.050 607.200 ;
        RECT 734.400 607.050 735.600 637.950 ;
        RECT 739.950 622.950 742.050 625.050 ;
        RECT 740.400 619.050 741.600 622.950 ;
        RECT 739.950 616.950 742.050 619.050 ;
        RECT 746.400 613.050 747.600 649.950 ;
        RECT 749.400 634.050 750.600 652.950 ;
        RECT 752.400 652.050 753.600 676.950 ;
        RECT 755.400 655.050 756.600 679.950 ;
        RECT 758.400 676.050 759.600 682.800 ;
        RECT 767.400 682.050 768.600 683.100 ;
        RECT 773.400 682.050 774.600 683.100 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 760.950 676.950 763.050 679.050 ;
        RECT 757.950 673.950 760.050 676.050 ;
        RECT 757.950 655.950 760.050 658.050 ;
        RECT 754.950 652.950 757.050 655.050 ;
        RECT 751.950 649.950 754.050 652.050 ;
        RECT 758.400 649.050 759.600 655.950 ;
        RECT 761.400 655.050 762.600 676.950 ;
        RECT 764.400 673.050 765.600 679.950 ;
        RECT 763.950 670.950 766.050 673.050 ;
        RECT 770.400 667.050 771.600 679.950 ;
        RECT 775.950 676.950 778.050 679.050 ;
        RECT 763.950 664.950 766.050 667.050 ;
        RECT 769.950 664.950 772.050 667.050 ;
        RECT 760.950 652.950 763.050 655.050 ;
        RECT 764.400 652.200 765.600 664.950 ;
        RECT 766.950 655.950 769.050 658.050 ;
        RECT 763.950 650.100 766.050 652.200 ;
        RECT 767.400 652.050 768.600 655.950 ;
        RECT 764.400 649.050 765.600 650.100 ;
        RECT 766.950 649.950 769.050 652.050 ;
        RECT 772.950 651.600 775.050 652.050 ;
        RECT 776.400 651.600 777.600 676.950 ;
        RECT 782.400 667.050 783.600 694.950 ;
        RECT 781.950 664.950 784.050 667.050 ;
        RECT 772.950 650.400 777.600 651.600 ;
        RECT 772.950 649.950 775.050 650.400 ;
        RECT 781.950 650.100 784.050 655.050 ;
        RECT 785.400 651.600 786.600 718.950 ;
        RECT 788.400 712.050 789.600 721.950 ;
        RECT 790.950 721.800 793.050 723.900 ;
        RECT 796.950 721.800 799.050 723.900 ;
        RECT 803.400 718.050 804.600 724.950 ;
        RECT 812.400 723.900 813.600 748.950 ;
        RECT 814.950 745.950 817.050 748.050 ;
        RECT 811.950 721.800 814.050 723.900 ;
        RECT 802.950 715.950 805.050 718.050 ;
        RECT 787.950 709.950 790.050 712.050 ;
        RECT 805.950 709.950 808.050 712.050 ;
        RECT 787.950 703.950 790.050 706.050 ;
        RECT 788.400 700.050 789.600 703.950 ;
        RECT 787.950 697.950 790.050 700.050 ;
        RECT 802.950 697.950 805.050 700.050 ;
        RECT 803.400 691.050 804.600 697.950 ;
        RECT 802.950 688.950 805.050 691.050 ;
        RECT 790.950 683.100 793.050 685.200 ;
        RECT 796.950 684.000 799.050 688.050 ;
        RECT 806.400 685.050 807.600 709.950 ;
        RECT 812.400 691.050 813.600 721.800 ;
        RECT 811.950 688.950 814.050 691.050 ;
        RECT 791.400 682.050 792.600 683.100 ;
        RECT 797.400 682.050 798.600 684.000 ;
        RECT 805.950 682.950 808.050 685.050 ;
        RECT 812.400 682.050 813.600 688.950 ;
        RECT 815.400 688.050 816.600 745.950 ;
        RECT 817.950 727.950 820.050 733.050 ;
        RECT 821.400 727.050 822.600 766.950 ;
        RECT 824.400 763.050 825.600 793.950 ;
        RECT 826.950 778.950 829.050 781.050 ;
        RECT 823.950 760.950 826.050 763.050 ;
        RECT 827.400 760.050 828.600 778.950 ;
        RECT 836.400 765.600 837.600 799.950 ;
        RECT 842.400 771.600 843.600 815.400 ;
        RECT 860.400 814.050 861.600 829.950 ;
        RECT 844.950 811.950 847.050 814.050 ;
        RECT 853.950 811.950 856.050 814.050 ;
        RECT 859.950 811.950 862.050 814.050 ;
        RECT 845.400 808.050 846.600 811.950 ;
        RECT 844.950 805.950 847.050 808.050 ;
        RECT 847.950 806.100 850.050 808.200 ;
        RECT 848.400 805.050 849.600 806.100 ;
        RECT 854.400 805.050 855.600 811.950 ;
        RECT 869.400 811.050 870.600 832.950 ;
        RECT 877.950 832.800 880.050 834.900 ;
        RECT 889.950 832.950 892.050 835.050 ;
        RECT 874.950 826.950 877.050 829.050 ;
        RECT 875.400 822.600 876.600 826.950 ;
        RECT 914.400 823.050 915.600 877.950 ;
        RECT 875.400 821.400 879.600 822.600 ;
        RECT 871.950 816.600 874.050 820.050 ;
        RECT 871.950 816.000 876.600 816.600 ;
        RECT 872.400 815.400 876.600 816.000 ;
        RECT 862.950 808.950 865.050 811.050 ;
        RECT 847.950 802.950 850.050 805.050 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 856.950 802.950 859.050 805.050 ;
        RECT 851.400 796.050 852.600 802.950 ;
        RECT 850.950 793.950 853.050 796.050 ;
        RECT 857.400 793.050 858.600 802.950 ;
        RECT 859.950 799.950 862.050 802.050 ;
        RECT 856.950 790.950 859.050 793.050 ;
        RECT 860.400 781.050 861.600 799.950 ;
        RECT 863.400 790.050 864.600 808.950 ;
        RECT 868.950 807.000 871.050 811.050 ;
        RECT 875.400 808.050 876.600 815.400 ;
        RECT 869.400 805.050 870.600 807.000 ;
        RECT 874.950 805.950 877.050 808.050 ;
        RECT 868.950 802.950 871.050 805.050 ;
        RECT 871.950 802.950 874.050 805.050 ;
        RECT 872.400 801.900 873.600 802.950 ;
        RECT 878.400 802.050 879.600 821.400 ;
        RECT 898.950 820.950 901.050 823.050 ;
        RECT 913.950 820.950 916.050 823.050 ;
        RECT 892.950 811.950 895.050 814.050 ;
        RECT 893.400 805.050 894.600 811.950 ;
        RECT 889.950 802.950 892.050 805.050 ;
        RECT 892.950 802.950 895.050 805.050 ;
        RECT 871.950 799.800 874.050 801.900 ;
        RECT 877.950 799.950 880.050 802.050 ;
        RECT 890.400 801.900 891.600 802.950 ;
        RECT 889.950 799.800 892.050 801.900 ;
        RECT 862.950 787.950 865.050 790.050 ;
        RECT 859.950 778.950 862.050 781.050 ;
        RECT 850.950 775.950 853.050 778.050 ;
        RECT 851.400 772.050 852.600 775.950 ;
        RECT 842.400 770.400 846.600 771.600 ;
        RECT 841.950 766.950 844.050 769.050 ;
        RECT 833.400 764.400 837.600 765.600 ;
        RECT 833.400 760.050 834.600 764.400 ;
        RECT 826.950 757.950 829.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 832.950 757.950 835.050 760.050 ;
        RECT 835.950 757.950 838.050 760.050 ;
        RECT 830.400 756.900 831.600 757.950 ;
        RECT 836.400 756.900 837.600 757.950 ;
        RECT 842.400 756.900 843.600 766.950 ;
        RECT 829.950 754.800 832.050 756.900 ;
        RECT 835.950 754.800 838.050 756.900 ;
        RECT 841.950 754.800 844.050 756.900 ;
        RECT 830.400 747.600 831.600 754.800 ;
        RECT 830.400 746.400 834.600 747.600 ;
        RECT 826.950 728.100 829.050 730.200 ;
        RECT 833.400 730.050 834.600 746.400 ;
        RECT 838.950 739.950 841.050 742.050 ;
        RECT 835.950 730.950 838.050 733.050 ;
        RECT 827.400 727.050 828.600 728.100 ;
        RECT 832.950 727.950 835.050 730.050 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 823.950 724.950 826.050 727.050 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 829.950 724.950 832.050 727.050 ;
        RECT 817.950 721.950 820.050 724.050 ;
        RECT 824.400 723.900 825.600 724.950 ;
        RECT 814.950 685.950 817.050 688.050 ;
        RECT 818.400 685.200 819.600 721.950 ;
        RECT 823.950 721.800 826.050 723.900 ;
        RECT 820.950 703.950 823.050 706.050 ;
        RECT 817.950 683.100 820.050 685.200 ;
        RECT 821.400 685.050 822.600 703.950 ;
        RECT 830.400 697.050 831.600 724.950 ;
        RECT 832.950 721.950 835.050 724.050 ;
        RECT 833.400 706.050 834.600 721.950 ;
        RECT 832.950 703.950 835.050 706.050 ;
        RECT 829.950 694.950 832.050 697.050 ;
        RECT 836.400 694.050 837.600 730.950 ;
        RECT 839.400 730.050 840.600 739.950 ;
        RECT 842.400 733.050 843.600 754.800 ;
        RECT 845.400 736.050 846.600 770.400 ;
        RECT 850.950 769.950 853.050 772.050 ;
        RECT 877.950 769.950 880.050 772.050 ;
        RECT 851.400 760.050 852.600 769.950 ;
        RECT 878.400 763.200 879.600 769.950 ;
        RECT 899.400 769.050 900.600 820.950 ;
        RECT 917.400 808.050 918.600 892.950 ;
        RECT 916.950 805.950 919.050 808.050 ;
        RECT 907.950 802.950 910.050 805.050 ;
        RECT 908.400 795.600 909.600 802.950 ;
        RECT 916.950 799.950 919.050 802.050 ;
        RECT 905.400 794.400 909.600 795.600 ;
        RECT 905.400 781.050 906.600 794.400 ;
        RECT 904.950 778.950 907.050 781.050 ;
        RECT 898.950 766.950 901.050 769.050 ;
        RECT 913.950 766.950 916.050 769.050 ;
        RECT 856.950 761.100 859.050 763.200 ;
        RECT 877.950 761.100 880.050 763.200 ;
        RECT 883.950 762.000 886.050 766.050 ;
        RECT 895.950 765.600 900.000 766.050 ;
        RECT 895.950 763.950 900.600 765.600 ;
        RECT 857.400 760.050 858.600 761.100 ;
        RECT 878.400 760.050 879.600 761.100 ;
        RECT 884.400 760.050 885.600 762.000 ;
        RECT 899.400 760.050 900.600 763.950 ;
        RECT 904.950 761.100 907.050 763.200 ;
        RECT 910.950 761.100 913.050 763.200 ;
        RECT 905.400 760.050 906.600 761.100 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 856.950 757.950 859.050 760.050 ;
        RECT 859.950 757.950 862.050 760.050 ;
        RECT 877.950 757.950 880.050 760.050 ;
        RECT 880.950 757.950 883.050 760.050 ;
        RECT 883.950 757.950 886.050 760.050 ;
        RECT 886.950 757.950 889.050 760.050 ;
        RECT 895.950 757.950 898.050 760.050 ;
        RECT 898.950 757.950 901.050 760.050 ;
        RECT 901.950 757.950 904.050 760.050 ;
        RECT 904.950 757.950 907.050 760.050 ;
        RECT 854.400 756.900 855.600 757.950 ;
        RECT 853.950 754.800 856.050 756.900 ;
        RECT 860.400 751.050 861.600 757.950 ;
        RECT 881.400 751.050 882.600 757.950 ;
        RECT 887.400 756.600 888.600 757.950 ;
        RECT 896.400 756.900 897.600 757.950 ;
        RECT 887.400 756.000 891.600 756.600 ;
        RECT 887.400 755.400 892.050 756.000 ;
        RECT 889.950 751.950 892.050 755.400 ;
        RECT 895.950 754.800 898.050 756.900 ;
        RECT 859.950 748.950 862.050 751.050 ;
        RECT 874.950 748.950 877.050 751.050 ;
        RECT 880.950 748.950 883.050 751.050 ;
        RECT 886.950 748.950 889.050 751.050 ;
        RECT 847.950 745.950 850.050 748.050 ;
        RECT 856.950 745.950 859.050 748.050 ;
        RECT 844.950 733.950 847.050 736.050 ;
        RECT 841.950 730.950 844.050 733.050 ;
        RECT 838.950 727.950 841.050 730.050 ;
        RECT 842.400 727.050 843.600 730.950 ;
        RECT 848.400 727.050 849.600 745.950 ;
        RECT 857.400 739.050 858.600 745.950 ;
        RECT 856.950 736.950 859.050 739.050 ;
        RECT 862.950 736.950 865.050 739.050 ;
        RECT 856.950 733.800 859.050 735.900 ;
        RECT 841.950 724.950 844.050 727.050 ;
        RECT 844.950 724.950 847.050 727.050 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 845.400 723.900 846.600 724.950 ;
        RECT 844.950 721.800 847.050 723.900 ;
        RECT 845.400 718.050 846.600 721.800 ;
        RECT 851.400 721.050 852.600 724.950 ;
        RECT 850.950 720.600 853.050 721.050 ;
        RECT 848.400 719.400 853.050 720.600 ;
        RECT 844.950 715.950 847.050 718.050 ;
        RECT 848.400 703.050 849.600 719.400 ;
        RECT 850.950 718.950 853.050 719.400 ;
        RECT 847.950 700.950 850.050 703.050 ;
        RECT 844.950 697.950 847.050 700.050 ;
        RECT 857.400 699.600 858.600 733.800 ;
        RECT 863.400 733.050 864.600 736.950 ;
        RECT 862.950 730.950 865.050 733.050 ;
        RECT 875.400 732.600 876.600 748.950 ;
        RECT 875.400 732.000 879.600 732.600 ;
        RECT 875.400 731.400 880.050 732.000 ;
        RECT 865.950 728.100 868.050 730.200 ;
        RECT 871.950 728.100 874.050 730.200 ;
        RECT 866.400 727.050 867.600 728.100 ;
        RECT 872.400 727.050 873.600 728.100 ;
        RECT 877.950 727.950 880.050 731.400 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 871.950 724.950 874.050 727.050 ;
        RECT 874.950 724.950 877.050 727.050 ;
        RECT 862.950 718.950 865.050 724.050 ;
        RECT 869.400 718.050 870.600 724.950 ;
        RECT 875.400 723.900 876.600 724.950 ;
        RECT 874.950 721.800 877.050 723.900 ;
        RECT 868.950 715.950 871.050 718.050 ;
        RECT 854.400 698.400 858.600 699.600 ;
        RECT 826.950 691.950 829.050 694.050 ;
        RECT 835.950 691.950 838.050 694.050 ;
        RECT 818.400 682.050 819.600 683.100 ;
        RECT 820.950 682.950 823.050 685.050 ;
        RECT 823.950 682.950 826.050 685.050 ;
        RECT 790.950 679.950 793.050 682.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 796.950 679.950 799.050 682.050 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 808.950 679.950 811.050 682.050 ;
        RECT 811.950 679.950 814.050 682.050 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 787.950 676.950 790.050 679.050 ;
        RECT 788.400 673.050 789.600 676.950 ;
        RECT 787.950 670.950 790.050 673.050 ;
        RECT 790.950 655.950 793.050 658.050 ;
        RECT 785.400 650.400 789.600 651.600 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 757.950 646.950 760.050 649.050 ;
        RECT 760.950 646.950 763.050 649.050 ;
        RECT 763.950 646.950 766.050 649.050 ;
        RECT 751.950 643.950 754.050 646.050 ;
        RECT 748.950 631.950 751.050 634.050 ;
        RECT 752.400 619.050 753.600 643.950 ;
        RECT 755.400 637.050 756.600 646.950 ;
        RECT 757.950 637.950 760.050 640.050 ;
        RECT 754.950 634.950 757.050 637.050 ;
        RECT 758.400 628.050 759.600 637.950 ;
        RECT 757.950 625.950 760.050 628.050 ;
        RECT 761.400 622.050 762.600 646.950 ;
        RECT 763.950 640.950 766.050 643.050 ;
        RECT 760.950 619.950 763.050 622.050 ;
        RECT 751.950 616.950 754.050 619.050 ;
        RECT 742.800 609.300 744.900 611.400 ;
        RECT 745.950 610.950 748.050 613.050 ;
        RECT 752.400 610.500 754.500 612.600 ;
        RECT 760.950 610.950 763.050 613.050 ;
        RECT 725.400 604.050 726.600 605.100 ;
        RECT 733.950 604.950 736.050 607.050 ;
        RECT 740.400 604.050 741.600 606.600 ;
        RECT 724.950 601.950 727.050 604.050 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 740.400 601.950 742.500 604.050 ;
        RECT 724.950 595.950 727.050 598.050 ;
        RECT 718.950 589.950 721.050 592.050 ;
        RECT 725.400 571.050 726.600 595.950 ;
        RECT 728.400 595.050 729.600 601.950 ;
        RECT 736.950 598.950 739.050 601.050 ;
        RECT 743.700 600.300 744.600 609.300 ;
        RECT 746.100 605.700 748.200 607.800 ;
        RECT 749.400 606.900 750.600 609.450 ;
        RECT 747.300 603.300 748.200 605.700 ;
        RECT 749.100 604.800 751.200 606.900 ;
        RECT 753.000 603.300 754.050 610.500 ;
        RECT 747.300 602.100 754.050 603.300 ;
        RECT 750.150 600.300 752.250 601.200 ;
        RECT 743.700 599.100 752.250 600.300 ;
        RECT 727.950 592.950 730.050 595.050 ;
        RECT 730.950 589.950 733.050 592.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 724.950 568.950 727.050 571.050 ;
        RECT 722.400 567.600 723.600 568.950 ;
        RECT 719.400 566.400 723.600 567.600 ;
        RECT 715.950 544.950 718.050 547.050 ;
        RECT 719.400 541.050 720.600 566.400 ;
        RECT 718.950 538.950 721.050 541.050 ;
        RECT 709.950 536.400 712.050 538.500 ;
        RECT 724.950 537.300 727.050 539.400 ;
        RECT 703.950 532.950 706.050 535.050 ;
        RECT 700.950 526.950 703.050 529.050 ;
        RECT 704.400 526.050 705.600 532.950 ;
        RECT 703.950 523.950 706.050 526.050 ;
        RECT 698.400 521.400 702.600 522.600 ;
        RECT 694.950 517.950 697.050 520.050 ;
        RECT 688.950 514.500 691.050 516.600 ;
        RECT 685.950 505.950 688.050 508.050 ;
        RECT 682.950 496.950 685.050 499.050 ;
        RECT 686.400 496.200 687.600 505.950 ;
        RECT 685.950 494.100 688.050 496.200 ;
        RECT 691.950 495.000 694.050 499.050 ;
        RECT 686.400 493.050 687.600 494.100 ;
        RECT 692.400 493.050 693.600 495.000 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 688.950 490.950 691.050 493.050 ;
        RECT 691.950 490.950 694.050 493.050 ;
        RECT 694.950 490.950 697.050 493.050 ;
        RECT 682.950 487.950 685.050 490.050 ;
        RECT 689.400 489.900 690.600 490.950 ;
        RECT 683.400 484.050 684.600 487.950 ;
        RECT 688.950 487.800 691.050 489.900 ;
        RECT 695.400 484.050 696.600 490.950 ;
        RECT 682.950 481.950 685.050 484.050 ;
        RECT 694.950 481.950 697.050 484.050 ;
        RECT 701.400 481.050 702.600 521.400 ;
        RECT 703.950 517.950 706.050 520.050 ;
        RECT 704.400 484.050 705.600 517.950 ;
        RECT 710.100 516.600 711.300 536.400 ;
        RECT 725.850 533.700 727.050 537.300 ;
        RECT 724.950 531.600 727.050 533.700 ;
        RECT 712.950 527.400 715.050 529.500 ;
        RECT 713.400 526.050 714.600 527.400 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 722.400 522.600 723.600 523.950 ;
        RECT 719.400 521.400 723.600 522.600 ;
        RECT 719.400 517.050 720.600 521.400 ;
        RECT 709.950 514.500 712.050 516.600 ;
        RECT 718.950 514.950 721.050 517.050 ;
        RECT 725.850 516.600 727.050 531.600 ;
        RECT 724.950 514.500 727.050 516.600 ;
        RECT 721.950 508.950 724.050 511.050 ;
        RECT 731.400 510.600 732.600 589.950 ;
        RECT 737.400 589.050 738.600 598.950 ;
        RECT 745.200 597.300 747.300 599.100 ;
        RECT 749.100 596.100 751.200 598.200 ;
        RECT 753.150 596.700 754.050 602.100 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 755.400 599.400 756.600 601.950 ;
        RECT 736.950 586.950 739.050 589.050 ;
        RECT 733.950 580.950 736.050 583.050 ;
        RECT 734.400 573.600 735.600 580.950 ;
        RECT 749.400 577.050 750.600 596.100 ;
        RECT 752.400 594.600 754.500 596.700 ;
        RECT 751.950 586.950 754.050 589.050 ;
        RECT 752.400 580.050 753.600 586.950 ;
        RECT 761.400 583.050 762.600 610.950 ;
        RECT 764.400 600.900 765.600 640.950 ;
        RECT 773.400 637.050 774.600 649.950 ;
        RECT 782.400 649.050 783.600 650.100 ;
        RECT 778.950 646.950 781.050 649.050 ;
        RECT 781.950 646.950 784.050 649.050 ;
        RECT 775.950 643.950 778.050 646.050 ;
        RECT 772.950 634.950 775.050 637.050 ;
        RECT 776.400 634.050 777.600 643.950 ;
        RECT 775.950 631.950 778.050 634.050 ;
        RECT 779.400 610.050 780.600 646.950 ;
        RECT 788.400 643.050 789.600 650.400 ;
        RECT 791.400 646.050 792.600 655.950 ;
        RECT 794.400 655.050 795.600 679.950 ;
        RECT 800.400 670.050 801.600 679.950 ;
        RECT 802.950 676.950 805.050 679.050 ;
        RECT 799.950 667.950 802.050 670.050 ;
        RECT 793.950 652.950 796.050 655.050 ;
        RECT 799.950 650.100 802.050 652.200 ;
        RECT 803.400 652.050 804.600 676.950 ;
        RECT 809.400 676.050 810.600 679.950 ;
        RECT 808.950 673.950 811.050 676.050 ;
        RECT 815.400 675.600 816.600 679.950 ;
        RECT 820.950 676.950 823.050 679.050 ;
        RECT 812.400 674.400 816.600 675.600 ;
        RECT 805.950 670.950 808.050 673.050 ;
        RECT 800.400 649.050 801.600 650.100 ;
        RECT 802.950 649.950 805.050 652.050 ;
        RECT 796.950 646.950 799.050 649.050 ;
        RECT 799.950 646.950 802.050 649.050 ;
        RECT 790.950 643.950 793.050 646.050 ;
        RECT 797.400 645.900 798.600 646.950 ;
        RECT 796.950 643.800 799.050 645.900 ;
        RECT 802.950 643.950 805.050 646.050 ;
        RECT 787.950 640.950 790.050 643.050 ;
        RECT 797.400 637.050 798.600 643.800 ;
        RECT 796.950 634.950 799.050 637.050 ;
        RECT 803.400 619.050 804.600 643.950 ;
        RECT 806.400 631.050 807.600 670.950 ;
        RECT 809.400 667.050 810.600 673.950 ;
        RECT 808.950 664.950 811.050 667.050 ;
        RECT 812.400 652.200 813.600 674.400 ;
        RECT 821.400 673.050 822.600 676.950 ;
        RECT 820.950 670.950 823.050 673.050 ;
        RECT 811.950 650.100 814.050 652.200 ;
        RECT 817.950 650.100 820.050 652.200 ;
        RECT 824.400 652.050 825.600 682.950 ;
        RECT 827.400 670.050 828.600 691.950 ;
        RECT 832.950 688.950 835.050 691.050 ;
        RECT 833.400 682.050 834.600 688.950 ;
        RECT 841.950 683.100 844.050 685.200 ;
        RECT 845.400 685.050 846.600 697.950 ;
        RECT 847.950 691.950 850.050 694.050 ;
        RECT 842.400 682.050 843.600 683.100 ;
        RECT 844.950 682.950 847.050 685.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 841.950 679.950 844.050 682.050 ;
        RECT 829.950 673.950 832.050 676.050 ;
        RECT 832.950 673.950 835.050 676.050 ;
        RECT 826.950 667.950 829.050 670.050 ;
        RECT 812.400 649.050 813.600 650.100 ;
        RECT 818.400 649.050 819.600 650.100 ;
        RECT 823.950 649.950 826.050 652.050 ;
        RECT 826.950 649.950 829.050 652.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 817.950 646.950 820.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 805.950 628.950 808.050 631.050 ;
        RECT 815.400 622.050 816.600 646.950 ;
        RECT 821.400 645.900 822.600 646.950 ;
        RECT 820.950 643.800 823.050 645.900 ;
        RECT 820.950 640.650 823.050 642.750 ;
        RECT 808.950 619.950 811.050 622.050 ;
        RECT 814.950 619.950 817.050 622.050 ;
        RECT 781.950 616.950 784.050 619.050 ;
        RECT 802.950 616.950 805.050 619.050 ;
        RECT 766.950 604.950 769.050 610.050 ;
        RECT 772.950 606.000 775.050 610.050 ;
        RECT 778.950 607.950 781.050 610.050 ;
        RECT 773.400 604.050 774.600 606.000 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 763.950 598.800 766.050 600.900 ;
        RECT 766.950 598.950 769.050 601.050 ;
        RECT 770.400 600.900 771.600 601.950 ;
        RECT 767.400 595.050 768.600 598.950 ;
        RECT 769.950 598.800 772.050 600.900 ;
        RECT 766.950 592.950 769.050 595.050 ;
        RECT 763.950 589.950 766.050 592.050 ;
        RECT 764.400 586.050 765.600 589.950 ;
        RECT 782.400 589.050 783.600 616.950 ;
        RECT 787.950 605.100 790.050 607.200 ;
        RECT 793.950 606.000 796.050 610.050 ;
        RECT 805.950 607.950 808.050 610.050 ;
        RECT 788.400 604.050 789.600 605.100 ;
        RECT 794.400 604.050 795.600 606.000 ;
        RECT 787.950 601.950 790.050 604.050 ;
        RECT 790.950 601.950 793.050 604.050 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 784.950 598.950 787.050 601.050 ;
        RECT 781.950 586.950 784.050 589.050 ;
        RECT 763.950 583.950 766.050 586.050 ;
        RECT 760.950 580.950 763.050 583.050 ;
        RECT 785.400 580.050 786.600 598.950 ;
        RECT 791.400 595.050 792.600 601.950 ;
        RECT 797.400 601.050 798.600 601.950 ;
        RECT 797.400 599.400 802.050 601.050 ;
        RECT 798.000 598.950 802.050 599.400 ;
        RECT 790.950 592.950 793.050 595.050 ;
        RECT 787.950 586.950 790.050 589.050 ;
        RECT 751.950 577.950 754.050 580.050 ;
        RECT 784.950 577.950 787.050 580.050 ;
        RECT 734.400 572.400 738.600 573.600 ;
        RECT 742.950 573.000 745.050 577.050 ;
        RECT 748.950 574.950 751.050 577.050 ;
        RECT 737.400 571.050 738.600 572.400 ;
        RECT 743.400 571.050 744.600 573.000 ;
        RECT 736.950 568.950 739.050 571.050 ;
        RECT 739.950 568.950 742.050 571.050 ;
        RECT 742.950 568.950 745.050 571.050 ;
        RECT 740.400 567.900 741.600 568.950 ;
        RECT 739.950 565.800 742.050 567.900 ;
        RECT 739.950 562.650 742.050 564.750 ;
        RECT 733.950 532.950 736.050 535.050 ;
        RECT 728.400 509.400 732.600 510.600 ;
        RECT 715.950 502.950 718.050 505.050 ;
        RECT 709.950 499.950 712.050 502.050 ;
        RECT 710.400 493.050 711.600 499.950 ;
        RECT 716.400 493.050 717.600 502.950 ;
        RECT 722.400 496.050 723.600 508.950 ;
        RECT 724.950 496.950 727.050 499.050 ;
        RECT 721.950 493.950 724.050 496.050 ;
        RECT 709.950 490.950 712.050 493.050 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 715.950 490.950 718.050 493.050 ;
        RECT 718.950 490.950 721.050 493.050 ;
        RECT 713.400 489.900 714.600 490.950 ;
        RECT 719.400 490.050 720.600 490.950 ;
        RECT 712.950 487.800 715.050 489.900 ;
        RECT 719.400 488.400 724.050 490.050 ;
        RECT 720.000 487.950 724.050 488.400 ;
        RECT 725.400 486.600 726.600 496.950 ;
        RECT 722.400 485.400 726.600 486.600 ;
        RECT 703.950 481.950 706.050 484.050 ;
        RECT 715.950 481.950 718.050 484.050 ;
        RECT 700.950 478.950 703.050 481.050 ;
        RECT 712.950 478.950 715.050 481.050 ;
        RECT 697.950 460.950 700.050 463.050 ;
        RECT 691.950 458.400 694.050 460.500 ;
        RECT 685.950 449.400 688.050 451.500 ;
        RECT 686.400 448.050 687.600 449.400 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 682.950 442.950 685.050 445.050 ;
        RECT 683.400 439.050 684.600 442.950 ;
        RECT 682.950 436.950 685.050 439.050 ;
        RECT 692.100 438.600 693.300 458.400 ;
        RECT 694.950 454.950 697.050 457.050 ;
        RECT 695.400 448.050 696.600 454.950 ;
        RECT 698.400 451.050 699.600 460.950 ;
        RECT 706.950 459.300 709.050 461.400 ;
        RECT 707.850 455.700 709.050 459.300 ;
        RECT 706.950 453.600 709.050 455.700 ;
        RECT 697.950 448.950 700.050 451.050 ;
        RECT 694.950 445.950 697.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 697.950 442.950 700.050 445.050 ;
        RECT 704.400 444.600 705.600 445.950 ;
        RECT 701.400 443.400 706.050 444.600 ;
        RECT 691.950 436.500 694.050 438.600 ;
        RECT 679.950 433.950 682.050 436.050 ;
        RECT 680.400 427.050 681.600 433.950 ;
        RECT 688.950 427.950 691.050 430.050 ;
        RECT 679.950 424.950 682.050 427.050 ;
        RECT 676.950 421.950 679.050 424.050 ;
        RECT 682.950 421.950 685.050 424.050 ;
        RECT 667.950 415.950 670.050 418.050 ;
        RECT 676.950 416.100 679.050 418.200 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 656.400 411.900 657.600 412.950 ;
        RECT 655.950 409.800 658.050 411.900 ;
        RECT 662.400 408.600 663.600 412.950 ;
        RECT 659.400 407.400 663.600 408.600 ;
        RECT 659.400 388.050 660.600 407.400 ;
        RECT 661.950 403.950 664.050 406.050 ;
        RECT 649.950 385.950 652.050 388.050 ;
        RECT 658.950 385.950 661.050 388.050 ;
        RECT 658.950 382.800 661.050 384.900 ;
        RECT 646.950 379.950 649.050 382.050 ;
        RECT 654.000 375.600 658.050 376.050 ;
        RECT 653.400 373.950 658.050 375.600 ;
        RECT 653.400 370.050 654.600 373.950 ;
        RECT 659.400 373.050 660.600 382.800 ;
        RECT 658.950 370.950 661.050 373.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 650.400 366.900 651.600 367.950 ;
        RECT 656.400 366.900 657.600 367.950 ;
        RECT 649.950 366.600 652.050 366.900 ;
        RECT 640.950 350.400 645.600 352.050 ;
        RECT 647.400 365.400 652.050 366.600 ;
        RECT 640.950 349.950 645.000 350.400 ;
        RECT 616.950 346.950 619.050 349.050 ;
        RECT 622.950 346.950 625.050 349.050 ;
        RECT 628.950 346.950 631.050 349.050 ;
        RECT 643.950 346.950 646.050 349.050 ;
        RECT 613.950 340.950 616.050 343.050 ;
        RECT 610.950 337.950 613.050 340.050 ;
        RECT 617.400 337.050 618.600 346.950 ;
        RECT 623.400 337.050 624.600 346.950 ;
        RECT 616.950 334.950 619.050 337.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 610.950 331.950 613.050 334.050 ;
        RECT 620.400 333.900 621.600 334.950 ;
        RECT 611.400 319.050 612.600 331.950 ;
        RECT 619.950 331.800 622.050 333.900 ;
        RECT 610.950 316.950 613.050 319.050 ;
        RECT 620.400 300.600 621.600 331.800 ;
        RECT 622.950 301.950 625.050 304.050 ;
        RECT 617.400 299.400 621.600 300.600 ;
        RECT 617.400 292.050 618.600 299.400 ;
        RECT 623.400 292.050 624.600 301.950 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 616.950 289.950 619.050 292.050 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 622.950 289.950 625.050 292.050 ;
        RECT 614.400 288.900 615.600 289.950 ;
        RECT 613.950 286.800 616.050 288.900 ;
        RECT 595.950 277.800 598.050 279.900 ;
        RECT 607.950 277.950 610.050 280.050 ;
        RECT 587.400 263.400 591.600 264.600 ;
        RECT 590.400 262.200 591.600 263.400 ;
        RECT 568.950 259.950 571.050 262.050 ;
        RECT 574.950 260.100 577.050 262.200 ;
        RECT 583.950 260.100 586.050 262.200 ;
        RECT 589.950 260.100 592.050 262.200 ;
        RECT 596.400 262.050 597.600 277.800 ;
        RECT 607.950 274.800 610.050 276.900 ;
        RECT 598.950 268.950 601.050 271.050 ;
        RECT 575.400 259.050 576.600 260.100 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 568.950 253.950 571.050 256.050 ;
        RECT 569.400 229.050 570.600 253.950 ;
        RECT 572.400 241.050 573.600 256.950 ;
        RECT 578.400 255.900 579.600 256.950 ;
        RECT 577.950 253.800 580.050 255.900 ;
        RECT 584.400 249.600 585.600 260.100 ;
        RECT 590.400 259.050 591.600 260.100 ;
        RECT 595.950 259.950 598.050 262.050 ;
        RECT 589.950 256.950 592.050 259.050 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 586.950 253.950 589.050 256.050 ;
        RECT 581.400 248.400 585.600 249.600 ;
        RECT 571.950 238.950 574.050 241.050 ;
        RECT 577.950 238.950 580.050 241.050 ;
        RECT 568.950 226.950 571.050 229.050 ;
        RECT 565.950 215.100 568.050 217.200 ;
        RECT 571.950 215.100 574.050 217.200 ;
        RECT 572.400 214.050 573.600 215.100 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 571.950 211.950 574.050 214.050 ;
        RECT 565.950 205.950 568.050 208.050 ;
        RECT 566.400 184.050 567.600 205.950 ;
        RECT 569.400 205.050 570.600 211.950 ;
        RECT 578.400 205.050 579.600 238.950 ;
        RECT 568.950 202.950 571.050 205.050 ;
        RECT 577.950 202.950 580.050 205.050 ;
        RECT 581.400 202.050 582.600 248.400 ;
        RECT 587.400 244.050 588.600 253.950 ;
        RECT 586.950 241.950 589.050 244.050 ;
        RECT 593.400 220.050 594.600 256.950 ;
        RECT 595.950 253.950 598.050 256.050 ;
        RECT 592.950 217.950 595.050 220.050 ;
        RECT 596.400 217.200 597.600 253.950 ;
        RECT 589.950 215.100 592.050 217.200 ;
        RECT 595.950 215.100 598.050 217.200 ;
        RECT 599.400 216.600 600.600 268.950 ;
        RECT 608.400 265.050 609.600 274.800 ;
        RECT 610.950 268.950 613.050 271.050 ;
        RECT 620.400 270.600 621.600 289.950 ;
        RECT 620.400 269.400 624.600 270.600 ;
        RECT 607.950 262.950 610.050 265.050 ;
        RECT 604.950 260.100 607.050 262.200 ;
        RECT 605.400 259.050 606.600 260.100 ;
        RECT 611.400 259.050 612.600 268.950 ;
        RECT 619.950 265.950 622.050 268.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 610.950 256.950 613.050 259.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 608.400 255.900 609.600 256.950 ;
        RECT 607.950 253.800 610.050 255.900 ;
        RECT 614.400 255.000 615.600 256.950 ;
        RECT 620.400 255.900 621.600 265.950 ;
        RECT 623.400 262.050 624.600 269.400 ;
        RECT 629.400 265.050 630.600 346.950 ;
        RECT 631.950 340.950 634.050 343.050 ;
        RECT 632.400 313.050 633.600 340.950 ;
        RECT 637.950 338.100 640.050 343.050 ;
        RECT 638.400 337.050 639.600 338.100 ;
        RECT 644.400 337.050 645.600 346.950 ;
        RECT 647.400 340.050 648.600 365.400 ;
        RECT 649.950 364.800 652.050 365.400 ;
        RECT 655.950 364.800 658.050 366.900 ;
        RECT 658.950 364.950 661.050 367.050 ;
        RECT 662.400 366.900 663.600 403.950 ;
        RECT 668.400 394.050 669.600 415.950 ;
        RECT 677.400 415.050 678.600 416.100 ;
        RECT 683.400 415.050 684.600 421.950 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 682.950 412.950 685.050 415.050 ;
        RECT 667.950 391.950 670.050 394.050 ;
        RECT 674.400 385.050 675.600 412.950 ;
        RECT 685.950 409.950 688.050 412.050 ;
        RECT 686.400 406.050 687.600 409.950 ;
        RECT 685.950 403.950 688.050 406.050 ;
        RECT 673.950 382.950 676.050 385.050 ;
        RECT 667.950 379.950 670.050 382.050 ;
        RECT 668.400 373.200 669.600 379.950 ;
        RECT 673.950 376.950 676.050 379.050 ;
        RECT 667.950 371.100 670.050 373.200 ;
        RECT 668.400 370.050 669.600 371.100 ;
        RECT 674.400 370.050 675.600 376.950 ;
        RECT 689.400 376.200 690.600 427.950 ;
        RECT 698.400 424.050 699.600 442.950 ;
        RECT 701.400 432.600 702.600 443.400 ;
        RECT 703.950 442.500 706.050 443.400 ;
        RECT 707.850 438.600 709.050 453.600 ;
        RECT 706.950 436.500 709.050 438.600 ;
        RECT 701.400 431.400 705.600 432.600 ;
        RECT 700.950 427.950 703.050 430.050 ;
        RECT 697.950 421.950 700.050 424.050 ;
        RECT 701.400 415.050 702.600 427.950 ;
        RECT 704.400 418.050 705.600 431.400 ;
        RECT 713.400 430.050 714.600 478.950 ;
        RECT 712.950 427.950 715.050 430.050 ;
        RECT 716.400 427.050 717.600 481.950 ;
        RECT 718.950 466.950 721.050 469.050 ;
        RECT 719.400 451.050 720.600 466.950 ;
        RECT 718.950 448.950 721.050 451.050 ;
        RECT 722.400 448.050 723.600 485.400 ;
        RECT 728.400 466.050 729.600 509.400 ;
        RECT 734.400 505.050 735.600 532.950 ;
        RECT 740.400 526.050 741.600 562.650 ;
        RECT 752.400 562.050 753.600 577.950 ;
        RECT 754.950 574.950 757.050 577.050 ;
        RECT 751.950 559.950 754.050 562.050 ;
        RECT 755.400 553.050 756.600 574.950 ;
        RECT 763.950 572.100 766.050 574.200 ;
        RECT 764.400 571.050 765.600 572.100 ;
        RECT 760.950 568.950 763.050 571.050 ;
        RECT 763.950 568.950 766.050 571.050 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 781.950 568.950 784.050 571.050 ;
        RECT 757.950 565.950 760.050 568.050 ;
        RECT 754.950 550.950 757.050 553.050 ;
        RECT 751.950 547.950 754.050 550.050 ;
        RECT 752.400 544.050 753.600 547.950 ;
        RECT 751.950 541.950 754.050 544.050 ;
        RECT 758.400 543.600 759.600 565.950 ;
        RECT 761.400 556.050 762.600 568.950 ;
        RECT 770.400 567.600 771.600 568.950 ;
        RECT 770.400 566.400 774.600 567.600 ;
        RECT 769.950 559.950 772.050 562.050 ;
        RECT 760.950 553.950 763.050 556.050 ;
        RECT 755.400 542.400 759.600 543.600 ;
        RECT 745.950 536.400 748.050 538.500 ;
        RECT 739.950 523.950 742.050 526.050 ;
        RECT 746.100 516.600 747.300 536.400 ;
        RECT 752.400 534.600 753.600 541.950 ;
        RECT 749.400 533.400 753.600 534.600 ;
        RECT 749.400 529.500 750.600 533.400 ;
        RECT 748.950 527.400 751.050 529.500 ;
        RECT 755.400 529.050 756.600 542.400 ;
        RECT 760.950 537.300 763.050 539.400 ;
        RECT 761.850 533.700 763.050 537.300 ;
        RECT 760.950 531.600 763.050 533.700 ;
        RECT 766.950 532.950 769.050 535.050 ;
        RECT 749.400 526.050 750.600 527.400 ;
        RECT 754.950 526.950 757.050 529.050 ;
        RECT 748.950 523.950 751.050 526.050 ;
        RECT 757.950 523.950 760.050 526.050 ;
        RECT 751.800 520.950 753.900 523.050 ;
        RECT 758.400 522.600 759.600 523.950 ;
        RECT 755.400 521.400 760.050 522.600 ;
        RECT 745.950 514.500 748.050 516.600 ;
        RECT 752.400 510.600 753.600 520.950 ;
        RECT 749.400 509.400 753.600 510.600 ;
        RECT 733.950 502.950 736.050 505.050 ;
        RECT 730.950 493.950 733.050 499.050 ;
        RECT 736.950 495.000 739.050 499.050 ;
        RECT 737.400 493.050 738.600 495.000 ;
        RECT 745.950 493.950 748.050 496.050 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 734.400 489.600 735.600 490.950 ;
        RECT 740.400 489.900 741.600 490.950 ;
        RECT 731.400 488.400 735.600 489.600 ;
        RECT 731.400 478.050 732.600 488.400 ;
        RECT 739.950 484.950 742.050 489.900 ;
        RECT 746.400 489.600 747.600 493.950 ;
        RECT 743.400 488.400 747.600 489.600 ;
        RECT 743.400 478.050 744.600 488.400 ;
        RECT 745.950 484.950 748.050 487.050 ;
        RECT 730.950 475.950 733.050 478.050 ;
        RECT 742.950 475.950 745.050 478.050 ;
        RECT 733.950 472.950 736.050 475.050 ;
        RECT 739.950 472.950 742.050 475.050 ;
        RECT 727.950 463.950 730.050 466.050 ;
        RECT 727.950 458.400 730.050 460.500 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 728.100 438.600 729.300 458.400 ;
        RECT 730.950 454.950 733.050 457.050 ;
        RECT 731.400 451.500 732.600 454.950 ;
        RECT 734.400 454.050 735.600 472.950 ;
        RECT 736.950 466.950 739.050 469.050 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 730.950 449.400 733.050 451.500 ;
        RECT 731.400 448.050 732.600 449.400 ;
        RECT 730.950 445.950 733.050 448.050 ;
        RECT 733.950 442.800 736.050 444.900 ;
        RECT 727.950 436.500 730.050 438.600 ;
        RECT 734.400 436.050 735.600 442.800 ;
        RECT 733.950 433.950 736.050 436.050 ;
        RECT 724.950 427.950 727.050 430.050 ;
        RECT 709.950 424.950 712.050 427.050 ;
        RECT 715.950 424.950 718.050 427.050 ;
        RECT 706.950 421.950 709.050 424.050 ;
        RECT 703.950 415.950 706.050 418.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 698.400 411.900 699.600 412.950 ;
        RECT 697.950 409.800 700.050 411.900 ;
        RECT 703.950 409.950 706.050 412.050 ;
        RECT 704.400 396.600 705.600 409.950 ;
        RECT 707.400 397.050 708.600 421.950 ;
        RECT 701.400 395.400 705.600 396.600 ;
        RECT 694.950 391.950 697.050 394.050 ;
        RECT 691.950 388.950 694.050 391.050 ;
        RECT 692.400 382.050 693.600 388.950 ;
        RECT 691.950 379.950 694.050 382.050 ;
        RECT 695.400 379.050 696.600 391.950 ;
        RECT 694.950 376.950 697.050 379.050 ;
        RECT 682.950 373.950 685.050 376.050 ;
        RECT 688.950 374.100 691.050 376.200 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 670.950 367.950 673.050 370.050 ;
        RECT 673.950 367.950 676.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 671.400 366.900 672.600 367.950 ;
        RECT 652.950 361.950 655.050 364.050 ;
        RECT 653.400 358.050 654.600 361.950 ;
        RECT 652.950 355.950 655.050 358.050 ;
        RECT 649.950 352.950 652.050 355.050 ;
        RECT 646.950 337.950 649.050 340.050 ;
        RECT 637.950 334.950 640.050 337.050 ;
        RECT 640.950 334.950 643.050 337.050 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 641.400 333.900 642.600 334.950 ;
        RECT 640.950 331.800 643.050 333.900 ;
        RECT 650.400 316.050 651.600 352.950 ;
        RECT 653.400 340.050 654.600 355.950 ;
        RECT 652.950 337.950 655.050 340.050 ;
        RECT 659.400 337.050 660.600 364.950 ;
        RECT 661.950 364.800 664.050 366.900 ;
        RECT 670.950 364.800 673.050 366.900 ;
        RECT 680.400 352.050 681.600 367.950 ;
        RECT 670.950 349.950 673.050 352.050 ;
        RECT 679.950 349.950 682.050 352.050 ;
        RECT 664.950 338.100 667.050 340.200 ;
        RECT 671.400 339.600 672.600 349.950 ;
        RECT 676.950 344.400 679.050 346.500 ;
        RECT 671.400 338.400 675.600 339.600 ;
        RECT 665.400 337.050 666.600 338.100 ;
        RECT 674.400 337.050 675.600 338.400 ;
        RECT 655.950 334.950 658.050 337.050 ;
        RECT 658.950 334.950 661.050 337.050 ;
        RECT 661.950 334.950 664.050 337.050 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 656.400 325.050 657.600 334.950 ;
        RECT 655.950 322.950 658.050 325.050 ;
        RECT 649.950 313.950 652.050 316.050 ;
        RECT 662.400 313.050 663.600 334.950 ;
        RECT 668.400 319.050 669.600 334.950 ;
        RECT 670.950 331.950 673.050 334.050 ;
        RECT 667.950 316.950 670.050 319.050 ;
        RECT 631.950 310.950 634.050 313.050 ;
        RECT 661.950 310.950 664.050 313.050 ;
        RECT 671.400 304.050 672.600 331.950 ;
        RECT 677.850 329.400 679.050 344.400 ;
        RECT 676.950 327.300 679.050 329.400 ;
        RECT 677.850 323.700 679.050 327.300 ;
        RECT 676.950 321.600 679.050 323.700 ;
        RECT 673.950 316.950 676.050 319.050 ;
        RECT 670.950 301.950 673.050 304.050 ;
        RECT 637.950 300.600 640.050 301.050 ;
        RECT 632.400 299.400 640.050 300.600 ;
        RECT 632.400 295.050 633.600 299.400 ;
        RECT 637.950 298.950 640.050 299.400 ;
        RECT 646.950 298.950 649.050 301.050 ;
        RECT 631.950 292.950 634.050 295.050 ;
        RECT 640.950 293.100 643.050 295.200 ;
        RECT 647.400 295.050 648.600 298.950 ;
        RECT 670.950 298.800 673.050 300.900 ;
        RECT 641.400 292.050 642.600 293.100 ;
        RECT 646.950 292.950 649.050 295.050 ;
        RECT 658.950 293.100 661.050 295.200 ;
        RECT 664.950 293.100 667.050 295.200 ;
        RECT 659.400 292.050 660.600 293.100 ;
        RECT 665.400 292.050 666.600 293.100 ;
        RECT 637.950 289.950 640.050 292.050 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 655.950 289.950 658.050 292.050 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 638.400 288.900 639.600 289.950 ;
        RECT 637.950 286.800 640.050 288.900 ;
        RECT 644.400 283.050 645.600 289.950 ;
        RECT 646.950 286.950 649.050 289.050 ;
        RECT 631.950 280.950 634.050 283.050 ;
        RECT 643.950 280.950 646.050 283.050 ;
        RECT 628.950 262.950 631.050 265.050 ;
        RECT 622.950 259.950 625.050 262.050 ;
        RECT 632.400 261.600 633.600 280.950 ;
        RECT 640.950 277.950 643.050 280.050 ;
        RECT 629.400 260.400 633.600 261.600 ;
        RECT 629.400 259.050 630.600 260.400 ;
        RECT 625.950 256.950 628.050 259.050 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 604.950 250.950 607.050 253.050 ;
        RECT 613.950 250.950 616.050 255.000 ;
        RECT 619.950 253.800 622.050 255.900 ;
        RECT 622.950 253.950 625.050 256.050 ;
        RECT 626.400 255.900 627.600 256.950 ;
        RECT 599.400 215.400 603.600 216.600 ;
        RECT 590.400 214.050 591.600 215.100 ;
        RECT 596.400 214.050 597.600 215.100 ;
        RECT 586.950 211.950 589.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 595.950 211.950 598.050 214.050 ;
        RECT 587.400 210.900 588.600 211.950 ;
        RECT 586.950 208.800 589.050 210.900 ;
        RECT 580.950 199.950 583.050 202.050 ;
        RECT 587.400 199.050 588.600 208.800 ;
        RECT 593.400 205.050 594.600 211.950 ;
        RECT 592.950 202.950 595.050 205.050 ;
        RECT 586.950 196.950 589.050 199.050 ;
        RECT 602.400 190.050 603.600 215.400 ;
        RECT 605.400 210.900 606.600 250.950 ;
        RECT 623.400 250.050 624.600 253.950 ;
        RECT 625.950 253.800 628.050 255.900 ;
        RECT 635.400 255.000 636.600 256.950 ;
        RECT 634.950 250.950 637.050 255.000 ;
        RECT 622.950 247.950 625.050 250.050 ;
        RECT 625.950 226.950 628.050 229.050 ;
        RECT 610.950 215.100 613.050 217.200 ;
        RECT 619.950 215.100 622.050 217.200 ;
        RECT 611.400 214.050 612.600 215.100 ;
        RECT 620.400 214.050 621.600 215.100 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 619.950 211.950 622.050 214.050 ;
        RECT 614.400 210.900 615.600 211.950 ;
        RECT 604.950 208.800 607.050 210.900 ;
        RECT 613.950 208.800 616.050 210.900 ;
        RECT 626.400 193.050 627.600 226.950 ;
        RECT 641.400 223.050 642.600 277.950 ;
        RECT 647.400 274.050 648.600 286.950 ;
        RECT 649.950 283.950 652.050 288.900 ;
        RECT 656.400 288.000 657.600 289.950 ;
        RECT 655.950 283.950 658.050 288.000 ;
        RECT 662.400 280.050 663.600 289.950 ;
        RECT 664.950 283.950 667.050 286.050 ;
        RECT 661.950 277.950 664.050 280.050 ;
        RECT 646.950 271.950 649.050 274.050 ;
        RECT 643.950 262.950 646.050 265.050 ;
        RECT 644.400 235.050 645.600 262.950 ;
        RECT 652.950 260.100 655.050 262.200 ;
        RECT 653.400 259.050 654.600 260.100 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 650.400 244.050 651.600 256.950 ;
        RECT 652.950 247.950 655.050 250.050 ;
        RECT 649.950 241.950 652.050 244.050 ;
        RECT 653.400 238.050 654.600 247.950 ;
        RECT 656.400 241.050 657.600 256.950 ;
        RECT 665.400 253.050 666.600 283.950 ;
        RECT 671.400 280.050 672.600 298.800 ;
        RECT 674.400 286.050 675.600 316.950 ;
        RECT 683.400 304.050 684.600 373.950 ;
        RECT 688.950 370.950 691.050 373.050 ;
        RECT 689.400 370.050 690.600 370.950 ;
        RECT 695.400 370.050 696.600 376.950 ;
        RECT 701.400 373.050 702.600 395.400 ;
        RECT 706.950 394.950 709.050 397.050 ;
        RECT 710.400 393.600 711.600 424.950 ;
        RECT 721.950 421.950 724.050 424.050 ;
        RECT 715.950 416.100 718.050 418.200 ;
        RECT 716.400 415.050 717.600 416.100 ;
        RECT 722.400 415.050 723.600 421.950 ;
        RECT 725.400 418.050 726.600 427.950 ;
        RECT 730.950 422.400 733.050 424.500 ;
        RECT 737.400 424.050 738.600 466.950 ;
        RECT 740.400 445.050 741.600 472.950 ;
        RECT 746.400 463.050 747.600 484.950 ;
        RECT 749.400 484.050 750.600 509.400 ;
        RECT 755.400 505.050 756.600 521.400 ;
        RECT 757.950 520.500 760.050 521.400 ;
        RECT 761.850 516.600 763.050 531.600 ;
        RECT 760.950 514.500 763.050 516.600 ;
        RECT 760.950 508.950 763.050 511.050 ;
        RECT 754.950 502.950 757.050 505.050 ;
        RECT 761.400 493.050 762.600 508.950 ;
        RECT 757.950 490.950 760.050 493.050 ;
        RECT 760.950 490.950 763.050 493.050 ;
        RECT 751.950 484.950 754.050 490.050 ;
        RECT 748.950 481.950 751.050 484.050 ;
        RECT 754.950 481.950 757.050 484.050 ;
        RECT 745.950 460.950 748.050 463.050 ;
        RECT 746.400 457.050 747.600 460.950 ;
        RECT 745.950 454.950 748.050 457.050 ;
        RECT 751.950 454.950 754.050 457.050 ;
        RECT 742.950 448.950 745.050 451.050 ;
        RECT 748.800 449.100 750.900 451.200 ;
        RECT 752.400 451.050 753.600 454.950 ;
        RECT 739.950 442.950 742.050 445.050 ;
        RECT 724.950 415.950 727.050 418.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 712.950 409.950 715.050 412.050 ;
        RECT 707.400 392.400 711.600 393.600 ;
        RECT 700.950 370.950 703.050 373.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 691.950 367.950 694.050 370.050 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 697.950 367.950 700.050 370.050 ;
        RECT 692.400 342.600 693.600 367.950 ;
        RECT 698.400 366.900 699.600 367.950 ;
        RECT 697.950 364.800 700.050 366.900 ;
        RECT 698.400 358.050 699.600 364.800 ;
        RECT 707.400 364.050 708.600 392.400 ;
        RECT 713.400 385.050 714.600 409.950 ;
        RECT 719.400 406.050 720.600 412.950 ;
        RECT 724.950 409.950 727.050 412.050 ;
        RECT 728.400 411.000 729.600 412.950 ;
        RECT 721.950 406.950 724.050 409.050 ;
        RECT 718.950 403.950 721.050 406.050 ;
        RECT 722.400 403.050 723.600 406.950 ;
        RECT 721.950 400.950 724.050 403.050 ;
        RECT 712.950 382.950 715.050 385.050 ;
        RECT 715.950 371.100 718.050 373.200 ;
        RECT 722.400 373.050 723.600 400.950 ;
        RECT 725.400 376.050 726.600 409.950 ;
        RECT 727.950 406.950 730.050 411.000 ;
        RECT 731.700 402.600 732.900 422.400 ;
        RECT 736.950 421.950 739.050 424.050 ;
        RECT 736.950 412.950 739.050 415.050 ;
        RECT 737.400 411.600 738.600 412.950 ;
        RECT 736.950 409.500 739.050 411.600 ;
        RECT 743.400 409.050 744.600 448.950 ;
        RECT 749.400 448.050 750.600 449.100 ;
        RECT 751.950 448.950 754.050 451.050 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 745.950 442.950 748.050 445.050 ;
        RECT 742.950 406.950 745.050 409.050 ;
        RECT 746.400 405.600 747.600 442.950 ;
        RECT 755.400 442.050 756.600 481.950 ;
        RECT 758.400 469.050 759.600 490.950 ;
        RECT 763.950 487.950 766.050 490.050 ;
        RECT 764.400 475.050 765.600 487.950 ;
        RECT 763.950 472.950 766.050 475.050 ;
        RECT 767.400 471.600 768.600 532.950 ;
        RECT 770.400 511.050 771.600 559.950 ;
        RECT 773.400 559.050 774.600 566.400 ;
        RECT 772.950 556.950 775.050 559.050 ;
        RECT 772.950 550.950 775.050 553.050 ;
        RECT 773.400 529.050 774.600 550.950 ;
        RECT 782.400 544.050 783.600 568.950 ;
        RECT 788.400 568.050 789.600 586.950 ;
        RECT 790.950 583.950 793.050 586.050 ;
        RECT 791.400 577.050 792.600 583.950 ;
        RECT 793.950 580.950 796.050 583.050 ;
        RECT 790.950 574.950 793.050 577.050 ;
        RECT 787.950 565.950 790.050 568.050 ;
        RECT 791.400 564.600 792.600 574.950 ;
        RECT 788.400 563.400 792.600 564.600 ;
        RECT 788.400 550.050 789.600 563.400 ;
        RECT 787.950 547.950 790.050 550.050 ;
        RECT 781.950 541.950 784.050 544.050 ;
        RECT 787.950 541.950 790.050 544.050 ;
        RECT 781.950 536.400 784.050 538.500 ;
        RECT 772.950 526.950 775.050 529.050 ;
        RECT 777.000 528.600 781.050 529.050 ;
        RECT 776.400 526.950 781.050 528.600 ;
        RECT 776.400 526.050 777.600 526.950 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 772.950 520.950 775.050 523.050 ;
        RECT 769.950 508.950 772.050 511.050 ;
        RECT 769.950 502.950 772.050 505.050 ;
        RECT 770.400 481.050 771.600 502.950 ;
        RECT 773.400 499.050 774.600 520.950 ;
        RECT 782.100 516.600 783.300 536.400 ;
        RECT 788.400 528.600 789.600 541.950 ;
        RECT 794.400 535.050 795.600 580.950 ;
        RECT 806.400 574.050 807.600 607.950 ;
        RECT 809.400 607.050 810.600 619.950 ;
        RECT 821.400 616.050 822.600 640.650 ;
        RECT 827.400 628.050 828.600 649.950 ;
        RECT 830.400 645.900 831.600 673.950 ;
        RECT 833.400 652.050 834.600 673.950 ;
        RECT 836.400 670.050 837.600 679.950 ;
        RECT 844.950 676.950 847.050 679.050 ;
        RECT 835.950 667.950 838.050 670.050 ;
        RECT 845.400 664.050 846.600 676.950 ;
        RECT 838.950 661.950 841.050 664.050 ;
        RECT 844.950 661.950 847.050 664.050 ;
        RECT 832.950 649.950 835.050 652.050 ;
        RECT 839.400 649.050 840.600 661.950 ;
        RECT 844.950 655.950 847.050 658.050 ;
        RECT 845.400 649.050 846.600 655.950 ;
        RECT 848.400 655.050 849.600 691.950 ;
        RECT 847.950 652.950 850.050 655.050 ;
        RECT 835.950 646.950 838.050 649.050 ;
        RECT 838.950 646.950 841.050 649.050 ;
        RECT 841.950 646.950 844.050 649.050 ;
        RECT 844.950 646.950 847.050 649.050 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 836.400 645.900 837.600 646.950 ;
        RECT 829.950 643.800 832.050 645.900 ;
        RECT 835.950 643.800 838.050 645.900 ;
        RECT 842.400 645.000 843.600 646.950 ;
        RECT 841.950 640.950 844.050 645.000 ;
        RECT 844.950 640.950 847.050 643.050 ;
        RECT 832.950 634.950 835.050 637.050 ;
        RECT 826.950 625.950 829.050 628.050 ;
        RECT 829.950 619.950 832.050 622.050 ;
        RECT 820.950 613.950 823.050 616.050 ;
        RECT 814.800 609.300 816.900 611.400 ;
        RECT 824.400 610.500 826.500 612.600 ;
        RECT 808.950 604.950 811.050 607.050 ;
        RECT 812.400 604.050 813.600 606.600 ;
        RECT 808.950 601.800 811.050 603.900 ;
        RECT 812.400 601.950 814.500 604.050 ;
        RECT 805.950 571.950 808.050 574.050 ;
        RECT 796.950 562.950 799.050 565.050 ;
        RECT 793.950 532.950 796.050 535.050 ;
        RECT 785.400 527.400 789.600 528.600 ;
        RECT 785.400 526.050 786.600 527.400 ;
        RECT 784.950 523.950 787.050 526.050 ;
        RECT 787.950 520.950 790.050 523.050 ;
        RECT 781.950 514.500 784.050 516.600 ;
        RECT 788.400 511.050 789.600 520.950 ;
        RECT 787.950 508.950 790.050 511.050 ;
        RECT 787.950 505.800 790.050 507.900 ;
        RECT 781.950 499.950 784.050 502.050 ;
        RECT 772.950 496.950 775.050 499.050 ;
        RECT 782.400 493.050 783.600 499.950 ;
        RECT 788.400 493.050 789.600 505.800 ;
        RECT 797.400 502.050 798.600 562.950 ;
        RECT 809.400 529.050 810.600 601.800 ;
        RECT 815.700 600.300 816.600 609.300 ;
        RECT 818.100 605.700 820.200 607.800 ;
        RECT 821.400 606.900 822.600 609.450 ;
        RECT 819.300 603.300 820.200 605.700 ;
        RECT 821.100 604.800 823.200 606.900 ;
        RECT 825.000 603.300 826.050 610.500 ;
        RECT 830.400 610.050 831.600 619.950 ;
        RECT 829.950 607.950 832.050 610.050 ;
        RECT 833.400 604.050 834.600 634.950 ;
        RECT 835.950 625.950 838.050 628.050 ;
        RECT 819.300 602.100 826.050 603.300 ;
        RECT 822.150 600.300 824.250 601.200 ;
        RECT 815.700 599.100 824.250 600.300 ;
        RECT 817.200 597.300 819.300 599.100 ;
        RECT 821.100 596.100 823.200 598.200 ;
        RECT 825.150 596.700 826.050 602.100 ;
        RECT 826.950 601.950 829.050 604.050 ;
        RECT 832.950 601.950 835.050 604.050 ;
        RECT 827.400 599.400 828.600 601.950 ;
        RECT 821.400 580.050 822.600 596.100 ;
        RECT 824.400 594.600 826.500 596.700 ;
        RECT 811.950 577.950 814.050 580.050 ;
        RECT 820.950 577.950 823.050 580.050 ;
        RECT 829.950 577.950 832.050 580.050 ;
        RECT 812.400 562.050 813.600 577.950 ;
        RECT 817.950 572.100 820.050 574.200 ;
        RECT 823.950 573.000 826.050 577.050 ;
        RECT 826.950 574.050 829.050 574.200 ;
        RECT 830.400 574.050 831.600 577.950 ;
        RECT 818.400 571.050 819.600 572.100 ;
        RECT 824.400 571.050 825.600 573.000 ;
        RECT 826.950 572.100 831.600 574.050 ;
        RECT 836.400 573.600 837.600 625.950 ;
        RECT 841.950 610.950 844.050 613.050 ;
        RECT 842.400 607.050 843.600 610.950 ;
        RECT 841.950 604.950 844.050 607.050 ;
        RECT 845.400 604.050 846.600 640.950 ;
        RECT 848.400 634.050 849.600 646.950 ;
        RECT 847.950 631.950 850.050 634.050 ;
        RECT 854.400 610.050 855.600 698.400 ;
        RECT 875.400 697.050 876.600 721.800 ;
        RECT 883.950 697.950 886.050 700.050 ;
        RECT 856.950 694.950 859.050 697.050 ;
        RECT 874.950 694.950 877.050 697.050 ;
        RECT 857.400 688.050 858.600 694.950 ;
        RECT 862.500 688.500 864.600 690.600 ;
        RECT 856.950 685.950 859.050 688.050 ;
        RECT 859.950 679.950 862.050 682.050 ;
        RECT 862.950 681.300 864.000 688.500 ;
        RECT 866.400 684.900 867.600 687.450 ;
        RECT 872.100 687.300 874.200 689.400 ;
        RECT 865.800 682.800 867.900 684.900 ;
        RECT 868.800 683.700 870.900 685.800 ;
        RECT 868.800 681.300 869.700 683.700 ;
        RECT 862.950 680.100 869.700 681.300 ;
        RECT 860.400 677.400 861.600 679.950 ;
        RECT 856.950 673.950 859.050 676.050 ;
        RECT 862.950 674.700 863.850 680.100 ;
        RECT 864.750 678.300 866.850 679.200 ;
        RECT 872.400 678.300 873.300 687.300 ;
        RECT 884.400 685.050 885.600 697.950 ;
        RECT 887.400 694.050 888.600 748.950 ;
        RECT 902.400 739.050 903.600 757.950 ;
        RECT 911.400 751.050 912.600 761.100 ;
        RECT 914.400 754.050 915.600 766.950 ;
        RECT 913.950 751.950 916.050 754.050 ;
        RECT 910.950 748.950 913.050 751.050 ;
        RECT 901.950 736.950 904.050 739.050 ;
        RECT 899.400 732.900 900.600 735.450 ;
        RECT 895.200 729.900 897.300 731.700 ;
        RECT 899.100 730.800 901.200 732.900 ;
        RECT 902.400 732.300 904.500 734.400 ;
        RECT 893.700 728.700 902.250 729.900 ;
        RECT 890.400 724.950 892.500 727.050 ;
        RECT 890.400 722.400 891.600 724.950 ;
        RECT 893.700 719.700 894.600 728.700 ;
        RECT 900.150 727.800 902.250 728.700 ;
        RECT 903.150 726.900 904.050 732.300 ;
        RECT 913.950 729.600 916.050 730.050 ;
        RECT 917.400 729.600 918.600 799.950 ;
        RECT 919.950 733.950 922.050 736.050 ;
        RECT 905.400 727.050 906.600 729.600 ;
        RECT 913.950 728.400 918.600 729.600 ;
        RECT 913.950 727.950 916.050 728.400 ;
        RECT 897.300 725.700 904.050 726.900 ;
        RECT 897.300 723.300 898.200 725.700 ;
        RECT 896.100 721.200 898.200 723.300 ;
        RECT 899.100 722.100 901.200 724.200 ;
        RECT 892.800 717.600 894.900 719.700 ;
        RECT 899.400 719.550 900.600 722.100 ;
        RECT 903.000 718.500 904.050 725.700 ;
        RECT 904.950 724.950 907.050 727.050 ;
        RECT 910.950 724.950 913.050 727.050 ;
        RECT 911.400 720.600 912.600 724.950 ;
        RECT 908.400 719.400 912.600 720.600 ;
        RECT 902.400 716.400 904.500 718.500 ;
        RECT 908.400 715.050 909.600 719.400 ;
        RECT 907.950 712.950 910.050 715.050 ;
        RECT 898.950 706.950 901.050 709.050 ;
        RECT 886.950 691.950 889.050 694.050 ;
        RECT 899.400 688.050 900.600 706.950 ;
        RECT 914.400 700.050 915.600 727.950 ;
        RECT 913.950 697.950 916.050 700.050 ;
        RECT 920.400 688.050 921.600 733.950 ;
        RECT 898.950 685.950 901.050 688.050 ;
        RECT 919.950 685.950 922.050 688.050 ;
        RECT 875.400 682.050 876.600 684.600 ;
        RECT 883.950 682.950 886.050 685.050 ;
        RECT 889.950 683.100 892.050 685.200 ;
        RECT 899.400 683.400 906.600 684.600 ;
        RECT 890.400 682.050 891.600 683.100 ;
        RECT 874.500 679.950 876.600 682.050 ;
        RECT 886.950 679.950 889.050 682.050 ;
        RECT 889.950 679.950 892.050 682.050 ;
        RECT 892.950 679.950 895.050 682.050 ;
        RECT 864.750 677.100 873.300 678.300 ;
        RECT 857.400 667.050 858.600 673.950 ;
        RECT 862.500 672.600 864.600 674.700 ;
        RECT 865.800 674.100 867.900 676.200 ;
        RECT 869.700 675.300 871.800 677.100 ;
        RECT 883.950 676.950 886.050 679.050 ;
        RECT 887.400 678.900 888.600 679.950 ;
        RECT 856.950 664.950 859.050 667.050 ;
        RECT 866.400 661.050 867.600 674.100 ;
        RECT 884.400 673.050 885.600 676.950 ;
        RECT 886.950 676.800 889.050 678.900 ;
        RECT 883.950 670.950 886.050 673.050 ;
        RECT 871.950 664.950 874.050 667.050 ;
        RECT 856.950 658.950 859.050 661.050 ;
        RECT 865.950 658.950 868.050 661.050 ;
        RECT 857.400 652.050 858.600 658.950 ;
        RECT 856.950 649.950 859.050 652.050 ;
        RECT 859.950 651.000 862.050 655.050 ;
        RECT 860.400 649.050 861.600 651.000 ;
        RECT 865.950 650.100 868.050 652.200 ;
        RECT 872.400 652.050 873.600 664.950 ;
        RECT 887.400 655.050 888.600 676.800 ;
        RECT 893.400 664.050 894.600 679.950 ;
        RECT 895.950 676.950 898.050 679.050 ;
        RECT 892.950 661.950 895.050 664.050 ;
        RECT 889.950 655.950 892.050 658.050 ;
        RECT 886.950 652.950 889.050 655.050 ;
        RECT 866.400 649.050 867.600 650.100 ;
        RECT 871.950 649.950 874.050 652.050 ;
        RECT 880.950 649.950 883.050 652.050 ;
        RECT 859.950 646.950 862.050 649.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 856.950 643.950 859.050 646.050 ;
        RECT 863.400 645.000 864.600 646.950 ;
        RECT 869.400 645.000 870.600 646.950 ;
        RECT 853.950 607.950 856.050 610.050 ;
        RECT 854.400 606.600 855.600 607.950 ;
        RECT 851.400 605.400 855.600 606.600 ;
        RECT 851.400 604.050 852.600 605.400 ;
        RECT 844.950 601.950 847.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 850.950 601.950 853.050 604.050 ;
        RECT 844.950 580.950 847.050 583.050 ;
        RECT 838.950 577.950 841.050 580.050 ;
        RECT 828.000 571.950 831.600 572.100 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 811.950 559.950 814.050 562.050 ;
        RECT 821.400 559.050 822.600 568.950 ;
        RECT 826.950 559.950 829.050 562.050 ;
        RECT 820.950 556.950 823.050 559.050 ;
        RECT 799.950 528.600 804.000 529.050 ;
        RECT 799.950 526.950 804.600 528.600 ;
        RECT 808.950 526.950 811.050 529.050 ;
        RECT 820.950 528.000 823.050 532.050 ;
        RECT 803.400 526.050 804.600 526.950 ;
        RECT 821.400 526.050 822.600 528.000 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 799.950 520.950 802.050 523.050 ;
        RECT 800.400 508.050 801.600 520.950 ;
        RECT 818.400 514.050 819.600 523.950 ;
        RECT 823.950 517.950 826.050 520.050 ;
        RECT 817.950 511.950 820.050 514.050 ;
        RECT 814.950 508.950 817.050 511.050 ;
        RECT 799.950 505.950 802.050 508.050 ;
        RECT 796.950 499.950 799.050 502.050 ;
        RECT 796.950 494.100 799.050 496.200 ;
        RECT 815.400 496.050 816.600 508.950 ;
        RECT 817.950 505.950 820.050 508.050 ;
        RECT 797.400 493.050 798.600 494.100 ;
        RECT 814.950 493.950 817.050 496.050 ;
        RECT 818.400 493.050 819.600 505.950 ;
        RECT 824.400 499.200 825.600 517.950 ;
        RECT 827.400 511.050 828.600 559.950 ;
        RECT 830.400 532.050 831.600 571.950 ;
        RECT 833.400 572.400 837.600 573.600 ;
        RECT 833.400 541.050 834.600 572.400 ;
        RECT 839.400 571.050 840.600 577.950 ;
        RECT 845.400 571.050 846.600 580.950 ;
        RECT 848.400 577.050 849.600 601.950 ;
        RECT 857.400 580.050 858.600 643.950 ;
        RECT 859.950 640.950 862.050 643.050 ;
        RECT 862.950 640.950 865.050 645.000 ;
        RECT 868.950 640.950 871.050 645.000 ;
        RECT 881.400 643.050 882.600 649.950 ;
        RECT 890.400 649.050 891.600 655.950 ;
        RECT 896.400 652.050 897.600 676.950 ;
        RECT 899.400 670.050 900.600 683.400 ;
        RECT 905.400 682.050 906.600 683.400 ;
        RECT 910.950 683.100 913.050 685.200 ;
        RECT 911.400 682.050 912.600 683.100 ;
        RECT 919.950 682.800 922.050 684.900 ;
        RECT 904.950 679.950 907.050 682.050 ;
        RECT 907.950 679.950 910.050 682.050 ;
        RECT 910.950 679.950 913.050 682.050 ;
        RECT 913.950 679.950 916.050 682.050 ;
        RECT 908.400 678.900 909.600 679.950 ;
        RECT 907.950 676.800 910.050 678.900 ;
        RECT 914.400 673.050 915.600 679.950 ;
        RECT 916.950 676.950 919.050 679.050 ;
        RECT 913.950 670.950 916.050 673.050 ;
        RECT 898.950 667.950 901.050 670.050 ;
        RECT 913.950 667.800 916.050 669.900 ;
        RECT 901.950 661.950 904.050 664.050 ;
        RECT 895.950 649.950 898.050 652.050 ;
        RECT 902.400 649.050 903.600 661.950 ;
        RECT 910.950 655.950 913.050 658.050 ;
        RECT 886.950 646.950 889.050 649.050 ;
        RECT 889.950 646.950 892.050 649.050 ;
        RECT 892.950 646.950 895.050 649.050 ;
        RECT 901.950 646.950 904.050 649.050 ;
        RECT 904.950 646.950 907.050 649.050 ;
        RECT 883.950 643.950 886.050 646.050 ;
        RECT 887.400 645.000 888.600 646.950 ;
        RECT 880.950 640.950 883.050 643.050 ;
        RECT 860.400 607.050 861.600 640.950 ;
        RECT 869.400 619.050 870.600 640.950 ;
        RECT 884.400 625.050 885.600 643.950 ;
        RECT 886.950 640.950 889.050 645.000 ;
        RECT 883.950 622.950 886.050 625.050 ;
        RECT 862.950 616.950 865.050 619.050 ;
        RECT 868.950 616.950 871.050 619.050 ;
        RECT 863.400 613.050 864.600 616.950 ;
        RECT 868.950 613.800 871.050 615.900 ;
        RECT 862.950 610.950 865.050 613.050 ;
        RECT 859.950 604.950 862.050 607.050 ;
        RECT 862.950 606.000 865.050 609.900 ;
        RECT 869.400 607.200 870.600 613.800 ;
        RECT 887.400 610.200 888.600 640.950 ;
        RECT 893.400 637.050 894.600 646.950 ;
        RECT 895.950 643.950 898.050 646.050 ;
        RECT 892.950 634.950 895.050 637.050 ;
        RECT 892.950 616.950 895.050 619.050 ;
        RECT 886.950 608.100 889.050 610.200 ;
        RECT 863.400 604.050 864.600 606.000 ;
        RECT 868.950 605.100 871.050 607.200 ;
        RECT 869.400 604.050 870.600 605.100 ;
        RECT 886.950 604.950 889.050 607.050 ;
        RECT 887.400 604.050 888.600 604.950 ;
        RECT 893.400 604.050 894.600 616.950 ;
        RECT 896.400 607.050 897.600 643.950 ;
        RECT 905.400 637.050 906.600 646.950 ;
        RECT 904.950 636.600 907.050 637.050 ;
        RECT 902.400 635.400 907.050 636.600 ;
        RECT 898.950 607.950 901.050 610.050 ;
        RECT 895.950 604.950 898.050 607.050 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 868.950 601.950 871.050 604.050 ;
        RECT 883.950 601.950 886.050 604.050 ;
        RECT 886.950 601.950 889.050 604.050 ;
        RECT 889.950 601.950 892.050 604.050 ;
        RECT 892.950 601.950 895.050 604.050 ;
        RECT 859.950 598.950 862.050 601.050 ;
        RECT 850.950 577.950 853.050 580.050 ;
        RECT 856.950 577.950 859.050 580.050 ;
        RECT 847.950 574.950 850.050 577.050 ;
        RECT 851.400 574.050 852.600 577.950 ;
        RECT 860.400 574.050 861.600 598.950 ;
        RECT 866.400 595.050 867.600 601.950 ;
        RECT 871.950 598.950 874.050 601.050 ;
        RECT 880.950 598.950 883.050 601.050 ;
        RECT 865.950 592.950 868.050 595.050 ;
        RECT 868.950 580.950 871.050 583.050 ;
        RECT 865.950 577.950 868.050 580.050 ;
        RECT 850.950 571.950 853.050 574.050 ;
        RECT 859.950 571.950 862.050 574.050 ;
        RECT 866.400 571.050 867.600 577.950 ;
        RECT 869.400 577.050 870.600 580.950 ;
        RECT 868.950 574.950 871.050 577.050 ;
        RECT 872.400 574.050 873.600 598.950 ;
        RECT 881.400 595.050 882.600 598.950 ;
        RECT 880.950 592.950 883.050 595.050 ;
        RECT 884.400 580.050 885.600 601.950 ;
        RECT 890.400 595.050 891.600 601.950 ;
        RECT 889.950 592.950 892.050 595.050 ;
        RECT 874.950 577.950 877.050 580.050 ;
        RECT 883.950 577.950 886.050 580.050 ;
        RECT 889.950 577.950 892.050 580.050 ;
        RECT 871.950 571.950 874.050 574.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 844.950 568.950 847.050 571.050 ;
        RECT 847.950 568.950 850.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 865.950 568.950 868.050 571.050 ;
        RECT 868.950 568.950 871.050 571.050 ;
        RECT 835.950 565.950 838.050 568.050 ;
        RECT 842.400 567.900 843.600 568.950 ;
        RECT 832.950 538.950 835.050 541.050 ;
        RECT 836.400 538.050 837.600 565.950 ;
        RECT 841.950 562.950 844.050 567.900 ;
        RECT 848.400 562.050 849.600 568.950 ;
        RECT 859.950 565.950 862.050 568.050 ;
        RECT 863.400 567.000 864.600 568.950 ;
        RECT 869.400 567.900 870.600 568.950 ;
        RECT 847.950 559.950 850.050 562.050 ;
        RECT 838.950 547.950 841.050 550.050 ;
        RECT 835.950 535.950 838.050 538.050 ;
        RECT 829.950 526.950 832.050 532.050 ;
        RECT 839.400 526.050 840.600 547.950 ;
        RECT 860.400 544.050 861.600 565.950 ;
        RECT 862.950 562.950 865.050 567.000 ;
        RECT 868.950 565.800 871.050 567.900 ;
        RECT 865.950 562.950 868.050 565.050 ;
        RECT 859.950 541.950 862.050 544.050 ;
        RECT 856.950 538.950 859.050 541.050 ;
        RECT 857.400 532.050 858.600 538.950 ;
        RECT 856.950 529.950 859.050 532.050 ;
        RECT 866.400 529.200 867.600 562.950 ;
        RECT 868.950 562.650 871.050 564.750 ;
        RECT 869.400 538.050 870.600 562.650 ;
        RECT 868.950 535.950 871.050 538.050 ;
        RECT 859.950 527.100 862.050 529.200 ;
        RECT 865.950 527.100 868.050 529.200 ;
        RECT 860.400 526.050 861.600 527.100 ;
        RECT 866.400 526.050 867.600 527.100 ;
        RECT 871.950 526.950 874.050 529.050 ;
        RECT 835.950 523.950 838.050 526.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 856.950 523.950 859.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 865.950 523.950 868.050 526.050 ;
        RECT 829.950 520.950 832.050 523.050 ;
        RECT 836.400 522.900 837.600 523.950 ;
        RECT 826.950 508.950 829.050 511.050 ;
        RECT 823.950 497.100 826.050 499.200 ;
        RECT 830.400 496.050 831.600 520.950 ;
        RECT 835.950 520.800 838.050 522.900 ;
        RECT 838.950 517.950 841.050 520.050 ;
        RECT 832.950 508.950 835.050 511.050 ;
        RECT 823.950 493.950 826.050 496.050 ;
        RECT 829.950 493.950 832.050 496.050 ;
        RECT 824.400 493.050 825.600 493.950 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 802.950 490.950 805.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 823.950 490.950 826.050 493.050 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 769.950 478.950 772.050 481.050 ;
        RECT 779.400 478.050 780.600 490.950 ;
        RECT 785.400 484.050 786.600 490.950 ;
        RECT 803.400 489.900 804.600 490.950 ;
        RECT 821.400 489.900 822.600 490.950 ;
        RECT 827.400 489.900 828.600 490.950 ;
        RECT 802.950 487.800 805.050 489.900 ;
        RECT 820.950 487.800 823.050 489.900 ;
        RECT 826.950 487.800 829.050 489.900 ;
        RECT 829.950 487.950 832.050 490.050 ;
        RECT 784.950 481.950 787.050 484.050 ;
        RECT 790.950 481.950 793.050 484.050 ;
        RECT 805.950 481.950 808.050 484.050 ;
        RECT 778.950 475.950 781.050 478.050 ;
        RECT 764.400 470.400 768.600 471.600 ;
        RECT 757.950 466.950 760.050 469.050 ;
        RECT 760.950 463.950 763.050 466.050 ;
        RECT 757.950 457.950 760.050 460.050 ;
        RECT 754.950 439.950 757.050 442.050 ;
        RECT 743.400 405.000 747.600 405.600 ;
        RECT 742.950 404.400 747.600 405.000 ;
        RECT 751.950 422.400 754.050 424.500 ;
        RECT 751.950 407.400 753.150 422.400 ;
        RECT 758.400 421.050 759.600 457.950 ;
        RECT 761.400 439.050 762.600 463.950 ;
        RECT 760.950 436.950 763.050 439.050 ;
        RECT 754.950 419.400 759.600 421.050 ;
        RECT 754.950 418.950 759.000 419.400 ;
        RECT 760.950 417.600 763.050 418.050 ;
        RECT 755.400 416.400 763.050 417.600 ;
        RECT 755.400 415.050 756.600 416.400 ;
        RECT 760.950 415.950 763.050 416.400 ;
        RECT 754.950 412.950 757.050 415.050 ;
        RECT 760.950 412.800 763.050 414.900 ;
        RECT 757.950 409.950 760.050 412.050 ;
        RECT 751.950 405.300 754.050 407.400 ;
        RECT 730.950 400.500 733.050 402.600 ;
        RECT 736.950 400.950 739.050 403.050 ;
        RECT 742.950 400.950 745.050 404.400 ;
        RECT 751.950 401.700 753.150 405.300 ;
        RECT 724.950 373.950 727.050 376.050 ;
        RECT 716.400 370.050 717.600 371.100 ;
        RECT 721.950 370.950 724.050 373.050 ;
        RECT 730.950 372.000 733.050 376.050 ;
        RECT 731.400 370.050 732.600 372.000 ;
        RECT 737.400 370.050 738.600 400.950 ;
        RECT 751.950 399.600 754.050 401.700 ;
        RECT 742.950 394.950 745.050 397.050 ;
        RECT 739.950 388.950 742.050 391.050 ;
        RECT 740.400 372.600 741.600 388.950 ;
        RECT 743.400 375.600 744.600 394.950 ;
        RECT 746.400 386.400 753.600 387.600 ;
        RECT 746.400 382.050 747.600 386.400 ;
        RECT 748.950 382.950 751.050 385.050 ;
        RECT 745.950 379.950 748.050 382.050 ;
        RECT 743.400 374.400 747.600 375.600 ;
        RECT 740.400 371.400 744.600 372.600 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 715.950 367.950 718.050 370.050 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 709.950 364.950 712.050 367.050 ;
        RECT 713.400 366.000 714.600 367.950 ;
        RECT 706.950 361.950 709.050 364.050 ;
        RECT 697.950 355.950 700.050 358.050 ;
        RECT 706.950 349.950 709.050 352.050 ;
        RECT 697.950 344.400 700.050 346.500 ;
        RECT 692.400 342.000 696.600 342.600 ;
        RECT 692.400 341.400 697.050 342.000 ;
        RECT 685.950 338.100 688.050 340.200 ;
        RECT 686.400 333.600 687.600 338.100 ;
        RECT 694.950 337.950 697.050 341.400 ;
        RECT 691.950 334.950 694.050 337.050 ;
        RECT 692.400 333.600 693.600 334.950 ;
        RECT 686.400 332.400 690.600 333.600 ;
        RECT 689.400 325.050 690.600 332.400 ;
        RECT 691.950 331.500 694.050 333.600 ;
        RECT 688.950 322.950 691.050 325.050 ;
        RECT 698.100 324.600 699.300 344.400 ;
        RECT 700.950 334.950 703.050 337.050 ;
        RECT 701.400 333.600 702.600 334.950 ;
        RECT 707.400 333.600 708.600 349.950 ;
        RECT 701.400 332.400 708.600 333.600 ;
        RECT 697.950 322.500 700.050 324.600 ;
        RECT 691.950 319.950 694.050 322.050 ;
        RECT 692.400 316.050 693.600 319.950 ;
        RECT 691.950 313.950 694.050 316.050 ;
        RECT 706.950 313.950 709.050 316.050 ;
        RECT 688.950 310.950 691.050 313.050 ;
        RECT 679.950 300.600 682.050 304.050 ;
        RECT 682.950 301.950 685.050 304.050 ;
        RECT 679.950 300.000 684.600 300.600 ;
        RECT 680.400 299.400 684.600 300.000 ;
        RECT 679.950 294.000 682.050 298.050 ;
        RECT 683.400 297.600 684.600 299.400 ;
        RECT 685.950 297.600 688.050 298.050 ;
        RECT 683.400 296.400 688.050 297.600 ;
        RECT 685.950 295.950 688.050 296.400 ;
        RECT 680.400 292.050 681.600 294.000 ;
        RECT 686.400 292.050 687.600 295.950 ;
        RECT 689.400 295.050 690.600 310.950 ;
        RECT 707.400 307.050 708.600 313.950 ;
        RECT 706.950 304.950 709.050 307.050 ;
        RECT 691.950 301.950 694.050 304.050 ;
        RECT 688.950 292.950 691.050 295.050 ;
        RECT 679.950 289.950 682.050 292.050 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 683.400 288.900 684.600 289.950 ;
        RECT 682.950 286.800 685.050 288.900 ;
        RECT 688.950 286.950 691.050 289.050 ;
        RECT 673.950 283.950 676.050 286.050 ;
        RECT 679.950 283.950 682.050 286.050 ;
        RECT 676.950 280.950 679.050 283.050 ;
        RECT 670.950 277.950 673.050 280.050 ;
        RECT 670.950 271.950 673.050 274.050 ;
        RECT 671.400 259.050 672.600 271.950 ;
        RECT 677.400 262.200 678.600 280.950 ;
        RECT 676.950 260.100 679.050 262.200 ;
        RECT 680.400 262.050 681.600 283.950 ;
        RECT 682.950 280.950 685.050 283.050 ;
        RECT 677.400 259.050 678.600 260.100 ;
        RECT 679.950 259.950 682.050 262.050 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 674.400 255.000 675.600 256.950 ;
        RECT 661.950 250.950 664.050 253.050 ;
        RECT 664.950 250.950 667.050 253.050 ;
        RECT 655.950 238.950 658.050 241.050 ;
        RECT 652.950 235.950 655.050 238.050 ;
        RECT 643.950 232.950 646.050 235.050 ;
        RECT 662.400 226.050 663.600 250.950 ;
        RECT 670.950 249.600 673.050 253.050 ;
        RECT 673.950 250.950 676.050 255.000 ;
        RECT 676.950 249.600 679.050 250.050 ;
        RECT 670.950 249.000 679.050 249.600 ;
        RECT 671.400 248.400 679.050 249.000 ;
        RECT 676.950 247.950 679.050 248.400 ;
        RECT 683.400 241.050 684.600 280.950 ;
        RECT 689.400 265.050 690.600 286.950 ;
        RECT 692.400 280.050 693.600 301.950 ;
        RECT 710.400 298.050 711.600 364.950 ;
        RECT 712.950 361.950 715.050 366.000 ;
        RECT 721.950 364.950 724.050 367.050 ;
        RECT 722.400 352.050 723.600 364.950 ;
        RECT 721.950 349.950 724.050 352.050 ;
        RECT 721.950 346.800 724.050 348.900 ;
        RECT 715.950 338.100 718.050 340.200 ;
        RECT 716.400 337.050 717.600 338.100 ;
        RECT 722.400 337.050 723.600 346.800 ;
        RECT 725.400 340.200 726.600 367.950 ;
        RECT 730.950 340.950 733.050 343.050 ;
        RECT 724.950 338.100 727.050 340.200 ;
        RECT 727.950 337.950 730.050 340.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 719.400 325.050 720.600 334.950 ;
        RECT 728.400 328.050 729.600 337.950 ;
        RECT 727.950 325.950 730.050 328.050 ;
        RECT 718.950 322.950 721.050 325.050 ;
        RECT 724.950 319.950 727.050 322.050 ;
        RECT 712.950 307.950 715.050 310.050 ;
        RECT 694.950 295.950 697.050 298.050 ;
        RECT 709.950 295.950 712.050 298.050 ;
        RECT 695.400 283.050 696.600 295.950 ;
        RECT 697.950 292.950 700.050 295.050 ;
        RECT 703.950 293.100 706.050 295.200 ;
        RECT 694.950 280.950 697.050 283.050 ;
        RECT 691.950 277.950 694.050 280.050 ;
        RECT 694.950 271.950 697.050 274.050 ;
        RECT 688.950 262.950 691.050 265.050 ;
        RECT 695.400 259.050 696.600 271.950 ;
        RECT 698.400 265.050 699.600 292.950 ;
        RECT 704.400 292.050 705.600 293.100 ;
        RECT 703.950 289.950 706.050 292.050 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 703.950 265.950 706.050 268.050 ;
        RECT 697.950 262.950 700.050 265.050 ;
        RECT 688.950 256.950 691.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 689.400 255.900 690.600 256.950 ;
        RECT 688.800 253.800 690.900 255.900 ;
        RECT 691.950 253.950 694.050 256.050 ;
        RECT 688.950 250.650 691.050 252.750 ;
        RECT 682.950 238.950 685.050 241.050 ;
        RECT 646.950 223.950 649.050 226.050 ;
        RECT 661.950 223.950 664.050 226.050 ;
        RECT 628.950 220.950 631.050 223.050 ;
        RECT 640.950 220.950 643.050 223.050 ;
        RECT 625.950 190.950 628.050 193.050 ;
        RECT 583.950 187.950 586.050 190.050 ;
        RECT 592.950 187.950 595.050 190.050 ;
        RECT 601.950 189.600 604.050 190.050 ;
        RECT 601.950 188.400 606.600 189.600 ;
        RECT 601.950 187.950 604.050 188.400 ;
        RECT 565.950 181.950 568.050 184.050 ;
        RECT 571.950 182.100 574.050 184.200 ;
        RECT 577.950 182.100 580.050 184.200 ;
        RECT 572.400 181.050 573.600 182.100 ;
        RECT 578.400 181.050 579.600 182.100 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 571.950 178.950 574.050 181.050 ;
        RECT 574.950 178.950 577.050 181.050 ;
        RECT 577.950 178.950 580.050 181.050 ;
        RECT 569.400 178.050 570.600 178.950 ;
        RECT 565.950 176.400 570.600 178.050 ;
        RECT 575.400 177.000 576.600 178.950 ;
        RECT 565.950 175.950 570.000 176.400 ;
        RECT 568.950 172.950 571.050 175.050 ;
        RECT 574.950 172.950 577.050 177.000 ;
        RECT 584.400 175.050 585.600 187.950 ;
        RECT 593.400 181.050 594.600 187.950 ;
        RECT 598.950 182.100 601.050 184.200 ;
        RECT 599.400 181.050 600.600 182.100 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 595.950 178.950 598.050 181.050 ;
        RECT 598.950 178.950 601.050 181.050 ;
        RECT 590.400 177.900 591.600 178.950 ;
        RECT 596.400 177.900 597.600 178.950 ;
        RECT 605.400 177.900 606.600 188.400 ;
        RECT 616.950 187.950 619.050 190.050 ;
        RECT 607.950 181.950 610.050 184.050 ;
        RECT 583.950 172.950 586.050 175.050 ;
        RECT 589.950 172.950 592.050 177.900 ;
        RECT 595.950 175.800 598.050 177.900 ;
        RECT 604.950 175.800 607.050 177.900 ;
        RECT 563.400 158.400 567.600 159.600 ;
        RECT 562.950 154.950 565.050 157.050 ;
        RECT 550.950 148.950 553.050 151.050 ;
        RECT 547.950 141.600 550.050 142.050 ;
        RECT 545.400 140.400 550.050 141.600 ;
        RECT 545.400 136.050 546.600 140.400 ;
        RECT 547.950 139.950 550.050 140.400 ;
        RECT 551.400 136.050 552.600 148.950 ;
        RECT 556.950 138.000 559.050 142.050 ;
        RECT 563.400 139.050 564.600 154.950 ;
        RECT 557.400 136.050 558.600 138.000 ;
        RECT 562.950 136.950 565.050 139.050 ;
        RECT 484.950 133.950 487.050 136.050 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 508.950 133.950 511.050 136.050 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 535.950 133.950 538.050 136.050 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 544.950 133.950 547.050 136.050 ;
        RECT 550.950 133.950 553.050 136.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 556.950 133.950 559.050 136.050 ;
        RECT 559.950 133.950 562.050 136.050 ;
        RECT 475.950 130.800 478.050 132.900 ;
        RECT 485.400 118.050 486.600 133.950 ;
        RECT 491.400 132.900 492.600 133.950 ;
        RECT 506.400 132.900 507.600 133.950 ;
        RECT 490.950 127.950 493.050 132.900 ;
        RECT 499.950 127.950 502.050 132.900 ;
        RECT 505.950 130.800 508.050 132.900 ;
        RECT 475.950 115.950 478.050 118.050 ;
        RECT 484.950 115.950 487.050 118.050 ;
        RECT 476.400 106.050 477.600 115.950 ;
        RECT 512.400 112.050 513.600 133.950 ;
        RECT 530.400 132.900 531.600 133.950 ;
        RECT 536.400 132.900 537.600 133.950 ;
        RECT 554.400 132.900 555.600 133.950 ;
        RECT 517.950 130.800 520.050 132.900 ;
        RECT 529.950 130.800 532.050 132.900 ;
        RECT 535.950 130.800 538.050 132.900 ;
        RECT 553.950 130.800 556.050 132.900 ;
        RECT 481.950 109.950 484.050 112.050 ;
        RECT 487.950 109.950 490.050 112.050 ;
        RECT 502.950 109.950 505.050 112.050 ;
        RECT 511.950 109.950 514.050 112.050 ;
        RECT 475.950 103.950 478.050 106.050 ;
        RECT 482.400 103.050 483.600 109.950 ;
        RECT 488.400 103.050 489.600 109.950 ;
        RECT 503.400 103.050 504.600 109.950 ;
        RECT 508.950 104.100 511.050 106.200 ;
        RECT 509.400 103.050 510.600 104.100 ;
        RECT 514.950 103.950 517.050 106.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 463.950 100.950 466.050 103.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 481.950 100.950 484.050 103.050 ;
        RECT 484.950 100.950 487.050 103.050 ;
        RECT 487.950 100.950 490.050 103.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 499.950 100.950 502.050 103.050 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 508.950 100.950 511.050 103.050 ;
        RECT 455.400 99.900 456.600 100.950 ;
        RECT 448.950 97.800 451.050 99.900 ;
        RECT 454.950 97.800 457.050 99.900 ;
        RECT 445.950 88.950 448.050 91.050 ;
        RECT 442.950 85.950 445.050 88.050 ;
        RECT 424.950 64.950 427.050 67.050 ;
        RECT 427.950 64.950 430.050 67.050 ;
        RECT 418.950 61.950 421.050 64.050 ;
        RECT 407.400 58.050 408.600 60.000 ;
        RECT 412.950 59.100 415.050 61.200 ;
        RECT 413.400 58.050 414.600 59.100 ;
        RECT 425.400 58.050 426.600 64.950 ;
        RECT 430.950 60.000 433.050 64.050 ;
        RECT 431.400 58.050 432.600 60.000 ;
        RECT 446.400 58.050 447.600 88.950 ;
        RECT 461.400 67.050 462.600 100.950 ;
        RECT 467.400 85.050 468.600 100.950 ;
        RECT 469.950 97.950 472.050 100.050 ;
        RECT 475.950 99.900 480.000 100.050 ;
        RECT 485.400 99.900 486.600 100.950 ;
        RECT 475.950 97.950 481.050 99.900 ;
        RECT 470.400 91.050 471.600 97.950 ;
        RECT 478.950 97.800 481.050 97.950 ;
        RECT 484.950 97.800 487.050 99.900 ;
        RECT 491.400 94.050 492.600 100.950 ;
        RECT 500.400 94.050 501.600 100.950 ;
        RECT 490.950 91.950 493.050 94.050 ;
        RECT 499.950 91.950 502.050 94.050 ;
        RECT 506.400 91.050 507.600 100.950 ;
        RECT 515.400 97.050 516.600 103.950 ;
        RECT 514.950 94.950 517.050 97.050 ;
        RECT 518.400 91.050 519.600 130.800 ;
        RECT 526.950 124.950 529.050 127.050 ;
        RECT 527.400 103.050 528.600 124.950 ;
        RECT 560.400 124.050 561.600 133.950 ;
        RECT 532.950 121.950 535.050 124.050 ;
        RECT 538.950 121.950 541.050 124.050 ;
        RECT 559.950 121.950 562.050 124.050 ;
        RECT 533.400 112.050 534.600 121.950 ;
        RECT 532.950 109.950 535.050 112.050 ;
        RECT 533.400 103.050 534.600 109.950 ;
        RECT 523.950 100.950 526.050 103.050 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 524.400 91.050 525.600 100.950 ;
        RECT 530.400 99.900 531.600 100.950 ;
        RECT 539.400 100.050 540.600 121.950 ;
        RECT 544.950 115.950 547.050 118.050 ;
        RECT 541.950 109.950 544.050 112.050 ;
        RECT 542.400 106.050 543.600 109.950 ;
        RECT 541.950 103.950 544.050 106.050 ;
        RECT 545.400 103.050 546.600 115.950 ;
        RECT 550.950 105.000 553.050 109.050 ;
        RECT 559.950 106.950 562.050 109.050 ;
        RECT 551.400 103.050 552.600 105.000 ;
        RECT 544.950 100.950 547.050 103.050 ;
        RECT 547.950 100.950 550.050 103.050 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 529.950 97.800 532.050 99.900 ;
        RECT 538.950 97.950 541.050 100.050 ;
        RECT 548.400 99.900 549.600 100.950 ;
        RECT 554.400 99.900 555.600 100.950 ;
        RECT 547.950 97.800 550.050 99.900 ;
        RECT 553.950 97.800 556.050 99.900 ;
        RECT 556.950 97.950 559.050 100.050 ;
        RECT 560.400 99.900 561.600 106.950 ;
        RECT 562.950 103.950 565.050 106.050 ;
        RECT 563.400 100.050 564.600 103.950 ;
        RECT 566.400 103.050 567.600 158.400 ;
        RECT 569.400 118.050 570.600 172.950 ;
        RECT 592.950 169.950 595.050 175.050 ;
        RECT 592.950 160.950 595.050 163.050 ;
        RECT 574.950 145.950 577.050 148.050 ;
        RECT 575.400 136.050 576.600 145.950 ;
        RECT 580.950 137.100 583.050 139.200 ;
        RECT 581.400 136.050 582.600 137.100 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 577.950 133.950 580.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 578.400 132.900 579.600 133.950 ;
        RECT 584.400 132.900 585.600 133.950 ;
        RECT 593.400 133.050 594.600 160.950 ;
        RECT 604.950 142.950 607.050 145.050 ;
        RECT 598.950 137.100 601.050 139.200 ;
        RECT 605.400 139.050 606.600 142.950 ;
        RECT 608.400 139.200 609.600 181.950 ;
        RECT 617.400 181.050 618.600 187.950 ;
        RECT 622.950 182.100 625.050 184.200 ;
        RECT 623.400 181.050 624.600 182.100 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 616.950 178.950 619.050 181.050 ;
        RECT 619.950 178.950 622.050 181.050 ;
        RECT 622.950 178.950 625.050 181.050 ;
        RECT 614.400 172.050 615.600 178.950 ;
        RECT 620.400 177.000 621.600 178.950 ;
        RECT 619.950 172.950 622.050 177.000 ;
        RECT 629.400 172.050 630.600 220.950 ;
        RECT 637.950 215.100 640.050 220.050 ;
        RECT 647.400 216.600 648.600 223.950 ;
        RECT 644.400 215.400 648.600 216.600 ;
        RECT 655.950 216.000 658.050 220.050 ;
        RECT 638.400 214.050 639.600 215.100 ;
        RECT 644.400 214.050 645.600 215.400 ;
        RECT 656.400 214.050 657.600 216.000 ;
        RECT 662.400 214.050 663.600 223.950 ;
        RECT 679.950 215.100 682.050 217.200 ;
        RECT 689.400 217.050 690.600 250.650 ;
        RECT 680.400 214.050 681.600 215.100 ;
        RECT 688.950 214.950 691.050 217.050 ;
        RECT 634.950 211.950 637.050 214.050 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 640.950 211.950 643.050 214.050 ;
        RECT 643.950 211.950 646.050 214.050 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 658.950 211.950 661.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 676.950 211.950 679.050 214.050 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 635.400 187.050 636.600 211.950 ;
        RECT 641.400 205.050 642.600 211.950 ;
        RECT 659.400 205.050 660.600 211.950 ;
        RECT 665.400 210.900 666.600 211.950 ;
        RECT 664.950 208.800 667.050 210.900 ;
        RECT 670.950 210.600 673.050 211.050 ;
        RECT 677.400 210.600 678.600 211.950 ;
        RECT 683.400 210.900 684.600 211.950 ;
        RECT 670.950 209.400 678.600 210.600 ;
        RECT 670.950 208.950 673.050 209.400 ;
        RECT 682.950 208.800 685.050 210.900 ;
        RECT 688.950 208.950 691.050 211.050 ;
        RECT 673.950 205.950 676.050 208.050 ;
        RECT 640.950 202.950 643.050 205.050 ;
        RECT 658.950 202.950 661.050 205.050 ;
        RECT 649.950 190.950 652.050 193.050 ;
        RECT 634.950 184.950 637.050 187.050 ;
        RECT 631.950 181.950 634.050 184.050 ;
        RECT 640.950 182.100 643.050 184.200 ;
        RECT 613.950 169.950 616.050 172.050 ;
        RECT 628.950 169.950 631.050 172.050 ;
        RECT 632.400 148.050 633.600 181.950 ;
        RECT 641.400 181.050 642.600 182.100 ;
        RECT 637.950 178.950 640.050 181.050 ;
        RECT 640.950 178.950 643.050 181.050 ;
        RECT 643.950 178.950 646.050 181.050 ;
        RECT 631.950 145.950 634.050 148.050 ;
        RECT 632.400 142.050 633.600 145.950 ;
        RECT 638.400 145.050 639.600 178.950 ;
        RECT 644.400 163.050 645.600 178.950 ;
        RECT 650.400 169.050 651.600 190.950 ;
        RECT 663.000 186.600 667.050 187.050 ;
        RECT 662.400 184.950 667.050 186.600 ;
        RECT 670.950 184.950 673.050 187.050 ;
        RECT 662.400 181.050 663.600 184.950 ;
        RECT 658.950 178.950 661.050 181.050 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 664.950 178.950 667.050 181.050 ;
        RECT 659.400 177.900 660.600 178.950 ;
        RECT 665.400 177.900 666.600 178.950 ;
        RECT 658.950 175.800 661.050 177.900 ;
        RECT 664.950 175.800 667.050 177.900 ;
        RECT 664.950 169.950 667.050 172.050 ;
        RECT 649.950 166.950 652.050 169.050 ;
        RECT 643.950 160.950 646.050 163.050 ;
        RECT 644.400 154.050 645.600 160.950 ;
        RECT 649.950 157.950 652.050 160.050 ;
        RECT 643.950 151.950 646.050 154.050 ;
        RECT 650.400 145.050 651.600 157.950 ;
        RECT 655.950 145.950 658.050 148.050 ;
        RECT 637.950 142.950 640.050 145.050 ;
        RECT 649.950 142.950 652.050 145.050 ;
        RECT 599.400 136.050 600.600 137.100 ;
        RECT 604.950 136.950 607.050 139.050 ;
        RECT 607.950 137.100 610.050 139.200 ;
        RECT 616.950 137.100 619.050 139.200 ;
        RECT 622.950 138.000 625.050 142.050 ;
        RECT 631.950 139.950 634.050 142.050 ;
        RECT 643.950 141.600 646.050 142.200 ;
        RECT 638.400 140.400 646.050 141.600 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 577.950 130.800 580.050 132.900 ;
        RECT 583.950 130.800 586.050 132.900 ;
        RECT 592.950 130.950 595.050 133.050 ;
        RECT 602.400 132.900 603.600 133.950 ;
        RECT 608.400 132.900 609.600 137.100 ;
        RECT 617.400 136.050 618.600 137.100 ;
        RECT 623.400 136.050 624.600 138.000 ;
        RECT 628.950 136.950 631.050 139.050 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 614.400 132.900 615.600 133.950 ;
        RECT 601.950 130.800 604.050 132.900 ;
        RECT 607.800 130.800 609.900 132.900 ;
        RECT 613.950 132.600 616.050 132.900 ;
        RECT 611.400 132.000 616.050 132.600 ;
        RECT 610.950 131.400 616.050 132.000 ;
        RECT 610.950 127.950 613.050 131.400 ;
        RECT 613.950 130.800 616.050 131.400 ;
        RECT 607.950 121.950 610.050 124.050 ;
        RECT 568.950 115.950 571.050 118.050 ;
        RECT 601.950 112.950 604.050 115.050 ;
        RECT 577.950 109.950 580.050 112.050 ;
        RECT 571.950 104.100 574.050 106.200 ;
        RECT 572.400 103.050 573.600 104.100 ;
        RECT 578.400 103.050 579.600 109.950 ;
        RECT 586.950 106.950 589.050 109.050 ;
        RECT 565.950 100.950 568.050 103.050 ;
        RECT 571.950 100.950 574.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 577.950 100.950 580.050 103.050 ;
        RECT 580.950 100.950 583.050 103.050 ;
        RECT 469.950 88.950 472.050 91.050 ;
        RECT 505.950 88.950 508.050 91.050 ;
        RECT 517.950 88.950 520.050 91.050 ;
        RECT 523.950 88.950 526.050 91.050 ;
        RECT 506.400 85.050 507.600 88.950 ;
        RECT 466.950 82.950 469.050 85.050 ;
        RECT 505.950 82.950 508.050 85.050 ;
        RECT 505.950 76.950 508.050 79.050 ;
        RECT 553.950 76.950 556.050 79.050 ;
        RECT 478.950 67.950 481.050 70.050 ;
        RECT 490.950 67.950 493.050 70.050 ;
        RECT 451.950 64.950 454.050 67.050 ;
        RECT 460.950 64.950 463.050 67.050 ;
        RECT 452.400 58.050 453.600 64.950 ;
        RECT 457.950 60.000 460.050 64.050 ;
        RECT 472.950 60.000 475.050 64.050 ;
        RECT 458.400 58.050 459.600 60.000 ;
        RECT 473.400 58.050 474.600 60.000 ;
        RECT 479.400 58.050 480.600 67.950 ;
        RECT 481.950 64.950 484.050 67.050 ;
        RECT 482.400 61.050 483.600 64.950 ;
        RECT 487.950 61.950 490.050 64.050 ;
        RECT 481.950 58.950 484.050 61.050 ;
        RECT 484.950 59.100 487.050 61.200 ;
        RECT 403.950 55.950 406.050 58.050 ;
        RECT 406.950 55.950 409.050 58.050 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 430.950 55.950 433.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 445.950 55.950 448.050 58.050 ;
        RECT 451.950 55.950 454.050 58.050 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 469.950 55.950 472.050 58.050 ;
        RECT 472.950 55.950 475.050 58.050 ;
        RECT 475.950 55.950 478.050 58.050 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 397.950 52.950 400.050 55.050 ;
        RECT 404.400 54.900 405.600 55.950 ;
        RECT 410.400 54.900 411.600 55.950 ;
        RECT 403.950 52.800 406.050 54.900 ;
        RECT 409.950 52.800 412.050 54.900 ;
        RECT 419.400 52.050 420.600 55.950 ;
        RECT 428.400 54.900 429.600 55.950 ;
        RECT 427.950 52.800 430.050 54.900 ;
        RECT 412.950 49.950 415.050 52.050 ;
        RECT 418.950 49.950 421.050 52.050 ;
        RECT 406.950 43.950 409.050 46.050 ;
        RECT 400.950 31.950 403.050 34.050 ;
        RECT 394.950 28.950 397.050 31.050 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 386.400 21.000 387.600 22.950 ;
        RECT 392.400 21.900 393.600 22.950 ;
        RECT 401.400 21.900 402.600 31.950 ;
        RECT 407.400 25.050 408.600 43.950 ;
        RECT 413.400 25.050 414.600 49.950 ;
        RECT 424.950 46.950 427.050 49.050 ;
        RECT 421.950 40.950 424.050 43.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 415.950 22.950 418.050 25.050 ;
        RECT 410.400 21.900 411.600 22.950 ;
        RECT 379.950 16.950 382.050 19.050 ;
        RECT 385.950 16.950 388.050 21.000 ;
        RECT 391.950 16.950 394.050 21.900 ;
        RECT 400.950 19.800 403.050 21.900 ;
        RECT 409.950 19.800 412.050 21.900 ;
        RECT 416.400 21.000 417.600 22.950 ;
        RECT 415.950 16.950 418.050 21.000 ;
        RECT 367.950 13.950 370.050 16.050 ;
        RECT 422.400 10.050 423.600 40.950 ;
        RECT 425.400 31.050 426.600 46.950 ;
        RECT 434.400 43.050 435.600 55.950 ;
        RECT 455.400 54.900 456.600 55.950 ;
        RECT 454.950 52.800 457.050 54.900 ;
        RECT 461.400 54.000 462.600 55.950 ;
        RECT 470.400 54.000 471.600 55.950 ;
        RECT 460.950 49.950 463.050 54.000 ;
        RECT 469.950 49.950 472.050 54.000 ;
        RECT 476.400 49.050 477.600 55.950 ;
        RECT 485.400 55.050 486.600 59.100 ;
        RECT 481.950 49.950 484.050 55.050 ;
        RECT 484.950 52.950 487.050 55.050 ;
        RECT 475.950 46.950 478.050 49.050 ;
        RECT 484.950 46.950 487.050 51.900 ;
        RECT 488.400 46.050 489.600 61.950 ;
        RECT 491.400 61.050 492.600 67.950 ;
        RECT 490.950 58.950 493.050 61.050 ;
        RECT 493.950 60.000 496.050 64.050 ;
        RECT 494.400 58.050 495.600 60.000 ;
        RECT 506.400 58.050 507.600 76.950 ;
        RECT 554.400 73.050 555.600 76.950 ;
        RECT 520.950 70.950 523.050 73.050 ;
        RECT 553.950 70.950 556.050 73.050 ;
        RECT 511.950 59.100 514.050 61.200 ;
        RECT 512.400 58.050 513.600 59.100 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 496.950 55.950 499.050 58.050 ;
        RECT 505.950 55.950 508.050 58.050 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 497.400 49.050 498.600 55.950 ;
        RECT 509.400 54.900 510.600 55.950 ;
        RECT 508.950 52.800 511.050 54.900 ;
        RECT 515.400 49.050 516.600 55.950 ;
        RECT 521.400 54.900 522.600 70.950 ;
        RECT 535.950 67.950 538.050 70.050 ;
        RECT 529.950 60.000 532.050 64.050 ;
        RECT 530.400 58.050 531.600 60.000 ;
        RECT 536.400 58.050 537.600 67.950 ;
        RECT 544.950 61.950 547.050 64.050 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 520.950 52.800 523.050 54.900 ;
        RECT 496.950 46.950 499.050 49.050 ;
        RECT 502.950 46.950 505.050 49.050 ;
        RECT 514.950 46.950 517.050 49.050 ;
        RECT 454.950 43.950 457.050 46.050 ;
        RECT 487.950 43.950 490.050 46.050 ;
        RECT 433.950 40.950 436.050 43.050 ;
        RECT 424.950 28.950 427.050 31.050 ;
        RECT 436.950 28.950 442.050 31.050 ;
        RECT 425.400 21.900 426.600 28.950 ;
        RECT 455.400 28.200 456.600 43.950 ;
        RECT 484.950 42.600 487.050 43.050 ;
        RECT 490.950 42.600 493.050 43.050 ;
        RECT 484.950 41.400 493.050 42.600 ;
        RECT 484.950 40.950 487.050 41.400 ;
        RECT 490.950 40.950 493.050 41.400 ;
        RECT 481.950 37.950 484.050 40.050 ;
        RECT 487.950 37.950 490.050 40.050 ;
        RECT 433.950 26.100 436.050 28.200 ;
        RECT 441.000 27.600 445.050 28.050 ;
        RECT 434.400 25.050 435.600 26.100 ;
        RECT 440.400 25.950 445.050 27.600 ;
        RECT 445.950 25.950 448.050 28.050 ;
        RECT 454.950 26.100 457.050 28.200 ;
        RECT 460.950 26.100 463.050 28.200 ;
        RECT 440.400 25.050 441.600 25.950 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 431.400 21.900 432.600 22.950 ;
        RECT 437.400 21.900 438.600 22.950 ;
        RECT 446.400 21.900 447.600 25.950 ;
        RECT 455.400 25.050 456.600 26.100 ;
        RECT 461.400 25.050 462.600 26.100 ;
        RECT 469.950 25.950 472.050 28.050 ;
        RECT 451.950 22.950 454.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 424.950 19.800 427.050 21.900 ;
        RECT 430.950 19.800 433.050 21.900 ;
        RECT 436.950 19.800 439.050 21.900 ;
        RECT 445.950 19.800 448.050 21.900 ;
        RECT 448.950 19.950 451.050 22.050 ;
        RECT 452.400 21.900 453.600 22.950 ;
        RECT 458.400 21.900 459.600 22.950 ;
        RECT 470.400 21.900 471.600 25.950 ;
        RECT 482.400 25.050 483.600 37.950 ;
        RECT 488.400 25.050 489.600 37.950 ;
        RECT 503.400 25.200 504.600 46.950 ;
        RECT 526.950 43.950 529.050 46.050 ;
        RECT 511.950 34.950 514.050 37.050 ;
        RECT 505.950 31.950 508.050 34.050 ;
        RECT 506.400 28.050 507.600 31.950 ;
        RECT 505.950 25.950 508.050 28.050 ;
        RECT 512.400 25.200 513.600 34.950 ;
        RECT 472.950 22.950 475.050 25.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 487.950 22.950 490.050 25.050 ;
        RECT 502.950 23.100 505.050 25.200 ;
        RECT 508.950 23.100 511.050 25.200 ;
        RECT 511.950 23.100 514.050 25.200 ;
        RECT 517.950 23.100 520.050 25.200 ;
        RECT 449.400 16.050 450.600 19.950 ;
        RECT 451.950 19.800 454.050 21.900 ;
        RECT 457.950 19.800 460.050 21.900 ;
        RECT 469.950 19.800 472.050 21.900 ;
        RECT 473.400 16.050 474.600 22.950 ;
        RECT 479.400 21.900 480.600 22.950 ;
        RECT 485.400 21.900 486.600 22.950 ;
        RECT 509.400 22.050 510.600 23.100 ;
        RECT 478.950 19.800 481.050 21.900 ;
        RECT 484.950 19.800 487.050 21.900 ;
        RECT 508.950 19.950 511.050 22.050 ;
        RECT 448.950 13.950 451.050 16.050 ;
        RECT 472.950 13.950 475.050 16.050 ;
        RECT 479.400 13.050 480.600 19.800 ;
        RECT 478.950 10.950 481.050 13.050 ;
        RECT 361.950 7.950 364.050 10.050 ;
        RECT 421.950 7.950 424.050 10.050 ;
        RECT 509.400 7.050 510.600 19.950 ;
        RECT 518.400 7.050 519.600 23.100 ;
        RECT 527.400 22.050 528.600 43.950 ;
        RECT 533.400 43.050 534.600 55.950 ;
        RECT 539.400 52.050 540.600 55.950 ;
        RECT 545.400 54.900 546.600 61.950 ;
        RECT 554.400 58.050 555.600 70.950 ;
        RECT 557.400 64.050 558.600 97.950 ;
        RECT 559.950 97.800 562.050 99.900 ;
        RECT 562.950 97.950 565.050 100.050 ;
        RECT 575.400 99.900 576.600 100.950 ;
        RECT 565.950 94.950 568.050 97.050 ;
        RECT 574.950 94.950 577.050 99.900 ;
        RECT 566.400 70.050 567.600 94.950 ;
        RECT 581.400 94.050 582.600 100.950 ;
        RECT 587.400 94.050 588.600 106.950 ;
        RECT 595.950 105.000 598.050 109.050 ;
        RECT 596.400 103.050 597.600 105.000 ;
        RECT 602.400 103.050 603.600 112.950 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 598.950 100.950 601.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 593.400 99.000 594.600 100.950 ;
        RECT 599.400 99.900 600.600 100.950 ;
        RECT 592.950 94.950 595.050 99.000 ;
        RECT 598.950 97.800 601.050 99.900 ;
        RECT 580.950 91.950 583.050 94.050 ;
        RECT 586.950 91.950 589.050 94.050 ;
        RECT 565.950 67.950 568.050 70.050 ;
        RECT 571.950 64.950 574.050 67.050 ;
        RECT 595.950 64.950 598.050 67.050 ;
        RECT 556.950 61.950 559.050 64.050 ;
        RECT 562.950 59.100 565.050 61.200 ;
        RECT 550.950 55.950 553.050 58.050 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 551.400 54.900 552.600 55.950 ;
        RECT 544.950 52.800 547.050 54.900 ;
        RECT 550.950 52.800 553.050 54.900 ;
        RECT 539.400 50.400 544.050 52.050 ;
        RECT 552.000 51.750 556.050 52.050 ;
        RECT 540.000 49.950 544.050 50.400 ;
        RECT 550.950 49.950 556.050 51.750 ;
        RECT 550.950 49.650 553.050 49.950 ;
        RECT 563.400 49.050 564.600 59.100 ;
        RECT 572.400 58.050 573.600 64.950 ;
        RECT 577.950 59.100 580.050 61.200 ;
        RECT 589.950 59.100 592.050 61.200 ;
        RECT 578.400 58.050 579.600 59.100 ;
        RECT 590.400 58.050 591.600 59.100 ;
        RECT 596.400 58.050 597.600 64.950 ;
        RECT 604.950 58.950 607.050 61.050 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 547.950 46.950 550.050 49.050 ;
        RECT 562.950 46.950 565.050 49.050 ;
        RECT 535.950 43.950 538.050 46.050 ;
        RECT 532.950 40.950 535.050 43.050 ;
        RECT 529.950 34.950 532.050 37.050 ;
        RECT 526.950 19.950 529.050 22.050 ;
        RECT 530.400 19.050 531.600 34.950 ;
        RECT 532.950 31.950 535.050 34.050 ;
        RECT 533.400 28.050 534.600 31.950 ;
        RECT 532.950 25.950 535.050 28.050 ;
        RECT 536.400 25.050 537.600 43.950 ;
        RECT 541.950 26.100 544.050 28.200 ;
        RECT 548.400 28.050 549.600 46.950 ;
        RECT 569.400 40.050 570.600 55.950 ;
        RECT 575.400 54.000 576.600 55.950 ;
        RECT 593.400 54.000 594.600 55.950 ;
        RECT 599.400 54.900 600.600 55.950 ;
        RECT 574.950 49.950 577.050 54.000 ;
        RECT 592.950 49.950 595.050 54.000 ;
        RECT 598.950 52.800 601.050 54.900 ;
        RECT 589.950 46.950 592.050 49.050 ;
        RECT 568.950 37.950 571.050 40.050 ;
        RECT 559.950 31.950 562.050 34.050 ;
        RECT 574.950 31.950 577.050 34.050 ;
        RECT 542.400 25.050 543.600 26.100 ;
        RECT 547.950 25.950 550.050 28.050 ;
        RECT 560.400 25.050 561.600 31.950 ;
        RECT 565.950 26.100 568.050 28.200 ;
        RECT 566.400 25.050 567.600 26.100 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 544.950 22.950 547.050 25.050 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 568.950 22.950 571.050 25.050 ;
        RECT 539.400 21.000 540.600 22.950 ;
        RECT 545.400 21.900 546.600 22.950 ;
        RECT 529.950 16.950 532.050 19.050 ;
        RECT 538.950 16.950 541.050 21.000 ;
        RECT 544.950 19.800 547.050 21.900 ;
        RECT 554.400 16.050 555.600 22.950 ;
        RECT 553.950 13.950 556.050 16.050 ;
        RECT 563.400 7.050 564.600 22.950 ;
        RECT 569.400 21.900 570.600 22.950 ;
        RECT 575.400 22.050 576.600 31.950 ;
        RECT 586.200 29.100 588.300 31.200 ;
        RECT 590.400 30.900 591.600 46.950 ;
        RECT 605.400 34.050 606.600 58.950 ;
        RECT 608.400 49.050 609.600 121.950 ;
        RECT 613.950 115.950 616.050 118.050 ;
        RECT 610.950 109.950 613.050 112.050 ;
        RECT 611.400 99.900 612.600 109.950 ;
        RECT 610.950 97.800 613.050 99.900 ;
        RECT 614.400 91.050 615.600 115.950 ;
        RECT 620.400 112.050 621.600 133.950 ;
        RECT 629.400 133.050 630.600 136.950 ;
        RECT 638.400 136.050 639.600 140.400 ;
        RECT 643.950 140.100 646.050 140.400 ;
        RECT 643.950 136.950 646.050 139.050 ;
        RECT 644.400 136.050 645.600 136.950 ;
        RECT 634.950 133.950 637.050 136.050 ;
        RECT 637.950 133.950 640.050 136.050 ;
        RECT 640.950 133.950 643.050 136.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 628.950 130.950 631.050 133.050 ;
        RECT 635.400 132.000 636.600 133.950 ;
        RECT 641.400 132.900 642.600 133.950 ;
        RECT 650.400 133.050 651.600 142.950 ;
        RECT 656.400 139.050 657.600 145.950 ;
        RECT 658.950 141.600 663.000 142.050 ;
        RECT 658.950 139.950 663.600 141.600 ;
        RECT 655.950 136.950 658.050 139.050 ;
        RECT 662.400 136.050 663.600 139.950 ;
        RECT 665.400 138.600 666.600 169.950 ;
        RECT 671.400 169.050 672.600 184.950 ;
        RECT 674.400 184.050 675.600 205.950 ;
        RECT 673.950 181.950 676.050 184.050 ;
        RECT 676.950 183.000 679.050 187.050 ;
        RECT 677.400 181.050 678.600 183.000 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 680.400 177.900 681.600 178.950 ;
        RECT 679.950 175.800 682.050 177.900 ;
        RECT 667.800 166.950 669.900 169.050 ;
        RECT 670.950 166.950 673.050 169.050 ;
        RECT 668.400 159.600 669.600 166.950 ;
        RECT 668.400 158.400 672.600 159.600 ;
        RECT 665.400 137.400 669.600 138.600 ;
        RECT 658.950 133.950 661.050 136.050 ;
        RECT 661.950 133.950 664.050 136.050 ;
        RECT 634.950 127.950 637.050 132.000 ;
        RECT 640.950 130.800 643.050 132.900 ;
        RECT 649.950 130.950 652.050 133.050 ;
        RECT 659.400 132.900 660.600 133.950 ;
        RECT 658.950 130.800 661.050 132.900 ;
        RECT 668.400 121.050 669.600 137.400 ;
        RECT 667.950 118.950 670.050 121.050 ;
        RECT 646.950 115.950 649.050 118.050 ;
        RECT 637.950 112.950 640.050 115.050 ;
        RECT 619.950 109.950 622.050 112.050 ;
        RECT 638.400 109.050 639.600 112.950 ;
        RECT 637.950 106.950 640.050 109.050 ;
        RECT 628.950 104.250 631.050 106.350 ;
        RECT 629.400 103.200 630.600 104.250 ;
        RECT 638.400 103.200 639.600 106.950 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 622.950 101.100 625.050 103.200 ;
        RECT 628.950 101.100 631.050 103.200 ;
        RECT 631.950 101.100 634.050 103.200 ;
        RECT 637.950 101.100 640.050 103.200 ;
        RECT 613.950 88.950 616.050 91.050 ;
        RECT 617.400 79.050 618.600 100.950 ;
        RECT 623.400 88.050 624.600 101.100 ;
        RECT 632.400 100.050 633.600 101.100 ;
        RECT 632.400 98.400 637.050 100.050 ;
        RECT 647.400 99.900 648.600 115.950 ;
        RECT 671.400 112.050 672.600 158.400 ;
        RECT 673.950 151.950 676.050 154.050 ;
        RECT 674.400 139.050 675.600 151.950 ;
        RECT 680.400 141.600 681.600 175.800 ;
        RECT 682.950 157.950 685.050 160.050 ;
        RECT 677.400 140.400 681.600 141.600 ;
        RECT 673.950 136.950 676.050 139.050 ;
        RECT 677.400 136.050 678.600 140.400 ;
        RECT 683.400 136.050 684.600 157.950 ;
        RECT 689.400 157.050 690.600 208.950 ;
        RECT 692.400 205.050 693.600 253.950 ;
        RECT 698.400 250.050 699.600 256.950 ;
        RECT 700.950 253.950 703.050 256.050 ;
        RECT 697.950 247.950 700.050 250.050 ;
        RECT 697.950 235.950 700.050 238.050 ;
        RECT 694.950 220.950 697.050 223.050 ;
        RECT 695.400 210.900 696.600 220.950 ;
        RECT 698.400 217.050 699.600 235.950 ;
        RECT 701.400 219.600 702.600 253.950 ;
        RECT 704.400 223.050 705.600 265.950 ;
        RECT 707.400 265.050 708.600 289.950 ;
        RECT 709.950 286.950 712.050 289.050 ;
        RECT 706.950 262.950 709.050 265.050 ;
        RECT 710.400 259.050 711.600 286.950 ;
        RECT 713.400 265.050 714.600 307.950 ;
        RECT 718.950 293.100 721.050 295.200 ;
        RECT 719.400 292.050 720.600 293.100 ;
        RECT 725.400 292.050 726.600 319.950 ;
        RECT 731.400 304.050 732.600 340.950 ;
        RECT 734.400 340.050 735.600 367.950 ;
        RECT 743.400 361.050 744.600 371.400 ;
        RECT 742.950 358.950 745.050 361.050 ;
        RECT 736.950 355.950 739.050 358.050 ;
        RECT 733.950 337.950 736.050 340.050 ;
        RECT 737.400 337.050 738.600 355.950 ;
        RECT 746.400 355.050 747.600 374.400 ;
        RECT 749.400 373.050 750.600 382.950 ;
        RECT 752.400 375.600 753.600 386.400 ;
        RECT 758.400 376.050 759.600 409.950 ;
        RECT 761.400 391.050 762.600 412.800 ;
        RECT 764.400 412.050 765.600 470.400 ;
        RECT 766.950 463.950 769.050 466.050 ;
        RECT 767.400 454.050 768.600 463.950 ;
        RECT 791.400 454.050 792.600 481.950 ;
        RECT 799.950 472.950 802.050 475.050 ;
        RECT 806.400 474.600 807.600 481.950 ;
        RECT 814.950 475.950 817.050 478.050 ;
        RECT 806.400 473.400 810.600 474.600 ;
        RECT 766.950 451.950 769.050 454.050 ;
        RECT 778.950 451.950 781.050 454.050 ;
        RECT 790.950 451.950 793.050 454.050 ;
        RECT 769.950 439.950 775.050 442.050 ;
        RECT 766.950 436.950 769.050 439.050 ;
        RECT 767.400 418.050 768.600 436.950 ;
        RECT 772.950 433.950 775.050 436.050 ;
        RECT 769.950 427.950 772.050 430.050 ;
        RECT 766.950 415.950 769.050 418.050 ;
        RECT 770.400 415.050 771.600 427.950 ;
        RECT 773.400 421.050 774.600 433.950 ;
        RECT 779.400 433.050 780.600 451.950 ;
        RECT 791.400 448.050 792.600 451.950 ;
        RECT 800.400 451.050 801.600 472.950 ;
        RECT 802.950 469.950 805.050 472.050 ;
        RECT 803.400 453.600 804.600 469.950 ;
        RECT 809.400 457.050 810.600 473.400 ;
        RECT 808.950 454.950 811.050 457.050 ;
        RECT 803.400 453.000 807.600 453.600 ;
        RECT 803.400 452.400 808.050 453.000 ;
        RECT 799.950 448.950 802.050 451.050 ;
        RECT 805.950 448.950 808.050 452.400 ;
        RECT 809.400 448.050 810.600 454.950 ;
        RECT 784.950 445.950 787.050 448.050 ;
        RECT 790.950 445.950 793.050 448.050 ;
        RECT 802.950 445.950 805.050 448.050 ;
        RECT 808.950 445.950 811.050 448.050 ;
        RECT 785.400 444.900 786.600 445.950 ;
        RECT 784.950 442.800 787.050 444.900 ;
        RECT 799.950 442.950 802.050 445.050 ;
        RECT 803.400 444.900 804.600 445.950 ;
        RECT 781.950 439.950 784.050 442.050 ;
        RECT 778.950 430.950 781.050 433.050 ;
        RECT 775.950 421.800 778.050 423.900 ;
        RECT 772.950 418.950 775.050 421.050 ;
        RECT 776.400 415.050 777.600 421.800 ;
        RECT 782.400 418.050 783.600 439.950 ;
        RECT 784.950 430.950 787.050 433.050 ;
        RECT 781.950 415.950 784.050 418.050 ;
        RECT 769.950 412.950 772.050 415.050 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 775.950 412.950 778.050 415.050 ;
        RECT 778.950 412.950 781.050 415.050 ;
        RECT 763.950 409.950 766.050 412.050 ;
        RECT 773.400 411.900 774.600 412.950 ;
        RECT 772.950 409.800 775.050 411.900 ;
        RECT 763.950 406.800 766.050 408.900 ;
        RECT 766.950 406.950 769.050 409.050 ;
        RECT 760.950 388.950 763.050 391.050 ;
        RECT 752.400 374.400 756.600 375.600 ;
        RECT 748.950 370.950 751.050 373.050 ;
        RECT 755.400 370.050 756.600 374.400 ;
        RECT 757.950 373.950 760.050 376.050 ;
        RECT 760.950 371.100 763.050 373.200 ;
        RECT 764.400 373.050 765.600 406.800 ;
        RECT 761.400 370.050 762.600 371.100 ;
        RECT 763.950 370.950 766.050 373.050 ;
        RECT 751.950 367.950 754.050 370.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 748.950 364.950 751.050 367.050 ;
        RECT 745.950 352.950 748.050 355.050 ;
        RECT 749.400 352.050 750.600 364.950 ;
        RECT 748.950 349.950 751.050 352.050 ;
        RECT 745.950 340.950 748.050 343.050 ;
        RECT 736.950 334.950 739.050 337.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 740.400 316.050 741.600 334.950 ;
        RECT 739.950 313.950 742.050 316.050 ;
        RECT 730.950 301.950 733.050 304.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 722.400 288.900 723.600 289.950 ;
        RECT 721.950 286.800 724.050 288.900 ;
        RECT 724.950 283.950 727.050 286.050 ;
        RECT 715.950 274.950 718.050 277.050 ;
        RECT 712.950 262.950 715.050 265.050 ;
        RECT 716.400 259.050 717.600 274.950 ;
        RECT 725.400 262.050 726.600 283.950 ;
        RECT 731.400 274.050 732.600 301.950 ;
        RECT 746.400 298.050 747.600 340.950 ;
        RECT 749.400 339.600 750.600 349.950 ;
        RECT 752.400 343.050 753.600 367.950 ;
        RECT 758.400 366.900 759.600 367.950 ;
        RECT 757.950 364.800 760.050 366.900 ;
        RECT 763.950 364.950 766.050 367.050 ;
        RECT 760.950 358.950 763.050 361.050 ;
        RECT 757.950 349.950 760.050 352.050 ;
        RECT 751.950 340.950 754.050 343.050 ;
        RECT 758.400 340.050 759.600 349.950 ;
        RECT 761.400 349.050 762.600 358.950 ;
        RECT 764.400 349.050 765.600 364.950 ;
        RECT 767.400 358.050 768.600 406.950 ;
        RECT 779.400 406.050 780.600 412.950 ;
        RECT 778.950 403.950 781.050 406.050 ;
        RECT 785.400 394.050 786.600 430.950 ;
        RECT 787.950 421.950 790.050 424.050 ;
        RECT 788.400 418.050 789.600 421.950 ;
        RECT 787.950 415.950 790.050 418.050 ;
        RECT 793.950 416.100 796.050 418.200 ;
        RECT 800.400 418.050 801.600 442.950 ;
        RECT 802.950 442.800 805.050 444.900 ;
        RECT 811.950 442.950 814.050 445.050 ;
        RECT 812.400 436.050 813.600 442.950 ;
        RECT 811.950 433.950 814.050 436.050 ;
        RECT 802.950 430.950 805.050 433.050 ;
        RECT 803.400 421.050 804.600 430.950 ;
        RECT 802.950 418.950 805.050 421.050 ;
        RECT 812.400 418.050 813.600 433.950 ;
        RECT 815.400 424.050 816.600 475.950 ;
        RECT 826.950 457.950 829.050 460.050 ;
        RECT 817.950 454.950 820.050 457.050 ;
        RECT 814.950 421.950 817.050 424.050 ;
        RECT 818.400 421.050 819.600 454.950 ;
        RECT 820.950 448.950 823.050 451.050 ;
        RECT 821.400 427.050 822.600 448.950 ;
        RECT 827.400 448.050 828.600 457.950 ;
        RECT 830.400 451.050 831.600 487.950 ;
        RECT 833.400 478.050 834.600 508.950 ;
        RECT 835.950 502.950 838.050 505.050 ;
        RECT 836.400 496.050 837.600 502.950 ;
        RECT 839.400 498.600 840.600 517.950 ;
        RECT 842.400 502.050 843.600 523.950 ;
        RECT 844.950 520.950 847.050 523.050 ;
        RECT 845.400 505.050 846.600 520.950 ;
        RECT 857.400 514.050 858.600 523.950 ;
        RECT 863.400 522.900 864.600 523.950 ;
        RECT 862.950 520.800 865.050 522.900 ;
        RECT 868.950 520.800 871.050 522.900 ;
        RECT 856.950 511.950 859.050 514.050 ;
        RECT 865.950 511.950 868.050 514.050 ;
        RECT 856.950 505.950 859.050 508.050 ;
        RECT 862.950 505.950 865.050 508.050 ;
        RECT 844.950 502.950 847.050 505.050 ;
        RECT 857.400 502.050 858.600 505.950 ;
        RECT 841.950 499.950 844.050 502.050 ;
        RECT 856.950 499.950 859.050 502.050 ;
        RECT 863.400 499.050 864.600 505.950 ;
        RECT 839.400 497.400 843.600 498.600 ;
        RECT 835.950 493.950 838.050 496.050 ;
        RECT 842.400 493.050 843.600 497.400 ;
        RECT 862.950 496.950 865.050 499.050 ;
        RECT 866.400 493.050 867.600 511.950 ;
        RECT 869.400 496.050 870.600 520.800 ;
        RECT 868.950 493.950 871.050 496.050 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 844.950 490.950 847.050 493.050 ;
        RECT 862.950 490.950 865.050 493.050 ;
        RECT 865.950 490.950 868.050 493.050 ;
        RECT 835.950 487.950 838.050 490.050 ;
        RECT 832.950 475.950 835.050 478.050 ;
        RECT 836.400 472.050 837.600 487.950 ;
        RECT 839.400 481.050 840.600 490.950 ;
        RECT 845.400 484.050 846.600 490.950 ;
        RECT 844.950 481.950 847.050 484.050 ;
        RECT 838.950 478.950 841.050 481.050 ;
        RECT 847.950 475.950 850.050 478.050 ;
        RECT 835.950 469.950 838.050 472.050 ;
        RECT 832.950 463.950 835.050 466.050 ;
        RECT 833.400 460.050 834.600 463.950 ;
        RECT 832.950 457.950 835.050 460.050 ;
        RECT 848.400 451.050 849.600 475.950 ;
        RECT 863.400 475.050 864.600 490.950 ;
        RECT 868.950 487.950 871.050 490.050 ;
        RECT 869.400 478.050 870.600 487.950 ;
        RECT 872.400 487.050 873.600 526.950 ;
        RECT 875.400 514.050 876.600 577.950 ;
        RECT 880.950 576.600 885.000 577.050 ;
        RECT 880.950 574.950 885.600 576.600 ;
        RECT 884.400 574.200 885.600 574.950 ;
        RECT 883.950 572.100 886.050 574.200 ;
        RECT 890.400 574.050 891.600 577.950 ;
        RECT 899.400 574.050 900.600 607.950 ;
        RECT 902.400 607.050 903.600 635.400 ;
        RECT 904.950 634.950 907.050 635.400 ;
        RECT 904.950 616.950 907.050 619.050 ;
        RECT 901.950 604.950 904.050 607.050 ;
        RECT 905.400 604.050 906.600 616.950 ;
        RECT 911.400 610.200 912.600 655.950 ;
        RECT 914.400 613.050 915.600 667.800 ;
        RECT 917.400 664.050 918.600 676.950 ;
        RECT 916.950 661.950 919.050 664.050 ;
        RECT 913.950 610.950 916.050 613.050 ;
        RECT 910.950 608.100 913.050 610.200 ;
        RECT 910.950 604.950 913.050 607.050 ;
        RECT 917.400 606.600 918.600 661.950 ;
        RECT 920.400 610.050 921.600 682.800 ;
        RECT 919.950 607.950 922.050 610.050 ;
        RECT 917.400 605.400 921.600 606.600 ;
        RECT 911.400 604.050 912.600 604.950 ;
        RECT 904.950 601.950 907.050 604.050 ;
        RECT 907.950 601.950 910.050 604.050 ;
        RECT 910.950 601.950 913.050 604.050 ;
        RECT 913.950 601.950 916.050 604.050 ;
        RECT 901.950 598.950 904.050 601.050 ;
        RECT 908.400 600.900 909.600 601.950 ;
        RECT 902.400 583.050 903.600 598.950 ;
        RECT 907.950 598.800 910.050 600.900 ;
        RECT 904.950 595.950 907.050 598.050 ;
        RECT 901.950 580.950 904.050 583.050 ;
        RECT 905.400 577.050 906.600 595.950 ;
        RECT 914.400 589.050 915.600 601.950 ;
        RECT 920.400 595.050 921.600 605.400 ;
        RECT 919.950 594.600 922.050 595.050 ;
        RECT 917.400 593.400 922.050 594.600 ;
        RECT 907.950 586.950 910.050 589.050 ;
        RECT 913.950 586.950 916.050 589.050 ;
        RECT 904.950 576.600 907.050 577.050 ;
        RECT 902.400 575.400 907.050 576.600 ;
        RECT 884.400 571.050 885.600 572.100 ;
        RECT 889.950 571.950 892.050 574.050 ;
        RECT 892.950 571.950 895.050 574.050 ;
        RECT 898.950 571.950 901.050 574.050 ;
        RECT 880.950 568.950 883.050 571.050 ;
        RECT 883.950 568.950 886.050 571.050 ;
        RECT 886.950 568.950 889.050 571.050 ;
        RECT 877.950 565.950 880.050 568.050 ;
        RECT 881.400 567.000 882.600 568.950 ;
        RECT 878.400 562.050 879.600 565.950 ;
        RECT 880.950 562.950 883.050 567.000 ;
        RECT 887.400 562.050 888.600 568.950 ;
        RECT 889.950 565.950 892.050 568.050 ;
        RECT 877.950 559.950 880.050 562.050 ;
        RECT 886.950 559.950 889.050 562.050 ;
        RECT 880.950 547.950 883.050 550.050 ;
        RECT 877.950 541.950 880.050 544.050 ;
        RECT 874.950 511.950 877.050 514.050 ;
        RECT 878.400 508.050 879.600 541.950 ;
        RECT 881.400 529.050 882.600 547.950 ;
        RECT 890.400 541.050 891.600 565.950 ;
        RECT 889.950 538.950 892.050 541.050 ;
        RECT 883.950 532.950 886.050 535.050 ;
        RECT 880.950 526.950 883.050 529.050 ;
        RECT 884.400 526.050 885.600 532.950 ;
        RECT 890.400 526.050 891.600 538.950 ;
        RECT 893.400 529.050 894.600 571.950 ;
        RECT 902.400 571.050 903.600 575.400 ;
        RECT 904.950 574.950 907.050 575.400 ;
        RECT 908.400 574.050 909.600 586.950 ;
        RECT 910.950 580.950 913.050 583.050 ;
        RECT 907.950 571.950 910.050 574.050 ;
        RECT 901.950 568.950 904.050 571.050 ;
        RECT 904.950 568.950 907.050 571.050 ;
        RECT 901.950 550.950 904.050 553.050 ;
        RECT 902.400 529.050 903.600 550.950 ;
        RECT 905.400 547.050 906.600 568.950 ;
        RECT 907.950 565.950 910.050 568.050 ;
        RECT 904.950 544.950 907.050 547.050 ;
        RECT 908.400 534.600 909.600 565.950 ;
        RECT 911.400 535.050 912.600 580.950 ;
        RECT 913.950 574.950 916.050 577.050 ;
        RECT 914.400 550.050 915.600 574.950 ;
        RECT 917.400 553.050 918.600 593.400 ;
        RECT 919.950 592.950 922.050 593.400 ;
        RECT 919.950 586.950 922.050 589.050 ;
        RECT 916.950 550.950 919.050 553.050 ;
        RECT 913.950 547.950 916.050 550.050 ;
        RECT 916.950 544.950 919.050 547.050 ;
        RECT 913.950 538.950 916.050 541.050 ;
        RECT 905.400 534.000 909.600 534.600 ;
        RECT 904.950 533.400 909.600 534.000 ;
        RECT 904.950 529.950 907.050 533.400 ;
        RECT 910.950 532.950 913.050 535.050 ;
        RECT 911.400 531.600 912.600 532.950 ;
        RECT 908.400 530.400 912.600 531.600 ;
        RECT 892.950 526.950 895.050 529.050 ;
        RECT 898.950 526.950 901.050 529.050 ;
        RECT 901.950 526.950 904.050 529.050 ;
        RECT 883.950 523.950 886.050 526.050 ;
        RECT 886.950 523.950 889.050 526.050 ;
        RECT 889.950 523.950 892.050 526.050 ;
        RECT 880.950 520.950 883.050 523.050 ;
        RECT 877.950 505.950 880.050 508.050 ;
        RECT 881.400 502.050 882.600 520.950 ;
        RECT 887.400 517.050 888.600 523.950 ;
        RECT 892.950 520.950 895.050 523.050 ;
        RECT 889.950 517.950 892.050 520.050 ;
        RECT 886.950 514.950 889.050 517.050 ;
        RECT 874.950 499.950 877.050 502.050 ;
        RECT 880.950 499.950 883.050 502.050 ;
        RECT 871.950 484.950 874.050 487.050 ;
        RECT 868.950 475.950 871.050 478.050 ;
        RECT 862.950 472.950 865.050 475.050 ;
        RECT 862.950 463.950 865.050 466.050 ;
        RECT 829.950 448.950 832.050 451.050 ;
        RECT 841.950 448.950 844.050 451.050 ;
        RECT 847.950 448.950 850.050 451.050 ;
        RECT 853.950 449.100 856.050 451.200 ;
        RECT 826.950 445.950 829.050 448.050 ;
        RECT 832.950 445.950 835.050 448.050 ;
        RECT 833.400 444.900 834.600 445.950 ;
        RECT 832.950 442.800 835.050 444.900 ;
        RECT 838.950 439.950 841.050 445.050 ;
        RECT 842.400 433.050 843.600 448.950 ;
        RECT 854.400 448.050 855.600 449.100 ;
        RECT 850.950 445.950 853.050 448.050 ;
        RECT 853.950 445.950 856.050 448.050 ;
        RECT 829.950 430.950 832.050 433.050 ;
        RECT 841.950 430.950 844.050 433.050 ;
        RECT 830.400 427.050 831.600 430.950 ;
        RECT 842.400 427.050 843.600 430.950 ;
        RECT 851.400 427.050 852.600 445.950 ;
        RECT 863.400 436.050 864.600 463.950 ;
        RECT 868.950 457.950 871.050 460.050 ;
        RECT 869.400 448.050 870.600 457.950 ;
        RECT 875.400 451.050 876.600 499.950 ;
        RECT 890.400 499.050 891.600 517.950 ;
        RECT 893.400 499.050 894.600 520.950 ;
        RECT 883.950 495.000 886.050 499.050 ;
        RECT 889.800 496.950 891.900 499.050 ;
        RECT 892.950 496.950 895.050 499.050 ;
        RECT 891.000 495.900 894.000 496.050 ;
        RECT 891.000 495.600 895.050 495.900 ;
        RECT 884.400 493.050 885.600 495.000 ;
        RECT 890.400 493.950 895.050 495.600 ;
        RECT 890.400 493.050 891.600 493.950 ;
        RECT 892.950 493.800 895.050 493.950 ;
        RECT 880.950 490.950 883.050 493.050 ;
        RECT 883.950 490.950 886.050 493.050 ;
        RECT 886.950 490.950 889.050 493.050 ;
        RECT 889.950 490.950 892.050 493.050 ;
        RECT 881.400 489.000 882.600 490.950 ;
        RECT 880.950 484.950 883.050 489.000 ;
        RECT 883.950 481.950 886.050 484.050 ;
        RECT 880.950 475.950 883.050 478.050 ;
        RECT 877.950 466.950 880.050 469.050 ;
        RECT 874.950 448.950 877.050 451.050 ;
        RECT 868.950 445.950 871.050 448.050 ;
        RECT 871.950 445.950 874.050 448.050 ;
        RECT 872.400 439.050 873.600 445.950 ;
        RECT 874.950 442.950 877.050 445.050 ;
        RECT 871.950 436.950 874.050 439.050 ;
        RECT 862.950 433.950 865.050 436.050 ;
        RECT 820.950 424.950 823.050 427.050 ;
        RECT 829.950 424.950 832.050 427.050 ;
        RECT 832.950 421.950 835.050 427.050 ;
        RECT 841.950 424.950 844.050 427.050 ;
        RECT 850.950 424.950 853.050 427.050 ;
        RECT 856.950 424.950 859.050 427.050 ;
        RECT 847.950 421.950 850.050 424.050 ;
        RECT 794.400 415.050 795.600 416.100 ;
        RECT 799.950 415.950 802.050 418.050 ;
        RECT 802.950 415.800 805.050 417.900 ;
        RECT 811.950 415.950 814.050 418.050 ;
        RECT 814.950 417.000 817.050 420.900 ;
        RECT 817.950 418.950 820.050 421.050 ;
        RECT 790.950 412.950 793.050 415.050 ;
        RECT 793.950 412.950 796.050 415.050 ;
        RECT 796.950 412.950 799.050 415.050 ;
        RECT 787.950 409.950 790.050 412.050 ;
        RECT 769.950 391.950 772.050 394.050 ;
        RECT 784.950 391.950 787.050 394.050 ;
        RECT 770.400 373.050 771.600 391.950 ;
        RECT 788.400 390.600 789.600 409.950 ;
        RECT 791.400 408.600 792.600 412.950 ;
        RECT 797.400 411.900 798.600 412.950 ;
        RECT 796.950 409.800 799.050 411.900 ;
        RECT 799.950 409.950 802.050 412.050 ;
        RECT 796.950 408.600 799.050 408.750 ;
        RECT 791.400 407.400 799.050 408.600 ;
        RECT 796.950 406.650 799.050 407.400 ;
        RECT 785.400 389.400 789.600 390.600 ;
        RECT 781.950 382.950 784.050 385.050 ;
        RECT 775.950 376.950 778.050 379.050 ;
        RECT 769.950 370.950 772.050 373.050 ;
        RECT 776.400 370.050 777.600 376.950 ;
        RECT 772.950 367.950 775.050 370.050 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 769.950 364.950 772.050 367.050 ;
        RECT 773.400 366.900 774.600 367.950 ;
        RECT 766.950 355.950 769.050 358.050 ;
        RECT 760.950 346.950 763.050 349.050 ;
        RECT 763.950 346.950 766.050 349.050 ;
        RECT 766.950 346.950 769.050 352.050 ;
        RECT 760.950 340.950 763.050 343.050 ;
        RECT 749.400 338.400 753.600 339.600 ;
        RECT 752.400 337.050 753.600 338.400 ;
        RECT 757.950 337.950 760.050 340.050 ;
        RECT 751.950 334.950 754.050 337.050 ;
        RECT 754.950 334.950 757.050 337.050 ;
        RECT 755.400 333.900 756.600 334.950 ;
        RECT 754.950 331.800 757.050 333.900 ;
        RECT 761.400 333.600 762.600 340.950 ;
        RECT 764.400 337.050 765.600 346.950 ;
        RECT 770.400 339.600 771.600 364.950 ;
        RECT 772.950 364.800 775.050 366.900 ;
        RECT 782.400 357.600 783.600 382.950 ;
        RECT 779.400 356.400 783.600 357.600 ;
        RECT 772.950 346.950 775.050 349.050 ;
        RECT 767.400 338.400 771.600 339.600 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 758.400 332.400 762.600 333.600 ;
        RECT 754.950 325.950 757.050 328.050 ;
        RECT 733.950 295.950 736.050 298.050 ;
        RECT 745.950 295.950 748.050 298.050 ;
        RECT 751.950 295.950 754.050 298.050 ;
        RECT 730.950 271.950 733.050 274.050 ;
        RECT 734.400 273.600 735.600 295.950 ;
        RECT 739.950 293.100 742.050 295.200 ;
        RECT 740.400 292.050 741.600 293.100 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 742.950 286.950 745.050 289.050 ;
        RECT 739.950 283.950 742.050 286.050 ;
        RECT 734.400 272.400 738.600 273.600 ;
        RECT 730.950 266.400 733.050 268.500 ;
        RECT 724.950 259.950 727.050 262.050 ;
        RECT 727.950 261.000 730.050 265.050 ;
        RECT 728.400 259.050 729.600 261.000 ;
        RECT 709.950 256.950 712.050 259.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 727.950 256.950 730.050 259.050 ;
        RECT 713.400 229.050 714.600 256.950 ;
        RECT 719.400 255.900 720.600 256.950 ;
        RECT 718.950 253.800 721.050 255.900 ;
        RECT 724.950 253.950 727.050 256.050 ;
        RECT 725.400 235.050 726.600 253.950 ;
        RECT 731.850 251.400 733.050 266.400 ;
        RECT 730.950 249.300 733.050 251.400 ;
        RECT 731.850 245.700 733.050 249.300 ;
        RECT 730.950 243.600 733.050 245.700 ;
        RECT 724.950 232.950 727.050 235.050 ;
        RECT 712.950 226.950 715.050 229.050 ;
        RECT 733.950 223.950 736.050 226.050 ;
        RECT 703.950 220.950 706.050 223.050 ;
        RECT 701.400 218.400 705.600 219.600 ;
        RECT 697.950 214.950 700.050 217.050 ;
        RECT 704.400 214.050 705.600 218.400 ;
        RECT 709.950 216.000 712.050 220.050 ;
        RECT 718.950 217.950 721.050 220.050 ;
        RECT 710.400 214.050 711.600 216.000 ;
        RECT 715.950 214.950 718.050 217.050 ;
        RECT 700.950 211.950 703.050 214.050 ;
        RECT 703.950 211.950 706.050 214.050 ;
        RECT 706.950 211.950 709.050 214.050 ;
        RECT 709.950 211.950 712.050 214.050 ;
        RECT 701.400 210.900 702.600 211.950 ;
        RECT 694.950 208.800 697.050 210.900 ;
        RECT 700.950 208.800 703.050 210.900 ;
        RECT 691.950 202.950 694.050 205.050 ;
        RECT 701.400 202.050 702.600 208.800 ;
        RECT 700.950 199.950 703.050 202.050 ;
        RECT 707.400 196.050 708.600 211.950 ;
        RECT 706.950 193.950 709.050 196.050 ;
        RECT 709.950 188.400 712.050 190.500 ;
        RECT 700.950 182.100 703.050 184.200 ;
        RECT 706.950 182.400 709.050 184.500 ;
        RECT 701.400 181.050 702.600 182.100 ;
        RECT 707.400 181.050 708.600 182.400 ;
        RECT 700.950 178.950 703.050 181.050 ;
        RECT 706.950 178.950 709.050 181.050 ;
        RECT 710.850 173.400 712.050 188.400 ;
        RECT 716.400 184.500 717.600 214.950 ;
        RECT 719.400 211.050 720.600 217.950 ;
        RECT 727.950 215.100 730.050 217.200 ;
        RECT 728.400 214.050 729.600 215.100 ;
        RECT 734.400 214.050 735.600 223.950 ;
        RECT 737.400 220.050 738.600 272.400 ;
        RECT 740.400 255.600 741.600 283.950 ;
        RECT 743.400 262.050 744.600 286.950 ;
        RECT 746.400 274.050 747.600 289.950 ;
        RECT 752.400 274.050 753.600 295.950 ;
        RECT 745.950 271.950 748.050 274.050 ;
        RECT 751.950 271.950 754.050 274.050 ;
        RECT 755.400 273.600 756.600 325.950 ;
        RECT 758.400 286.050 759.600 332.400 ;
        RECT 767.400 316.050 768.600 338.400 ;
        RECT 773.400 337.050 774.600 346.950 ;
        RECT 779.400 337.050 780.600 356.400 ;
        RECT 785.400 354.600 786.600 389.400 ;
        RECT 800.400 385.050 801.600 409.950 ;
        RECT 803.400 406.050 804.600 415.800 ;
        RECT 815.400 415.050 816.600 417.000 ;
        RECT 820.950 416.100 823.050 418.200 ;
        RECT 826.950 417.000 829.050 421.050 ;
        RECT 832.950 418.800 835.050 420.900 ;
        RECT 821.400 415.050 822.600 416.100 ;
        RECT 827.400 415.050 828.600 417.000 ;
        RECT 805.950 412.950 808.050 415.050 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 817.950 412.950 820.050 415.050 ;
        RECT 820.950 412.950 823.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 806.400 409.050 807.600 412.950 ;
        RECT 811.950 409.950 814.050 412.050 ;
        RECT 805.950 406.950 808.050 409.050 ;
        RECT 802.950 403.950 805.050 406.050 ;
        RECT 799.950 382.950 802.050 385.050 ;
        RECT 805.950 382.950 808.050 385.050 ;
        RECT 787.950 379.950 790.050 382.050 ;
        RECT 788.400 364.050 789.600 379.950 ;
        RECT 793.950 371.100 796.050 373.200 ;
        RECT 799.950 371.100 802.050 373.200 ;
        RECT 806.400 373.050 807.600 382.950 ;
        RECT 812.400 373.050 813.600 409.950 ;
        RECT 818.400 397.050 819.600 412.950 ;
        RECT 824.400 411.900 825.600 412.950 ;
        RECT 823.950 406.950 826.050 411.900 ;
        RECT 829.950 409.950 832.050 412.050 ;
        RECT 833.400 411.900 834.600 418.800 ;
        RECT 841.950 417.000 844.050 421.050 ;
        RECT 842.400 415.050 843.600 417.000 ;
        RECT 838.950 412.950 841.050 415.050 ;
        RECT 841.950 412.950 844.050 415.050 ;
        RECT 817.950 394.950 820.050 397.050 ;
        RECT 830.400 393.600 831.600 409.950 ;
        RECT 832.950 409.800 835.050 411.900 ;
        RECT 839.400 411.000 840.600 412.950 ;
        RECT 838.950 406.950 841.050 411.000 ;
        RECT 848.400 400.050 849.600 421.950 ;
        RECT 857.400 415.050 858.600 424.950 ;
        RECT 875.400 424.050 876.600 442.950 ;
        RECT 878.400 439.050 879.600 466.950 ;
        RECT 881.400 457.050 882.600 475.950 ;
        RECT 884.400 469.050 885.600 481.950 ;
        RECT 887.400 481.050 888.600 490.950 ;
        RECT 892.950 487.950 895.050 490.050 ;
        RECT 889.950 484.950 892.050 487.050 ;
        RECT 886.950 478.950 889.050 481.050 ;
        RECT 883.950 466.950 886.050 469.050 ;
        RECT 883.950 463.800 886.050 465.900 ;
        RECT 880.950 454.950 883.050 457.050 ;
        RECT 884.400 448.050 885.600 463.800 ;
        RECT 890.400 462.600 891.600 484.950 ;
        RECT 887.400 461.400 891.600 462.600 ;
        RECT 887.400 454.050 888.600 461.400 ;
        RECT 889.950 457.950 892.050 460.050 ;
        RECT 886.950 451.950 889.050 454.050 ;
        RECT 890.400 448.050 891.600 457.950 ;
        RECT 893.400 451.050 894.600 487.950 ;
        RECT 899.400 484.050 900.600 526.950 ;
        RECT 908.400 526.050 909.600 530.400 ;
        RECT 914.400 526.050 915.600 538.950 ;
        RECT 917.400 529.050 918.600 544.950 ;
        RECT 916.950 526.950 919.050 529.050 ;
        RECT 904.950 523.950 907.050 526.050 ;
        RECT 907.950 523.950 910.050 526.050 ;
        RECT 910.950 523.950 913.050 526.050 ;
        RECT 913.950 523.950 916.050 526.050 ;
        RECT 901.950 505.950 904.050 508.050 ;
        RECT 902.400 496.050 903.600 505.950 ;
        RECT 905.400 499.050 906.600 523.950 ;
        RECT 911.400 522.900 912.600 523.950 ;
        RECT 910.950 520.800 913.050 522.900 ;
        RECT 907.950 499.950 910.050 502.050 ;
        RECT 916.950 499.950 919.050 502.050 ;
        RECT 904.950 496.950 907.050 499.050 ;
        RECT 901.950 493.950 904.050 496.050 ;
        RECT 908.400 493.050 909.600 499.950 ;
        RECT 904.950 490.950 907.050 493.050 ;
        RECT 907.950 490.950 910.050 493.050 ;
        RECT 910.950 490.950 913.050 493.050 ;
        RECT 901.950 487.950 904.050 490.050 ;
        RECT 905.400 489.000 906.600 490.950 ;
        RECT 898.950 481.950 901.050 484.050 ;
        RECT 898.950 472.950 901.050 475.050 ;
        RECT 892.950 448.950 895.050 451.050 ;
        RECT 883.950 445.950 886.050 448.050 ;
        RECT 886.950 445.950 889.050 448.050 ;
        RECT 889.950 445.950 892.050 448.050 ;
        RECT 883.950 439.950 886.050 442.050 ;
        RECT 877.950 436.950 880.050 439.050 ;
        RECT 880.950 436.950 883.050 439.050 ;
        RECT 881.400 430.050 882.600 436.950 ;
        RECT 880.950 427.950 883.050 430.050 ;
        RECT 868.950 421.950 871.050 424.050 ;
        RECT 874.950 421.950 877.050 424.050 ;
        RECT 862.950 417.000 865.050 421.050 ;
        RECT 869.400 418.050 870.600 421.950 ;
        RECT 884.400 421.200 885.600 439.950 ;
        RECT 887.400 430.050 888.600 445.950 ;
        RECT 892.950 442.950 895.050 445.050 ;
        RECT 889.950 436.950 892.050 439.050 ;
        RECT 886.950 427.950 889.050 430.050 ;
        RECT 871.950 418.950 874.050 421.050 ;
        RECT 883.950 419.100 886.050 421.200 ;
        RECT 863.400 415.050 864.600 417.000 ;
        RECT 868.950 415.950 871.050 418.050 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 865.950 412.950 868.050 415.050 ;
        RECT 854.400 411.000 855.600 412.950 ;
        RECT 853.950 406.950 856.050 411.000 ;
        RECT 838.950 397.950 841.050 400.050 ;
        RECT 847.950 397.950 850.050 400.050 ;
        RECT 827.400 392.400 831.600 393.600 ;
        RECT 814.950 379.950 817.050 382.050 ;
        RECT 794.400 370.050 795.600 371.100 ;
        RECT 800.400 370.050 801.600 371.100 ;
        RECT 805.950 370.950 808.050 373.050 ;
        RECT 811.950 370.950 814.050 373.050 ;
        RECT 815.400 370.050 816.600 379.950 ;
        RECT 823.950 372.000 826.050 376.050 ;
        RECT 827.400 373.050 828.600 392.400 ;
        RECT 829.950 382.950 832.050 385.050 ;
        RECT 824.400 370.050 825.600 372.000 ;
        RECT 826.950 370.950 829.050 373.050 ;
        RECT 793.950 367.950 796.050 370.050 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 799.950 367.950 802.050 370.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 814.950 367.950 817.050 370.050 ;
        RECT 817.950 367.950 820.050 370.050 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 790.950 364.950 793.050 367.050 ;
        RECT 797.400 366.000 798.600 367.950 ;
        RECT 803.400 366.900 804.600 367.950 ;
        RECT 818.400 366.900 819.600 367.950 ;
        RECT 830.400 367.050 831.600 382.950 ;
        RECT 832.950 373.950 835.050 376.050 ;
        RECT 787.950 361.950 790.050 364.050 ;
        RECT 787.950 355.950 790.050 358.050 ;
        RECT 782.400 353.400 786.600 354.600 ;
        RECT 782.400 343.050 783.600 353.400 ;
        RECT 788.400 352.050 789.600 355.950 ;
        RECT 787.950 351.600 790.050 352.050 ;
        RECT 785.400 350.400 790.050 351.600 ;
        RECT 781.950 340.950 784.050 343.050 ;
        RECT 772.950 334.950 775.050 337.050 ;
        RECT 775.950 334.950 778.050 337.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 769.950 328.950 772.050 334.050 ;
        RECT 766.950 313.950 769.050 316.050 ;
        RECT 760.950 307.950 763.050 310.050 ;
        RECT 761.400 295.050 762.600 307.950 ;
        RECT 776.400 301.050 777.600 334.950 ;
        RECT 775.950 298.950 778.050 301.050 ;
        RECT 760.950 292.950 763.050 295.050 ;
        RECT 763.950 294.000 766.050 298.050 ;
        RECT 764.400 292.050 765.600 294.000 ;
        RECT 778.950 293.100 781.050 295.200 ;
        RECT 779.400 292.050 780.600 293.100 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 775.950 289.950 778.050 292.050 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 767.400 288.900 768.600 289.950 ;
        RECT 766.950 286.800 769.050 288.900 ;
        RECT 757.950 283.950 760.050 286.050 ;
        RECT 763.950 283.950 766.050 286.050 ;
        RECT 776.400 285.600 777.600 289.950 ;
        RECT 776.400 284.400 780.600 285.600 ;
        RECT 760.950 274.950 763.050 277.050 ;
        RECT 755.400 272.400 759.600 273.600 ;
        RECT 746.400 268.050 747.600 271.950 ;
        RECT 745.950 265.950 748.050 268.050 ;
        RECT 751.950 266.400 754.050 268.500 ;
        RECT 742.950 259.950 745.050 262.050 ;
        RECT 745.950 256.950 748.050 259.050 ;
        RECT 740.400 254.400 744.600 255.600 ;
        RECT 739.950 250.950 742.050 253.050 ;
        RECT 736.950 217.950 739.050 220.050 ;
        RECT 740.400 217.050 741.600 250.950 ;
        RECT 743.400 229.050 744.600 254.400 ;
        RECT 746.400 247.050 747.600 256.950 ;
        RECT 745.950 244.950 748.050 247.050 ;
        RECT 752.100 246.600 753.300 266.400 ;
        RECT 758.400 262.050 759.600 272.400 ;
        RECT 757.950 259.950 760.050 262.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 755.400 255.000 756.600 256.950 ;
        RECT 754.950 250.950 757.050 255.000 ;
        RECT 757.950 253.950 760.050 256.050 ;
        RECT 751.950 244.500 754.050 246.600 ;
        RECT 742.950 226.950 745.050 229.050 ;
        RECT 754.950 226.950 757.050 229.050 ;
        RECT 742.950 223.800 745.050 225.900 ;
        RECT 739.950 214.950 742.050 217.050 ;
        RECT 727.950 211.950 730.050 214.050 ;
        RECT 730.950 211.950 733.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 736.950 211.950 739.050 214.050 ;
        RECT 718.950 208.950 721.050 211.050 ;
        RECT 731.400 210.900 732.600 211.950 ;
        RECT 730.950 208.800 733.050 210.900 ;
        RECT 737.400 205.050 738.600 211.950 ;
        RECT 739.950 208.950 742.050 211.050 ;
        RECT 736.950 202.950 739.050 205.050 ;
        RECT 718.950 199.950 721.050 202.050 ;
        RECT 715.950 182.400 718.050 184.500 ;
        RECT 709.950 171.300 712.050 173.400 ;
        RECT 719.400 172.050 720.600 199.950 ;
        RECT 721.950 193.950 724.050 196.050 ;
        RECT 722.400 184.050 723.600 193.950 ;
        RECT 730.950 188.400 733.050 190.500 ;
        RECT 721.950 181.950 724.050 184.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 725.400 178.050 726.600 178.950 ;
        RECT 721.950 176.400 726.600 178.050 ;
        RECT 721.950 175.950 726.000 176.400 ;
        RECT 700.800 166.950 702.900 169.050 ;
        RECT 710.850 167.700 712.050 171.300 ;
        RECT 718.950 169.950 721.050 172.050 ;
        RECT 731.100 168.600 732.300 188.400 ;
        RECT 733.950 178.950 736.050 181.050 ;
        RECT 734.400 177.600 735.600 178.950 ;
        RECT 740.400 177.600 741.600 208.950 ;
        RECT 743.400 208.050 744.600 223.800 ;
        RECT 745.950 217.950 748.050 220.050 ;
        RECT 742.950 205.950 745.050 208.050 ;
        RECT 742.950 199.950 745.050 202.050 ;
        RECT 733.950 176.400 741.600 177.600 ;
        RECT 733.950 175.500 736.050 176.400 ;
        RECT 688.950 154.950 691.050 157.050 ;
        RECT 691.950 148.950 694.050 151.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 679.950 133.950 682.050 136.050 ;
        RECT 682.950 133.950 685.050 136.050 ;
        RECT 685.950 133.950 688.050 136.050 ;
        RECT 680.400 132.900 681.600 133.950 ;
        RECT 686.400 132.900 687.600 133.950 ;
        RECT 679.950 130.800 682.050 132.900 ;
        RECT 685.950 130.800 688.050 132.900 ;
        RECT 686.400 118.050 687.600 130.800 ;
        RECT 692.400 124.050 693.600 148.950 ;
        RECT 701.400 145.050 702.600 166.950 ;
        RECT 709.950 165.600 712.050 167.700 ;
        RECT 730.950 166.500 733.050 168.600 ;
        RECT 712.950 160.950 715.050 163.050 ;
        RECT 700.950 142.950 703.050 145.050 ;
        RECT 706.950 142.950 709.050 145.050 ;
        RECT 694.950 137.100 697.050 139.200 ;
        RECT 700.950 137.100 703.050 139.200 ;
        RECT 695.400 133.050 696.600 137.100 ;
        RECT 701.400 136.050 702.600 137.100 ;
        RECT 707.400 136.050 708.600 142.950 ;
        RECT 700.950 133.950 703.050 136.050 ;
        RECT 703.950 133.950 706.050 136.050 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 694.950 130.950 697.050 133.050 ;
        RECT 704.400 132.900 705.600 133.950 ;
        RECT 713.400 133.050 714.600 160.950 ;
        RECT 724.950 148.950 727.050 151.050 ;
        RECT 715.950 145.950 718.050 148.050 ;
        RECT 703.950 130.800 706.050 132.900 ;
        RECT 712.950 130.950 715.050 133.050 ;
        RECT 716.400 127.050 717.600 145.950 ;
        RECT 725.400 136.050 726.600 148.950 ;
        RECT 730.950 137.100 733.050 139.200 ;
        RECT 731.400 136.050 732.600 137.100 ;
        RECT 721.950 133.950 724.050 136.050 ;
        RECT 724.950 133.950 727.050 136.050 ;
        RECT 727.950 133.950 730.050 136.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 722.400 127.050 723.600 133.950 ;
        RECT 694.950 124.950 697.050 127.050 ;
        RECT 715.950 124.950 718.050 127.050 ;
        RECT 721.950 124.950 724.050 127.050 ;
        RECT 691.950 121.950 694.050 124.050 ;
        RECT 685.950 115.950 688.050 118.050 ;
        RECT 670.950 109.950 673.050 112.050 ;
        RECT 685.950 109.950 688.050 112.050 ;
        RECT 649.950 105.600 652.050 109.050 ;
        RECT 649.950 105.000 654.600 105.600 ;
        RECT 650.400 104.400 654.600 105.000 ;
        RECT 653.400 103.050 654.600 104.400 ;
        RECT 658.950 104.100 661.050 106.200 ;
        RECT 659.400 103.050 660.600 104.100 ;
        RECT 667.950 103.950 670.050 106.050 ;
        RECT 673.950 104.100 676.050 106.200 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 633.000 97.950 637.050 98.400 ;
        RECT 646.950 97.800 649.050 99.900 ;
        RECT 622.950 85.950 625.050 88.050 ;
        RECT 616.950 76.950 619.050 79.050 ;
        RECT 623.400 67.050 624.600 85.950 ;
        RECT 656.400 79.050 657.600 100.950 ;
        RECT 662.400 99.900 663.600 100.950 ;
        RECT 661.950 97.800 664.050 99.900 ;
        RECT 668.400 94.050 669.600 103.950 ;
        RECT 674.400 103.050 675.600 104.100 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 670.950 97.950 673.050 100.050 ;
        RECT 677.400 99.000 678.600 100.950 ;
        RECT 667.950 91.950 670.050 94.050 ;
        RECT 671.400 88.050 672.600 97.950 ;
        RECT 676.950 94.950 679.050 99.000 ;
        RECT 670.950 85.950 673.050 88.050 ;
        RECT 686.400 82.050 687.600 109.950 ;
        RECT 695.400 103.050 696.600 124.950 ;
        RECT 709.950 118.950 712.050 121.050 ;
        RECT 703.950 106.950 706.050 109.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 692.400 94.050 693.600 100.950 ;
        RECT 698.400 99.000 699.600 100.950 ;
        RECT 697.950 94.950 700.050 99.000 ;
        RECT 691.950 91.950 694.050 94.050 ;
        RECT 688.950 88.950 691.050 91.050 ;
        RECT 689.400 85.050 690.600 88.950 ;
        RECT 688.950 82.950 691.050 85.050 ;
        RECT 685.950 79.950 688.050 82.050 ;
        RECT 655.950 76.950 658.050 79.050 ;
        RECT 673.950 73.950 676.050 76.050 ;
        RECT 646.950 70.950 649.050 73.050 ;
        RECT 622.950 64.950 625.050 67.050 ;
        RECT 616.950 59.100 619.050 61.200 ;
        RECT 631.950 59.100 634.050 61.200 ;
        RECT 617.400 58.050 618.600 59.100 ;
        RECT 632.400 58.050 633.600 59.100 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 628.950 55.950 631.050 58.050 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 607.950 46.950 610.050 49.050 ;
        RECT 614.400 40.050 615.600 55.950 ;
        RECT 629.400 54.900 630.600 55.950 ;
        RECT 635.400 54.900 636.600 55.950 ;
        RECT 647.400 55.050 648.600 70.950 ;
        RECT 652.950 67.950 655.050 70.050 ;
        RECT 653.400 58.050 654.600 67.950 ;
        RECT 658.950 60.000 661.050 64.050 ;
        RECT 659.400 58.050 660.600 60.000 ;
        RECT 664.950 59.100 667.050 61.200 ;
        RECT 665.400 58.050 666.600 59.100 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 628.950 52.800 631.050 54.900 ;
        RECT 634.950 52.800 637.050 54.900 ;
        RECT 646.950 52.950 649.050 55.050 ;
        RECT 656.400 49.050 657.600 55.950 ;
        RECT 662.400 54.000 663.600 55.950 ;
        RECT 674.400 54.600 675.600 73.950 ;
        RECT 691.950 69.300 694.050 71.400 ;
        RECT 692.850 65.700 694.050 69.300 ;
        RECT 691.950 63.600 694.050 65.700 ;
        RECT 679.950 59.100 682.050 61.200 ;
        RECT 680.400 58.050 681.600 59.100 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 683.400 54.900 684.600 55.950 ;
        RECT 661.950 49.950 664.050 54.000 ;
        RECT 674.400 53.400 678.600 54.600 ;
        RECT 655.950 46.950 658.050 49.050 ;
        RECT 613.950 37.950 616.050 40.050 ;
        RECT 652.950 37.950 655.050 40.050 ;
        RECT 604.950 31.950 607.050 34.050 ;
        RECT 584.400 25.200 585.600 27.600 ;
        RECT 583.950 23.100 586.050 25.200 ;
        RECT 586.950 24.000 587.850 29.100 ;
        RECT 589.500 28.800 591.600 30.900 ;
        RECT 596.250 29.400 598.350 31.500 ;
        RECT 593.700 27.000 595.800 27.900 ;
        RECT 588.750 25.800 595.800 27.000 ;
        RECT 588.750 24.900 590.850 25.800 ;
        RECT 593.700 24.000 595.800 24.900 ;
        RECT 586.950 23.100 595.800 24.000 ;
        RECT 568.950 19.800 571.050 21.900 ;
        RECT 574.950 19.950 577.050 22.050 ;
        RECT 586.950 16.500 587.850 23.100 ;
        RECT 593.700 22.800 595.800 23.100 ;
        RECT 589.500 20.100 591.600 22.200 ;
        RECT 590.400 17.550 591.600 20.100 ;
        RECT 596.700 16.800 597.600 29.400 ;
        RECT 598.500 23.100 600.600 25.200 ;
        RECT 599.400 20.550 600.600 23.100 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 586.800 14.400 588.900 16.500 ;
        RECT 595.800 14.700 597.900 16.800 ;
        RECT 602.400 10.050 603.600 22.950 ;
        RECT 605.400 21.900 606.600 31.950 ;
        RECT 613.950 26.100 616.050 28.200 ;
        RECT 614.400 25.050 615.600 26.100 ;
        RECT 619.950 25.950 622.050 31.050 ;
        RECT 622.950 26.100 625.050 28.200 ;
        RECT 631.950 26.100 634.050 28.200 ;
        RECT 637.950 26.100 640.050 28.200 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 611.400 21.900 612.600 22.950 ;
        RECT 604.950 19.800 607.050 21.900 ;
        RECT 610.950 19.800 613.050 21.900 ;
        RECT 611.400 13.050 612.600 19.800 ;
        RECT 617.400 16.050 618.600 22.950 ;
        RECT 623.400 16.050 624.600 26.100 ;
        RECT 632.400 25.050 633.600 26.100 ;
        RECT 638.400 25.050 639.600 26.100 ;
        RECT 646.950 25.950 649.050 28.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 637.950 22.950 640.050 25.050 ;
        RECT 629.400 21.900 630.600 22.950 ;
        RECT 635.400 21.900 636.600 22.950 ;
        RECT 628.950 19.800 631.050 21.900 ;
        RECT 634.950 19.800 637.050 21.900 ;
        RECT 647.400 19.050 648.600 25.950 ;
        RECT 653.400 25.050 654.600 37.950 ;
        RECT 658.950 26.100 661.050 28.200 ;
        RECT 664.950 26.100 667.050 28.200 ;
        RECT 667.950 27.600 672.000 28.050 ;
        RECT 659.400 25.050 660.600 26.100 ;
        RECT 652.950 22.950 655.050 25.050 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 658.950 22.950 661.050 25.050 ;
        RECT 656.400 21.900 657.600 22.950 ;
        RECT 655.950 19.800 658.050 21.900 ;
        RECT 616.950 13.950 619.050 16.050 ;
        RECT 622.950 13.950 625.050 16.050 ;
        RECT 631.950 13.950 634.050 19.050 ;
        RECT 646.950 16.950 649.050 19.050 ;
        RECT 661.950 16.950 664.050 22.050 ;
        RECT 665.400 16.050 666.600 26.100 ;
        RECT 667.950 25.950 672.600 27.600 ;
        RECT 671.400 25.050 672.600 25.950 ;
        RECT 677.400 25.050 678.600 53.400 ;
        RECT 682.950 52.800 685.050 54.900 ;
        RECT 689.400 54.600 690.600 55.950 ;
        RECT 683.400 28.200 684.600 52.800 ;
        RECT 688.950 52.500 691.050 54.600 ;
        RECT 692.850 48.600 694.050 63.600 ;
        RECT 704.400 60.600 705.600 106.950 ;
        RECT 710.400 88.050 711.600 118.950 ;
        RECT 721.950 115.950 724.050 118.050 ;
        RECT 715.950 105.000 718.050 109.050 ;
        RECT 716.400 103.050 717.600 105.000 ;
        RECT 722.400 103.050 723.600 115.950 ;
        RECT 728.400 106.050 729.600 133.950 ;
        RECT 737.400 109.050 738.600 176.400 ;
        RECT 743.400 175.050 744.600 199.950 ;
        RECT 742.950 172.950 745.050 175.050 ;
        RECT 743.400 160.050 744.600 172.950 ;
        RECT 742.950 157.950 745.050 160.050 ;
        RECT 742.950 148.050 745.050 151.050 ;
        RECT 739.950 147.000 745.050 148.050 ;
        RECT 739.950 146.400 744.600 147.000 ;
        RECT 739.950 145.950 744.000 146.400 ;
        RECT 742.950 142.950 745.050 145.050 ;
        RECT 743.400 136.050 744.600 142.950 ;
        RECT 746.400 142.050 747.600 217.950 ;
        RECT 755.400 214.050 756.600 226.950 ;
        RECT 758.400 220.050 759.600 253.950 ;
        RECT 761.400 247.050 762.600 274.950 ;
        RECT 760.950 244.950 763.050 247.050 ;
        RECT 757.950 217.950 760.050 220.050 ;
        RECT 751.950 211.950 754.050 214.050 ;
        RECT 754.950 211.950 757.050 214.050 ;
        RECT 757.950 211.950 760.050 214.050 ;
        RECT 752.400 210.000 753.600 211.950 ;
        RECT 751.950 205.950 754.050 210.000 ;
        RECT 758.400 205.050 759.600 211.950 ;
        RECT 760.950 208.950 763.050 211.050 ;
        RECT 757.950 202.950 760.050 205.050 ;
        RECT 757.950 181.950 760.050 184.050 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 752.400 177.900 753.600 178.950 ;
        RECT 751.950 175.800 754.050 177.900 ;
        RECT 748.950 157.950 751.050 160.050 ;
        RECT 745.950 139.950 748.050 142.050 ;
        RECT 749.400 139.200 750.600 157.950 ;
        RECT 758.400 145.050 759.600 181.950 ;
        RECT 757.950 142.950 760.050 145.050 ;
        RECT 761.400 142.050 762.600 208.950 ;
        RECT 764.400 151.050 765.600 283.950 ;
        RECT 775.950 277.950 778.050 280.050 ;
        RECT 766.950 268.950 769.050 271.050 ;
        RECT 767.400 223.050 768.600 268.950 ;
        RECT 776.400 259.050 777.600 277.950 ;
        RECT 779.400 277.050 780.600 284.400 ;
        RECT 778.950 274.950 781.050 277.050 ;
        RECT 785.400 268.050 786.600 350.400 ;
        RECT 787.950 349.950 790.050 350.400 ;
        RECT 791.400 349.050 792.600 364.950 ;
        RECT 796.950 364.050 799.050 366.000 ;
        RECT 802.950 364.800 805.050 366.900 ;
        RECT 817.800 364.800 819.900 366.900 ;
        RECT 820.950 364.950 823.050 367.050 ;
        RECT 829.950 364.950 832.050 367.050 ;
        RECT 796.800 363.000 799.050 364.050 ;
        RECT 796.800 361.950 798.900 363.000 ;
        RECT 799.950 361.950 802.050 364.050 ;
        RECT 793.950 352.950 796.050 355.050 ;
        RECT 790.950 346.950 793.050 349.050 ;
        RECT 794.400 337.050 795.600 352.950 ;
        RECT 800.400 340.050 801.600 361.950 ;
        RECT 821.400 352.050 822.600 364.950 ;
        RECT 833.400 364.050 834.600 373.950 ;
        RECT 839.400 370.050 840.600 397.950 ;
        RECT 860.400 378.600 861.600 412.950 ;
        RECT 862.950 385.950 865.050 388.050 ;
        RECT 857.400 377.400 861.600 378.600 ;
        RECT 857.400 373.050 858.600 377.400 ;
        RECT 863.400 375.600 864.600 385.950 ;
        RECT 866.400 382.050 867.600 412.950 ;
        RECT 872.400 412.050 873.600 418.950 ;
        RECT 883.950 415.950 886.050 418.050 ;
        RECT 884.400 415.050 885.600 415.950 ;
        RECT 880.950 412.950 883.050 415.050 ;
        RECT 883.950 412.950 886.050 415.050 ;
        RECT 868.950 409.950 871.050 412.050 ;
        RECT 871.950 409.950 874.050 412.050 ;
        RECT 881.400 411.900 882.600 412.950 ;
        RECT 865.950 379.950 868.050 382.050 ;
        RECT 869.400 376.050 870.600 409.950 ;
        RECT 872.400 397.050 873.600 409.950 ;
        RECT 880.950 409.800 883.050 411.900 ;
        RECT 886.950 409.950 889.050 412.050 ;
        RECT 871.950 394.950 874.050 397.050 ;
        RECT 887.400 394.050 888.600 409.950 ;
        RECT 886.950 391.950 889.050 394.050 ;
        RECT 880.950 388.950 883.050 391.050 ;
        RECT 874.950 382.950 877.050 385.050 ;
        RECT 863.400 374.400 867.600 375.600 ;
        RECT 856.950 370.950 859.050 373.050 ;
        RECT 866.400 370.050 867.600 374.400 ;
        RECT 868.950 373.950 871.050 376.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 865.950 367.950 868.050 370.050 ;
        RECT 868.950 367.950 871.050 370.050 ;
        RECT 842.400 366.900 843.600 367.950 ;
        RECT 841.950 364.800 844.050 366.900 ;
        RECT 850.950 364.950 853.050 367.050 ;
        RECT 832.950 361.950 835.050 364.050 ;
        RECT 838.950 361.950 841.050 364.050 ;
        RECT 823.950 352.950 826.050 355.050 ;
        RECT 802.950 349.950 805.050 352.050 ;
        RECT 820.950 349.950 823.050 352.050 ;
        RECT 799.950 337.950 802.050 340.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 791.400 330.600 792.600 334.950 ;
        RECT 791.400 329.400 795.600 330.600 ;
        RECT 787.950 310.950 790.050 313.050 ;
        RECT 784.950 265.950 787.050 268.050 ;
        RECT 784.950 262.800 787.050 264.900 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 778.950 256.950 781.050 259.050 ;
        RECT 773.400 250.050 774.600 256.950 ;
        RECT 772.950 247.950 775.050 250.050 ;
        RECT 775.950 232.950 778.050 235.050 ;
        RECT 769.950 226.950 772.050 229.050 ;
        RECT 766.950 220.950 769.050 223.050 ;
        RECT 770.400 214.050 771.600 226.950 ;
        RECT 776.400 217.200 777.600 232.950 ;
        RECT 779.400 232.050 780.600 256.950 ;
        RECT 781.950 253.950 784.050 256.050 ;
        RECT 778.950 229.950 781.050 232.050 ;
        RECT 778.950 220.950 781.050 223.050 ;
        RECT 775.950 215.100 778.050 217.200 ;
        RECT 779.400 217.050 780.600 220.950 ;
        RECT 776.400 214.050 777.600 215.100 ;
        RECT 778.950 214.950 781.050 217.050 ;
        RECT 769.950 211.950 772.050 214.050 ;
        RECT 772.950 211.950 775.050 214.050 ;
        RECT 775.950 211.950 778.050 214.050 ;
        RECT 773.400 190.050 774.600 211.950 ;
        RECT 772.950 187.950 775.050 190.050 ;
        RECT 782.400 186.600 783.600 253.950 ;
        RECT 785.400 241.050 786.600 262.800 ;
        RECT 788.400 262.050 789.600 310.950 ;
        RECT 794.400 310.050 795.600 329.400 ;
        RECT 793.950 307.950 796.050 310.050 ;
        RECT 797.400 298.050 798.600 334.950 ;
        RECT 799.950 331.950 802.050 334.050 ;
        RECT 800.400 328.050 801.600 331.950 ;
        RECT 799.950 325.950 802.050 328.050 ;
        RECT 803.400 313.050 804.600 349.950 ;
        RECT 824.400 348.600 825.600 352.950 ;
        RECT 839.400 352.050 840.600 361.950 ;
        RECT 838.950 349.950 841.050 352.050 ;
        RECT 847.950 349.950 850.050 352.050 ;
        RECT 821.400 347.400 825.600 348.600 ;
        RECT 814.950 338.100 817.050 340.200 ;
        RECT 815.400 337.050 816.600 338.100 ;
        RECT 821.400 337.050 822.600 347.400 ;
        RECT 835.950 346.950 838.050 349.050 ;
        RECT 836.400 343.050 837.600 346.950 ;
        RECT 835.950 340.950 838.050 343.050 ;
        RECT 826.950 338.100 829.050 340.200 ;
        RECT 832.950 338.100 835.050 340.200 ;
        RECT 838.950 338.100 841.050 340.200 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 814.950 334.950 817.050 337.050 ;
        RECT 817.950 334.950 820.050 337.050 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 812.400 330.600 813.600 334.950 ;
        RECT 818.400 333.900 819.600 334.950 ;
        RECT 817.950 331.800 820.050 333.900 ;
        RECT 809.400 329.400 813.600 330.600 ;
        RECT 805.950 313.950 808.050 316.050 ;
        RECT 802.950 310.950 805.050 313.050 ;
        RECT 796.950 295.950 799.050 298.050 ;
        RECT 793.950 293.100 796.050 295.200 ;
        RECT 799.950 293.100 802.050 295.200 ;
        RECT 806.400 295.050 807.600 313.950 ;
        RECT 809.400 310.050 810.600 329.400 ;
        RECT 827.400 328.050 828.600 338.100 ;
        RECT 833.400 337.050 834.600 338.100 ;
        RECT 839.400 337.050 840.600 338.100 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 835.950 334.950 838.050 337.050 ;
        RECT 838.950 334.950 841.050 337.050 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 836.400 333.900 837.600 334.950 ;
        RECT 835.950 331.800 838.050 333.900 ;
        RECT 838.950 328.950 841.050 331.050 ;
        RECT 811.950 325.950 814.050 328.050 ;
        RECT 826.950 325.950 829.050 328.050 ;
        RECT 812.400 319.050 813.600 325.950 ;
        RECT 814.950 322.950 817.050 325.050 ;
        RECT 811.950 316.950 814.050 319.050 ;
        RECT 808.950 307.950 811.050 310.050 ;
        RECT 808.950 298.950 811.050 301.050 ;
        RECT 794.400 292.050 795.600 293.100 ;
        RECT 800.400 292.050 801.600 293.100 ;
        RECT 805.950 292.950 808.050 295.050 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 796.950 289.950 799.050 292.050 ;
        RECT 799.950 289.950 802.050 292.050 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 797.400 286.050 798.600 289.950 ;
        RECT 803.400 288.900 804.600 289.950 ;
        RECT 802.950 286.800 805.050 288.900 ;
        RECT 805.950 286.950 808.050 289.050 ;
        RECT 790.950 283.950 793.050 286.050 ;
        RECT 796.950 283.950 799.050 286.050 ;
        RECT 791.400 265.050 792.600 283.950 ;
        RECT 797.400 271.050 798.600 283.950 ;
        RECT 806.400 277.050 807.600 286.950 ;
        RECT 805.950 274.950 808.050 277.050 ;
        RECT 796.950 268.950 799.050 271.050 ;
        RECT 809.400 268.050 810.600 298.950 ;
        RECT 812.400 289.050 813.600 316.950 ;
        RECT 815.400 295.050 816.600 322.950 ;
        RECT 835.950 313.950 838.050 316.050 ;
        RECT 836.400 310.050 837.600 313.950 ;
        RECT 835.950 307.950 838.050 310.050 ;
        RECT 817.950 301.950 820.050 304.050 ;
        RECT 814.950 292.950 817.050 295.050 ;
        RECT 818.400 292.050 819.600 301.950 ;
        RECT 823.950 293.100 826.050 295.200 ;
        RECT 829.950 294.000 832.050 298.050 ;
        RECT 824.400 292.050 825.600 293.100 ;
        RECT 830.400 292.050 831.600 294.000 ;
        RECT 832.950 292.950 835.050 298.050 ;
        RECT 817.950 289.950 820.050 292.050 ;
        RECT 820.950 289.950 823.050 292.050 ;
        RECT 823.950 289.950 826.050 292.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 811.800 286.950 813.900 289.050 ;
        RECT 821.400 288.900 822.600 289.950 ;
        RECT 827.400 288.900 828.600 289.950 ;
        RECT 836.400 288.900 837.600 307.950 ;
        RECT 839.400 298.050 840.600 328.950 ;
        RECT 838.950 295.950 841.050 298.050 ;
        RECT 842.400 295.050 843.600 334.950 ;
        RECT 848.400 325.050 849.600 349.950 ;
        RECT 847.950 322.950 850.050 325.050 ;
        RECT 851.400 310.050 852.600 364.950 ;
        RECT 863.400 345.600 864.600 367.950 ;
        RECT 869.400 366.900 870.600 367.950 ;
        RECT 868.950 364.800 871.050 366.900 ;
        RECT 871.950 364.950 874.050 367.050 ;
        RECT 875.400 366.900 876.600 382.950 ;
        RECT 877.950 373.950 880.050 376.050 ;
        RECT 863.400 344.400 867.600 345.600 ;
        RECT 866.400 340.050 867.600 344.400 ;
        RECT 865.950 337.950 868.050 340.050 ;
        RECT 872.400 339.600 873.600 364.950 ;
        RECT 874.950 364.800 877.050 366.900 ;
        RECT 878.400 349.050 879.600 373.950 ;
        RECT 881.400 373.050 882.600 388.950 ;
        RECT 886.950 385.950 889.050 388.050 ;
        RECT 880.950 370.950 883.050 373.050 ;
        RECT 887.400 370.050 888.600 385.950 ;
        RECT 890.400 376.050 891.600 436.950 ;
        RECT 893.400 430.050 894.600 442.950 ;
        RECT 899.400 442.050 900.600 472.950 ;
        RECT 902.400 451.050 903.600 487.950 ;
        RECT 904.950 484.950 907.050 489.000 ;
        RECT 904.950 481.800 907.050 483.900 ;
        RECT 905.400 460.050 906.600 481.800 ;
        RECT 911.400 475.050 912.600 490.950 ;
        RECT 913.950 484.950 916.050 487.050 ;
        RECT 910.950 472.950 913.050 475.050 ;
        RECT 904.950 457.950 907.050 460.050 ;
        RECT 907.950 454.950 910.050 457.050 ;
        RECT 901.950 448.950 904.050 451.050 ;
        RECT 908.400 448.050 909.600 454.950 ;
        RECT 914.400 454.050 915.600 484.950 ;
        RECT 917.400 481.050 918.600 499.950 ;
        RECT 916.950 478.950 919.050 481.050 ;
        RECT 916.950 472.950 919.050 475.050 ;
        RECT 913.950 451.950 916.050 454.050 ;
        RECT 917.400 450.600 918.600 472.950 ;
        RECT 920.400 460.050 921.600 586.950 ;
        RECT 919.950 457.950 922.050 460.050 ;
        RECT 919.950 451.950 922.050 454.050 ;
        RECT 914.400 449.400 918.600 450.600 ;
        RECT 914.400 448.050 915.600 449.400 ;
        RECT 904.950 445.950 907.050 448.050 ;
        RECT 907.950 445.950 910.050 448.050 ;
        RECT 910.950 445.950 913.050 448.050 ;
        RECT 913.950 445.950 916.050 448.050 ;
        RECT 901.950 442.950 904.050 445.050 ;
        RECT 898.950 439.950 901.050 442.050 ;
        RECT 892.950 427.950 895.050 430.050 ;
        RECT 902.400 424.050 903.600 442.950 ;
        RECT 905.400 436.050 906.600 445.950 ;
        RECT 911.400 444.900 912.600 445.950 ;
        RECT 920.400 444.900 921.600 451.950 ;
        RECT 910.950 442.800 913.050 444.900 ;
        RECT 919.950 442.800 922.050 444.900 ;
        RECT 913.950 439.950 916.050 442.050 ;
        RECT 904.950 433.950 907.050 436.050 ;
        RECT 901.950 421.950 904.050 424.050 ;
        RECT 907.950 421.950 910.050 424.050 ;
        RECT 901.950 412.950 904.050 415.050 ;
        RECT 902.400 411.900 903.600 412.950 ;
        RECT 901.950 409.800 904.050 411.900 ;
        RECT 902.400 400.050 903.600 409.800 ;
        RECT 901.950 397.950 904.050 400.050 ;
        RECT 901.950 391.950 904.050 394.050 ;
        RECT 898.950 385.950 901.050 388.050 ;
        RECT 889.950 373.950 892.050 376.050 ;
        RECT 899.400 373.050 900.600 385.950 ;
        RECT 902.400 376.050 903.600 391.950 ;
        RECT 908.400 388.050 909.600 421.950 ;
        RECT 910.950 397.950 913.050 400.050 ;
        RECT 907.950 385.950 910.050 388.050 ;
        RECT 907.950 379.950 910.050 382.050 ;
        RECT 901.950 373.950 904.050 376.050 ;
        RECT 898.950 370.950 901.050 373.050 ;
        RECT 902.400 370.050 903.600 373.950 ;
        RECT 908.400 370.050 909.600 379.950 ;
        RECT 911.400 373.050 912.600 397.950 ;
        RECT 910.950 370.950 913.050 373.050 ;
        RECT 883.950 367.950 886.050 370.050 ;
        RECT 886.950 367.950 889.050 370.050 ;
        RECT 901.950 367.950 904.050 370.050 ;
        RECT 904.950 367.950 907.050 370.050 ;
        RECT 907.950 367.950 910.050 370.050 ;
        RECT 880.950 364.950 883.050 367.050 ;
        RECT 877.950 346.950 880.050 349.050 ;
        RECT 869.400 338.400 873.600 339.600 ;
        RECT 881.400 339.600 882.600 364.950 ;
        RECT 884.400 361.050 885.600 367.950 ;
        RECT 892.950 364.950 895.050 367.050 ;
        RECT 898.950 364.950 901.050 367.050 ;
        RECT 883.950 358.950 886.050 361.050 ;
        RECT 893.400 349.050 894.600 364.950 ;
        RECT 895.950 352.950 898.050 355.050 ;
        RECT 886.950 346.950 889.050 349.050 ;
        RECT 892.950 346.950 895.050 349.050 ;
        RECT 887.400 340.050 888.600 346.950 ;
        RECT 881.400 338.400 885.600 339.600 ;
        RECT 859.950 334.950 862.050 337.050 ;
        RECT 860.400 328.050 861.600 334.950 ;
        RECT 859.950 325.950 862.050 328.050 ;
        RECT 865.950 316.950 868.050 319.050 ;
        RECT 850.950 307.950 853.050 310.050 ;
        RECT 866.400 304.050 867.600 316.950 ;
        RECT 865.950 301.950 868.050 304.050 ;
        RECT 844.950 295.950 847.050 301.050 ;
        RECT 850.950 298.950 856.050 301.050 ;
        RECT 865.950 298.800 868.050 300.900 ;
        RECT 841.950 292.950 844.050 295.050 ;
        RECT 847.950 293.100 850.050 295.200 ;
        RECT 853.950 294.000 856.050 297.900 ;
        RECT 862.950 295.950 865.050 298.050 ;
        RECT 848.400 292.050 849.600 293.100 ;
        RECT 854.400 292.050 855.600 294.000 ;
        RECT 859.950 293.100 862.050 295.200 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 844.950 289.950 847.050 292.050 ;
        RECT 847.950 289.950 850.050 292.050 ;
        RECT 850.950 289.950 853.050 292.050 ;
        RECT 853.950 289.950 856.050 292.050 ;
        RECT 814.950 286.800 817.050 288.900 ;
        RECT 820.950 286.800 823.050 288.900 ;
        RECT 826.950 286.800 829.050 288.900 ;
        RECT 835.950 286.800 838.050 288.900 ;
        RECT 802.950 265.950 805.050 268.050 ;
        RECT 808.950 265.950 811.050 268.050 ;
        RECT 787.950 259.950 790.050 262.050 ;
        RECT 790.950 261.000 793.050 265.050 ;
        RECT 796.950 261.000 799.050 265.050 ;
        RECT 791.400 259.050 792.600 261.000 ;
        RECT 797.400 259.050 798.600 261.000 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 796.950 256.950 799.050 259.050 ;
        RECT 794.400 250.050 795.600 256.950 ;
        RECT 803.400 255.600 804.600 265.950 ;
        RECT 808.950 261.000 811.050 264.900 ;
        RECT 815.400 262.050 816.600 286.800 ;
        RECT 817.950 283.950 820.050 286.050 ;
        RECT 818.400 280.050 819.600 283.950 ;
        RECT 839.400 283.050 840.600 289.950 ;
        RECT 841.950 283.950 844.050 289.050 ;
        RECT 820.950 280.950 823.050 283.050 ;
        RECT 838.800 280.950 840.900 283.050 ;
        RECT 817.950 277.950 820.050 280.050 ;
        RECT 809.400 259.050 810.600 261.000 ;
        RECT 814.950 259.950 817.050 262.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 800.400 254.400 804.600 255.600 ;
        RECT 793.950 247.950 796.050 250.050 ;
        RECT 790.950 241.950 793.050 244.050 ;
        RECT 784.950 238.950 787.050 241.050 ;
        RECT 791.400 232.050 792.600 241.950 ;
        RECT 790.950 229.950 793.050 232.050 ;
        RECT 796.950 229.950 799.050 232.050 ;
        RECT 784.800 214.950 786.900 217.050 ;
        RECT 779.400 185.400 783.600 186.600 ;
        RECT 769.950 175.950 772.050 178.050 ;
        RECT 763.950 148.950 766.050 151.050 ;
        RECT 763.950 142.950 766.050 145.050 ;
        RECT 757.800 139.800 759.900 141.900 ;
        RECT 760.950 139.950 763.050 142.050 ;
        RECT 748.950 137.100 751.050 139.200 ;
        RECT 749.400 136.050 750.600 137.100 ;
        RECT 754.950 136.950 757.050 139.050 ;
        RECT 742.950 133.950 745.050 136.050 ;
        RECT 745.950 133.950 748.050 136.050 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 746.400 132.900 747.600 133.950 ;
        RECT 755.400 132.900 756.600 136.950 ;
        RECT 745.950 130.800 748.050 132.900 ;
        RECT 754.950 130.800 757.050 132.900 ;
        RECT 755.400 127.050 756.600 130.800 ;
        RECT 754.950 124.950 757.050 127.050 ;
        RECT 736.950 106.950 739.050 109.050 ;
        RECT 727.800 103.950 729.900 106.050 ;
        RECT 730.950 104.100 733.050 106.200 ;
        RECT 739.950 104.100 742.050 106.200 ;
        RECT 745.950 105.000 748.050 109.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 718.950 100.950 721.050 103.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 724.950 100.950 727.050 103.050 ;
        RECT 719.400 93.600 720.600 100.950 ;
        RECT 725.400 99.900 726.600 100.950 ;
        RECT 724.950 97.800 727.050 99.900 ;
        RECT 727.950 97.950 730.050 100.050 ;
        RECT 721.950 93.600 724.050 97.050 ;
        RECT 719.400 93.000 724.050 93.600 ;
        RECT 719.400 92.400 723.600 93.000 ;
        RECT 709.950 85.950 712.050 88.050 ;
        RECT 712.950 68.400 715.050 70.500 ;
        RECT 701.400 59.400 705.600 60.600 ;
        RECT 706.950 60.000 709.050 64.050 ;
        RECT 701.400 49.050 702.600 59.400 ;
        RECT 707.400 58.050 708.600 60.000 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 691.950 46.500 694.050 48.600 ;
        RECT 700.950 46.950 703.050 49.050 ;
        RECT 713.100 48.600 714.300 68.400 ;
        RECT 715.950 59.400 718.050 61.500 ;
        RECT 716.400 58.050 717.600 59.400 ;
        RECT 715.950 55.950 718.050 58.050 ;
        RECT 722.400 52.050 723.600 92.400 ;
        RECT 728.400 61.500 729.600 97.950 ;
        RECT 731.400 97.050 732.600 104.100 ;
        RECT 740.400 103.050 741.600 104.100 ;
        RECT 746.400 103.050 747.600 105.000 ;
        RECT 754.950 103.950 757.050 106.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 742.950 100.950 745.050 103.050 ;
        RECT 745.950 100.950 748.050 103.050 ;
        RECT 748.950 100.950 751.050 103.050 ;
        RECT 737.400 99.600 738.600 100.950 ;
        RECT 734.400 98.400 738.600 99.600 ;
        RECT 730.950 94.950 733.050 97.050 ;
        RECT 727.950 59.400 730.050 61.500 ;
        RECT 721.950 49.950 724.050 52.050 ;
        RECT 712.950 46.500 715.050 48.600 ;
        RECT 712.950 32.400 715.050 34.500 ;
        RECT 682.950 26.100 685.050 28.200 ;
        RECT 694.950 26.100 697.050 28.200 ;
        RECT 695.400 25.050 696.600 26.100 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 673.950 22.950 676.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 694.950 22.950 697.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 674.400 21.900 675.600 22.950 ;
        RECT 673.950 19.800 676.050 21.900 ;
        RECT 710.400 21.600 711.600 22.950 ;
        RECT 709.950 19.500 712.050 21.600 ;
        RECT 664.950 13.950 667.050 16.050 ;
        RECT 610.950 10.950 613.050 13.050 ;
        RECT 713.700 12.600 714.900 32.400 ;
        RECT 724.950 31.950 727.050 34.050 ;
        RECT 718.950 22.950 721.050 25.050 ;
        RECT 719.400 21.600 720.600 22.950 ;
        RECT 725.400 21.600 726.600 31.950 ;
        RECT 728.400 21.600 729.600 59.400 ;
        RECT 734.400 58.050 735.600 98.400 ;
        RECT 733.950 55.950 736.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 737.400 40.050 738.600 55.950 ;
        RECT 736.950 37.950 739.050 40.050 ;
        RECT 733.950 32.400 736.050 34.500 ;
        RECT 743.400 34.050 744.600 100.950 ;
        RECT 745.950 91.950 748.050 94.050 ;
        RECT 746.400 73.050 747.600 91.950 ;
        RECT 749.400 88.050 750.600 100.950 ;
        RECT 748.950 85.950 751.050 88.050 ;
        RECT 751.950 82.950 754.050 85.050 ;
        RECT 745.950 70.950 748.050 73.050 ;
        RECT 752.400 58.050 753.600 82.950 ;
        RECT 755.400 64.050 756.600 103.950 ;
        RECT 758.400 97.050 759.600 139.800 ;
        RECT 764.400 139.050 765.600 142.950 ;
        RECT 770.400 142.050 771.600 175.950 ;
        RECT 772.950 145.950 775.050 148.050 ;
        RECT 766.800 141.000 768.900 142.050 ;
        RECT 766.800 139.950 769.050 141.000 ;
        RECT 769.950 139.950 772.050 142.050 ;
        RECT 760.950 136.800 763.050 138.900 ;
        RECT 763.950 136.950 766.050 139.050 ;
        RECT 766.950 138.000 769.050 139.950 ;
        RECT 761.400 112.050 762.600 136.800 ;
        RECT 767.400 136.050 768.600 138.000 ;
        RECT 773.400 136.050 774.600 145.950 ;
        RECT 779.400 145.050 780.600 185.400 ;
        RECT 785.400 183.600 786.600 214.950 ;
        RECT 791.400 214.050 792.600 229.950 ;
        RECT 797.400 217.050 798.600 229.950 ;
        RECT 796.950 214.950 799.050 217.050 ;
        RECT 790.950 211.950 793.050 214.050 ;
        RECT 793.950 211.950 796.050 214.050 ;
        RECT 787.950 208.950 790.050 211.050 ;
        RECT 788.400 186.600 789.600 208.950 ;
        RECT 794.400 205.050 795.600 211.950 ;
        RECT 793.950 202.950 796.050 205.050 ;
        RECT 788.400 185.400 792.600 186.600 ;
        RECT 782.400 182.400 786.600 183.600 ;
        RECT 782.400 175.050 783.600 182.400 ;
        RECT 791.400 181.050 792.600 185.400 ;
        RECT 796.800 182.100 798.900 184.200 ;
        RECT 800.400 184.050 801.600 254.400 ;
        RECT 805.950 253.950 808.050 256.050 ;
        RECT 802.950 250.950 805.050 253.050 ;
        RECT 803.400 217.050 804.600 250.950 ;
        RECT 806.400 228.600 807.600 253.950 ;
        RECT 806.400 227.400 810.600 228.600 ;
        RECT 805.950 223.950 808.050 226.050 ;
        RECT 802.950 214.950 805.050 217.050 ;
        RECT 806.400 214.050 807.600 223.950 ;
        RECT 809.400 220.050 810.600 227.400 ;
        RECT 812.400 226.050 813.600 256.950 ;
        RECT 814.950 253.950 817.050 256.050 ;
        RECT 815.400 232.050 816.600 253.950 ;
        RECT 814.950 229.950 817.050 232.050 ;
        RECT 811.950 223.950 814.050 226.050 ;
        RECT 818.400 223.050 819.600 277.950 ;
        RECT 821.400 255.600 822.600 280.950 ;
        RECT 841.950 280.800 844.050 282.900 ;
        RECT 842.400 268.050 843.600 280.800 ;
        RECT 845.400 277.050 846.600 289.950 ;
        RECT 851.400 288.900 852.600 289.950 ;
        RECT 850.950 286.800 853.050 288.900 ;
        RECT 856.950 280.950 859.050 286.050 ;
        RECT 860.400 280.050 861.600 293.100 ;
        RECT 863.400 289.050 864.600 295.950 ;
        RECT 866.400 294.600 867.600 298.800 ;
        RECT 869.400 298.050 870.600 338.400 ;
        RECT 877.950 334.950 880.050 337.050 ;
        RECT 871.950 331.950 874.050 334.050 ;
        RECT 868.950 295.950 871.050 298.050 ;
        RECT 872.400 297.600 873.600 331.950 ;
        RECT 878.400 316.050 879.600 334.950 ;
        RECT 877.950 313.950 880.050 316.050 ;
        RECT 872.400 296.400 876.600 297.600 ;
        RECT 866.400 293.400 870.600 294.600 ;
        RECT 869.400 292.050 870.600 293.400 ;
        RECT 875.400 292.050 876.600 296.400 ;
        RECT 877.950 292.950 880.050 298.050 ;
        RECT 880.950 292.950 883.050 295.050 ;
        RECT 868.950 289.950 871.050 292.050 ;
        RECT 871.950 289.950 874.050 292.050 ;
        RECT 874.950 289.950 877.050 292.050 ;
        RECT 862.950 286.950 865.050 289.050 ;
        RECT 865.950 283.950 871.050 286.050 ;
        RECT 859.950 277.950 862.050 280.050 ;
        RECT 844.950 274.950 847.050 277.050 ;
        RECT 853.950 274.950 856.050 277.050 ;
        RECT 845.400 271.050 846.600 274.950 ;
        RECT 844.950 268.950 847.050 271.050 ;
        RECT 823.950 265.950 826.050 268.050 ;
        RECT 841.950 265.950 844.050 268.050 ;
        RECT 824.400 262.050 825.600 265.950 ;
        RECT 823.950 259.950 826.050 262.050 ;
        RECT 826.950 260.100 829.050 262.200 ;
        RECT 832.950 260.100 835.050 265.050 ;
        RECT 827.400 259.050 828.600 260.100 ;
        RECT 833.400 259.050 834.600 260.100 ;
        RECT 826.950 256.950 829.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 838.950 258.000 841.050 262.200 ;
        RECT 821.400 254.400 825.600 255.600 ;
        RECT 820.950 250.950 823.050 253.050 ;
        RECT 821.400 244.050 822.600 250.950 ;
        RECT 820.950 241.950 823.050 244.050 ;
        RECT 817.950 220.950 820.050 223.050 ;
        RECT 824.400 220.050 825.600 254.400 ;
        RECT 830.400 247.050 831.600 256.950 ;
        RECT 839.400 256.050 840.600 258.000 ;
        RECT 847.950 257.100 850.050 259.200 ;
        RECT 848.400 256.050 849.600 257.100 ;
        RECT 838.950 253.950 841.050 256.050 ;
        RECT 847.950 253.950 850.050 256.050 ;
        RECT 835.950 250.950 838.050 253.050 ;
        RECT 829.950 244.950 832.050 247.050 ;
        RECT 808.950 217.950 811.050 220.050 ;
        RECT 823.950 217.950 826.050 220.050 ;
        RECT 811.950 215.100 814.050 217.200 ;
        RECT 812.400 214.050 813.600 215.100 ;
        RECT 820.950 214.950 823.050 217.050 ;
        RECT 829.950 214.950 832.050 217.050 ;
        RECT 805.950 211.950 808.050 214.050 ;
        RECT 808.950 211.950 811.050 214.050 ;
        RECT 811.950 211.950 814.050 214.050 ;
        RECT 814.950 211.950 817.050 214.050 ;
        RECT 821.400 213.900 822.600 214.950 ;
        RECT 830.400 213.900 831.600 214.950 ;
        RECT 836.400 213.900 837.600 250.950 ;
        RECT 854.400 247.050 855.600 274.950 ;
        RECT 872.400 274.050 873.600 289.950 ;
        RECT 881.400 286.050 882.600 292.950 ;
        RECT 880.950 283.950 883.050 286.050 ;
        RECT 877.950 280.950 880.050 283.050 ;
        RECT 878.400 274.050 879.600 280.950 ;
        RECT 884.400 274.050 885.600 338.400 ;
        RECT 886.950 337.950 889.050 340.050 ;
        RECT 896.400 337.050 897.600 352.950 ;
        RECT 899.400 343.050 900.600 364.950 ;
        RECT 901.950 358.950 904.050 361.050 ;
        RECT 902.400 354.600 903.600 358.950 ;
        RECT 905.400 358.050 906.600 367.950 ;
        RECT 910.950 364.950 913.050 367.050 ;
        RECT 907.950 358.950 910.050 361.050 ;
        RECT 904.950 355.950 907.050 358.050 ;
        RECT 902.400 353.400 906.600 354.600 ;
        RECT 901.950 346.950 904.050 349.050 ;
        RECT 898.950 340.950 901.050 343.050 ;
        RECT 902.400 340.050 903.600 346.950 ;
        RECT 901.950 337.950 904.050 340.050 ;
        RECT 889.950 334.950 892.050 337.050 ;
        RECT 895.950 334.950 898.050 337.050 ;
        RECT 898.950 334.950 901.050 337.050 ;
        RECT 886.950 331.950 889.050 334.050 ;
        RECT 887.400 295.050 888.600 331.950 ;
        RECT 890.400 310.050 891.600 334.950 ;
        RECT 889.950 307.950 892.050 310.050 ;
        RECT 892.950 301.950 895.050 304.050 ;
        RECT 886.950 292.950 889.050 295.050 ;
        RECT 893.400 292.050 894.600 301.950 ;
        RECT 899.400 292.050 900.600 334.950 ;
        RECT 901.950 331.950 904.050 334.050 ;
        RECT 902.400 294.600 903.600 331.950 ;
        RECT 905.400 304.050 906.600 353.400 ;
        RECT 908.400 349.050 909.600 358.950 ;
        RECT 907.950 346.950 910.050 349.050 ;
        RECT 907.950 340.950 910.050 343.050 ;
        RECT 904.950 301.950 907.050 304.050 ;
        RECT 902.400 293.400 906.600 294.600 ;
        RECT 889.950 289.950 892.050 292.050 ;
        RECT 892.950 289.950 895.050 292.050 ;
        RECT 895.950 289.950 898.050 292.050 ;
        RECT 898.950 289.950 901.050 292.050 ;
        RECT 886.950 286.950 889.050 289.050 ;
        RECT 890.400 288.900 891.600 289.950 ;
        RECT 887.400 277.050 888.600 286.950 ;
        RECT 889.950 286.800 892.050 288.900 ;
        RECT 896.400 283.050 897.600 289.950 ;
        RECT 895.950 280.950 898.050 283.050 ;
        RECT 886.950 274.950 889.050 277.050 ;
        RECT 892.950 276.600 895.050 277.050 ;
        RECT 892.950 275.400 900.600 276.600 ;
        RECT 892.950 274.950 895.050 275.400 ;
        RECT 871.950 271.950 874.050 274.050 ;
        RECT 877.950 271.950 880.050 274.050 ;
        RECT 883.950 271.950 886.050 274.050 ;
        RECT 895.950 271.950 898.050 274.050 ;
        RECT 859.950 266.400 862.050 268.500 ;
        RECT 856.950 262.950 859.050 265.050 ;
        RECT 857.400 253.050 858.600 262.950 ;
        RECT 856.950 250.950 859.050 253.050 ;
        RECT 860.850 249.600 862.050 266.400 ;
        RECT 859.950 247.500 862.050 249.600 ;
        RECT 853.950 244.950 856.050 247.050 ;
        RECT 860.850 242.700 862.050 247.500 ;
        RECT 862.950 266.400 865.050 268.500 ;
        RECT 865.950 266.400 868.050 268.500 ;
        RECT 868.950 266.400 871.050 268.500 ;
        RECT 874.950 266.400 877.050 268.500 ;
        RECT 883.950 266.400 886.050 268.500 ;
        RECT 886.950 266.400 889.050 268.500 ;
        RECT 889.950 266.400 892.050 268.500 ;
        RECT 862.950 245.700 864.150 266.400 ;
        RECT 865.950 249.600 867.450 266.400 ;
        RECT 869.850 254.700 871.050 266.400 ;
        RECT 875.250 254.700 876.450 266.400 ;
        RECT 877.950 259.950 880.050 262.050 ;
        RECT 878.400 258.900 879.600 259.950 ;
        RECT 877.950 256.800 880.050 258.900 ;
        RECT 868.950 252.600 871.050 254.700 ;
        RECT 874.950 252.600 877.050 254.700 ;
        RECT 865.950 247.500 868.050 249.600 ;
        RECT 859.950 240.600 862.050 242.700 ;
        RECT 863.100 242.700 864.150 245.700 ;
        RECT 866.100 242.700 867.300 247.500 ;
        RECT 869.850 245.700 871.050 252.600 ;
        RECT 875.850 247.200 877.050 252.600 ;
        RECT 868.950 243.600 871.050 245.700 ;
        RECT 874.950 245.100 877.050 247.200 ;
        RECT 883.950 245.400 885.150 266.400 ;
        RECT 886.950 250.800 888.150 266.400 ;
        RECT 886.950 248.700 889.050 250.800 ;
        RECT 887.400 245.400 888.600 248.700 ;
        RECT 890.400 245.400 891.600 266.400 ;
        RECT 896.400 262.050 897.600 271.950 ;
        RECT 895.950 259.950 898.050 262.050 ;
        RECT 899.400 259.050 900.600 275.400 ;
        RECT 898.950 256.950 901.050 259.050 ;
        RECT 905.400 258.600 906.600 293.400 ;
        RECT 908.400 261.600 909.600 340.950 ;
        RECT 911.400 288.900 912.600 364.950 ;
        RECT 914.400 361.050 915.600 439.950 ;
        RECT 916.950 436.950 919.050 439.050 ;
        RECT 913.950 358.950 916.050 361.050 ;
        RECT 913.950 352.950 916.050 355.050 ;
        RECT 910.950 286.800 913.050 288.900 ;
        RECT 908.400 260.400 912.600 261.600 ;
        RECT 905.400 257.400 909.600 258.600 ;
        RECT 901.950 253.950 904.050 256.050 ;
        RECT 895.950 247.950 898.050 250.050 ;
        RECT 883.950 243.300 886.050 245.400 ;
        RECT 886.950 243.300 889.050 245.400 ;
        RECT 889.950 243.300 892.050 245.400 ;
        RECT 863.100 240.600 865.200 242.700 ;
        RECT 866.100 240.600 868.200 242.700 ;
        RECT 856.950 235.950 859.050 238.050 ;
        RECT 841.950 228.300 844.050 230.400 ;
        RECT 842.850 223.500 844.050 228.300 ;
        RECT 845.100 228.300 847.200 230.400 ;
        RECT 848.100 228.300 850.200 230.400 ;
        RECT 857.400 229.050 858.600 235.950 ;
        RECT 845.100 225.300 846.150 228.300 ;
        RECT 841.950 221.400 844.050 223.500 ;
        RECT 838.950 217.950 841.050 220.050 ;
        RECT 802.950 208.950 805.050 211.050 ;
        RECT 809.400 210.900 810.600 211.950 ;
        RECT 797.400 181.050 798.600 182.100 ;
        RECT 799.950 181.950 802.050 184.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 793.950 178.950 796.050 181.050 ;
        RECT 796.950 178.950 799.050 181.050 ;
        RECT 788.400 177.000 789.600 178.950 ;
        RECT 794.400 177.000 795.600 178.950 ;
        RECT 781.950 172.950 784.050 175.050 ;
        RECT 787.950 172.950 790.050 177.000 ;
        RECT 793.950 172.950 796.050 177.000 ;
        RECT 790.950 169.950 793.050 172.050 ;
        RECT 781.950 154.950 784.050 157.050 ;
        RECT 778.950 142.950 781.050 145.050 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 763.950 130.950 766.050 133.050 ;
        RECT 764.400 121.050 765.600 130.950 ;
        RECT 770.400 126.600 771.600 133.950 ;
        RECT 776.400 132.900 777.600 133.950 ;
        RECT 775.950 127.950 778.050 132.900 ;
        RECT 778.950 130.950 781.050 133.050 ;
        RECT 782.400 132.900 783.600 154.950 ;
        RECT 791.400 141.600 792.600 169.950 ;
        RECT 803.400 169.050 804.600 208.950 ;
        RECT 808.950 208.800 811.050 210.900 ;
        RECT 811.950 187.950 814.050 190.050 ;
        RECT 815.400 189.600 816.600 211.950 ;
        RECT 820.950 211.800 823.050 213.900 ;
        RECT 829.950 211.800 832.050 213.900 ;
        RECT 835.950 211.800 838.050 213.900 ;
        RECT 821.400 205.050 822.600 211.800 ;
        RECT 823.950 208.950 826.050 211.050 ;
        RECT 820.950 202.950 823.050 205.050 ;
        RECT 820.950 190.950 823.050 193.050 ;
        RECT 815.400 188.400 819.600 189.600 ;
        RECT 805.950 181.950 808.050 184.050 ;
        RECT 806.400 178.050 807.600 181.950 ;
        RECT 812.400 181.050 813.600 187.950 ;
        RECT 818.400 184.050 819.600 188.400 ;
        RECT 817.950 181.950 820.050 184.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 814.950 178.950 817.050 181.050 ;
        RECT 805.950 175.950 808.050 178.050 ;
        RECT 815.400 177.900 816.600 178.950 ;
        RECT 821.400 178.050 822.600 190.950 ;
        RECT 814.950 175.800 817.050 177.900 ;
        RECT 817.950 175.950 820.050 178.050 ;
        RECT 820.950 175.950 823.050 178.050 ;
        RECT 802.950 166.950 805.050 169.050 ;
        RECT 815.400 151.050 816.600 175.800 ;
        RECT 818.400 157.050 819.600 175.950 ;
        RECT 824.400 157.050 825.600 208.950 ;
        RECT 829.950 205.950 832.050 208.050 ;
        RECT 830.400 196.050 831.600 205.950 ;
        RECT 832.950 202.950 835.050 205.050 ;
        RECT 829.950 193.950 832.050 196.050 ;
        RECT 833.400 193.050 834.600 202.950 ;
        RECT 836.400 199.050 837.600 211.800 ;
        RECT 839.400 208.050 840.600 217.950 ;
        RECT 838.950 205.950 841.050 208.050 ;
        RECT 842.850 204.600 844.050 221.400 ;
        RECT 841.950 202.500 844.050 204.600 ;
        RECT 844.950 204.600 846.150 225.300 ;
        RECT 848.100 223.500 849.300 228.300 ;
        RECT 850.950 225.300 853.050 227.400 ;
        RECT 856.950 226.950 859.050 229.050 ;
        RECT 847.950 221.400 850.050 223.500 ;
        RECT 847.950 204.600 849.450 221.400 ;
        RECT 851.850 218.400 853.050 225.300 ;
        RECT 856.950 223.800 859.050 225.900 ;
        RECT 857.850 218.400 859.050 223.800 ;
        RECT 850.950 216.300 853.050 218.400 ;
        RECT 856.950 216.300 859.050 218.400 ;
        RECT 865.950 225.600 868.050 227.700 ;
        RECT 868.950 225.600 871.050 227.700 ;
        RECT 871.950 225.600 874.050 227.700 ;
        RECT 892.950 226.950 895.050 229.050 ;
        RECT 851.850 204.600 853.050 216.300 ;
        RECT 857.250 204.600 858.450 216.300 ;
        RECT 859.950 212.100 862.050 214.200 ;
        RECT 860.400 211.050 861.600 212.100 ;
        RECT 859.950 208.950 862.050 211.050 ;
        RECT 865.950 204.600 867.150 225.600 ;
        RECT 869.400 222.300 870.600 225.600 ;
        RECT 868.950 220.200 871.050 222.300 ;
        RECT 868.950 204.600 870.150 220.200 ;
        RECT 872.400 204.600 873.600 225.600 ;
        RECT 889.950 220.950 892.050 223.050 ;
        RECT 877.950 214.950 880.050 217.050 ;
        RECT 878.400 213.900 879.600 214.950 ;
        RECT 877.950 211.800 880.050 213.900 ;
        RECT 844.950 202.500 847.050 204.600 ;
        RECT 847.950 202.500 850.050 204.600 ;
        RECT 850.950 202.500 853.050 204.600 ;
        RECT 856.950 202.500 859.050 204.600 ;
        RECT 865.950 202.500 868.050 204.600 ;
        RECT 868.950 202.500 871.050 204.600 ;
        RECT 871.950 202.500 874.050 204.600 ;
        RECT 835.950 196.950 838.050 199.050 ;
        RECT 850.950 196.950 853.050 199.050 ;
        RECT 856.950 196.950 859.050 199.050 ;
        RECT 832.950 190.950 835.050 193.050 ;
        RECT 826.950 182.100 829.050 187.050 ;
        RECT 832.950 182.100 835.050 184.200 ;
        RECT 833.400 181.050 834.600 182.100 ;
        RECT 851.400 181.200 852.600 196.950 ;
        RECT 853.950 193.950 856.050 196.050 ;
        RECT 854.400 184.050 855.600 193.950 ;
        RECT 853.950 181.950 856.050 184.050 ;
        RECT 857.400 183.600 858.600 196.950 ;
        RECT 878.400 196.050 879.600 211.800 ;
        RECT 890.400 205.050 891.600 220.950 ;
        RECT 889.950 202.950 892.050 205.050 ;
        RECT 893.400 202.050 894.600 226.950 ;
        RECT 892.950 199.950 895.050 202.050 ;
        RECT 896.400 199.050 897.600 247.950 ;
        RECT 902.400 217.200 903.600 253.950 ;
        RECT 904.950 250.950 907.050 253.050 ;
        RECT 905.400 220.050 906.600 250.950 ;
        RECT 908.400 223.050 909.600 257.400 ;
        RECT 911.400 229.050 912.600 260.400 ;
        RECT 910.950 226.950 913.050 229.050 ;
        RECT 907.950 220.950 910.050 223.050 ;
        RECT 904.950 217.950 907.050 220.050 ;
        RECT 910.950 217.950 913.050 220.050 ;
        RECT 901.950 215.100 904.050 217.200 ;
        RECT 902.400 214.050 903.600 215.100 ;
        RECT 901.950 211.950 904.050 214.050 ;
        RECT 907.950 208.950 910.050 211.050 ;
        RECT 898.950 202.950 901.050 205.050 ;
        RECT 895.950 196.950 898.050 199.050 ;
        RECT 877.950 193.950 880.050 196.050 ;
        RECT 862.950 188.400 865.050 190.500 ;
        RECT 857.400 182.400 861.600 183.600 ;
        RECT 829.950 178.950 832.050 181.050 ;
        RECT 832.950 178.950 835.050 181.050 ;
        RECT 841.950 179.100 844.050 181.200 ;
        RECT 850.950 179.100 853.050 181.200 ;
        RECT 856.950 179.100 859.050 181.200 ;
        RECT 830.400 177.900 831.600 178.950 ;
        RECT 842.400 178.050 843.600 179.100 ;
        RECT 851.400 178.050 852.600 179.100 ;
        RECT 829.950 177.600 832.050 177.900 ;
        RECT 827.400 177.000 832.050 177.600 ;
        RECT 826.950 176.400 832.050 177.000 ;
        RECT 826.950 172.950 829.050 176.400 ;
        RECT 829.950 175.800 832.050 176.400 ;
        RECT 841.950 175.950 844.050 178.050 ;
        RECT 850.950 175.950 853.050 178.050 ;
        RECT 857.400 174.600 858.600 179.100 ;
        RECT 860.400 175.050 861.600 182.400 ;
        RECT 854.400 173.400 858.600 174.600 ;
        RECT 826.950 166.950 829.050 169.050 ;
        RECT 817.950 154.950 820.050 157.050 ;
        RECT 823.950 154.950 826.050 157.050 ;
        RECT 808.950 148.950 811.050 151.050 ;
        RECT 814.950 148.950 817.050 151.050 ;
        RECT 823.950 148.950 826.050 151.050 ;
        RECT 791.400 140.400 795.600 141.600 ;
        RECT 794.400 139.200 795.600 140.400 ;
        RECT 802.950 139.950 805.050 142.050 ;
        RECT 784.950 138.600 789.000 139.050 ;
        RECT 784.950 136.950 789.600 138.600 ;
        RECT 793.950 137.100 796.050 139.200 ;
        RECT 788.400 136.050 789.600 136.950 ;
        RECT 794.400 136.050 795.600 137.100 ;
        RECT 787.950 133.950 790.050 136.050 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 791.400 132.900 792.600 133.950 ;
        RECT 779.400 126.600 780.600 130.950 ;
        RECT 781.950 130.800 784.050 132.900 ;
        RECT 790.950 130.800 793.050 132.900 ;
        RECT 770.400 125.400 780.600 126.600 ;
        RECT 763.950 118.950 766.050 121.050 ;
        RECT 784.950 118.950 787.050 121.050 ;
        RECT 760.950 109.950 763.050 112.050 ;
        RECT 769.950 109.950 772.050 112.050 ;
        RECT 763.950 105.000 766.050 109.050 ;
        RECT 764.400 103.050 765.600 105.000 ;
        RECT 770.400 103.050 771.600 109.950 ;
        RECT 785.400 103.050 786.600 118.950 ;
        RECT 791.400 118.050 792.600 130.800 ;
        RECT 790.950 115.950 793.050 118.050 ;
        RECT 791.400 112.050 792.600 115.950 ;
        RECT 790.950 109.950 793.050 112.050 ;
        RECT 797.400 106.200 798.600 133.950 ;
        RECT 803.400 133.050 804.600 139.950 ;
        RECT 809.400 136.050 810.600 148.950 ;
        RECT 816.000 138.600 820.050 139.050 ;
        RECT 815.400 136.950 820.050 138.600 ;
        RECT 815.400 136.050 816.600 136.950 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 802.950 130.950 805.050 133.050 ;
        RECT 812.400 132.900 813.600 133.950 ;
        RECT 811.950 130.800 814.050 132.900 ;
        RECT 817.950 127.950 820.050 133.050 ;
        RECT 821.400 106.200 822.600 133.950 ;
        RECT 790.950 104.100 793.050 106.200 ;
        RECT 796.950 104.100 799.050 106.200 ;
        RECT 808.950 104.100 811.050 106.200 ;
        RECT 814.950 104.100 817.050 106.200 ;
        RECT 820.950 104.100 823.050 106.200 ;
        RECT 791.400 103.050 792.600 104.100 ;
        RECT 809.400 103.050 810.600 104.100 ;
        RECT 815.400 103.050 816.600 104.100 ;
        RECT 763.950 100.950 766.050 103.050 ;
        RECT 766.950 100.950 769.050 103.050 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 808.950 100.950 811.050 103.050 ;
        RECT 811.950 100.950 814.050 103.050 ;
        RECT 814.950 100.950 817.050 103.050 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 767.400 99.900 768.600 100.950 ;
        RECT 766.950 97.800 769.050 99.900 ;
        RECT 757.950 94.950 760.050 97.050 ;
        RECT 757.950 64.950 760.050 67.050 ;
        RECT 754.950 61.950 757.050 64.050 ;
        RECT 758.400 58.050 759.600 64.950 ;
        RECT 763.950 59.100 766.050 61.200 ;
        RECT 767.400 60.600 768.600 97.800 ;
        RECT 773.400 76.050 774.600 100.950 ;
        RECT 782.400 94.050 783.600 100.950 ;
        RECT 788.400 99.900 789.600 100.950 ;
        RECT 787.950 97.800 790.050 99.900 ;
        RECT 806.400 99.000 807.600 100.950 ;
        RECT 781.950 91.950 784.050 94.050 ;
        RECT 788.400 91.050 789.600 97.800 ;
        RECT 805.950 94.950 808.050 99.000 ;
        RECT 787.950 88.950 790.050 91.050 ;
        RECT 812.400 76.050 813.600 100.950 ;
        RECT 818.400 88.050 819.600 100.950 ;
        RECT 817.950 85.950 820.050 88.050 ;
        RECT 824.400 85.050 825.600 148.950 ;
        RECT 827.400 121.050 828.600 166.950 ;
        RECT 838.950 163.950 841.050 166.050 ;
        RECT 832.950 138.000 835.050 142.050 ;
        RECT 833.400 136.050 834.600 138.000 ;
        RECT 839.400 136.050 840.600 163.950 ;
        RECT 854.400 147.600 855.600 173.400 ;
        RECT 859.950 172.950 862.050 175.050 ;
        RECT 856.950 169.950 859.050 172.050 ;
        RECT 863.850 171.600 865.050 188.400 ;
        RECT 857.400 151.050 858.600 169.950 ;
        RECT 862.950 169.500 865.050 171.600 ;
        RECT 863.850 164.700 865.050 169.500 ;
        RECT 865.950 188.400 868.050 190.500 ;
        RECT 868.950 188.400 871.050 190.500 ;
        RECT 871.950 188.400 874.050 190.500 ;
        RECT 877.950 188.400 880.050 190.500 ;
        RECT 886.950 188.400 889.050 190.500 ;
        RECT 889.950 188.400 892.050 190.500 ;
        RECT 892.950 188.400 895.050 190.500 ;
        RECT 865.950 167.700 867.150 188.400 ;
        RECT 868.950 171.600 870.450 188.400 ;
        RECT 872.850 176.700 874.050 188.400 ;
        RECT 878.250 176.700 879.450 188.400 ;
        RECT 880.950 181.950 883.050 184.050 ;
        RECT 881.400 180.900 882.600 181.950 ;
        RECT 880.950 178.800 883.050 180.900 ;
        RECT 871.950 174.600 874.050 176.700 ;
        RECT 877.950 174.600 880.050 176.700 ;
        RECT 868.950 169.500 871.050 171.600 ;
        RECT 862.950 162.600 865.050 164.700 ;
        RECT 866.100 164.700 867.150 167.700 ;
        RECT 869.100 164.700 870.300 169.500 ;
        RECT 872.850 167.700 874.050 174.600 ;
        RECT 878.850 169.200 880.050 174.600 ;
        RECT 871.950 165.600 874.050 167.700 ;
        RECT 877.950 167.100 880.050 169.200 ;
        RECT 886.950 167.400 888.150 188.400 ;
        RECT 889.950 172.800 891.150 188.400 ;
        RECT 889.950 170.700 892.050 172.800 ;
        RECT 890.400 167.400 891.600 170.700 ;
        RECT 893.400 167.400 894.600 188.400 ;
        RECT 899.400 184.050 900.600 202.950 ;
        RECT 901.950 199.950 904.050 202.050 ;
        RECT 898.950 181.950 901.050 184.050 ;
        RECT 902.400 181.050 903.600 199.950 ;
        RECT 908.400 184.050 909.600 208.950 ;
        RECT 907.950 181.950 910.050 184.050 ;
        RECT 911.400 181.050 912.600 217.950 ;
        RECT 914.400 195.600 915.600 352.950 ;
        RECT 917.400 351.600 918.600 436.950 ;
        RECT 919.950 427.950 922.050 430.050 ;
        RECT 920.400 391.050 921.600 427.950 ;
        RECT 919.950 388.950 922.050 391.050 ;
        RECT 919.950 379.950 922.050 382.050 ;
        RECT 920.400 355.050 921.600 379.950 ;
        RECT 919.950 352.950 922.050 355.050 ;
        RECT 917.400 350.400 921.600 351.600 ;
        RECT 916.950 346.950 919.050 349.050 ;
        RECT 917.400 211.050 918.600 346.950 ;
        RECT 916.950 208.950 919.050 211.050 ;
        RECT 914.400 194.400 918.600 195.600 ;
        RECT 913.950 190.950 916.050 193.050 ;
        RECT 901.950 178.950 904.050 181.050 ;
        RECT 910.950 178.950 913.050 181.050 ;
        RECT 904.950 175.950 907.050 178.050 ;
        RECT 914.400 177.600 915.600 190.950 ;
        RECT 911.400 176.400 915.600 177.600 ;
        RECT 905.400 174.600 906.600 175.950 ;
        RECT 911.400 174.600 912.600 176.400 ;
        RECT 905.400 173.400 912.600 174.600 ;
        RECT 913.950 172.950 916.050 175.050 ;
        RECT 910.950 169.950 913.050 172.050 ;
        RECT 886.950 165.300 889.050 167.400 ;
        RECT 889.950 165.300 892.050 167.400 ;
        RECT 892.950 165.300 895.050 167.400 ;
        RECT 907.950 166.950 910.050 169.050 ;
        RECT 866.100 162.600 868.200 164.700 ;
        RECT 869.100 162.600 871.200 164.700 ;
        RECT 889.950 160.950 892.050 163.050 ;
        RECT 856.950 148.950 859.050 151.050 ;
        RECT 871.950 148.950 874.050 151.050 ;
        RECT 854.400 147.000 858.600 147.600 ;
        RECT 854.400 146.400 859.050 147.000 ;
        RECT 854.400 142.200 855.600 146.400 ;
        RECT 856.950 142.950 859.050 146.400 ;
        RECT 847.950 139.950 850.050 142.050 ;
        RECT 853.950 140.100 856.050 142.200 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 826.950 118.950 829.050 121.050 ;
        RECT 836.400 112.050 837.600 133.950 ;
        RECT 842.400 132.000 843.600 133.950 ;
        RECT 841.950 127.950 844.050 132.000 ;
        RECT 844.950 114.600 847.050 115.050 ;
        RECT 839.400 113.400 847.050 114.600 ;
        RECT 832.800 109.950 834.900 112.050 ;
        RECT 835.950 109.950 838.050 112.050 ;
        RECT 833.400 103.050 834.600 109.950 ;
        RECT 839.400 103.050 840.600 113.400 ;
        RECT 844.950 112.950 847.050 113.400 ;
        RECT 841.950 109.950 844.050 112.050 ;
        RECT 848.400 111.600 849.600 139.950 ;
        RECT 859.950 133.950 862.050 136.050 ;
        RECT 860.400 132.000 861.600 133.950 ;
        RECT 859.950 127.950 862.050 132.000 ;
        RECT 856.950 112.950 859.050 115.050 ;
        RECT 845.400 110.400 849.600 111.600 ;
        RECT 842.400 106.050 843.600 109.950 ;
        RECT 841.950 103.950 844.050 106.050 ;
        RECT 829.950 100.950 832.050 103.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 830.400 99.900 831.600 100.950 ;
        RECT 829.950 97.800 832.050 99.900 ;
        RECT 836.400 91.050 837.600 100.950 ;
        RECT 835.950 88.950 838.050 91.050 ;
        RECT 823.950 82.950 826.050 85.050 ;
        RECT 772.950 73.950 775.050 76.050 ;
        RECT 805.950 73.950 808.050 76.050 ;
        RECT 811.950 73.950 814.050 76.050 ;
        RECT 845.400 75.600 846.600 110.400 ;
        RECT 847.950 106.950 850.050 109.050 ;
        RECT 848.400 91.050 849.600 106.950 ;
        RECT 857.400 103.050 858.600 112.950 ;
        RECT 862.950 105.000 865.050 109.050 ;
        RECT 863.400 103.050 864.600 105.000 ;
        RECT 853.950 100.950 856.050 103.050 ;
        RECT 856.950 100.950 859.050 103.050 ;
        RECT 859.950 100.950 862.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 865.950 100.950 868.050 103.050 ;
        RECT 850.950 97.950 853.050 100.050 ;
        RECT 847.950 88.950 850.050 91.050 ;
        RECT 842.400 74.400 846.600 75.600 ;
        RECT 851.400 75.600 852.600 97.950 ;
        RECT 854.400 82.050 855.600 100.950 ;
        RECT 856.950 82.950 859.050 85.050 ;
        RECT 853.950 79.950 856.050 82.050 ;
        RECT 851.400 74.400 855.600 75.600 ;
        RECT 790.950 69.300 793.050 71.400 ;
        RECT 772.950 64.950 775.050 67.050 ;
        RECT 791.850 65.700 793.050 69.300 ;
        RECT 767.400 59.400 771.600 60.600 ;
        RECT 764.400 58.050 765.600 59.100 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 755.400 54.900 756.600 55.950 ;
        RECT 754.950 52.800 757.050 54.900 ;
        RECT 761.400 54.000 762.600 55.950 ;
        RECT 760.950 49.950 763.050 54.000 ;
        RECT 770.400 52.050 771.600 59.400 ;
        RECT 769.950 49.950 772.050 52.050 ;
        RECT 773.400 40.050 774.600 64.950 ;
        RECT 790.950 63.600 793.050 65.700 ;
        RECT 778.950 59.100 781.050 61.200 ;
        RECT 779.400 58.050 780.600 59.100 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 787.950 55.950 790.050 58.050 ;
        RECT 751.950 37.950 754.050 40.050 ;
        RECT 772.950 37.950 775.050 40.050 ;
        RECT 778.950 37.950 781.050 40.050 ;
        RECT 718.950 19.500 721.050 21.600 ;
        RECT 724.800 19.500 726.900 21.600 ;
        RECT 727.950 19.500 730.050 21.600 ;
        RECT 733.950 17.400 735.150 32.400 ;
        RECT 742.950 31.950 745.050 34.050 ;
        RECT 736.950 26.400 739.050 28.500 ;
        RECT 752.400 28.200 753.600 37.950 ;
        RECT 769.950 32.400 772.050 34.500 ;
        RECT 737.400 25.050 738.600 26.400 ;
        RECT 751.950 26.100 754.050 28.200 ;
        RECT 752.400 25.050 753.600 26.100 ;
        RECT 736.950 22.950 739.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 767.400 21.600 768.600 22.950 ;
        RECT 766.950 19.500 769.050 21.600 ;
        RECT 733.950 15.300 736.050 17.400 ;
        RECT 712.950 10.500 715.050 12.600 ;
        RECT 733.950 11.700 735.150 15.300 ;
        RECT 770.700 12.600 771.900 32.400 ;
        RECT 779.400 27.600 780.600 37.950 ;
        RECT 782.400 34.050 783.600 55.950 ;
        RECT 788.400 54.600 789.600 55.950 ;
        RECT 787.950 52.500 790.050 54.600 ;
        RECT 791.850 48.600 793.050 63.600 ;
        RECT 806.400 58.050 807.600 73.950 ;
        RECT 838.950 70.950 841.050 73.050 ;
        RECT 811.950 68.400 814.050 70.500 ;
        RECT 826.950 68.400 829.050 70.500 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 812.100 48.600 813.300 68.400 ;
        RECT 814.950 60.000 817.050 64.050 ;
        RECT 823.950 60.000 826.050 64.050 ;
        RECT 815.400 58.050 816.600 60.000 ;
        RECT 824.400 58.050 825.600 60.000 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 827.700 48.600 828.900 68.400 ;
        RECT 832.950 67.950 835.050 70.050 ;
        RECT 833.400 58.050 834.600 67.950 ;
        RECT 839.400 58.050 840.600 70.950 ;
        RECT 842.400 64.050 843.600 74.400 ;
        RECT 847.950 69.300 850.050 71.400 ;
        RECT 847.950 65.700 849.150 69.300 ;
        RECT 841.950 61.950 844.050 64.050 ;
        RECT 847.950 63.600 850.050 65.700 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 838.950 55.950 841.050 58.050 ;
        RECT 790.950 46.500 793.050 48.600 ;
        RECT 811.950 46.500 814.050 48.600 ;
        RECT 826.950 46.500 829.050 48.600 ;
        RECT 781.950 31.950 784.050 34.050 ;
        RECT 790.950 32.400 793.050 34.500 ;
        RECT 779.400 26.400 783.600 27.600 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 776.400 21.600 777.600 22.950 ;
        RECT 782.400 21.600 783.600 26.400 ;
        RECT 775.950 19.500 778.050 21.600 ;
        RECT 781.950 19.500 784.050 21.600 ;
        RECT 790.950 17.400 792.150 32.400 ;
        RECT 805.950 31.950 808.050 34.050 ;
        RECT 793.950 26.400 796.050 28.500 ;
        RECT 806.400 28.200 807.600 31.950 ;
        RECT 839.400 28.200 840.600 55.950 ;
        RECT 847.950 48.600 849.150 63.600 ;
        RECT 854.400 61.050 855.600 74.400 ;
        RECT 853.950 58.950 856.050 61.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 851.400 54.600 852.600 55.950 ;
        RECT 850.950 53.400 855.600 54.600 ;
        RECT 850.950 52.500 853.050 53.400 ;
        RECT 847.950 46.500 850.050 48.600 ;
        RECT 794.400 25.050 795.600 26.400 ;
        RECT 805.950 26.100 808.050 28.200 ;
        RECT 826.950 26.100 829.050 28.200 ;
        RECT 838.950 26.100 841.050 28.200 ;
        RECT 854.400 27.600 855.600 53.400 ;
        RECT 857.400 46.050 858.600 82.950 ;
        RECT 860.400 70.050 861.600 100.950 ;
        RECT 866.400 99.000 867.600 100.950 ;
        RECT 865.950 94.950 868.050 99.000 ;
        RECT 868.950 97.950 871.050 100.050 ;
        RECT 865.950 78.600 868.050 82.050 ;
        RECT 863.400 78.000 868.050 78.600 ;
        RECT 863.400 77.400 867.600 78.000 ;
        RECT 859.950 67.950 862.050 70.050 ;
        RECT 863.400 58.050 864.600 77.400 ;
        RECT 865.950 73.950 868.050 76.050 ;
        RECT 866.400 63.600 867.600 73.950 ;
        RECT 869.400 73.050 870.600 97.950 ;
        RECT 868.950 70.950 871.050 73.050 ;
        RECT 872.400 64.050 873.600 148.950 ;
        RECT 877.950 142.950 880.050 145.050 ;
        RECT 878.400 136.050 879.600 142.950 ;
        RECT 877.950 133.950 880.050 136.050 ;
        RECT 886.950 118.950 889.050 121.050 ;
        RECT 874.950 105.600 879.000 106.050 ;
        RECT 874.950 103.950 879.600 105.600 ;
        RECT 878.400 103.050 879.600 103.950 ;
        RECT 877.950 100.950 880.050 103.050 ;
        RECT 880.950 100.950 883.050 103.050 ;
        RECT 881.400 88.050 882.600 100.950 ;
        RECT 880.950 85.950 883.050 88.050 ;
        RECT 887.400 64.050 888.600 118.950 ;
        RECT 890.400 82.050 891.600 160.950 ;
        RECT 904.950 154.950 907.050 157.050 ;
        RECT 895.950 104.100 898.050 106.200 ;
        RECT 896.400 103.050 897.600 104.100 ;
        RECT 895.950 100.950 898.050 103.050 ;
        RECT 898.950 100.950 901.050 103.050 ;
        RECT 899.400 99.000 900.600 100.950 ;
        RECT 898.950 94.950 901.050 99.000 ;
        RECT 889.950 79.950 892.050 82.050 ;
        RECT 901.950 73.950 904.050 76.050 ;
        RECT 889.950 64.950 892.050 67.050 ;
        RECT 866.400 62.400 870.600 63.600 ;
        RECT 869.400 58.050 870.600 62.400 ;
        RECT 871.950 61.950 874.050 64.050 ;
        RECT 877.950 61.950 880.050 64.050 ;
        RECT 880.950 61.950 883.050 64.050 ;
        RECT 886.950 61.950 889.050 64.050 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 865.950 55.950 868.050 58.050 ;
        RECT 868.950 55.950 871.050 58.050 ;
        RECT 871.950 55.950 874.050 58.050 ;
        RECT 866.400 54.900 867.600 55.950 ;
        RECT 865.950 52.800 868.050 54.900 ;
        RECT 872.400 46.050 873.600 55.950 ;
        RECT 856.950 43.950 859.050 46.050 ;
        RECT 865.950 43.950 868.050 46.050 ;
        RECT 871.950 43.950 874.050 46.050 ;
        RECT 854.400 26.400 858.600 27.600 ;
        RECT 806.400 25.050 807.600 26.100 ;
        RECT 827.400 25.050 828.600 26.100 ;
        RECT 857.400 25.050 858.600 26.400 ;
        RECT 866.400 25.050 867.600 43.950 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 856.950 22.950 859.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 878.400 21.900 879.600 61.950 ;
        RECT 881.400 54.900 882.600 61.950 ;
        RECT 890.400 58.050 891.600 64.950 ;
        RECT 895.950 59.100 898.050 61.200 ;
        RECT 896.400 58.050 897.600 59.100 ;
        RECT 886.950 55.950 889.050 58.050 ;
        RECT 889.950 55.950 892.050 58.050 ;
        RECT 892.950 55.950 895.050 58.050 ;
        RECT 895.950 55.950 898.050 58.050 ;
        RECT 887.400 54.900 888.600 55.950 ;
        RECT 880.950 52.800 883.050 54.900 ;
        RECT 886.950 52.800 889.050 54.900 ;
        RECT 893.400 51.600 894.600 55.950 ;
        RECT 893.400 50.400 897.600 51.600 ;
        RECT 892.950 46.950 895.050 49.050 ;
        RECT 893.400 25.050 894.600 46.950 ;
        RECT 896.400 43.050 897.600 50.400 ;
        RECT 902.400 49.050 903.600 73.950 ;
        RECT 905.400 54.900 906.600 154.950 ;
        RECT 904.950 52.800 907.050 54.900 ;
        RECT 901.950 46.950 904.050 49.050 ;
        RECT 908.400 43.050 909.600 166.950 ;
        RECT 911.400 67.050 912.600 169.950 ;
        RECT 910.950 64.950 913.050 67.050 ;
        RECT 895.950 40.950 898.050 43.050 ;
        RECT 907.950 40.950 910.050 43.050 ;
        RECT 889.950 22.950 892.050 25.050 ;
        RECT 892.950 22.950 895.050 25.050 ;
        RECT 895.950 22.950 898.050 25.050 ;
        RECT 890.400 21.900 891.600 22.950 ;
        RECT 877.950 19.800 880.050 21.900 ;
        RECT 889.950 19.800 892.050 21.900 ;
        RECT 896.400 21.000 897.600 22.950 ;
        RECT 790.950 15.300 793.050 17.400 ;
        RECT 895.950 16.950 898.050 21.000 ;
        RECT 911.400 19.050 912.600 64.950 ;
        RECT 914.400 61.200 915.600 172.950 ;
        RECT 917.400 76.050 918.600 194.400 ;
        RECT 920.400 169.050 921.600 350.400 ;
        RECT 919.950 166.950 922.050 169.050 ;
        RECT 919.950 160.950 922.050 163.050 ;
        RECT 916.950 73.950 919.050 76.050 ;
        RECT 913.950 59.100 916.050 61.200 ;
        RECT 920.400 46.050 921.600 160.950 ;
        RECT 919.950 43.950 922.050 46.050 ;
        RECT 910.950 16.950 913.050 19.050 ;
        RECT 601.950 7.950 604.050 10.050 ;
        RECT 733.950 9.600 736.050 11.700 ;
        RECT 769.950 10.500 772.050 12.600 ;
        RECT 790.950 11.700 792.150 15.300 ;
        RECT 790.950 9.600 793.050 11.700 ;
        RECT 112.950 4.950 115.050 7.050 ;
        RECT 199.950 4.950 202.050 7.050 ;
        RECT 319.950 4.950 322.050 7.050 ;
        RECT 415.950 4.950 421.050 7.050 ;
        RECT 424.950 4.950 430.050 7.050 ;
        RECT 508.950 4.950 511.050 7.050 ;
        RECT 517.950 4.950 520.050 7.050 ;
        RECT 562.950 4.950 565.050 7.050 ;
      LAYER metal3 ;
        RECT 664.950 936.600 667.050 937.050 ;
        RECT 847.950 936.600 850.050 937.050 ;
        RECT 664.950 935.400 744.600 936.600 ;
        RECT 664.950 934.950 667.050 935.400 ;
        RECT 43.950 933.600 46.050 934.050 ;
        RECT 97.950 933.600 100.050 934.050 ;
        RECT 136.950 933.600 139.050 934.050 ;
        RECT 43.950 932.400 139.050 933.600 ;
        RECT 43.950 931.950 46.050 932.400 ;
        RECT 97.950 931.950 100.050 932.400 ;
        RECT 136.950 931.950 139.050 932.400 ;
        RECT 652.950 933.600 655.050 934.050 ;
        RECT 739.950 933.600 742.050 934.050 ;
        RECT 652.950 932.400 742.050 933.600 ;
        RECT 743.400 933.600 744.600 935.400 ;
        RECT 770.400 935.400 850.050 936.600 ;
        RECT 770.400 933.600 771.600 935.400 ;
        RECT 847.950 934.950 850.050 935.400 ;
        RECT 743.400 932.400 771.600 933.600 ;
        RECT 652.950 931.950 655.050 932.400 ;
        RECT 739.950 931.950 742.050 932.400 ;
        RECT 112.950 930.600 115.050 931.050 ;
        RECT 214.950 930.600 217.050 931.050 ;
        RECT 298.950 930.600 301.050 931.050 ;
        RECT 310.950 930.600 313.050 931.050 ;
        RECT 112.950 929.400 313.050 930.600 ;
        RECT 112.950 928.950 115.050 929.400 ;
        RECT 214.950 928.950 217.050 929.400 ;
        RECT 298.950 928.950 301.050 929.400 ;
        RECT 310.950 928.950 313.050 929.400 ;
        RECT 334.950 930.600 337.050 931.050 ;
        RECT 334.950 929.400 357.600 930.600 ;
        RECT 334.950 928.950 337.050 929.400 ;
        RECT 356.400 928.050 357.600 929.400 ;
        RECT 76.950 927.600 79.050 928.050 ;
        RECT 109.950 927.600 112.050 928.050 ;
        RECT 76.950 926.400 112.050 927.600 ;
        RECT 76.950 925.950 79.050 926.400 ;
        RECT 109.950 925.950 112.050 926.400 ;
        RECT 304.950 927.600 307.050 928.050 ;
        RECT 337.950 927.600 340.050 928.050 ;
        RECT 304.950 926.400 340.050 927.600 ;
        RECT 304.950 925.950 307.050 926.400 ;
        RECT 337.950 925.950 340.050 926.400 ;
        RECT 355.950 927.600 358.050 928.050 ;
        RECT 370.950 927.600 373.050 928.050 ;
        RECT 355.950 926.400 373.050 927.600 ;
        RECT 355.950 925.950 358.050 926.400 ;
        RECT 370.950 925.950 373.050 926.400 ;
        RECT 463.950 927.600 466.050 928.050 ;
        RECT 505.950 927.600 508.050 928.050 ;
        RECT 463.950 926.400 508.050 927.600 ;
        RECT 463.950 925.950 466.050 926.400 ;
        RECT 505.950 925.950 508.050 926.400 ;
        RECT 841.950 927.600 844.050 928.050 ;
        RECT 874.950 927.600 877.050 928.050 ;
        RECT 841.950 926.400 877.050 927.600 ;
        RECT 841.950 925.950 844.050 926.400 ;
        RECT 874.950 925.950 877.050 926.400 ;
        RECT 13.950 924.600 16.050 925.050 ;
        RECT 37.950 924.600 40.050 925.050 ;
        RECT 58.950 924.600 61.050 925.050 ;
        RECT 13.950 923.400 61.050 924.600 ;
        RECT 13.950 922.950 16.050 923.400 ;
        RECT 37.950 922.950 40.050 923.400 ;
        RECT 58.950 922.950 61.050 923.400 ;
        RECT 130.950 924.600 133.050 925.050 ;
        RECT 163.950 924.600 166.050 925.050 ;
        RECT 130.950 923.400 166.050 924.600 ;
        RECT 130.950 922.950 133.050 923.400 ;
        RECT 163.950 922.950 166.050 923.400 ;
        RECT 178.950 924.600 181.050 925.050 ;
        RECT 205.950 924.600 208.050 925.050 ;
        RECT 178.950 923.400 208.050 924.600 ;
        RECT 178.950 922.950 181.050 923.400 ;
        RECT 205.950 922.950 208.050 923.400 ;
        RECT 247.950 924.600 250.050 925.050 ;
        RECT 265.950 924.600 268.050 925.050 ;
        RECT 280.950 924.600 283.050 925.050 ;
        RECT 247.950 923.400 283.050 924.600 ;
        RECT 247.950 922.950 250.050 923.400 ;
        RECT 265.950 922.950 268.050 923.400 ;
        RECT 280.950 922.950 283.050 923.400 ;
        RECT 415.950 924.600 418.050 925.050 ;
        RECT 427.950 924.600 430.050 925.050 ;
        RECT 415.950 923.400 430.050 924.600 ;
        RECT 415.950 922.950 418.050 923.400 ;
        RECT 427.950 922.950 430.050 923.400 ;
        RECT 556.950 924.600 559.050 925.050 ;
        RECT 571.950 924.600 574.050 925.050 ;
        RECT 556.950 923.400 574.050 924.600 ;
        RECT 556.950 922.950 559.050 923.400 ;
        RECT 571.950 922.950 574.050 923.400 ;
        RECT 583.950 924.600 586.050 925.050 ;
        RECT 601.950 924.600 604.050 925.050 ;
        RECT 583.950 923.400 604.050 924.600 ;
        RECT 583.950 922.950 586.050 923.400 ;
        RECT 601.950 922.950 604.050 923.400 ;
        RECT 643.950 924.600 646.050 925.050 ;
        RECT 658.950 924.600 661.050 925.050 ;
        RECT 718.950 924.600 721.050 925.050 ;
        RECT 745.950 924.600 748.050 925.050 ;
        RECT 643.950 923.400 748.050 924.600 ;
        RECT 643.950 922.950 646.050 923.400 ;
        RECT 658.950 922.950 661.050 923.400 ;
        RECT 718.950 922.950 721.050 923.400 ;
        RECT 745.950 922.950 748.050 923.400 ;
        RECT 790.950 924.600 793.050 925.050 ;
        RECT 838.950 924.600 841.050 925.050 ;
        RECT 790.950 923.400 841.050 924.600 ;
        RECT 790.950 922.950 793.050 923.400 ;
        RECT 838.950 922.950 841.050 923.400 ;
        RECT 88.950 921.600 91.050 922.050 ;
        RECT 112.950 921.600 115.050 922.050 ;
        RECT 88.950 920.400 115.050 921.600 ;
        RECT 88.950 919.950 91.050 920.400 ;
        RECT 112.950 919.950 115.050 920.400 ;
        RECT 118.950 921.600 121.050 922.050 ;
        RECT 127.950 921.600 130.050 922.050 ;
        RECT 118.950 920.400 130.050 921.600 ;
        RECT 118.950 919.950 121.050 920.400 ;
        RECT 127.950 919.950 130.050 920.400 ;
        RECT 493.950 921.600 496.050 922.050 ;
        RECT 499.950 921.600 502.050 922.050 ;
        RECT 493.950 920.400 502.050 921.600 ;
        RECT 493.950 919.950 496.050 920.400 ;
        RECT 499.950 919.950 502.050 920.400 ;
        RECT 751.950 921.600 754.050 922.050 ;
        RECT 781.950 921.600 784.050 922.050 ;
        RECT 751.950 920.400 784.050 921.600 ;
        RECT 751.950 919.950 754.050 920.400 ;
        RECT 781.950 919.950 784.050 920.400 ;
        RECT 814.950 921.600 817.050 922.050 ;
        RECT 820.950 921.600 823.050 922.050 ;
        RECT 814.950 920.400 823.050 921.600 ;
        RECT 814.950 919.950 817.050 920.400 ;
        RECT 820.950 919.950 823.050 920.400 ;
        RECT 826.950 921.600 829.050 922.050 ;
        RECT 832.950 921.600 835.050 922.050 ;
        RECT 826.950 920.400 835.050 921.600 ;
        RECT 826.950 919.950 829.050 920.400 ;
        RECT 832.950 919.950 835.050 920.400 ;
        RECT 25.950 918.750 28.050 919.200 ;
        RECT 31.950 918.750 34.050 919.200 ;
        RECT 25.950 917.550 34.050 918.750 ;
        RECT 43.800 918.600 45.900 919.050 ;
        RECT 25.950 917.100 28.050 917.550 ;
        RECT 31.950 917.100 34.050 917.550 ;
        RECT 38.400 917.400 45.900 918.600 ;
        RECT 38.400 915.600 39.600 917.400 ;
        RECT 43.800 916.950 45.900 917.400 ;
        RECT 46.950 918.750 49.050 919.200 ;
        RECT 52.950 918.750 55.050 919.200 ;
        RECT 46.950 917.550 55.050 918.750 ;
        RECT 46.950 917.100 49.050 917.550 ;
        RECT 52.950 917.100 55.050 917.550 ;
        RECT 76.950 918.600 79.050 919.200 ;
        RECT 76.950 917.400 96.600 918.600 ;
        RECT 76.950 917.100 79.050 917.400 ;
        RECT 35.400 914.400 39.600 915.600 ;
        RECT 95.400 915.600 96.600 917.400 ;
        RECT 103.950 917.100 106.050 919.200 ;
        RECT 142.950 918.750 145.050 919.200 ;
        RECT 151.950 918.750 154.050 919.200 ;
        RECT 142.950 917.550 154.050 918.750 ;
        RECT 142.950 917.100 145.050 917.550 ;
        RECT 151.950 917.100 154.050 917.550 ;
        RECT 169.950 918.600 172.050 919.200 ;
        RECT 184.950 918.600 187.050 919.200 ;
        RECT 169.950 917.400 187.050 918.600 ;
        RECT 169.950 917.100 172.050 917.400 ;
        RECT 184.950 917.100 187.050 917.400 ;
        RECT 199.950 917.100 202.050 919.200 ;
        RECT 220.950 918.600 223.050 919.200 ;
        RECT 212.400 917.400 223.050 918.600 ;
        RECT 95.400 914.400 102.600 915.600 ;
        RECT 35.400 912.900 36.600 914.400 ;
        RECT 34.950 910.800 37.050 912.900 ;
        RECT 40.950 912.600 43.050 912.900 ;
        RECT 46.950 912.600 49.050 913.050 ;
        RECT 40.950 911.400 49.050 912.600 ;
        RECT 40.950 910.800 43.050 911.400 ;
        RECT 46.950 910.950 49.050 911.400 ;
        RECT 61.950 912.450 64.050 912.900 ;
        RECT 70.950 912.450 73.050 912.900 ;
        RECT 61.950 911.250 73.050 912.450 ;
        RECT 61.950 910.800 64.050 911.250 ;
        RECT 70.950 910.800 73.050 911.250 ;
        RECT 88.950 912.600 91.050 913.050 ;
        RECT 101.400 912.900 102.600 914.400 ;
        RECT 94.950 912.600 97.050 912.900 ;
        RECT 88.950 911.400 97.050 912.600 ;
        RECT 88.950 910.950 91.050 911.400 ;
        RECT 94.950 910.800 97.050 911.400 ;
        RECT 100.950 910.800 103.050 912.900 ;
        RECT 104.400 912.600 105.600 917.100 ;
        RECT 130.950 915.600 133.050 916.050 ;
        RECT 125.400 914.400 133.050 915.600 ;
        RECT 115.950 912.600 118.050 912.900 ;
        RECT 104.400 911.400 118.050 912.600 ;
        RECT 115.950 910.800 118.050 911.400 ;
        RECT 121.950 912.600 124.050 912.900 ;
        RECT 125.400 912.600 126.600 914.400 ;
        RECT 130.950 913.950 133.050 914.400 ;
        RECT 121.950 911.400 126.600 912.600 ;
        RECT 139.950 912.600 142.050 912.900 ;
        RECT 166.950 912.600 169.050 912.900 ;
        RECT 200.400 912.600 201.600 917.100 ;
        RECT 139.950 911.400 169.050 912.600 ;
        RECT 121.950 910.800 124.050 911.400 ;
        RECT 139.950 910.800 142.050 911.400 ;
        RECT 166.950 910.800 169.050 911.400 ;
        RECT 185.400 911.400 201.600 912.600 ;
        RECT 127.950 909.600 130.050 910.050 ;
        RECT 185.400 909.600 186.600 911.400 ;
        RECT 127.950 908.400 186.600 909.600 ;
        RECT 187.950 909.600 190.050 910.050 ;
        RECT 199.950 909.600 202.050 910.050 ;
        RECT 212.400 909.600 213.600 917.400 ;
        RECT 220.950 917.100 223.050 917.400 ;
        RECT 226.950 918.750 229.050 919.200 ;
        RECT 235.950 918.750 238.050 919.200 ;
        RECT 226.950 917.550 238.050 918.750 ;
        RECT 226.950 917.100 229.050 917.550 ;
        RECT 235.950 917.100 238.050 917.550 ;
        RECT 259.950 918.750 262.050 919.200 ;
        RECT 271.950 918.750 274.050 919.200 ;
        RECT 259.950 917.550 274.050 918.750 ;
        RECT 259.950 917.100 262.050 917.550 ;
        RECT 271.950 917.100 274.050 917.550 ;
        RECT 286.950 918.750 289.050 919.200 ;
        RECT 292.950 918.750 295.050 919.200 ;
        RECT 286.950 917.550 295.050 918.750 ;
        RECT 286.950 917.100 289.050 917.550 ;
        RECT 292.950 917.100 295.050 917.550 ;
        RECT 316.950 918.750 319.050 919.200 ;
        RECT 325.950 918.750 328.050 919.200 ;
        RECT 316.950 917.550 328.050 918.750 ;
        RECT 316.950 917.100 319.050 917.550 ;
        RECT 325.950 917.100 328.050 917.550 ;
        RECT 340.950 916.950 343.050 919.050 ;
        RECT 367.950 918.750 370.050 919.200 ;
        RECT 385.950 918.750 388.050 919.200 ;
        RECT 367.950 917.550 388.050 918.750 ;
        RECT 367.950 917.100 370.050 917.550 ;
        RECT 385.950 917.100 388.050 917.550 ;
        RECT 409.950 918.750 412.050 919.200 ;
        RECT 415.950 918.750 418.050 919.200 ;
        RECT 409.950 917.550 418.050 918.750 ;
        RECT 409.950 917.100 412.050 917.550 ;
        RECT 415.950 917.100 418.050 917.550 ;
        RECT 421.950 917.100 424.050 919.200 ;
        RECT 442.950 918.600 445.050 919.200 ;
        RECT 454.950 918.600 457.050 919.050 ;
        RECT 442.950 917.400 457.050 918.600 ;
        RECT 442.950 917.100 445.050 917.400 ;
        RECT 214.950 912.450 217.050 912.900 ;
        RECT 223.950 912.450 226.050 912.900 ;
        RECT 214.950 911.250 226.050 912.450 ;
        RECT 214.950 910.800 217.050 911.250 ;
        RECT 223.950 910.800 226.050 911.250 ;
        RECT 250.950 912.450 253.050 912.900 ;
        RECT 256.950 912.600 259.050 912.900 ;
        RECT 268.950 912.600 271.050 912.900 ;
        RECT 256.950 912.450 271.050 912.600 ;
        RECT 250.950 911.400 271.050 912.450 ;
        RECT 250.950 911.250 259.050 911.400 ;
        RECT 250.950 910.800 253.050 911.250 ;
        RECT 256.950 910.800 259.050 911.250 ;
        RECT 268.950 910.800 271.050 911.400 ;
        RECT 286.950 912.450 289.050 912.900 ;
        RECT 313.950 912.450 316.050 912.900 ;
        RECT 286.950 911.250 316.050 912.450 ;
        RECT 286.950 910.800 289.050 911.250 ;
        RECT 313.950 910.800 316.050 911.250 ;
        RECT 325.950 912.600 328.050 913.050 ;
        RECT 337.950 912.600 340.050 912.900 ;
        RECT 325.950 911.400 340.050 912.600 ;
        RECT 341.400 912.600 342.600 916.950 ;
        RECT 352.950 912.600 355.050 912.900 ;
        RECT 376.950 912.600 379.050 912.900 ;
        RECT 341.400 911.400 379.050 912.600 ;
        RECT 325.950 910.950 328.050 911.400 ;
        RECT 337.950 910.800 340.050 911.400 ;
        RECT 352.950 910.800 355.050 911.400 ;
        RECT 376.950 910.800 379.050 911.400 ;
        RECT 406.950 912.600 409.050 912.900 ;
        RECT 422.400 912.600 423.600 917.100 ;
        RECT 454.950 916.950 457.050 917.400 ;
        RECT 517.950 918.750 520.050 919.200 ;
        RECT 523.950 918.750 526.050 919.200 ;
        RECT 517.950 917.550 526.050 918.750 ;
        RECT 517.950 917.100 520.050 917.550 ;
        RECT 523.950 917.100 526.050 917.550 ;
        RECT 535.950 918.750 538.050 919.200 ;
        RECT 541.950 918.750 544.050 919.200 ;
        RECT 535.950 917.550 544.050 918.750 ;
        RECT 535.950 917.100 538.050 917.550 ;
        RECT 541.950 917.100 544.050 917.550 ;
        RECT 547.950 918.600 550.050 919.200 ;
        RECT 565.950 918.750 568.050 919.200 ;
        RECT 583.800 918.750 585.900 919.200 ;
        RECT 565.950 918.600 585.900 918.750 ;
        RECT 547.950 917.550 585.900 918.600 ;
        RECT 547.950 917.400 568.050 917.550 ;
        RECT 547.950 917.100 550.050 917.400 ;
        RECT 565.950 917.100 568.050 917.400 ;
        RECT 583.800 917.100 585.900 917.550 ;
        RECT 586.950 918.750 589.050 919.200 ;
        RECT 592.950 918.750 595.050 919.200 ;
        RECT 586.950 917.550 595.050 918.750 ;
        RECT 586.950 917.100 589.050 917.550 ;
        RECT 592.950 917.100 595.050 917.550 ;
        RECT 598.950 918.750 601.050 919.200 ;
        RECT 604.950 918.750 607.050 919.200 ;
        RECT 598.950 917.550 607.050 918.750 ;
        RECT 598.950 917.100 601.050 917.550 ;
        RECT 604.950 917.100 607.050 917.550 ;
        RECT 613.950 918.600 616.050 919.200 ;
        RECT 619.800 918.600 621.900 919.050 ;
        RECT 613.950 917.400 621.900 918.600 ;
        RECT 613.950 917.100 616.050 917.400 ;
        RECT 619.800 916.950 621.900 917.400 ;
        RECT 622.950 918.750 625.050 919.200 ;
        RECT 628.950 918.750 631.050 919.200 ;
        RECT 622.950 917.550 631.050 918.750 ;
        RECT 622.950 917.100 625.050 917.550 ;
        RECT 628.950 917.100 631.050 917.550 ;
        RECT 634.950 918.600 637.050 919.200 ;
        RECT 652.950 918.600 655.050 919.200 ;
        RECT 634.950 917.400 655.050 918.600 ;
        RECT 634.950 917.100 637.050 917.400 ;
        RECT 551.400 914.400 594.600 915.600 ;
        RECT 406.950 911.400 423.600 912.600 ;
        RECT 454.950 912.450 457.050 912.900 ;
        RECT 460.950 912.450 463.050 912.900 ;
        RECT 406.950 910.800 409.050 911.400 ;
        RECT 454.950 911.250 463.050 912.450 ;
        RECT 454.950 910.800 457.050 911.250 ;
        RECT 460.950 910.800 463.050 911.250 ;
        RECT 481.950 912.600 484.050 912.900 ;
        RECT 493.950 912.600 496.050 913.050 ;
        RECT 551.400 912.900 552.600 914.400 ;
        RECT 481.950 911.400 496.050 912.600 ;
        RECT 481.950 910.800 484.050 911.400 ;
        RECT 493.950 910.950 496.050 911.400 ;
        RECT 550.950 910.800 553.050 912.900 ;
        RECT 583.950 912.600 586.050 913.050 ;
        RECT 589.950 912.600 592.050 912.900 ;
        RECT 583.950 911.400 592.050 912.600 ;
        RECT 593.400 912.600 594.600 914.400 ;
        RECT 637.950 912.600 640.050 912.900 ;
        RECT 593.400 911.400 640.050 912.600 ;
        RECT 583.950 910.950 586.050 911.400 ;
        RECT 589.950 910.800 592.050 911.400 ;
        RECT 637.950 910.800 640.050 911.400 ;
        RECT 187.950 908.400 213.600 909.600 ;
        RECT 295.950 909.600 298.050 910.050 ;
        RECT 304.950 909.600 307.050 910.050 ;
        RECT 295.950 908.400 307.050 909.600 ;
        RECT 127.950 907.950 130.050 908.400 ;
        RECT 187.950 907.950 190.050 908.400 ;
        RECT 199.950 907.950 202.050 908.400 ;
        RECT 295.950 907.950 298.050 908.400 ;
        RECT 304.950 907.950 307.050 908.400 ;
        RECT 595.950 909.600 598.050 910.050 ;
        RECT 601.950 909.600 604.050 910.050 ;
        RECT 595.950 908.400 604.050 909.600 ;
        RECT 595.950 907.950 598.050 908.400 ;
        RECT 601.950 907.950 604.050 908.400 ;
        RECT 619.950 909.600 622.050 910.050 ;
        RECT 634.950 909.600 637.050 910.050 ;
        RECT 619.950 908.400 637.050 909.600 ;
        RECT 619.950 907.950 622.050 908.400 ;
        RECT 634.950 907.950 637.050 908.400 ;
        RECT 643.950 909.600 646.050 910.050 ;
        RECT 650.400 909.600 651.600 917.400 ;
        RECT 652.950 917.100 655.050 917.400 ;
        RECT 673.950 918.600 676.050 919.200 ;
        RECT 682.950 918.600 685.050 919.050 ;
        RECT 673.950 917.400 685.050 918.600 ;
        RECT 673.950 917.100 676.050 917.400 ;
        RECT 682.950 916.950 685.050 917.400 ;
        RECT 724.950 918.750 727.050 919.200 ;
        RECT 733.950 918.750 736.050 919.200 ;
        RECT 724.950 917.550 736.050 918.750 ;
        RECT 769.950 918.600 772.050 919.200 ;
        RECT 724.950 917.100 727.050 917.550 ;
        RECT 733.950 917.100 736.050 917.550 ;
        RECT 755.400 917.400 772.050 918.600 ;
        RECT 755.400 912.900 756.600 917.400 ;
        RECT 769.950 917.100 772.050 917.400 ;
        RECT 808.950 917.100 811.050 919.200 ;
        RECT 823.950 917.100 826.050 919.200 ;
        RECT 838.950 918.600 841.050 919.050 ;
        RECT 830.400 917.400 841.050 918.600 ;
        RECT 809.400 913.050 810.600 917.100 ;
        RECT 824.400 913.050 825.600 917.100 ;
        RECT 830.400 915.600 831.600 917.400 ;
        RECT 838.950 916.950 841.050 917.400 ;
        RECT 859.950 917.100 862.050 919.200 ;
        RECT 667.950 912.450 670.050 912.900 ;
        RECT 676.950 912.450 679.050 912.900 ;
        RECT 667.950 911.250 679.050 912.450 ;
        RECT 667.950 910.800 670.050 911.250 ;
        RECT 676.950 910.800 679.050 911.250 ;
        RECT 682.950 912.450 685.050 912.900 ;
        RECT 721.950 912.450 724.050 912.900 ;
        RECT 682.950 911.250 724.050 912.450 ;
        RECT 682.950 910.800 685.050 911.250 ;
        RECT 721.950 910.800 724.050 911.250 ;
        RECT 754.950 910.800 757.050 912.900 ;
        RECT 766.950 912.600 769.050 912.900 ;
        RECT 775.950 912.600 778.050 913.050 ;
        RECT 766.950 911.400 778.050 912.600 ;
        RECT 766.950 910.800 769.050 911.400 ;
        RECT 775.950 910.950 778.050 911.400 ;
        RECT 781.950 912.600 784.050 913.050 ;
        RECT 793.950 912.600 796.050 913.050 ;
        RECT 781.950 911.400 796.050 912.600 ;
        RECT 781.950 910.950 784.050 911.400 ;
        RECT 793.950 910.950 796.050 911.400 ;
        RECT 805.950 911.400 810.600 913.050 ;
        RECT 820.950 911.400 825.600 913.050 ;
        RECT 827.400 914.400 831.600 915.600 ;
        RECT 860.400 915.600 861.600 917.100 ;
        RECT 868.950 915.600 871.050 916.050 ;
        RECT 860.400 914.400 871.050 915.600 ;
        RECT 827.400 912.900 828.600 914.400 ;
        RECT 868.950 913.950 871.050 914.400 ;
        RECT 805.950 910.950 810.000 911.400 ;
        RECT 820.950 910.950 825.000 911.400 ;
        RECT 826.950 910.800 829.050 912.900 ;
        RECT 835.950 912.600 838.050 912.900 ;
        RECT 856.950 912.600 859.050 912.900 ;
        RECT 835.950 911.400 859.050 912.600 ;
        RECT 835.950 910.800 838.050 911.400 ;
        RECT 856.950 910.800 859.050 911.400 ;
        RECT 643.950 908.400 651.600 909.600 ;
        RECT 862.950 909.600 865.050 910.050 ;
        RECT 892.950 909.600 895.050 910.050 ;
        RECT 862.950 908.400 895.050 909.600 ;
        RECT 643.950 907.950 646.050 908.400 ;
        RECT 862.950 907.950 865.050 908.400 ;
        RECT 892.950 907.950 895.050 908.400 ;
        RECT 79.950 906.600 82.050 907.050 ;
        RECT 94.950 906.600 97.050 907.050 ;
        RECT 79.950 905.400 97.050 906.600 ;
        RECT 79.950 904.950 82.050 905.400 ;
        RECT 94.950 904.950 97.050 905.400 ;
        RECT 115.950 906.600 118.050 907.050 ;
        RECT 223.950 906.600 226.050 907.050 ;
        RECT 274.950 906.600 277.050 907.050 ;
        RECT 406.950 906.600 409.050 907.050 ;
        RECT 412.950 906.600 415.050 907.050 ;
        RECT 115.950 905.400 415.050 906.600 ;
        RECT 115.950 904.950 118.050 905.400 ;
        RECT 223.950 904.950 226.050 905.400 ;
        RECT 274.950 904.950 277.050 905.400 ;
        RECT 406.950 904.950 409.050 905.400 ;
        RECT 412.950 904.950 415.050 905.400 ;
        RECT 448.950 906.600 451.050 907.050 ;
        RECT 508.950 906.600 511.050 907.050 ;
        RECT 517.950 906.600 520.050 907.050 ;
        RECT 448.950 905.400 520.050 906.600 ;
        RECT 448.950 904.950 451.050 905.400 ;
        RECT 508.950 904.950 511.050 905.400 ;
        RECT 517.950 904.950 520.050 905.400 ;
        RECT 544.950 906.600 547.050 907.050 ;
        RECT 556.950 906.600 559.050 907.050 ;
        RECT 544.950 905.400 559.050 906.600 ;
        RECT 544.950 904.950 547.050 905.400 ;
        RECT 556.950 904.950 559.050 905.400 ;
        RECT 631.950 906.600 634.050 907.050 ;
        RECT 640.950 906.600 643.050 907.050 ;
        RECT 631.950 905.400 643.050 906.600 ;
        RECT 631.950 904.950 634.050 905.400 ;
        RECT 640.950 904.950 643.050 905.400 ;
        RECT 658.950 906.600 661.050 907.050 ;
        RECT 673.800 906.600 675.900 907.050 ;
        RECT 658.950 905.400 675.900 906.600 ;
        RECT 658.950 904.950 661.050 905.400 ;
        RECT 673.800 904.950 675.900 905.400 ;
        RECT 676.950 906.600 679.050 907.050 ;
        RECT 685.950 906.600 688.050 907.050 ;
        RECT 700.950 906.600 703.050 907.050 ;
        RECT 676.950 905.400 703.050 906.600 ;
        RECT 676.950 904.950 679.050 905.400 ;
        RECT 685.950 904.950 688.050 905.400 ;
        RECT 700.950 904.950 703.050 905.400 ;
        RECT 739.950 906.600 742.050 907.050 ;
        RECT 766.950 906.600 769.050 907.050 ;
        RECT 739.950 905.400 769.050 906.600 ;
        RECT 739.950 904.950 742.050 905.400 ;
        RECT 766.950 904.950 769.050 905.400 ;
        RECT 781.950 906.600 784.050 907.050 ;
        RECT 811.950 906.600 814.050 907.050 ;
        RECT 781.950 905.400 814.050 906.600 ;
        RECT 781.950 904.950 784.050 905.400 ;
        RECT 811.950 904.950 814.050 905.400 ;
        RECT 847.950 906.600 850.050 907.050 ;
        RECT 859.950 906.600 862.050 907.050 ;
        RECT 847.950 905.400 862.050 906.600 ;
        RECT 847.950 904.950 850.050 905.400 ;
        RECT 859.950 904.950 862.050 905.400 ;
        RECT 118.950 903.600 121.050 904.050 ;
        RECT 145.950 903.600 148.050 904.050 ;
        RECT 208.950 903.600 211.050 904.050 ;
        RECT 118.950 902.400 211.050 903.600 ;
        RECT 118.950 901.950 121.050 902.400 ;
        RECT 145.950 901.950 148.050 902.400 ;
        RECT 208.950 901.950 211.050 902.400 ;
        RECT 259.950 903.600 262.050 904.050 ;
        RECT 292.950 903.600 295.050 904.050 ;
        RECT 259.950 902.400 295.050 903.600 ;
        RECT 259.950 901.950 262.050 902.400 ;
        RECT 292.950 901.950 295.050 902.400 ;
        RECT 565.950 903.600 568.050 904.050 ;
        RECT 622.950 903.600 625.050 904.050 ;
        RECT 649.950 903.600 652.050 904.050 ;
        RECT 772.950 903.600 775.050 904.050 ;
        RECT 820.950 903.600 823.050 904.050 ;
        RECT 565.950 902.400 823.050 903.600 ;
        RECT 565.950 901.950 568.050 902.400 ;
        RECT 622.950 901.950 625.050 902.400 ;
        RECT 649.950 901.950 652.050 902.400 ;
        RECT 772.950 901.950 775.050 902.400 ;
        RECT 820.950 901.950 823.050 902.400 ;
        RECT 88.950 900.600 91.050 901.050 ;
        RECT 127.950 900.600 130.050 901.050 ;
        RECT 88.950 899.400 130.050 900.600 ;
        RECT 88.950 898.950 91.050 899.400 ;
        RECT 127.950 898.950 130.050 899.400 ;
        RECT 202.950 900.600 205.050 901.050 ;
        RECT 235.950 900.600 238.050 901.050 ;
        RECT 202.950 899.400 238.050 900.600 ;
        RECT 202.950 898.950 205.050 899.400 ;
        RECT 235.950 898.950 238.050 899.400 ;
        RECT 307.950 900.600 310.050 901.050 ;
        RECT 532.950 900.600 535.050 901.050 ;
        RECT 307.950 899.400 535.050 900.600 ;
        RECT 307.950 898.950 310.050 899.400 ;
        RECT 532.950 898.950 535.050 899.400 ;
        RECT 568.950 900.600 571.050 901.050 ;
        RECT 628.950 900.600 631.050 901.050 ;
        RECT 568.950 899.400 631.050 900.600 ;
        RECT 568.950 898.950 571.050 899.400 ;
        RECT 628.950 898.950 631.050 899.400 ;
        RECT 634.950 900.600 637.050 901.050 ;
        RECT 649.800 900.600 651.900 900.900 ;
        RECT 634.950 899.400 651.900 900.600 ;
        RECT 634.950 898.950 637.050 899.400 ;
        RECT 649.800 898.800 651.900 899.400 ;
        RECT 652.950 900.600 655.050 901.050 ;
        RECT 664.950 900.600 667.050 901.050 ;
        RECT 652.950 899.400 667.050 900.600 ;
        RECT 652.950 898.950 655.050 899.400 ;
        RECT 664.950 898.950 667.050 899.400 ;
        RECT 718.950 900.600 721.050 901.050 ;
        RECT 727.950 900.600 730.050 901.050 ;
        RECT 718.950 899.400 730.050 900.600 ;
        RECT 718.950 898.950 721.050 899.400 ;
        RECT 727.950 898.950 730.050 899.400 ;
        RECT 733.950 900.600 736.050 901.050 ;
        RECT 781.950 900.600 784.050 901.050 ;
        RECT 733.950 899.400 784.050 900.600 ;
        RECT 733.950 898.950 736.050 899.400 ;
        RECT 781.950 898.950 784.050 899.400 ;
        RECT 805.950 900.600 808.050 901.050 ;
        RECT 811.950 900.600 814.050 901.050 ;
        RECT 805.950 899.400 814.050 900.600 ;
        RECT 805.950 898.950 808.050 899.400 ;
        RECT 811.950 898.950 814.050 899.400 ;
        RECT 862.950 900.600 865.050 901.050 ;
        RECT 868.950 900.600 871.050 901.050 ;
        RECT 895.950 900.600 898.050 901.050 ;
        RECT 862.950 899.400 898.050 900.600 ;
        RECT 862.950 898.950 865.050 899.400 ;
        RECT 868.950 898.950 871.050 899.400 ;
        RECT 895.950 898.950 898.050 899.400 ;
        RECT 97.950 897.600 100.050 898.050 ;
        RECT 118.950 897.600 121.050 898.050 ;
        RECT 97.950 896.400 121.050 897.600 ;
        RECT 97.950 895.950 100.050 896.400 ;
        RECT 118.950 895.950 121.050 896.400 ;
        RECT 151.950 897.600 154.050 898.050 ;
        RECT 178.950 897.600 181.050 898.050 ;
        RECT 211.950 897.600 214.050 898.050 ;
        RECT 151.950 896.400 214.050 897.600 ;
        RECT 151.950 895.950 154.050 896.400 ;
        RECT 178.950 895.950 181.050 896.400 ;
        RECT 211.950 895.950 214.050 896.400 ;
        RECT 523.950 897.600 526.050 898.050 ;
        RECT 535.950 897.600 538.050 898.050 ;
        RECT 562.950 897.600 565.050 898.050 ;
        RECT 670.950 897.600 673.050 898.050 ;
        RECT 523.950 896.400 673.050 897.600 ;
        RECT 523.950 895.950 526.050 896.400 ;
        RECT 535.950 895.950 538.050 896.400 ;
        RECT 562.950 895.950 565.050 896.400 ;
        RECT 670.950 895.950 673.050 896.400 ;
        RECT 694.950 897.600 697.050 898.050 ;
        RECT 709.950 897.600 712.050 898.050 ;
        RECT 748.950 897.600 751.050 898.050 ;
        RECT 694.950 896.400 751.050 897.600 ;
        RECT 694.950 895.950 697.050 896.400 ;
        RECT 709.950 895.950 712.050 896.400 ;
        RECT 748.950 895.950 751.050 896.400 ;
        RECT 859.950 897.600 862.050 898.050 ;
        RECT 868.950 897.600 871.050 897.900 ;
        RECT 889.950 897.600 892.050 898.050 ;
        RECT 859.950 896.400 892.050 897.600 ;
        RECT 859.950 895.950 862.050 896.400 ;
        RECT 868.950 895.800 871.050 896.400 ;
        RECT 889.950 895.950 892.050 896.400 ;
        RECT 55.950 894.600 58.050 895.050 ;
        RECT 94.950 894.600 97.050 895.050 ;
        RECT 55.950 893.400 97.050 894.600 ;
        RECT 55.950 892.950 58.050 893.400 ;
        RECT 94.950 892.950 97.050 893.400 ;
        RECT 265.950 894.600 268.050 895.050 ;
        RECT 280.950 894.600 283.050 895.050 ;
        RECT 265.950 893.400 283.050 894.600 ;
        RECT 265.950 892.950 268.050 893.400 ;
        RECT 280.950 892.950 283.050 893.400 ;
        RECT 319.950 894.600 322.050 895.050 ;
        RECT 364.950 894.600 367.050 895.050 ;
        RECT 319.950 893.400 367.050 894.600 ;
        RECT 319.950 892.950 322.050 893.400 ;
        RECT 364.950 892.950 367.050 893.400 ;
        RECT 628.950 894.600 631.050 895.050 ;
        RECT 667.950 894.600 670.050 895.050 ;
        RECT 628.950 893.400 670.050 894.600 ;
        RECT 628.950 892.950 631.050 893.400 ;
        RECT 667.950 892.950 670.050 893.400 ;
        RECT 706.950 894.600 709.050 895.050 ;
        RECT 715.950 894.600 718.050 895.050 ;
        RECT 766.950 894.600 769.050 895.050 ;
        RECT 706.950 893.400 718.050 894.600 ;
        RECT 706.950 892.950 709.050 893.400 ;
        RECT 715.950 892.950 718.050 893.400 ;
        RECT 722.400 893.400 769.050 894.600 ;
        RECT 148.950 891.600 151.050 892.050 ;
        RECT 160.950 891.600 163.050 892.050 ;
        RECT 148.950 890.400 163.050 891.600 ;
        RECT 148.950 889.950 151.050 890.400 ;
        RECT 160.950 889.950 163.050 890.400 ;
        RECT 208.950 891.600 211.050 892.050 ;
        RECT 244.950 891.600 247.050 892.050 ;
        RECT 208.950 890.400 247.050 891.600 ;
        RECT 208.950 889.950 211.050 890.400 ;
        RECT 244.950 889.950 247.050 890.400 ;
        RECT 283.950 891.600 286.050 892.050 ;
        RECT 316.950 891.600 319.050 892.050 ;
        RECT 283.950 890.400 319.050 891.600 ;
        RECT 283.950 889.950 286.050 890.400 ;
        RECT 316.950 889.950 319.050 890.400 ;
        RECT 382.950 891.600 385.050 892.050 ;
        RECT 394.950 891.600 397.050 892.050 ;
        RECT 424.950 891.600 427.050 892.050 ;
        RECT 382.950 890.400 427.050 891.600 ;
        RECT 382.950 889.950 385.050 890.400 ;
        RECT 394.950 889.950 397.050 890.400 ;
        RECT 424.950 889.950 427.050 890.400 ;
        RECT 490.950 891.600 493.050 892.050 ;
        RECT 502.950 891.600 505.050 892.050 ;
        RECT 490.950 890.400 505.050 891.600 ;
        RECT 490.950 889.950 493.050 890.400 ;
        RECT 502.950 889.950 505.050 890.400 ;
        RECT 595.950 891.600 598.050 892.050 ;
        RECT 604.950 891.600 607.050 892.050 ;
        RECT 619.950 891.600 622.050 892.050 ;
        RECT 673.950 891.600 676.050 892.050 ;
        RECT 679.950 891.600 682.050 892.050 ;
        RECT 595.950 890.400 666.600 891.600 ;
        RECT 595.950 889.950 598.050 890.400 ;
        RECT 604.950 889.950 607.050 890.400 ;
        RECT 619.950 889.950 622.050 890.400 ;
        RECT 665.400 889.050 666.600 890.400 ;
        RECT 673.950 890.400 682.050 891.600 ;
        RECT 673.950 889.950 676.050 890.400 ;
        RECT 679.950 889.950 682.050 890.400 ;
        RECT 691.950 891.600 694.050 892.050 ;
        RECT 722.400 891.600 723.600 893.400 ;
        RECT 766.950 892.950 769.050 893.400 ;
        RECT 829.950 894.600 832.050 895.050 ;
        RECT 847.950 894.600 850.050 895.050 ;
        RECT 829.950 893.400 850.050 894.600 ;
        RECT 829.950 892.950 832.050 893.400 ;
        RECT 847.950 892.950 850.050 893.400 ;
        RECT 877.950 894.600 880.050 895.050 ;
        RECT 916.950 894.600 919.050 895.050 ;
        RECT 877.950 893.400 919.050 894.600 ;
        RECT 877.950 892.950 880.050 893.400 ;
        RECT 916.950 892.950 919.050 893.400 ;
        RECT 691.950 890.400 723.600 891.600 ;
        RECT 724.950 891.600 727.050 892.050 ;
        RECT 736.950 891.600 739.050 892.050 ;
        RECT 787.950 891.600 790.050 892.050 ;
        RECT 724.950 890.400 790.050 891.600 ;
        RECT 691.950 889.950 694.050 890.400 ;
        RECT 724.950 889.950 727.050 890.400 ;
        RECT 736.950 889.950 739.050 890.400 ;
        RECT 787.950 889.950 790.050 890.400 ;
        RECT 823.950 891.600 826.050 892.050 ;
        RECT 853.950 891.600 856.050 892.050 ;
        RECT 823.950 890.400 856.050 891.600 ;
        RECT 823.950 889.950 826.050 890.400 ;
        RECT 853.950 889.950 856.050 890.400 ;
        RECT 889.950 891.600 892.050 892.050 ;
        RECT 904.950 891.600 907.050 892.050 ;
        RECT 889.950 890.400 907.050 891.600 ;
        RECT 889.950 889.950 892.050 890.400 ;
        RECT 904.950 889.950 907.050 890.400 ;
        RECT 16.950 888.600 19.050 889.050 ;
        RECT 58.950 888.600 61.050 889.050 ;
        RECT 82.950 888.600 85.050 889.050 ;
        RECT 184.950 888.600 187.050 889.050 ;
        RECT 16.950 887.400 85.050 888.600 ;
        RECT 16.950 886.950 19.050 887.400 ;
        RECT 58.950 886.950 61.050 887.400 ;
        RECT 82.950 886.950 85.050 887.400 ;
        RECT 170.400 887.400 187.050 888.600 ;
        RECT 170.400 886.200 171.600 887.400 ;
        RECT 184.950 886.950 187.050 887.400 ;
        RECT 445.950 888.600 448.050 889.050 ;
        RECT 472.950 888.600 475.050 889.050 ;
        RECT 526.950 888.600 529.050 889.050 ;
        RECT 541.950 888.600 544.050 889.050 ;
        RECT 550.950 888.600 553.050 889.050 ;
        RECT 445.950 887.400 504.600 888.600 ;
        RECT 445.950 886.950 448.050 887.400 ;
        RECT 472.950 886.950 475.050 887.400 ;
        RECT 22.950 884.100 25.050 886.200 ;
        RECT 31.950 885.600 34.050 886.050 ;
        RECT 40.950 885.600 43.050 886.200 ;
        RECT 31.950 884.400 43.050 885.600 ;
        RECT 23.400 879.600 24.600 884.100 ;
        RECT 31.950 883.950 34.050 884.400 ;
        RECT 40.950 884.100 43.050 884.400 ;
        RECT 49.950 885.750 52.050 886.200 ;
        RECT 58.950 885.750 61.050 886.200 ;
        RECT 49.950 884.550 61.050 885.750 ;
        RECT 49.950 884.100 52.050 884.550 ;
        RECT 58.950 884.100 61.050 884.550 ;
        RECT 64.950 885.600 67.050 886.200 ;
        RECT 73.950 885.600 76.050 886.050 ;
        RECT 64.950 884.400 76.050 885.600 ;
        RECT 64.950 884.100 67.050 884.400 ;
        RECT 73.950 883.950 76.050 884.400 ;
        RECT 109.950 885.600 112.050 886.200 ;
        RECT 121.950 885.600 124.050 886.050 ;
        RECT 133.950 885.600 136.050 886.200 ;
        RECT 109.950 884.400 136.050 885.600 ;
        RECT 109.950 884.100 112.050 884.400 ;
        RECT 121.950 883.950 124.050 884.400 ;
        RECT 133.950 884.100 136.050 884.400 ;
        RECT 139.950 884.100 142.050 886.200 ;
        RECT 157.950 885.750 160.050 886.200 ;
        RECT 169.950 885.750 172.050 886.200 ;
        RECT 157.950 884.550 172.050 885.750 ;
        RECT 157.950 884.100 160.050 884.550 ;
        RECT 169.950 884.100 172.050 884.550 ;
        RECT 193.950 885.750 196.050 886.200 ;
        RECT 208.950 885.750 211.050 886.200 ;
        RECT 193.950 884.550 211.050 885.750 ;
        RECT 193.950 884.100 196.050 884.550 ;
        RECT 208.950 884.100 211.050 884.550 ;
        RECT 232.950 885.750 235.050 886.200 ;
        RECT 241.950 885.750 244.050 886.200 ;
        RECT 232.950 884.550 244.050 885.750 ;
        RECT 232.950 884.100 235.050 884.550 ;
        RECT 241.950 884.100 244.050 884.550 ;
        RECT 250.950 884.100 253.050 886.200 ;
        RECT 271.950 884.100 274.050 886.200 ;
        RECT 280.950 885.750 283.050 886.200 ;
        RECT 298.950 885.750 301.050 886.200 ;
        RECT 280.950 884.550 301.050 885.750 ;
        RECT 280.950 884.100 283.050 884.550 ;
        RECT 298.950 884.100 301.050 884.550 ;
        RECT 337.950 885.600 340.050 886.200 ;
        RECT 352.950 885.600 355.050 886.200 ;
        RECT 367.950 885.600 370.050 886.050 ;
        RECT 379.950 885.750 382.050 886.200 ;
        RECT 385.950 885.750 388.050 886.200 ;
        RECT 337.950 884.400 378.600 885.600 ;
        RECT 337.950 884.100 340.050 884.400 ;
        RECT 352.950 884.100 355.050 884.400 ;
        RECT 140.400 882.600 141.600 884.100 ;
        RECT 251.400 882.600 252.600 884.100 ;
        RECT 272.400 882.600 273.600 884.100 ;
        RECT 367.950 883.950 370.050 884.400 ;
        RECT 140.400 881.400 150.600 882.600 ;
        RECT 251.400 881.400 273.600 882.600 ;
        RECT 43.950 879.600 46.050 879.900 ;
        RECT 23.400 878.400 46.050 879.600 ;
        RECT 43.950 877.800 46.050 878.400 ;
        RECT 61.950 879.600 64.050 879.900 ;
        RECT 79.950 879.600 82.050 879.900 ;
        RECT 61.950 878.400 84.600 879.600 ;
        RECT 61.950 877.800 64.050 878.400 ;
        RECT 79.950 877.800 82.050 878.400 ;
        RECT 49.950 876.600 52.050 877.050 ;
        RECT 58.950 876.600 61.050 877.050 ;
        RECT 49.950 875.400 61.050 876.600 ;
        RECT 83.400 876.600 84.600 878.400 ;
        RECT 85.950 879.450 88.050 879.900 ;
        RECT 91.950 879.450 94.050 879.900 ;
        RECT 85.950 878.250 94.050 879.450 ;
        RECT 149.400 879.600 150.600 881.400 ;
        RECT 272.400 880.050 273.600 881.400 ;
        RECT 181.950 879.600 184.050 879.900 ;
        RECT 196.950 879.600 199.050 879.900 ;
        RECT 149.400 878.400 199.050 879.600 ;
        RECT 85.950 877.800 88.050 878.250 ;
        RECT 91.950 877.800 94.050 878.250 ;
        RECT 181.950 877.800 184.050 878.400 ;
        RECT 196.950 877.800 199.050 878.400 ;
        RECT 211.950 879.600 214.050 880.050 ;
        RECT 220.950 879.600 223.050 879.900 ;
        RECT 211.950 878.400 223.050 879.600 ;
        RECT 211.950 877.950 214.050 878.400 ;
        RECT 220.950 877.800 223.050 878.400 ;
        RECT 238.950 879.600 241.050 879.900 ;
        RECT 253.950 879.600 256.050 879.900 ;
        RECT 238.950 878.400 256.050 879.600 ;
        RECT 238.950 877.800 241.050 878.400 ;
        RECT 253.950 877.800 256.050 878.400 ;
        RECT 268.950 878.400 273.600 880.050 ;
        RECT 274.950 879.600 277.050 879.900 ;
        RECT 295.950 879.600 298.050 879.900 ;
        RECT 274.950 878.400 298.050 879.600 ;
        RECT 268.950 877.950 273.000 878.400 ;
        RECT 274.950 877.800 277.050 878.400 ;
        RECT 295.950 877.800 298.050 878.400 ;
        RECT 301.950 879.600 304.050 879.900 ;
        RECT 316.950 879.600 319.050 879.900 ;
        RECT 301.950 878.400 319.050 879.600 ;
        RECT 301.950 877.800 304.050 878.400 ;
        RECT 316.950 877.800 319.050 878.400 ;
        RECT 355.950 879.600 358.050 879.900 ;
        RECT 370.950 879.600 373.050 879.900 ;
        RECT 355.950 878.400 373.050 879.600 ;
        RECT 377.400 879.600 378.600 884.400 ;
        RECT 379.950 884.550 388.050 885.750 ;
        RECT 379.950 884.100 382.050 884.550 ;
        RECT 385.950 884.100 388.050 884.550 ;
        RECT 400.950 885.600 403.050 886.200 ;
        RECT 406.950 885.600 409.050 886.050 ;
        RECT 400.950 884.400 409.050 885.600 ;
        RECT 400.950 884.100 403.050 884.400 ;
        RECT 406.950 883.950 409.050 884.400 ;
        RECT 454.950 885.600 457.050 886.200 ;
        RECT 478.950 885.600 481.050 886.200 ;
        RECT 454.950 884.400 474.600 885.600 ;
        RECT 454.950 884.100 457.050 884.400 ;
        RECT 391.950 879.600 394.050 879.900 ;
        RECT 377.400 878.400 394.050 879.600 ;
        RECT 355.950 877.800 358.050 878.400 ;
        RECT 370.950 877.800 373.050 878.400 ;
        RECT 391.950 877.800 394.050 878.400 ;
        RECT 397.950 879.600 400.050 879.900 ;
        RECT 415.950 879.600 418.050 879.900 ;
        RECT 397.950 878.400 418.050 879.600 ;
        RECT 397.950 877.800 400.050 878.400 ;
        RECT 415.950 877.800 418.050 878.400 ;
        RECT 430.950 879.450 433.050 879.900 ;
        RECT 448.950 879.450 451.050 883.050 ;
        RECT 469.950 879.450 472.050 879.900 ;
        RECT 430.950 878.250 472.050 879.450 ;
        RECT 473.400 879.600 474.600 884.400 ;
        RECT 478.950 884.400 498.600 885.600 ;
        RECT 478.950 884.100 481.050 884.400 ;
        RECT 497.400 879.900 498.600 884.400 ;
        RECT 499.950 884.100 502.050 886.200 ;
        RECT 503.400 885.600 504.600 887.400 ;
        RECT 526.950 887.400 534.600 888.600 ;
        RECT 526.950 886.950 529.050 887.400 ;
        RECT 505.950 885.600 508.050 886.200 ;
        RECT 503.400 884.400 508.050 885.600 ;
        RECT 505.950 884.100 508.050 884.400 ;
        RECT 517.950 884.100 520.050 886.200 ;
        RECT 533.400 885.600 534.600 887.400 ;
        RECT 541.950 887.400 553.050 888.600 ;
        RECT 541.950 886.950 544.050 887.400 ;
        RECT 550.950 886.950 553.050 887.400 ;
        RECT 637.950 888.600 640.050 889.050 ;
        RECT 643.950 888.600 646.050 889.050 ;
        RECT 637.950 887.400 646.050 888.600 ;
        RECT 637.950 886.950 640.050 887.400 ;
        RECT 643.950 886.950 646.050 887.400 ;
        RECT 655.950 888.600 658.050 889.050 ;
        RECT 664.950 888.600 667.050 889.050 ;
        RECT 742.950 888.600 745.050 889.050 ;
        RECT 655.950 887.400 663.600 888.600 ;
        RECT 655.950 886.950 658.050 887.400 ;
        RECT 553.950 885.600 556.050 886.050 ;
        RECT 533.400 884.400 556.050 885.600 ;
        RECT 475.950 879.600 478.050 879.900 ;
        RECT 473.400 878.400 478.050 879.600 ;
        RECT 430.950 877.800 433.050 878.250 ;
        RECT 469.950 877.800 472.050 878.250 ;
        RECT 475.950 877.800 478.050 878.400 ;
        RECT 496.950 877.800 499.050 879.900 ;
        RECT 500.400 877.050 501.600 884.100 ;
        RECT 502.950 879.600 505.050 879.900 ;
        RECT 518.400 879.600 519.600 884.100 ;
        RECT 553.950 883.950 556.050 884.400 ;
        RECT 613.950 884.100 616.050 886.200 ;
        RECT 619.950 885.600 622.050 886.200 ;
        RECT 619.950 884.400 630.600 885.600 ;
        RECT 619.950 884.100 622.050 884.400 ;
        RECT 550.950 882.600 553.050 883.050 ;
        RECT 527.400 881.400 553.050 882.600 ;
        RECT 614.400 882.600 615.600 884.100 ;
        RECT 614.400 882.000 627.450 882.600 ;
        RECT 614.400 881.400 628.050 882.000 ;
        RECT 527.400 879.900 528.600 881.400 ;
        RECT 550.950 880.950 553.050 881.400 ;
        RECT 625.950 880.050 628.050 881.400 ;
        RECT 502.950 878.400 519.600 879.600 ;
        RECT 502.950 877.800 505.050 878.400 ;
        RECT 526.950 877.800 529.050 879.900 ;
        RECT 532.950 879.600 535.050 880.050 ;
        RECT 544.950 879.600 547.050 879.900 ;
        RECT 532.950 878.400 547.050 879.600 ;
        RECT 532.950 877.950 535.050 878.400 ;
        RECT 544.950 877.800 547.050 878.400 ;
        RECT 553.950 879.450 556.050 879.900 ;
        RECT 568.950 879.450 571.050 879.900 ;
        RECT 553.950 878.250 571.050 879.450 ;
        RECT 553.950 877.800 556.050 878.250 ;
        RECT 568.950 877.800 571.050 878.250 ;
        RECT 586.950 879.600 589.050 879.900 ;
        RECT 610.950 879.600 613.050 879.900 ;
        RECT 586.950 878.400 613.050 879.600 ;
        RECT 586.950 877.800 589.050 878.400 ;
        RECT 610.950 877.800 613.050 878.400 ;
        RECT 625.800 879.000 628.050 880.050 ;
        RECT 629.400 879.900 630.600 884.400 ;
        RECT 631.950 884.100 634.050 886.200 ;
        RECT 662.400 885.600 663.600 887.400 ;
        RECT 664.950 887.400 745.050 888.600 ;
        RECT 664.950 886.950 667.050 887.400 ;
        RECT 742.950 886.950 745.050 887.400 ;
        RECT 691.950 885.600 694.050 886.050 ;
        RECT 662.400 884.400 694.050 885.600 ;
        RECT 625.800 877.950 627.900 879.000 ;
        RECT 628.950 877.800 631.050 879.900 ;
        RECT 632.400 879.600 633.600 884.100 ;
        RECT 691.950 883.950 694.050 884.400 ;
        RECT 700.950 885.600 705.000 886.050 ;
        RECT 711.000 885.600 715.050 886.050 ;
        RECT 700.950 883.950 705.600 885.600 ;
        RECT 640.950 879.600 643.050 880.050 ;
        RECT 704.400 879.900 705.600 883.950 ;
        RECT 710.400 883.950 715.050 885.600 ;
        RECT 718.950 885.600 721.050 886.050 ;
        RECT 730.950 885.600 733.050 886.200 ;
        RECT 739.950 885.600 742.050 886.050 ;
        RECT 718.950 884.400 729.600 885.600 ;
        RECT 718.950 883.950 721.050 884.400 ;
        RECT 710.400 879.900 711.600 883.950 ;
        RECT 728.400 879.900 729.600 884.400 ;
        RECT 730.950 884.400 742.050 885.600 ;
        RECT 730.950 884.100 733.050 884.400 ;
        RECT 739.950 883.950 742.050 884.400 ;
        RECT 766.950 885.600 771.000 886.050 ;
        RECT 772.950 885.600 775.050 886.200 ;
        RECT 781.950 885.600 784.050 886.050 ;
        RECT 796.950 885.750 799.050 886.200 ;
        RECT 805.950 885.750 808.050 886.200 ;
        RECT 766.950 883.950 771.600 885.600 ;
        RECT 772.950 884.400 780.600 885.600 ;
        RECT 772.950 884.100 775.050 884.400 ;
        RECT 770.400 879.900 771.600 883.950 ;
        RECT 632.400 878.400 643.050 879.600 ;
        RECT 640.950 877.950 643.050 878.400 ;
        RECT 649.950 879.450 652.050 879.900 ;
        RECT 655.950 879.450 658.050 879.900 ;
        RECT 649.950 878.250 658.050 879.450 ;
        RECT 649.950 877.800 652.050 878.250 ;
        RECT 655.950 877.800 658.050 878.250 ;
        RECT 670.950 879.450 673.050 879.900 ;
        RECT 676.950 879.450 679.050 879.900 ;
        RECT 670.950 878.250 679.050 879.450 ;
        RECT 670.950 877.800 673.050 878.250 ;
        RECT 676.950 877.800 679.050 878.250 ;
        RECT 688.950 879.450 691.050 879.900 ;
        RECT 694.950 879.450 697.050 879.900 ;
        RECT 688.950 878.250 697.050 879.450 ;
        RECT 688.950 877.800 691.050 878.250 ;
        RECT 694.950 877.800 697.050 878.250 ;
        RECT 703.950 877.800 706.050 879.900 ;
        RECT 709.950 877.800 712.050 879.900 ;
        RECT 715.950 879.450 718.050 879.900 ;
        RECT 721.950 879.450 724.050 879.900 ;
        RECT 715.950 878.250 724.050 879.450 ;
        RECT 715.950 877.800 718.050 878.250 ;
        RECT 721.950 877.800 724.050 878.250 ;
        RECT 727.950 877.800 730.050 879.900 ;
        RECT 769.950 877.800 772.050 879.900 ;
        RECT 779.400 879.600 780.600 884.400 ;
        RECT 781.950 884.400 792.600 885.600 ;
        RECT 781.950 883.950 784.050 884.400 ;
        RECT 791.400 879.900 792.600 884.400 ;
        RECT 796.950 884.550 808.050 885.750 ;
        RECT 796.950 884.100 799.050 884.550 ;
        RECT 805.950 884.100 808.050 884.550 ;
        RECT 820.950 885.750 823.050 886.200 ;
        RECT 829.950 885.750 832.050 886.200 ;
        RECT 820.950 884.550 832.050 885.750 ;
        RECT 820.950 884.100 823.050 884.550 ;
        RECT 829.950 884.100 832.050 884.550 ;
        RECT 835.950 884.100 838.050 886.200 ;
        RECT 874.950 885.600 877.050 886.200 ;
        RECT 857.400 884.400 877.050 885.600 ;
        RECT 784.950 879.600 787.050 879.900 ;
        RECT 779.400 878.400 787.050 879.600 ;
        RECT 784.950 877.800 787.050 878.400 ;
        RECT 790.950 877.800 793.050 879.900 ;
        RECT 808.950 879.600 811.050 879.900 ;
        RECT 832.950 879.600 835.050 879.900 ;
        RECT 808.950 878.400 835.050 879.600 ;
        RECT 836.400 879.600 837.600 884.100 ;
        RECT 857.400 879.900 858.600 884.400 ;
        RECT 874.950 884.100 877.050 884.400 ;
        RECT 892.950 884.100 895.050 886.200 ;
        RECT 893.400 882.600 894.600 884.100 ;
        RECT 881.400 882.000 894.600 882.600 ;
        RECT 880.950 881.400 894.600 882.000 ;
        RECT 850.950 879.600 853.050 879.900 ;
        RECT 836.400 878.400 853.050 879.600 ;
        RECT 808.950 877.800 811.050 878.400 ;
        RECT 832.950 877.800 835.050 878.400 ;
        RECT 850.950 877.800 853.050 878.400 ;
        RECT 856.950 877.800 859.050 879.900 ;
        RECT 880.950 877.950 883.050 881.400 ;
        RECT 895.950 879.600 898.050 879.900 ;
        RECT 904.950 879.600 907.050 880.050 ;
        RECT 913.950 879.600 916.050 880.050 ;
        RECT 895.950 878.400 916.050 879.600 ;
        RECT 895.950 877.800 898.050 878.400 ;
        RECT 904.950 877.950 907.050 878.400 ;
        RECT 913.950 877.950 916.050 878.400 ;
        RECT 106.950 876.600 109.050 877.050 ;
        RECT 83.400 875.400 109.050 876.600 ;
        RECT 49.950 874.950 52.050 875.400 ;
        RECT 58.950 874.950 61.050 875.400 ;
        RECT 106.950 874.950 109.050 875.400 ;
        RECT 136.950 876.600 139.050 877.050 ;
        RECT 154.950 876.600 157.050 877.050 ;
        RECT 136.950 875.400 157.050 876.600 ;
        RECT 136.950 874.950 139.050 875.400 ;
        RECT 154.950 874.950 157.050 875.400 ;
        RECT 205.950 876.600 208.050 877.050 ;
        RECT 307.950 876.600 310.050 877.050 ;
        RECT 205.950 875.400 310.050 876.600 ;
        RECT 500.400 876.750 504.000 877.050 ;
        RECT 500.400 875.400 505.050 876.750 ;
        RECT 205.950 874.950 208.050 875.400 ;
        RECT 307.950 874.950 310.050 875.400 ;
        RECT 501.000 874.950 505.050 875.400 ;
        RECT 592.950 876.600 595.050 877.050 ;
        RECT 601.950 876.600 604.050 877.050 ;
        RECT 592.950 875.400 604.050 876.600 ;
        RECT 592.950 874.950 595.050 875.400 ;
        RECT 601.950 874.950 604.050 875.400 ;
        RECT 502.950 874.650 505.050 874.950 ;
        RECT 13.950 873.600 16.050 874.050 ;
        RECT 28.950 873.600 31.050 874.050 ;
        RECT 55.950 873.600 58.050 874.050 ;
        RECT 13.950 872.400 58.050 873.600 ;
        RECT 13.950 871.950 16.050 872.400 ;
        RECT 28.950 871.950 31.050 872.400 ;
        RECT 55.950 871.950 58.050 872.400 ;
        RECT 70.950 873.600 73.050 874.050 ;
        RECT 82.950 873.600 85.050 874.050 ;
        RECT 91.950 873.600 94.050 874.050 ;
        RECT 70.950 872.400 94.050 873.600 ;
        RECT 70.950 871.950 73.050 872.400 ;
        RECT 82.950 871.950 85.050 872.400 ;
        RECT 91.950 871.950 94.050 872.400 ;
        RECT 187.950 873.600 190.050 874.050 ;
        RECT 202.950 873.600 205.050 874.050 ;
        RECT 187.950 872.400 205.050 873.600 ;
        RECT 187.950 871.950 190.050 872.400 ;
        RECT 202.950 871.950 205.050 872.400 ;
        RECT 232.950 873.600 235.050 874.050 ;
        RECT 280.950 873.600 283.050 874.050 ;
        RECT 340.950 873.600 343.050 874.050 ;
        RECT 232.950 872.400 343.050 873.600 ;
        RECT 232.950 871.950 235.050 872.400 ;
        RECT 280.950 871.950 283.050 872.400 ;
        RECT 340.950 871.950 343.050 872.400 ;
        RECT 376.950 873.600 379.050 874.050 ;
        RECT 436.950 873.600 439.050 874.050 ;
        RECT 376.950 872.400 439.050 873.600 ;
        RECT 376.950 871.950 379.050 872.400 ;
        RECT 436.950 871.950 439.050 872.400 ;
        RECT 478.950 873.600 481.050 874.050 ;
        RECT 508.950 873.600 511.050 874.050 ;
        RECT 532.950 873.600 535.050 874.050 ;
        RECT 478.950 872.400 535.050 873.600 ;
        RECT 478.950 871.950 481.050 872.400 ;
        RECT 508.950 871.950 511.050 872.400 ;
        RECT 532.950 871.950 535.050 872.400 ;
        RECT 610.950 873.600 613.050 874.050 ;
        RECT 661.950 873.600 664.050 874.050 ;
        RECT 721.950 873.600 724.050 874.050 ;
        RECT 610.950 872.400 724.050 873.600 ;
        RECT 610.950 871.950 613.050 872.400 ;
        RECT 661.950 871.950 664.050 872.400 ;
        RECT 721.950 871.950 724.050 872.400 ;
        RECT 778.950 873.600 781.050 874.050 ;
        RECT 793.950 873.600 796.050 874.050 ;
        RECT 778.950 872.400 796.050 873.600 ;
        RECT 778.950 871.950 781.050 872.400 ;
        RECT 793.950 871.950 796.050 872.400 ;
        RECT 820.950 873.600 823.050 874.050 ;
        RECT 877.950 873.600 880.050 874.050 ;
        RECT 820.950 872.400 880.050 873.600 ;
        RECT 820.950 871.950 823.050 872.400 ;
        RECT 877.950 871.950 880.050 872.400 ;
        RECT 106.950 870.600 109.050 871.050 ;
        RECT 115.950 870.600 118.050 871.050 ;
        RECT 106.950 869.400 118.050 870.600 ;
        RECT 106.950 868.950 109.050 869.400 ;
        RECT 115.950 868.950 118.050 869.400 ;
        RECT 409.950 870.600 412.050 871.050 ;
        RECT 427.950 870.600 430.050 871.050 ;
        RECT 409.950 869.400 430.050 870.600 ;
        RECT 409.950 868.950 412.050 869.400 ;
        RECT 427.950 868.950 430.050 869.400 ;
        RECT 484.950 870.600 487.050 871.050 ;
        RECT 511.950 870.600 514.050 871.050 ;
        RECT 484.950 869.400 514.050 870.600 ;
        RECT 484.950 868.950 487.050 869.400 ;
        RECT 511.950 868.950 514.050 869.400 ;
        RECT 568.950 870.600 571.050 871.050 ;
        RECT 616.950 870.600 619.050 871.050 ;
        RECT 640.950 870.600 643.050 871.050 ;
        RECT 568.950 869.400 643.050 870.600 ;
        RECT 568.950 868.950 571.050 869.400 ;
        RECT 616.950 868.950 619.050 869.400 ;
        RECT 640.950 868.950 643.050 869.400 ;
        RECT 850.950 870.600 853.050 871.050 ;
        RECT 871.950 870.600 874.050 871.050 ;
        RECT 850.950 869.400 874.050 870.600 ;
        RECT 850.950 868.950 853.050 869.400 ;
        RECT 871.950 868.950 874.050 869.400 ;
        RECT 25.950 867.600 28.050 868.050 ;
        RECT 37.950 867.600 40.050 868.050 ;
        RECT 107.400 867.600 108.600 868.950 ;
        RECT 25.950 866.400 108.600 867.600 ;
        RECT 190.950 867.600 193.050 868.050 ;
        RECT 229.950 867.600 232.050 868.050 ;
        RECT 286.950 867.600 289.050 868.050 ;
        RECT 190.950 866.400 289.050 867.600 ;
        RECT 25.950 865.950 28.050 866.400 ;
        RECT 37.950 865.950 40.050 866.400 ;
        RECT 190.950 865.950 193.050 866.400 ;
        RECT 229.950 865.950 232.050 866.400 ;
        RECT 286.950 865.950 289.050 866.400 ;
        RECT 490.950 867.600 493.050 868.050 ;
        RECT 520.950 867.600 523.050 868.050 ;
        RECT 490.950 866.400 523.050 867.600 ;
        RECT 490.950 865.950 493.050 866.400 ;
        RECT 520.950 865.950 523.050 866.400 ;
        RECT 772.950 867.600 775.050 868.050 ;
        RECT 817.950 867.600 820.050 868.050 ;
        RECT 772.950 866.400 820.050 867.600 ;
        RECT 772.950 865.950 775.050 866.400 ;
        RECT 817.950 865.950 820.050 866.400 ;
        RECT 538.950 864.600 541.050 864.900 ;
        RECT 568.950 864.600 571.050 865.050 ;
        RECT 538.950 863.400 571.050 864.600 ;
        RECT 538.950 862.800 541.050 863.400 ;
        RECT 568.950 862.950 571.050 863.400 ;
        RECT 763.950 864.600 766.050 865.050 ;
        RECT 778.950 864.600 781.050 865.050 ;
        RECT 763.950 863.400 781.050 864.600 ;
        RECT 763.950 862.950 766.050 863.400 ;
        RECT 778.950 862.950 781.050 863.400 ;
        RECT 826.950 864.600 829.050 865.050 ;
        RECT 856.950 864.600 859.050 865.050 ;
        RECT 826.950 863.400 859.050 864.600 ;
        RECT 826.950 862.950 829.050 863.400 ;
        RECT 856.950 862.950 859.050 863.400 ;
        RECT 259.950 861.600 262.050 862.050 ;
        RECT 268.950 861.600 271.050 862.050 ;
        RECT 334.950 861.600 337.050 862.050 ;
        RECT 259.950 860.400 337.050 861.600 ;
        RECT 259.950 859.950 262.050 860.400 ;
        RECT 268.950 859.950 271.050 860.400 ;
        RECT 334.950 859.950 337.050 860.400 ;
        RECT 499.950 861.600 502.050 862.050 ;
        RECT 583.950 861.600 586.050 862.050 ;
        RECT 499.950 860.400 586.050 861.600 ;
        RECT 499.950 859.950 502.050 860.400 ;
        RECT 583.950 859.950 586.050 860.400 ;
        RECT 721.950 861.600 724.050 862.050 ;
        RECT 742.950 861.600 745.050 862.050 ;
        RECT 772.950 861.600 775.050 862.050 ;
        RECT 721.950 860.400 775.050 861.600 ;
        RECT 721.950 859.950 724.050 860.400 ;
        RECT 742.950 859.950 745.050 860.400 ;
        RECT 772.950 859.950 775.050 860.400 ;
        RECT 22.950 858.600 25.050 859.050 ;
        RECT 70.950 858.600 73.050 859.050 ;
        RECT 91.950 858.600 94.050 859.050 ;
        RECT 22.950 857.400 94.050 858.600 ;
        RECT 22.950 856.950 25.050 857.400 ;
        RECT 70.950 856.950 73.050 857.400 ;
        RECT 91.950 856.950 94.050 857.400 ;
        RECT 262.950 858.600 265.050 859.050 ;
        RECT 286.950 858.600 289.050 859.050 ;
        RECT 262.950 857.400 289.050 858.600 ;
        RECT 262.950 856.950 265.050 857.400 ;
        RECT 286.950 856.950 289.050 857.400 ;
        RECT 361.950 858.600 364.050 859.050 ;
        RECT 424.950 858.600 427.050 859.050 ;
        RECT 361.950 857.400 427.050 858.600 ;
        RECT 361.950 856.950 364.050 857.400 ;
        RECT 424.950 856.950 427.050 857.400 ;
        RECT 505.950 858.600 508.050 859.050 ;
        RECT 553.950 858.600 556.050 859.050 ;
        RECT 505.950 857.400 556.050 858.600 ;
        RECT 505.950 856.950 508.050 857.400 ;
        RECT 553.950 856.950 556.050 857.400 ;
        RECT 577.950 858.600 580.050 859.050 ;
        RECT 634.950 858.600 637.050 859.050 ;
        RECT 709.950 858.600 712.050 859.050 ;
        RECT 577.950 857.400 712.050 858.600 ;
        RECT 577.950 856.950 580.050 857.400 ;
        RECT 634.950 856.950 637.050 857.400 ;
        RECT 709.950 856.950 712.050 857.400 ;
        RECT 784.950 858.600 787.050 859.050 ;
        RECT 820.950 858.600 823.050 859.050 ;
        RECT 784.950 857.400 823.050 858.600 ;
        RECT 784.950 856.950 787.050 857.400 ;
        RECT 820.950 856.950 823.050 857.400 ;
        RECT 43.950 855.600 46.050 856.050 ;
        RECT 121.950 855.600 124.050 856.050 ;
        RECT 43.950 854.400 124.050 855.600 ;
        RECT 43.950 853.950 46.050 854.400 ;
        RECT 121.950 853.950 124.050 854.400 ;
        RECT 289.950 855.600 292.050 856.050 ;
        RECT 427.950 855.600 430.050 856.050 ;
        RECT 436.950 855.600 439.050 856.050 ;
        RECT 289.950 854.400 439.050 855.600 ;
        RECT 289.950 853.950 292.050 854.400 ;
        RECT 427.950 853.950 430.050 854.400 ;
        RECT 436.950 853.950 439.050 854.400 ;
        RECT 451.950 855.600 454.050 856.050 ;
        RECT 592.950 855.600 595.050 856.050 ;
        RECT 451.950 854.400 595.050 855.600 ;
        RECT 451.950 853.950 454.050 854.400 ;
        RECT 592.950 853.950 595.050 854.400 ;
        RECT 598.950 855.600 601.050 856.050 ;
        RECT 688.950 855.600 691.050 856.050 ;
        RECT 598.950 854.400 691.050 855.600 ;
        RECT 598.950 853.950 601.050 854.400 ;
        RECT 688.950 853.950 691.050 854.400 ;
        RECT 727.950 855.600 730.050 856.050 ;
        RECT 769.950 855.600 772.050 856.050 ;
        RECT 727.950 854.400 772.050 855.600 ;
        RECT 727.950 853.950 730.050 854.400 ;
        RECT 769.950 853.950 772.050 854.400 ;
        RECT 787.950 855.600 790.050 856.050 ;
        RECT 796.950 855.600 799.050 856.050 ;
        RECT 787.950 854.400 799.050 855.600 ;
        RECT 787.950 853.950 790.050 854.400 ;
        RECT 796.950 853.950 799.050 854.400 ;
        RECT 817.950 855.600 820.050 856.050 ;
        RECT 829.950 855.600 832.050 856.050 ;
        RECT 862.950 855.600 865.050 856.050 ;
        RECT 877.950 855.600 880.050 856.050 ;
        RECT 817.950 854.400 880.050 855.600 ;
        RECT 817.950 853.950 820.050 854.400 ;
        RECT 829.950 853.950 832.050 854.400 ;
        RECT 862.950 853.950 865.050 854.400 ;
        RECT 877.950 853.950 880.050 854.400 ;
        RECT 163.950 852.600 166.050 853.050 ;
        RECT 172.950 852.600 175.050 853.050 ;
        RECT 163.950 851.400 175.050 852.600 ;
        RECT 163.950 850.950 166.050 851.400 ;
        RECT 172.950 850.950 175.050 851.400 ;
        RECT 265.950 852.600 268.050 853.050 ;
        RECT 298.950 852.600 301.050 853.050 ;
        RECT 265.950 851.400 301.050 852.600 ;
        RECT 265.950 850.950 268.050 851.400 ;
        RECT 298.950 850.950 301.050 851.400 ;
        RECT 661.950 852.600 664.050 853.050 ;
        RECT 682.950 852.600 685.050 853.050 ;
        RECT 661.950 851.400 685.050 852.600 ;
        RECT 661.950 850.950 664.050 851.400 ;
        RECT 682.950 850.950 685.050 851.400 ;
        RECT 721.950 852.600 724.050 853.050 ;
        RECT 739.950 852.600 742.050 853.050 ;
        RECT 721.950 851.400 742.050 852.600 ;
        RECT 721.950 850.950 724.050 851.400 ;
        RECT 739.950 850.950 742.050 851.400 ;
        RECT 841.950 852.600 844.050 853.050 ;
        RECT 856.950 852.600 859.050 853.050 ;
        RECT 889.950 852.600 892.050 853.050 ;
        RECT 841.950 851.400 892.050 852.600 ;
        RECT 841.950 850.950 844.050 851.400 ;
        RECT 856.950 850.950 859.050 851.400 ;
        RECT 889.950 850.950 892.050 851.400 ;
        RECT 31.950 849.600 34.050 850.050 ;
        RECT 40.950 849.600 43.050 850.050 ;
        RECT 31.950 848.400 43.050 849.600 ;
        RECT 31.950 847.950 34.050 848.400 ;
        RECT 40.950 847.950 43.050 848.400 ;
        RECT 127.950 849.600 130.050 850.050 ;
        RECT 187.950 849.600 190.050 850.050 ;
        RECT 127.950 848.400 190.050 849.600 ;
        RECT 127.950 847.950 130.050 848.400 ;
        RECT 187.950 847.950 190.050 848.400 ;
        RECT 364.950 849.600 367.050 850.050 ;
        RECT 403.950 849.600 406.050 850.050 ;
        RECT 364.950 848.400 406.050 849.600 ;
        RECT 364.950 847.950 367.050 848.400 ;
        RECT 403.950 847.950 406.050 848.400 ;
        RECT 502.950 849.600 505.050 850.050 ;
        RECT 514.950 849.600 517.050 850.050 ;
        RECT 502.950 848.400 517.050 849.600 ;
        RECT 502.950 847.950 505.050 848.400 ;
        RECT 514.950 847.950 517.050 848.400 ;
        RECT 526.950 849.600 529.050 850.050 ;
        RECT 550.950 849.600 553.050 850.050 ;
        RECT 526.950 848.400 553.050 849.600 ;
        RECT 526.950 847.950 529.050 848.400 ;
        RECT 550.950 847.950 553.050 848.400 ;
        RECT 772.950 849.600 775.050 850.050 ;
        RECT 790.950 849.600 793.050 850.050 ;
        RECT 772.950 848.400 793.050 849.600 ;
        RECT 772.950 847.950 775.050 848.400 ;
        RECT 790.950 847.950 793.050 848.400 ;
        RECT 85.950 846.600 88.050 847.050 ;
        RECT 94.950 846.600 97.050 847.050 ;
        RECT 85.950 845.400 97.050 846.600 ;
        RECT 85.950 844.950 88.050 845.400 ;
        RECT 94.950 844.950 97.050 845.400 ;
        RECT 118.950 846.600 121.050 847.050 ;
        RECT 154.950 846.600 157.050 847.050 ;
        RECT 388.950 846.600 391.050 847.050 ;
        RECT 412.950 846.600 415.050 847.050 ;
        RECT 118.950 845.400 157.050 846.600 ;
        RECT 118.950 844.950 121.050 845.400 ;
        RECT 154.950 844.950 157.050 845.400 ;
        RECT 374.400 845.400 391.050 846.600 ;
        RECT 374.400 844.050 375.600 845.400 ;
        RECT 388.950 844.950 391.050 845.400 ;
        RECT 395.400 845.400 415.050 846.600 ;
        RECT 13.950 843.600 16.050 844.050 ;
        RECT 169.950 843.600 172.050 844.050 ;
        RECT 184.950 843.600 187.050 844.050 ;
        RECT 13.950 842.400 30.600 843.600 ;
        RECT 13.950 841.950 16.050 842.400 ;
        RECT 10.950 840.600 13.050 841.200 ;
        RECT 25.950 840.600 28.050 841.050 ;
        RECT 10.950 839.400 28.050 840.600 ;
        RECT 10.950 839.100 13.050 839.400 ;
        RECT 25.950 838.950 28.050 839.400 ;
        RECT 29.400 834.600 30.600 842.400 ;
        RECT 169.950 842.400 187.050 843.600 ;
        RECT 169.950 841.950 172.050 842.400 ;
        RECT 184.950 841.950 187.050 842.400 ;
        RECT 241.950 843.600 244.050 844.050 ;
        RECT 268.950 843.600 271.050 844.050 ;
        RECT 292.950 843.600 295.050 844.050 ;
        RECT 241.950 842.400 271.050 843.600 ;
        RECT 241.950 841.950 244.050 842.400 ;
        RECT 268.950 841.950 271.050 842.400 ;
        RECT 278.400 842.400 295.050 843.600 ;
        RECT 34.950 840.750 37.050 841.200 ;
        RECT 43.950 840.750 46.050 841.200 ;
        RECT 34.950 839.550 46.050 840.750 ;
        RECT 34.950 839.100 37.050 839.550 ;
        RECT 43.950 839.100 46.050 839.550 ;
        RECT 49.950 839.100 52.050 841.200 ;
        RECT 58.950 840.600 63.000 841.050 ;
        RECT 64.950 840.750 67.050 841.200 ;
        RECT 79.950 840.750 82.050 841.200 ;
        RECT 64.950 840.600 82.050 840.750 ;
        RECT 100.950 840.600 103.050 841.200 ;
        RECT 50.400 837.600 51.600 839.100 ;
        RECT 58.950 838.950 63.600 840.600 ;
        RECT 64.950 839.550 103.050 840.600 ;
        RECT 64.950 839.100 67.050 839.550 ;
        RECT 79.950 839.400 103.050 839.550 ;
        RECT 79.950 839.100 82.050 839.400 ;
        RECT 100.950 839.100 103.050 839.400 ;
        RECT 121.950 840.600 124.050 841.200 ;
        RECT 136.950 840.600 139.050 841.200 ;
        RECT 121.950 839.400 139.050 840.600 ;
        RECT 121.950 839.100 124.050 839.400 ;
        RECT 136.950 839.100 139.050 839.400 ;
        RECT 172.950 840.750 175.050 841.200 ;
        RECT 178.950 840.750 181.050 841.200 ;
        RECT 172.950 839.550 181.050 840.750 ;
        RECT 172.950 839.100 175.050 839.550 ;
        RECT 178.950 839.100 181.050 839.550 ;
        RECT 187.950 838.950 190.050 841.050 ;
        RECT 196.950 839.100 199.050 841.200 ;
        RECT 220.950 840.600 223.050 841.200 ;
        RECT 235.950 840.600 238.050 841.200 ;
        RECT 247.950 840.600 250.050 841.050 ;
        RECT 220.950 839.400 250.050 840.600 ;
        RECT 220.950 839.100 223.050 839.400 ;
        RECT 235.950 839.100 238.050 839.400 ;
        RECT 50.400 836.400 57.600 837.600 ;
        RECT 56.400 835.050 57.600 836.400 ;
        RECT 31.950 834.600 34.050 834.900 ;
        RECT 29.400 833.400 34.050 834.600 ;
        RECT 31.950 832.800 34.050 833.400 ;
        RECT 43.950 834.600 46.050 835.050 ;
        RECT 52.950 834.600 55.050 834.900 ;
        RECT 43.950 833.400 55.050 834.600 ;
        RECT 56.400 833.400 61.050 835.050 ;
        RECT 62.400 834.600 63.600 838.950 ;
        RECT 127.950 837.600 130.050 838.050 ;
        RECT 119.400 836.400 130.050 837.600 ;
        RECT 91.950 834.600 94.050 834.900 ;
        RECT 62.400 833.400 94.050 834.600 ;
        RECT 43.950 832.950 46.050 833.400 ;
        RECT 52.950 832.800 55.050 833.400 ;
        RECT 57.000 832.950 61.050 833.400 ;
        RECT 91.950 832.800 94.050 833.400 ;
        RECT 106.950 834.600 109.050 835.050 ;
        RECT 119.400 834.900 120.600 836.400 ;
        RECT 127.950 835.950 130.050 836.400 ;
        RECT 112.950 834.600 115.050 834.900 ;
        RECT 106.950 833.400 115.050 834.600 ;
        RECT 106.950 832.950 109.050 833.400 ;
        RECT 112.950 832.800 115.050 833.400 ;
        RECT 118.950 832.800 121.050 834.900 ;
        RECT 160.950 834.600 163.050 834.900 ;
        RECT 169.950 834.600 172.050 835.050 ;
        RECT 160.950 833.400 172.050 834.600 ;
        RECT 160.950 832.800 163.050 833.400 ;
        RECT 169.950 832.950 172.050 833.400 ;
        RECT 181.950 834.600 184.050 834.900 ;
        RECT 188.400 834.600 189.600 838.950 ;
        RECT 181.950 833.400 189.600 834.600 ;
        RECT 197.400 834.600 198.600 839.100 ;
        RECT 247.950 838.950 250.050 839.400 ;
        RECT 274.950 840.600 277.050 841.200 ;
        RECT 278.400 840.600 279.600 842.400 ;
        RECT 292.950 841.950 295.050 842.400 ;
        RECT 319.950 843.600 322.050 844.050 ;
        RECT 334.950 843.600 337.050 844.050 ;
        RECT 358.950 843.600 361.050 844.050 ;
        RECT 373.950 843.600 376.050 844.050 ;
        RECT 319.950 842.400 342.600 843.600 ;
        RECT 319.950 841.950 322.050 842.400 ;
        RECT 334.950 841.950 337.050 842.400 ;
        RECT 274.950 839.400 279.600 840.600 ;
        RECT 280.950 840.750 283.050 841.200 ;
        RECT 289.950 840.750 292.050 841.200 ;
        RECT 280.950 839.550 292.050 840.750 ;
        RECT 274.950 839.100 277.050 839.400 ;
        RECT 280.950 839.100 283.050 839.550 ;
        RECT 289.950 839.100 292.050 839.550 ;
        RECT 307.950 840.600 310.050 841.200 ;
        RECT 319.950 840.600 322.050 841.200 ;
        RECT 307.950 839.400 322.050 840.600 ;
        RECT 307.950 839.100 310.050 839.400 ;
        RECT 319.950 839.100 322.050 839.400 ;
        RECT 325.950 840.750 328.050 841.200 ;
        RECT 331.950 840.750 334.050 841.200 ;
        RECT 325.950 839.550 334.050 840.750 ;
        RECT 325.950 839.100 328.050 839.550 ;
        RECT 331.950 839.100 334.050 839.550 ;
        RECT 341.400 840.600 342.600 842.400 ;
        RECT 358.950 842.400 376.050 843.600 ;
        RECT 358.950 841.950 361.050 842.400 ;
        RECT 373.950 841.950 376.050 842.400 ;
        RECT 382.950 843.600 385.050 844.050 ;
        RECT 395.400 843.600 396.600 845.400 ;
        RECT 412.950 844.950 415.050 845.400 ;
        RECT 676.950 846.600 679.050 847.050 ;
        RECT 703.950 846.600 706.050 847.050 ;
        RECT 676.950 845.400 706.050 846.600 ;
        RECT 676.950 844.950 679.050 845.400 ;
        RECT 703.950 844.950 706.050 845.400 ;
        RECT 724.950 846.600 727.050 847.050 ;
        RECT 874.950 846.600 877.050 847.050 ;
        RECT 880.950 846.600 883.050 847.050 ;
        RECT 898.950 846.600 901.050 847.050 ;
        RECT 724.950 845.400 753.600 846.600 ;
        RECT 724.950 844.950 727.050 845.400 ;
        RECT 382.950 842.400 396.600 843.600 ;
        RECT 752.400 843.600 753.600 845.400 ;
        RECT 874.950 845.400 901.050 846.600 ;
        RECT 874.950 844.950 877.050 845.400 ;
        RECT 880.950 844.950 883.050 845.400 ;
        RECT 898.950 844.950 901.050 845.400 ;
        RECT 757.950 843.600 760.050 844.050 ;
        RECT 784.950 843.600 787.050 844.050 ;
        RECT 752.400 842.400 787.050 843.600 ;
        RECT 382.950 841.950 385.050 842.400 ;
        RECT 757.950 841.950 760.050 842.400 ;
        RECT 784.950 841.950 787.050 842.400 ;
        RECT 349.950 840.600 352.050 841.200 ;
        RECT 341.400 839.400 352.050 840.600 ;
        RECT 349.950 839.100 352.050 839.400 ;
        RECT 367.950 840.750 370.050 841.200 ;
        RECT 379.950 840.750 382.050 841.200 ;
        RECT 367.950 839.550 382.050 840.750 ;
        RECT 367.950 839.100 370.050 839.550 ;
        RECT 379.950 839.100 382.050 839.550 ;
        RECT 397.950 840.600 400.050 841.200 ;
        RECT 397.950 839.400 402.600 840.600 ;
        RECT 397.950 839.100 400.050 839.400 ;
        RECT 290.400 837.600 291.600 839.100 ;
        RECT 209.400 836.400 291.600 837.600 ;
        RECT 209.400 834.600 210.600 836.400 ;
        RECT 401.400 835.050 402.600 839.400 ;
        RECT 409.950 837.600 412.050 841.050 ;
        RECT 418.950 839.100 421.050 841.200 ;
        RECT 442.950 840.750 445.050 841.200 ;
        RECT 448.950 840.750 451.050 841.200 ;
        RECT 442.950 839.550 451.050 840.750 ;
        RECT 442.950 839.100 445.050 839.550 ;
        RECT 448.950 839.100 451.050 839.550 ;
        RECT 475.950 840.750 478.050 841.200 ;
        RECT 490.950 840.750 493.050 841.050 ;
        RECT 499.950 840.750 502.050 841.200 ;
        RECT 475.950 839.550 502.050 840.750 ;
        RECT 475.950 839.100 478.050 839.550 ;
        RECT 409.950 837.000 417.600 837.600 ;
        RECT 410.400 836.400 417.600 837.000 ;
        RECT 197.400 833.400 210.600 834.600 ;
        RECT 229.950 834.600 232.050 835.050 ;
        RECT 238.950 834.600 241.050 834.900 ;
        RECT 229.950 833.400 241.050 834.600 ;
        RECT 181.950 832.800 184.050 833.400 ;
        RECT 229.950 832.950 232.050 833.400 ;
        RECT 238.950 832.800 241.050 833.400 ;
        RECT 247.950 834.450 250.050 834.900 ;
        RECT 256.950 834.450 259.050 834.900 ;
        RECT 247.950 833.250 259.050 834.450 ;
        RECT 247.950 832.800 250.050 833.250 ;
        RECT 256.950 832.800 259.050 833.250 ;
        RECT 277.950 834.600 280.050 834.900 ;
        RECT 286.950 834.600 289.050 835.050 ;
        RECT 277.950 833.400 289.050 834.600 ;
        RECT 277.950 832.800 280.050 833.400 ;
        RECT 286.950 832.950 289.050 833.400 ;
        RECT 322.950 834.600 325.050 834.900 ;
        RECT 337.950 834.600 340.050 835.050 ;
        RECT 322.950 833.400 340.050 834.600 ;
        RECT 322.950 832.800 325.050 833.400 ;
        RECT 337.950 832.950 340.050 833.400 ;
        RECT 400.950 832.950 403.050 835.050 ;
        RECT 416.400 834.900 417.600 836.400 ;
        RECT 415.950 832.800 418.050 834.900 ;
        RECT 419.400 832.050 420.600 839.100 ;
        RECT 490.950 838.950 493.050 839.550 ;
        RECT 499.950 839.100 502.050 839.550 ;
        RECT 520.950 839.100 523.050 841.200 ;
        RECT 532.950 839.100 535.050 841.200 ;
        RECT 553.950 839.100 556.050 841.200 ;
        RECT 589.950 839.100 592.050 841.200 ;
        RECT 613.950 840.750 616.050 841.200 ;
        RECT 619.950 840.750 622.050 841.200 ;
        RECT 613.950 839.550 622.050 840.750 ;
        RECT 613.950 839.100 616.050 839.550 ;
        RECT 619.950 839.100 622.050 839.550 ;
        RECT 628.950 839.100 631.050 841.200 ;
        RECT 640.950 840.750 643.050 841.200 ;
        RECT 646.950 840.750 649.050 841.200 ;
        RECT 640.950 839.550 649.050 840.750 ;
        RECT 640.950 839.100 643.050 839.550 ;
        RECT 646.950 839.100 649.050 839.550 ;
        RECT 652.950 839.100 655.050 841.200 ;
        RECT 664.950 840.750 667.050 841.200 ;
        RECT 670.950 840.750 673.050 841.200 ;
        RECT 664.950 839.550 673.050 840.750 ;
        RECT 664.950 839.100 667.050 839.550 ;
        RECT 670.950 839.100 673.050 839.550 ;
        RECT 694.950 839.100 697.050 841.200 ;
        RECT 715.950 840.600 718.050 841.200 ;
        RECT 713.400 839.400 718.050 840.600 ;
        RECT 481.950 834.600 484.050 834.900 ;
        RECT 496.950 834.600 499.050 834.900 ;
        RECT 521.400 834.600 522.600 839.100 ;
        RECT 533.400 837.600 534.600 839.100 ;
        RECT 554.400 837.600 555.600 839.100 ;
        RECT 533.400 837.000 537.600 837.600 ;
        RECT 545.400 837.000 555.600 837.600 ;
        RECT 533.400 836.400 538.050 837.000 ;
        RECT 481.950 833.400 495.600 834.600 ;
        RECT 481.950 832.800 484.050 833.400 ;
        RECT 70.950 831.600 73.050 832.050 ;
        RECT 79.950 831.600 82.050 832.050 ;
        RECT 70.950 830.400 82.050 831.600 ;
        RECT 70.950 829.950 73.050 830.400 ;
        RECT 79.950 829.950 82.050 830.400 ;
        RECT 292.950 831.600 295.050 832.050 ;
        RECT 316.950 831.600 319.050 832.050 ;
        RECT 292.950 830.400 319.050 831.600 ;
        RECT 292.950 829.950 295.050 830.400 ;
        RECT 316.950 829.950 319.050 830.400 ;
        RECT 346.950 831.600 349.050 832.050 ;
        RECT 358.950 831.600 361.050 832.050 ;
        RECT 346.950 830.400 361.050 831.600 ;
        RECT 346.950 829.950 349.050 830.400 ;
        RECT 358.950 829.950 361.050 830.400 ;
        RECT 418.950 829.950 421.050 832.050 ;
        RECT 430.950 831.600 433.050 832.050 ;
        RECT 442.950 831.600 445.050 832.050 ;
        RECT 430.950 830.400 445.050 831.600 ;
        RECT 494.400 831.600 495.600 833.400 ;
        RECT 496.950 833.400 522.600 834.600 ;
        RECT 496.950 832.800 499.050 833.400 ;
        RECT 535.950 832.950 538.050 836.400 ;
        RECT 544.950 836.400 555.600 837.000 ;
        RECT 544.950 832.950 547.050 836.400 ;
        RECT 590.400 835.050 591.600 839.100 ;
        RECT 550.950 834.600 553.050 834.900 ;
        RECT 577.800 834.600 579.900 835.050 ;
        RECT 550.950 833.400 579.900 834.600 ;
        RECT 590.400 833.400 595.050 835.050 ;
        RECT 629.400 834.600 630.600 839.100 ;
        RECT 649.950 834.600 652.050 834.900 ;
        RECT 629.400 833.400 652.050 834.600 ;
        RECT 653.400 834.600 654.600 839.100 ;
        RECT 695.400 835.050 696.600 839.100 ;
        RECT 673.950 834.600 676.050 834.900 ;
        RECT 653.400 833.400 676.050 834.600 ;
        RECT 695.400 833.400 700.050 835.050 ;
        RECT 550.950 832.800 553.050 833.400 ;
        RECT 577.800 832.950 579.900 833.400 ;
        RECT 591.000 832.950 595.050 833.400 ;
        RECT 649.950 832.800 652.050 833.400 ;
        RECT 673.950 832.800 676.050 833.400 ;
        RECT 696.000 832.950 700.050 833.400 ;
        RECT 514.950 831.600 517.050 832.050 ;
        RECT 532.950 831.600 535.050 832.050 ;
        RECT 494.400 830.400 517.050 831.600 ;
        RECT 430.950 829.950 433.050 830.400 ;
        RECT 442.950 829.950 445.050 830.400 ;
        RECT 514.950 829.950 517.050 830.400 ;
        RECT 521.400 830.400 535.050 831.600 ;
        RECT 4.950 828.600 7.050 829.050 ;
        RECT 19.950 828.600 22.050 829.050 ;
        RECT 4.950 827.400 22.050 828.600 ;
        RECT 4.950 826.950 7.050 827.400 ;
        RECT 19.950 826.950 22.050 827.400 ;
        RECT 130.950 828.600 133.050 829.050 ;
        RECT 139.950 828.600 142.050 829.050 ;
        RECT 199.950 828.600 202.050 829.050 ;
        RECT 208.950 828.600 211.050 829.050 ;
        RECT 130.950 827.400 211.050 828.600 ;
        RECT 130.950 826.950 133.050 827.400 ;
        RECT 139.950 826.950 142.050 827.400 ;
        RECT 199.950 826.950 202.050 827.400 ;
        RECT 208.950 826.950 211.050 827.400 ;
        RECT 223.950 828.600 226.050 829.050 ;
        RECT 253.950 828.600 256.050 829.050 ;
        RECT 223.950 827.400 256.050 828.600 ;
        RECT 223.950 826.950 226.050 827.400 ;
        RECT 253.950 826.950 256.050 827.400 ;
        RECT 322.950 828.600 325.050 829.050 ;
        RECT 334.950 828.600 337.050 829.050 ;
        RECT 322.950 827.400 337.050 828.600 ;
        RECT 322.950 826.950 325.050 827.400 ;
        RECT 334.950 826.950 337.050 827.400 ;
        RECT 340.950 828.600 343.050 829.050 ;
        RECT 346.950 828.600 349.050 828.900 ;
        RECT 352.950 828.600 355.050 829.050 ;
        RECT 340.950 827.400 355.050 828.600 ;
        RECT 340.950 826.950 343.050 827.400 ;
        RECT 346.950 826.800 349.050 827.400 ;
        RECT 352.950 826.950 355.050 827.400 ;
        RECT 451.950 828.600 454.050 829.050 ;
        RECT 457.950 828.600 460.050 829.050 ;
        RECT 451.950 827.400 460.050 828.600 ;
        RECT 451.950 826.950 454.050 827.400 ;
        RECT 457.950 826.950 460.050 827.400 ;
        RECT 499.950 828.600 502.050 829.050 ;
        RECT 521.400 828.600 522.600 830.400 ;
        RECT 532.950 829.950 535.050 830.400 ;
        RECT 625.950 831.600 628.050 832.050 ;
        RECT 637.950 831.600 640.050 832.050 ;
        RECT 625.950 830.400 640.050 831.600 ;
        RECT 625.950 829.950 628.050 830.400 ;
        RECT 637.950 829.950 640.050 830.400 ;
        RECT 691.950 831.600 694.050 832.050 ;
        RECT 713.400 831.600 714.600 839.400 ;
        RECT 715.950 839.100 718.050 839.400 ;
        RECT 736.950 838.950 739.050 841.050 ;
        RECT 772.950 840.600 775.050 841.050 ;
        RECT 755.400 839.400 775.050 840.600 ;
        RECT 737.400 837.600 738.600 838.950 ;
        RECT 755.400 837.600 756.600 839.400 ;
        RECT 772.950 838.950 775.050 839.400 ;
        RECT 790.950 840.600 793.050 841.050 ;
        RECT 826.950 840.600 829.050 841.050 ;
        RECT 835.950 840.600 838.050 841.200 ;
        RECT 840.000 840.600 844.050 841.050 ;
        RECT 790.950 839.400 810.600 840.600 ;
        RECT 790.950 838.950 793.050 839.400 ;
        RECT 722.400 837.000 756.600 837.600 ;
        RECT 721.950 836.400 756.600 837.000 ;
        RECT 809.400 837.600 810.600 839.400 ;
        RECT 826.950 839.400 838.050 840.600 ;
        RECT 826.950 838.950 829.050 839.400 ;
        RECT 835.950 839.100 838.050 839.400 ;
        RECT 839.400 838.950 844.050 840.600 ;
        RECT 850.950 838.950 853.050 841.050 ;
        RECT 862.950 839.100 865.050 841.200 ;
        RECT 874.950 840.600 877.050 841.200 ;
        RECT 872.400 839.400 877.050 840.600 ;
        RECT 809.400 836.400 813.600 837.600 ;
        RECT 721.950 832.950 724.050 836.400 ;
        RECT 739.950 834.600 742.050 834.900 ;
        RECT 760.950 834.600 763.050 834.900 ;
        RECT 739.950 833.400 763.050 834.600 ;
        RECT 739.950 832.800 742.050 833.400 ;
        RECT 760.950 832.800 763.050 833.400 ;
        RECT 766.950 834.450 769.050 834.900 ;
        RECT 781.950 834.450 784.050 834.900 ;
        RECT 766.950 833.250 784.050 834.450 ;
        RECT 812.400 834.600 813.600 836.400 ;
        RECT 839.400 834.900 840.600 838.950 ;
        RECT 851.400 835.050 852.600 838.950 ;
        RECT 823.950 834.600 826.050 834.900 ;
        RECT 812.400 833.400 826.050 834.600 ;
        RECT 766.950 832.800 769.050 833.250 ;
        RECT 781.950 832.800 784.050 833.250 ;
        RECT 823.950 832.800 826.050 833.400 ;
        RECT 838.950 832.800 841.050 834.900 ;
        RECT 850.950 832.950 853.050 835.050 ;
        RECT 863.400 834.600 864.600 839.100 ;
        RECT 868.950 834.600 871.050 835.050 ;
        RECT 863.400 833.400 871.050 834.600 ;
        RECT 868.950 832.950 871.050 833.400 ;
        RECT 691.950 830.400 714.600 831.600 ;
        RECT 826.950 831.600 829.050 832.050 ;
        RECT 835.950 831.600 838.050 832.050 ;
        RECT 826.950 830.400 838.050 831.600 ;
        RECT 691.950 829.950 694.050 830.400 ;
        RECT 826.950 829.950 829.050 830.400 ;
        RECT 835.950 829.950 838.050 830.400 ;
        RECT 859.950 831.600 862.050 832.050 ;
        RECT 872.400 831.600 873.600 839.400 ;
        RECT 874.950 839.100 877.050 839.400 ;
        RECT 877.950 834.600 880.050 834.900 ;
        RECT 889.950 834.600 892.050 835.050 ;
        RECT 877.950 833.400 892.050 834.600 ;
        RECT 877.950 832.800 880.050 833.400 ;
        RECT 889.950 832.950 892.050 833.400 ;
        RECT 859.950 830.400 873.600 831.600 ;
        RECT 859.950 829.950 862.050 830.400 ;
        RECT 499.950 827.400 522.600 828.600 ;
        RECT 547.950 828.600 550.050 829.050 ;
        RECT 577.950 828.600 580.050 829.050 ;
        RECT 547.950 827.400 580.050 828.600 ;
        RECT 499.950 826.950 502.050 827.400 ;
        RECT 547.950 826.950 550.050 827.400 ;
        RECT 577.950 826.950 580.050 827.400 ;
        RECT 598.950 828.600 601.050 829.050 ;
        RECT 604.950 828.600 607.050 829.050 ;
        RECT 598.950 827.400 607.050 828.600 ;
        RECT 598.950 826.950 601.050 827.400 ;
        RECT 604.950 826.950 607.050 827.400 ;
        RECT 610.950 828.600 613.050 829.050 ;
        RECT 655.950 828.600 658.050 829.050 ;
        RECT 664.950 828.600 667.050 829.050 ;
        RECT 688.950 828.600 691.050 829.050 ;
        RECT 610.950 827.400 691.050 828.600 ;
        RECT 610.950 826.950 613.050 827.400 ;
        RECT 655.950 826.950 658.050 827.400 ;
        RECT 664.950 826.950 667.050 827.400 ;
        RECT 688.950 826.950 691.050 827.400 ;
        RECT 694.950 828.600 697.050 829.050 ;
        RECT 724.950 828.600 727.050 829.050 ;
        RECT 694.950 827.400 727.050 828.600 ;
        RECT 694.950 826.950 697.050 827.400 ;
        RECT 724.950 826.950 727.050 827.400 ;
        RECT 754.950 828.600 757.050 829.050 ;
        RECT 778.950 828.600 781.050 828.900 ;
        RECT 754.950 827.400 781.050 828.600 ;
        RECT 754.950 826.950 757.050 827.400 ;
        RECT 778.950 826.800 781.050 827.400 ;
        RECT 814.950 828.600 817.050 829.050 ;
        RECT 874.950 828.600 877.050 829.050 ;
        RECT 814.950 827.400 877.050 828.600 ;
        RECT 814.950 826.950 817.050 827.400 ;
        RECT 874.950 826.950 877.050 827.400 ;
        RECT 217.950 825.600 220.050 826.050 ;
        RECT 244.950 825.600 247.050 826.050 ;
        RECT 217.950 824.400 247.050 825.600 ;
        RECT 217.950 823.950 220.050 824.400 ;
        RECT 244.950 823.950 247.050 824.400 ;
        RECT 256.950 825.600 259.050 826.050 ;
        RECT 283.950 825.600 286.050 826.050 ;
        RECT 256.950 824.400 286.050 825.600 ;
        RECT 256.950 823.950 259.050 824.400 ;
        RECT 283.950 823.950 286.050 824.400 ;
        RECT 289.950 825.600 292.050 826.050 ;
        RECT 319.950 825.600 322.050 826.050 ;
        RECT 289.950 824.400 322.050 825.600 ;
        RECT 289.950 823.950 292.050 824.400 ;
        RECT 319.950 823.950 322.050 824.400 ;
        RECT 328.950 825.600 331.050 826.050 ;
        RECT 337.950 825.600 340.050 826.050 ;
        RECT 358.950 825.600 361.050 826.050 ;
        RECT 328.950 824.400 361.050 825.600 ;
        RECT 328.950 823.950 331.050 824.400 ;
        RECT 337.950 823.950 340.050 824.400 ;
        RECT 358.950 823.950 361.050 824.400 ;
        RECT 391.950 825.600 394.050 826.050 ;
        RECT 439.950 825.600 442.050 826.050 ;
        RECT 391.950 824.400 442.050 825.600 ;
        RECT 391.950 823.950 394.050 824.400 ;
        RECT 439.950 823.950 442.050 824.400 ;
        RECT 475.950 825.600 478.050 826.050 ;
        RECT 520.800 825.600 522.900 826.050 ;
        RECT 475.950 824.400 522.900 825.600 ;
        RECT 475.950 823.950 478.050 824.400 ;
        RECT 520.800 823.950 522.900 824.400 ;
        RECT 523.950 825.600 526.050 826.050 ;
        RECT 544.950 825.600 547.050 825.900 ;
        RECT 523.950 824.400 547.050 825.600 ;
        RECT 523.950 823.950 526.050 824.400 ;
        RECT 544.950 823.800 547.050 824.400 ;
        RECT 703.950 825.600 706.050 826.050 ;
        RECT 715.800 825.600 717.900 826.050 ;
        RECT 703.950 824.400 717.900 825.600 ;
        RECT 703.950 823.950 706.050 824.400 ;
        RECT 715.800 823.950 717.900 824.400 ;
        RECT 718.950 825.600 721.050 826.050 ;
        RECT 727.950 825.600 730.050 826.050 ;
        RECT 718.950 824.400 730.050 825.600 ;
        RECT 718.950 823.950 721.050 824.400 ;
        RECT 727.950 823.950 730.050 824.400 ;
        RECT 796.950 825.600 799.050 826.050 ;
        RECT 811.950 825.600 814.050 826.050 ;
        RECT 796.950 824.400 814.050 825.600 ;
        RECT 796.950 823.950 799.050 824.400 ;
        RECT 811.950 823.950 814.050 824.400 ;
        RECT 13.950 822.600 16.050 823.050 ;
        RECT 19.950 822.600 22.050 823.050 ;
        RECT 13.950 821.400 22.050 822.600 ;
        RECT 13.950 820.950 16.050 821.400 ;
        RECT 19.950 820.950 22.050 821.400 ;
        RECT 52.950 822.600 55.050 823.050 ;
        RECT 58.950 822.600 61.050 823.050 ;
        RECT 67.950 822.600 70.050 823.050 ;
        RECT 97.950 822.600 100.050 823.050 ;
        RECT 52.950 821.400 100.050 822.600 ;
        RECT 52.950 820.950 55.050 821.400 ;
        RECT 58.950 820.950 61.050 821.400 ;
        RECT 67.950 820.950 70.050 821.400 ;
        RECT 97.950 820.950 100.050 821.400 ;
        RECT 253.950 822.600 256.050 823.050 ;
        RECT 364.950 822.600 367.050 823.050 ;
        RECT 253.950 821.400 367.050 822.600 ;
        RECT 253.950 820.950 256.050 821.400 ;
        RECT 364.950 820.950 367.050 821.400 ;
        RECT 502.950 822.600 505.050 823.050 ;
        RECT 508.950 822.600 511.050 823.050 ;
        RECT 502.950 821.400 511.050 822.600 ;
        RECT 502.950 820.950 505.050 821.400 ;
        RECT 508.950 820.950 511.050 821.400 ;
        RECT 523.950 822.600 526.050 822.900 ;
        RECT 535.950 822.600 538.050 823.050 ;
        RECT 565.950 822.600 568.050 823.050 ;
        RECT 523.950 821.400 568.050 822.600 ;
        RECT 28.950 819.600 31.050 820.050 ;
        RECT 43.950 819.600 46.050 820.050 ;
        RECT 28.950 818.400 46.050 819.600 ;
        RECT 28.950 817.950 31.050 818.400 ;
        RECT 43.950 817.950 46.050 818.400 ;
        RECT 202.950 819.600 205.050 820.050 ;
        RECT 217.800 819.600 219.900 820.050 ;
        RECT 202.950 818.400 219.900 819.600 ;
        RECT 202.950 817.950 205.050 818.400 ;
        RECT 217.800 817.950 219.900 818.400 ;
        RECT 220.950 819.600 223.050 820.050 ;
        RECT 292.800 819.600 294.900 820.050 ;
        RECT 220.950 818.400 294.900 819.600 ;
        RECT 220.950 817.950 223.050 818.400 ;
        RECT 292.800 817.950 294.900 818.400 ;
        RECT 295.950 819.600 298.050 820.050 ;
        RECT 346.950 819.600 349.050 820.050 ;
        RECT 295.950 818.400 349.050 819.600 ;
        RECT 295.950 817.950 298.050 818.400 ;
        RECT 346.950 817.950 349.050 818.400 ;
        RECT 397.950 819.600 400.050 820.050 ;
        RECT 430.950 819.600 433.050 820.050 ;
        RECT 448.950 819.600 451.050 820.050 ;
        RECT 454.950 819.600 457.050 820.050 ;
        RECT 397.950 818.400 420.600 819.600 ;
        RECT 397.950 817.950 400.050 818.400 ;
        RECT 7.950 816.600 10.050 817.050 ;
        RECT 37.950 816.600 40.050 817.050 ;
        RECT 7.950 815.400 40.050 816.600 ;
        RECT 7.950 814.950 10.050 815.400 ;
        RECT 37.950 814.950 40.050 815.400 ;
        RECT 148.950 816.600 151.050 817.050 ;
        RECT 166.950 816.600 169.050 817.050 ;
        RECT 148.950 815.400 169.050 816.600 ;
        RECT 148.950 814.950 151.050 815.400 ;
        RECT 166.950 814.950 169.050 815.400 ;
        RECT 301.950 816.600 304.050 817.050 ;
        RECT 331.950 816.600 334.050 817.050 ;
        RECT 301.950 815.400 334.050 816.600 ;
        RECT 419.400 816.600 420.600 818.400 ;
        RECT 430.950 818.400 457.050 819.600 ;
        RECT 430.950 817.950 433.050 818.400 ;
        RECT 448.950 817.950 451.050 818.400 ;
        RECT 454.950 817.950 457.050 818.400 ;
        RECT 460.950 819.600 463.050 820.050 ;
        RECT 502.950 819.600 505.050 819.900 ;
        RECT 460.950 818.400 505.050 819.600 ;
        RECT 509.400 819.600 510.600 820.950 ;
        RECT 523.950 820.800 526.050 821.400 ;
        RECT 535.950 820.950 538.050 821.400 ;
        RECT 565.950 820.950 568.050 821.400 ;
        RECT 586.950 822.600 589.050 823.050 ;
        RECT 622.950 822.600 625.050 823.050 ;
        RECT 586.950 821.400 625.050 822.600 ;
        RECT 586.950 820.950 589.050 821.400 ;
        RECT 622.950 820.950 625.050 821.400 ;
        RECT 631.950 822.600 634.050 823.050 ;
        RECT 694.950 822.600 697.050 823.050 ;
        RECT 631.950 821.400 697.050 822.600 ;
        RECT 631.950 820.950 634.050 821.400 ;
        RECT 694.950 820.950 697.050 821.400 ;
        RECT 700.950 822.600 703.050 823.050 ;
        RECT 736.950 822.600 739.050 823.050 ;
        RECT 700.950 821.400 739.050 822.600 ;
        RECT 700.950 820.950 703.050 821.400 ;
        RECT 736.950 820.950 739.050 821.400 ;
        RECT 778.950 822.600 781.050 823.050 ;
        RECT 898.950 822.600 901.050 823.050 ;
        RECT 913.950 822.600 916.050 823.050 ;
        RECT 778.950 821.400 825.600 822.600 ;
        RECT 778.950 820.950 781.050 821.400 ;
        RECT 824.400 820.050 825.600 821.400 ;
        RECT 898.950 821.400 916.050 822.600 ;
        RECT 898.950 820.950 901.050 821.400 ;
        RECT 913.950 820.950 916.050 821.400 ;
        RECT 529.950 819.600 532.050 820.050 ;
        RECT 538.950 819.600 541.050 820.050 ;
        RECT 509.400 818.400 541.050 819.600 ;
        RECT 460.950 817.950 463.050 818.400 ;
        RECT 502.950 817.800 505.050 818.400 ;
        RECT 529.950 817.950 532.050 818.400 ;
        RECT 538.950 817.950 541.050 818.400 ;
        RECT 559.950 819.600 562.050 820.050 ;
        RECT 583.950 819.600 586.050 820.050 ;
        RECT 559.950 818.400 586.050 819.600 ;
        RECT 559.950 817.950 562.050 818.400 ;
        RECT 583.950 817.950 586.050 818.400 ;
        RECT 715.950 819.600 718.050 820.050 ;
        RECT 727.800 819.600 729.900 820.050 ;
        RECT 715.950 818.400 729.900 819.600 ;
        RECT 715.950 817.950 718.050 818.400 ;
        RECT 727.800 817.950 729.900 818.400 ;
        RECT 730.950 819.600 733.050 820.050 ;
        RECT 760.950 819.600 763.050 820.050 ;
        RECT 730.950 818.400 763.050 819.600 ;
        RECT 730.950 817.950 733.050 818.400 ;
        RECT 760.950 817.950 763.050 818.400 ;
        RECT 823.950 819.600 826.050 820.050 ;
        RECT 871.950 819.600 874.050 820.050 ;
        RECT 823.950 818.400 874.050 819.600 ;
        RECT 823.950 817.950 826.050 818.400 ;
        RECT 871.950 817.950 874.050 818.400 ;
        RECT 427.950 816.600 430.050 817.050 ;
        RECT 419.400 815.400 430.050 816.600 ;
        RECT 301.950 814.950 304.050 815.400 ;
        RECT 331.950 814.950 334.050 815.400 ;
        RECT 427.950 814.950 430.050 815.400 ;
        RECT 481.950 816.600 484.050 817.050 ;
        RECT 490.950 816.600 493.050 817.050 ;
        RECT 481.950 815.400 493.050 816.600 ;
        RECT 481.950 814.950 484.050 815.400 ;
        RECT 490.950 814.950 493.050 815.400 ;
        RECT 544.950 816.600 547.050 817.050 ;
        RECT 589.950 816.600 592.050 817.050 ;
        RECT 544.950 815.400 592.050 816.600 ;
        RECT 544.950 814.950 547.050 815.400 ;
        RECT 589.950 814.950 592.050 815.400 ;
        RECT 595.950 816.600 598.050 817.050 ;
        RECT 610.950 816.600 613.050 817.050 ;
        RECT 658.950 816.600 661.050 817.050 ;
        RECT 595.950 815.400 613.050 816.600 ;
        RECT 595.950 814.950 598.050 815.400 ;
        RECT 610.950 814.950 613.050 815.400 ;
        RECT 632.400 815.400 661.050 816.600 ;
        RECT 43.950 813.600 46.050 814.050 ;
        RECT 61.950 813.600 64.050 814.050 ;
        RECT 43.950 812.400 64.050 813.600 ;
        RECT 43.950 811.950 46.050 812.400 ;
        RECT 61.950 811.950 64.050 812.400 ;
        RECT 82.950 813.600 85.050 814.050 ;
        RECT 112.950 813.600 115.050 814.050 ;
        RECT 124.950 813.600 127.050 814.050 ;
        RECT 82.950 812.400 127.050 813.600 ;
        RECT 82.950 811.950 85.050 812.400 ;
        RECT 112.950 811.950 115.050 812.400 ;
        RECT 124.950 811.950 127.050 812.400 ;
        RECT 136.950 813.600 139.050 814.050 ;
        RECT 175.950 813.600 178.050 814.050 ;
        RECT 136.950 812.400 178.050 813.600 ;
        RECT 136.950 811.950 139.050 812.400 ;
        RECT 175.950 811.950 178.050 812.400 ;
        RECT 262.950 813.600 265.050 814.050 ;
        RECT 268.950 813.600 271.050 814.050 ;
        RECT 262.950 812.400 271.050 813.600 ;
        RECT 262.950 811.950 265.050 812.400 ;
        RECT 268.950 811.950 271.050 812.400 ;
        RECT 340.950 813.600 343.050 814.050 ;
        RECT 352.950 813.600 355.050 814.050 ;
        RECT 340.950 812.400 355.050 813.600 ;
        RECT 340.950 811.950 343.050 812.400 ;
        RECT 352.950 811.950 355.050 812.400 ;
        RECT 388.950 813.600 391.050 814.050 ;
        RECT 406.950 813.600 409.050 814.050 ;
        RECT 388.950 812.400 409.050 813.600 ;
        RECT 388.950 811.950 391.050 812.400 ;
        RECT 406.950 811.950 409.050 812.400 ;
        RECT 478.950 813.600 481.050 814.050 ;
        RECT 529.950 813.600 532.050 814.050 ;
        RECT 478.950 812.400 532.050 813.600 ;
        RECT 478.950 811.950 481.050 812.400 ;
        RECT 529.950 811.950 532.050 812.400 ;
        RECT 613.950 813.600 616.050 814.050 ;
        RECT 632.400 813.600 633.600 815.400 ;
        RECT 658.950 814.950 661.050 815.400 ;
        RECT 613.950 812.400 633.600 813.600 ;
        RECT 661.950 813.600 664.050 814.050 ;
        RECT 691.950 813.600 694.050 814.050 ;
        RECT 661.950 812.400 694.050 813.600 ;
        RECT 613.950 811.950 616.050 812.400 ;
        RECT 661.950 811.950 664.050 812.400 ;
        RECT 691.950 811.950 694.050 812.400 ;
        RECT 712.950 813.600 715.050 814.050 ;
        RECT 724.800 813.600 726.900 814.050 ;
        RECT 712.950 812.400 726.900 813.600 ;
        RECT 712.950 811.950 715.050 812.400 ;
        RECT 724.800 811.950 726.900 812.400 ;
        RECT 727.950 813.600 730.050 814.050 ;
        RECT 751.950 813.600 754.050 814.050 ;
        RECT 727.950 812.400 754.050 813.600 ;
        RECT 727.950 811.950 730.050 812.400 ;
        RECT 751.950 811.950 754.050 812.400 ;
        RECT 802.950 813.600 805.050 814.050 ;
        RECT 829.950 813.600 832.050 814.050 ;
        RECT 802.950 812.400 832.050 813.600 ;
        RECT 802.950 811.950 805.050 812.400 ;
        RECT 829.950 811.950 832.050 812.400 ;
        RECT 844.950 813.600 847.050 814.050 ;
        RECT 853.950 813.600 856.050 814.050 ;
        RECT 844.950 812.400 856.050 813.600 ;
        RECT 844.950 811.950 847.050 812.400 ;
        RECT 853.950 811.950 856.050 812.400 ;
        RECT 859.950 813.600 862.050 814.050 ;
        RECT 892.950 813.600 895.050 814.050 ;
        RECT 859.950 812.400 895.050 813.600 ;
        RECT 859.950 811.950 862.050 812.400 ;
        RECT 892.950 811.950 895.050 812.400 ;
        RECT 31.950 810.600 34.050 811.050 ;
        RECT 40.950 810.600 43.050 811.050 ;
        RECT 31.950 809.400 43.050 810.600 ;
        RECT 31.950 808.950 34.050 809.400 ;
        RECT 40.950 808.950 43.050 809.400 ;
        RECT 85.950 810.600 88.050 811.050 ;
        RECT 91.950 810.600 94.050 811.050 ;
        RECT 100.950 810.600 103.050 811.050 ;
        RECT 85.950 809.400 103.050 810.600 ;
        RECT 85.950 808.950 88.050 809.400 ;
        RECT 91.950 808.950 94.050 809.400 ;
        RECT 100.950 808.950 103.050 809.400 ;
        RECT 379.950 810.600 382.050 811.050 ;
        RECT 391.950 810.600 394.050 811.050 ;
        RECT 379.950 809.400 394.050 810.600 ;
        RECT 379.950 808.950 382.050 809.400 ;
        RECT 391.950 808.950 394.050 809.400 ;
        RECT 400.950 808.950 403.050 811.050 ;
        RECT 469.950 810.600 472.050 811.050 ;
        RECT 475.950 810.600 478.050 811.050 ;
        RECT 469.950 809.400 478.050 810.600 ;
        RECT 469.950 808.950 472.050 809.400 ;
        RECT 475.950 808.950 478.050 809.400 ;
        RECT 493.950 810.600 496.050 811.050 ;
        RECT 505.950 810.600 508.050 811.050 ;
        RECT 493.950 809.400 508.050 810.600 ;
        RECT 493.950 808.950 496.050 809.400 ;
        RECT 505.950 808.950 508.050 809.400 ;
        RECT 511.950 810.600 516.000 811.050 ;
        RECT 511.950 808.950 516.600 810.600 ;
        RECT 523.950 808.950 526.050 811.050 ;
        RECT 790.950 810.600 793.050 811.050 ;
        RECT 808.950 810.600 811.050 811.050 ;
        RECT 790.950 809.400 811.050 810.600 ;
        RECT 790.950 808.950 793.050 809.400 ;
        RECT 808.950 808.950 811.050 809.400 ;
        RECT 862.950 810.600 865.050 811.050 ;
        RECT 868.950 810.600 871.050 811.050 ;
        RECT 862.950 809.400 871.050 810.600 ;
        RECT 862.950 808.950 865.050 809.400 ;
        RECT 868.950 808.950 871.050 809.400 ;
        RECT 1.950 807.750 4.050 808.200 ;
        RECT 19.950 807.750 22.050 808.200 ;
        RECT 1.950 806.550 22.050 807.750 ;
        RECT 76.950 807.600 79.050 808.200 ;
        RECT 1.950 806.100 4.050 806.550 ;
        RECT 19.950 806.100 22.050 806.550 ;
        RECT 62.400 806.400 79.050 807.600 ;
        RECT 31.950 801.450 34.050 801.900 ;
        RECT 40.950 801.450 43.050 801.900 ;
        RECT 31.950 800.250 43.050 801.450 ;
        RECT 31.950 799.800 34.050 800.250 ;
        RECT 40.950 799.800 43.050 800.250 ;
        RECT 62.400 799.050 63.600 806.400 ;
        RECT 76.950 806.100 79.050 806.400 ;
        RECT 106.950 807.600 109.050 808.200 ;
        RECT 115.950 807.600 118.050 808.050 ;
        RECT 106.950 806.400 118.050 807.600 ;
        RECT 106.950 806.100 109.050 806.400 ;
        RECT 115.950 805.950 118.050 806.400 ;
        RECT 130.950 807.600 133.050 808.200 ;
        RECT 139.950 807.750 142.050 808.200 ;
        RECT 145.950 807.750 148.050 808.200 ;
        RECT 130.950 806.400 138.600 807.600 ;
        RECT 130.950 806.100 133.050 806.400 ;
        RECT 137.400 804.600 138.600 806.400 ;
        RECT 139.950 806.550 148.050 807.750 ;
        RECT 139.950 806.100 142.050 806.550 ;
        RECT 145.950 806.100 148.050 806.550 ;
        RECT 151.950 807.600 154.050 808.200 ;
        RECT 160.950 807.600 163.050 807.900 ;
        RECT 190.950 807.600 193.050 808.200 ;
        RECT 151.950 806.400 163.050 807.600 ;
        RECT 151.950 806.100 154.050 806.400 ;
        RECT 160.950 805.800 163.050 806.400 ;
        RECT 179.400 806.400 193.050 807.600 ;
        RECT 137.400 803.400 144.600 804.600 ;
        RECT 85.950 801.450 88.050 801.900 ;
        RECT 91.950 801.450 94.050 801.900 ;
        RECT 85.950 800.250 94.050 801.450 ;
        RECT 85.950 799.800 88.050 800.250 ;
        RECT 91.950 799.800 94.050 800.250 ;
        RECT 97.950 801.450 100.050 801.900 ;
        RECT 112.950 801.450 115.050 801.900 ;
        RECT 97.950 800.250 115.050 801.450 ;
        RECT 143.400 801.600 144.600 803.400 ;
        RECT 179.400 801.900 180.600 806.400 ;
        RECT 190.950 806.100 193.050 806.400 ;
        RECT 196.950 807.600 199.050 808.200 ;
        RECT 208.950 807.600 211.050 808.050 ;
        RECT 196.950 806.400 211.050 807.600 ;
        RECT 196.950 806.100 199.050 806.400 ;
        RECT 208.950 805.950 211.050 806.400 ;
        RECT 232.950 807.600 235.050 808.050 ;
        RECT 244.950 807.600 247.050 808.200 ;
        RECT 262.950 807.600 265.050 808.200 ;
        RECT 232.950 806.400 265.050 807.600 ;
        RECT 232.950 805.950 235.050 806.400 ;
        RECT 244.950 806.100 247.050 806.400 ;
        RECT 262.950 806.100 265.050 806.400 ;
        RECT 274.950 807.600 277.050 808.200 ;
        RECT 280.950 807.750 283.050 808.200 ;
        RECT 286.950 807.750 289.050 808.200 ;
        RECT 280.950 807.600 289.050 807.750 ;
        RECT 274.950 806.550 289.050 807.600 ;
        RECT 274.950 806.400 283.050 806.550 ;
        RECT 274.950 806.100 277.050 806.400 ;
        RECT 280.950 806.100 283.050 806.400 ;
        RECT 286.950 806.100 289.050 806.550 ;
        RECT 301.950 807.750 304.050 808.200 ;
        RECT 307.950 807.750 310.050 808.200 ;
        RECT 301.950 806.550 310.050 807.750 ;
        RECT 301.950 806.100 304.050 806.550 ;
        RECT 307.950 806.100 310.050 806.550 ;
        RECT 340.950 805.950 343.050 808.050 ;
        RECT 346.950 806.100 349.050 808.200 ;
        RECT 373.950 807.600 376.050 808.200 ;
        RECT 373.950 806.400 381.600 807.600 ;
        RECT 373.950 806.100 376.050 806.400 ;
        RECT 148.950 801.600 151.050 801.900 ;
        RECT 143.400 800.400 151.050 801.600 ;
        RECT 97.950 799.800 100.050 800.250 ;
        RECT 112.950 799.800 115.050 800.250 ;
        RECT 148.950 799.800 151.050 800.400 ;
        RECT 178.950 799.800 181.050 801.900 ;
        RECT 22.950 798.600 25.050 799.050 ;
        RECT 28.950 798.600 31.050 799.050 ;
        RECT 22.950 797.400 31.050 798.600 ;
        RECT 22.950 796.950 25.050 797.400 ;
        RECT 28.950 796.950 31.050 797.400 ;
        RECT 61.950 796.950 64.050 799.050 ;
        RECT 92.400 798.600 93.600 799.800 ;
        RECT 121.950 798.600 124.050 799.050 ;
        RECT 92.400 797.400 124.050 798.600 ;
        RECT 121.950 796.950 124.050 797.400 ;
        RECT 268.950 798.600 271.050 799.050 ;
        RECT 280.950 798.600 283.050 799.050 ;
        RECT 268.950 797.400 283.050 798.600 ;
        RECT 341.400 798.600 342.600 805.950 ;
        RECT 347.400 804.600 348.600 806.100 ;
        RECT 344.400 804.000 348.600 804.600 ;
        RECT 343.950 803.400 348.600 804.000 ;
        RECT 343.950 799.950 346.050 803.400 ;
        RECT 361.950 801.600 364.050 802.050 ;
        RECT 367.950 801.600 370.050 802.050 ;
        RECT 361.950 800.400 370.050 801.600 ;
        RECT 380.400 801.600 381.600 806.400 ;
        RECT 401.400 801.900 402.600 808.950 ;
        RECT 406.950 807.750 409.050 808.200 ;
        RECT 412.950 807.750 415.050 808.200 ;
        RECT 406.950 806.550 415.050 807.750 ;
        RECT 406.950 806.100 409.050 806.550 ;
        RECT 412.950 806.100 415.050 806.550 ;
        RECT 433.950 806.100 436.050 808.200 ;
        RECT 454.950 807.600 457.050 808.050 ;
        RECT 454.950 806.400 477.600 807.600 ;
        RECT 434.400 802.050 435.600 806.100 ;
        RECT 454.950 805.950 457.050 806.400 ;
        RECT 476.400 804.600 477.600 806.400 ;
        RECT 499.950 805.950 502.050 808.050 ;
        RECT 515.400 807.600 516.600 808.950 ;
        RECT 515.400 806.400 519.600 807.600 ;
        RECT 476.400 804.000 489.600 804.600 ;
        RECT 476.400 803.400 490.050 804.000 ;
        RECT 394.950 801.600 397.050 801.900 ;
        RECT 380.400 800.400 397.050 801.600 ;
        RECT 361.950 799.950 364.050 800.400 ;
        RECT 367.950 799.950 370.050 800.400 ;
        RECT 394.950 799.800 397.050 800.400 ;
        RECT 400.950 799.800 403.050 801.900 ;
        RECT 421.950 801.450 424.050 801.900 ;
        RECT 427.800 801.450 429.900 801.900 ;
        RECT 421.950 800.250 429.900 801.450 ;
        RECT 421.950 799.800 424.050 800.250 ;
        RECT 427.800 799.800 429.900 800.250 ;
        RECT 430.950 800.400 435.600 802.050 ;
        RECT 442.950 801.600 445.050 802.050 ;
        RECT 454.950 801.600 457.050 802.050 ;
        RECT 442.950 800.400 457.050 801.600 ;
        RECT 430.950 799.950 435.000 800.400 ;
        RECT 442.950 799.950 445.050 800.400 ;
        RECT 454.950 799.950 457.050 800.400 ;
        RECT 472.950 801.600 475.050 801.900 ;
        RECT 478.950 801.600 481.050 802.050 ;
        RECT 472.950 800.400 481.050 801.600 ;
        RECT 472.950 799.800 475.050 800.400 ;
        RECT 478.950 799.950 481.050 800.400 ;
        RECT 487.950 799.950 490.050 803.400 ;
        RECT 496.950 801.600 499.050 801.900 ;
        RECT 500.400 801.600 501.600 805.950 ;
        RECT 496.950 800.400 501.600 801.600 ;
        RECT 505.950 801.450 508.050 802.050 ;
        RECT 511.950 801.450 514.050 801.900 ;
        RECT 496.950 799.800 499.050 800.400 ;
        RECT 505.950 800.250 514.050 801.450 ;
        RECT 505.950 799.950 508.050 800.250 ;
        RECT 511.950 799.800 514.050 800.250 ;
        RECT 518.400 799.050 519.600 806.400 ;
        RECT 524.400 801.900 525.600 808.950 ;
        RECT 529.950 807.600 532.050 808.050 ;
        RECT 538.950 807.600 541.050 808.200 ;
        RECT 556.950 807.600 559.050 808.200 ;
        RECT 529.950 806.400 537.600 807.600 ;
        RECT 529.950 805.950 532.050 806.400 ;
        RECT 536.400 801.900 537.600 806.400 ;
        RECT 538.950 806.400 559.050 807.600 ;
        RECT 538.950 806.100 541.050 806.400 ;
        RECT 556.950 806.100 559.050 806.400 ;
        RECT 562.950 807.600 565.050 808.200 ;
        RECT 571.800 807.600 573.900 808.050 ;
        RECT 562.950 806.400 573.900 807.600 ;
        RECT 562.950 806.100 565.050 806.400 ;
        RECT 571.800 805.950 573.900 806.400 ;
        RECT 589.950 807.600 592.050 808.050 ;
        RECT 628.950 807.600 631.050 808.200 ;
        RECT 664.950 807.600 667.050 808.200 ;
        RECT 673.950 807.600 676.050 808.050 ;
        RECT 589.950 806.400 621.600 807.600 ;
        RECT 589.950 805.950 592.050 806.400 ;
        RECT 620.400 801.900 621.600 806.400 ;
        RECT 628.950 806.400 676.050 807.600 ;
        RECT 628.950 806.100 631.050 806.400 ;
        RECT 664.950 806.100 667.050 806.400 ;
        RECT 673.950 805.950 676.050 806.400 ;
        RECT 682.950 807.600 685.050 808.200 ;
        RECT 688.950 807.750 691.050 808.200 ;
        RECT 718.950 807.750 721.050 808.200 ;
        RECT 682.950 806.400 687.600 807.600 ;
        RECT 682.950 806.100 685.050 806.400 ;
        RECT 686.400 804.600 687.600 806.400 ;
        RECT 688.950 806.550 721.050 807.750 ;
        RECT 688.950 806.100 691.050 806.550 ;
        RECT 718.950 806.100 721.050 806.550 ;
        RECT 748.950 805.950 751.050 808.050 ;
        RECT 781.950 805.950 784.050 808.050 ;
        RECT 802.950 807.600 805.050 808.050 ;
        RECT 814.950 807.600 817.050 808.200 ;
        RECT 834.000 807.600 838.050 808.050 ;
        RECT 802.950 806.400 810.600 807.600 ;
        RECT 802.950 805.950 805.050 806.400 ;
        RECT 686.400 803.400 699.600 804.600 ;
        RECT 523.950 799.800 526.050 801.900 ;
        RECT 535.950 799.800 538.050 801.900 ;
        RECT 541.950 801.600 544.050 801.900 ;
        RECT 586.800 801.600 588.900 801.900 ;
        RECT 541.950 800.400 588.900 801.600 ;
        RECT 541.950 799.800 544.050 800.400 ;
        RECT 586.800 799.800 588.900 800.400 ;
        RECT 589.950 801.450 592.050 801.900 ;
        RECT 601.950 801.450 604.050 801.900 ;
        RECT 589.950 800.250 604.050 801.450 ;
        RECT 589.950 799.800 592.050 800.250 ;
        RECT 601.950 799.800 604.050 800.250 ;
        RECT 619.950 799.800 622.050 801.900 ;
        RECT 625.950 801.600 628.050 801.900 ;
        RECT 637.950 801.600 640.050 802.050 ;
        RECT 625.950 800.400 640.050 801.600 ;
        RECT 625.950 799.800 628.050 800.400 ;
        RECT 637.950 799.950 640.050 800.400 ;
        RECT 646.950 801.600 649.050 801.900 ;
        RECT 655.950 801.600 658.050 802.050 ;
        RECT 698.400 801.900 699.600 803.400 ;
        RECT 749.400 802.050 750.600 805.950 ;
        RECT 646.950 800.400 658.050 801.600 ;
        RECT 646.950 799.800 649.050 800.400 ;
        RECT 655.950 799.950 658.050 800.400 ;
        RECT 673.950 801.450 676.050 801.900 ;
        RECT 679.950 801.450 682.050 801.900 ;
        RECT 673.950 800.250 682.050 801.450 ;
        RECT 673.950 799.800 676.050 800.250 ;
        RECT 679.950 799.800 682.050 800.250 ;
        RECT 697.950 799.800 700.050 801.900 ;
        RECT 748.950 799.950 751.050 802.050 ;
        RECT 782.400 801.600 783.600 805.950 ;
        RECT 809.400 804.600 810.600 806.400 ;
        RECT 814.950 806.400 828.600 807.600 ;
        RECT 814.950 806.100 817.050 806.400 ;
        RECT 809.400 803.400 813.600 804.600 ;
        RECT 812.400 801.900 813.600 803.400 ;
        RECT 827.400 801.900 828.600 806.400 ;
        RECT 833.400 805.950 838.050 807.600 ;
        RECT 847.950 806.100 850.050 808.200 ;
        RECT 833.400 801.900 834.600 805.950 ;
        RECT 787.950 801.600 790.050 801.900 ;
        RECT 782.400 800.400 790.050 801.600 ;
        RECT 787.950 799.800 790.050 800.400 ;
        RECT 811.950 799.800 814.050 801.900 ;
        RECT 826.950 799.800 829.050 801.900 ;
        RECT 832.950 799.800 835.050 801.900 ;
        RECT 848.400 801.600 849.600 806.100 ;
        RECT 874.950 805.950 877.050 808.050 ;
        RECT 915.000 807.600 919.050 808.050 ;
        RECT 914.400 805.950 919.050 807.600 ;
        RECT 859.950 801.600 862.050 802.050 ;
        RECT 848.400 800.400 862.050 801.600 ;
        RECT 859.950 799.950 862.050 800.400 ;
        RECT 871.950 801.600 874.050 801.900 ;
        RECT 875.400 801.600 876.600 805.950 ;
        RECT 914.400 802.050 915.600 805.950 ;
        RECT 871.950 800.400 876.600 801.600 ;
        RECT 877.950 801.600 880.050 802.050 ;
        RECT 889.950 801.600 892.050 801.900 ;
        RECT 877.950 800.400 892.050 801.600 ;
        RECT 914.400 800.400 919.050 802.050 ;
        RECT 871.950 799.800 874.050 800.400 ;
        RECT 877.950 799.950 880.050 800.400 ;
        RECT 889.950 799.800 892.050 800.400 ;
        RECT 915.000 799.950 919.050 800.400 ;
        RECT 346.950 798.600 349.050 799.050 ;
        RECT 341.400 797.400 349.050 798.600 ;
        RECT 268.950 796.950 271.050 797.400 ;
        RECT 280.950 796.950 283.050 797.400 ;
        RECT 346.950 796.950 349.050 797.400 ;
        RECT 415.950 798.600 418.050 799.050 ;
        RECT 436.950 798.600 439.050 799.050 ;
        RECT 415.950 797.400 439.050 798.600 ;
        RECT 415.950 796.950 418.050 797.400 ;
        RECT 436.950 796.950 439.050 797.400 ;
        RECT 514.950 797.400 519.600 799.050 ;
        RECT 643.950 798.600 646.050 799.050 ;
        RECT 706.950 798.600 709.050 799.050 ;
        RECT 712.950 798.600 715.050 799.050 ;
        RECT 643.950 797.400 715.050 798.600 ;
        RECT 514.950 796.950 519.000 797.400 ;
        RECT 643.950 796.950 646.050 797.400 ;
        RECT 706.950 796.950 709.050 797.400 ;
        RECT 712.950 796.950 715.050 797.400 ;
        RECT 718.950 798.600 721.050 799.050 ;
        RECT 745.950 798.600 748.050 799.050 ;
        RECT 718.950 797.400 748.050 798.600 ;
        RECT 718.950 796.950 721.050 797.400 ;
        RECT 745.950 796.950 748.050 797.400 ;
        RECT 29.400 795.600 30.600 796.950 ;
        RECT 58.950 795.600 61.050 796.050 ;
        RECT 29.400 794.400 61.050 795.600 ;
        RECT 58.950 793.950 61.050 794.400 ;
        RECT 103.950 795.600 106.050 796.050 ;
        RECT 127.950 795.600 130.050 796.050 ;
        RECT 103.950 794.400 130.050 795.600 ;
        RECT 103.950 793.950 106.050 794.400 ;
        RECT 127.950 793.950 130.050 794.400 ;
        RECT 145.950 795.600 148.050 796.050 ;
        RECT 154.950 795.600 157.050 796.050 ;
        RECT 145.950 794.400 157.050 795.600 ;
        RECT 145.950 793.950 148.050 794.400 ;
        RECT 154.950 793.950 157.050 794.400 ;
        RECT 160.950 795.600 163.050 796.050 ;
        RECT 193.950 795.600 196.050 796.050 ;
        RECT 160.950 794.400 196.050 795.600 ;
        RECT 160.950 793.950 163.050 794.400 ;
        RECT 193.950 793.950 196.050 794.400 ;
        RECT 271.950 795.600 274.050 796.050 ;
        RECT 289.950 795.600 292.050 796.050 ;
        RECT 271.950 794.400 292.050 795.600 ;
        RECT 271.950 793.950 274.050 794.400 ;
        RECT 289.950 793.950 292.050 794.400 ;
        RECT 310.950 795.600 313.050 796.050 ;
        RECT 322.950 795.600 325.050 796.050 ;
        RECT 349.950 795.600 352.050 796.050 ;
        RECT 310.950 794.400 352.050 795.600 ;
        RECT 310.950 793.950 313.050 794.400 ;
        RECT 322.950 793.950 325.050 794.400 ;
        RECT 349.950 793.950 352.050 794.400 ;
        RECT 364.950 795.600 367.050 796.050 ;
        RECT 385.950 795.600 388.050 796.050 ;
        RECT 364.950 794.400 388.050 795.600 ;
        RECT 364.950 793.950 367.050 794.400 ;
        RECT 385.950 793.950 388.050 794.400 ;
        RECT 397.950 795.600 400.050 796.050 ;
        RECT 416.400 795.600 417.600 796.950 ;
        RECT 397.950 794.400 417.600 795.600 ;
        RECT 515.400 795.600 516.600 796.950 ;
        RECT 541.950 795.600 544.050 796.050 ;
        RECT 515.400 794.400 544.050 795.600 ;
        RECT 397.950 793.950 400.050 794.400 ;
        RECT 541.950 793.950 544.050 794.400 ;
        RECT 571.950 795.600 574.050 796.050 ;
        RECT 598.950 795.600 601.050 796.050 ;
        RECT 571.950 794.400 601.050 795.600 ;
        RECT 571.950 793.950 574.050 794.400 ;
        RECT 598.950 793.950 601.050 794.400 ;
        RECT 610.950 795.600 613.050 796.050 ;
        RECT 631.950 795.600 634.050 796.050 ;
        RECT 610.950 794.400 634.050 795.600 ;
        RECT 610.950 793.950 613.050 794.400 ;
        RECT 631.950 793.950 634.050 794.400 ;
        RECT 652.950 795.600 655.050 796.050 ;
        RECT 667.950 795.600 670.050 796.050 ;
        RECT 652.950 794.400 670.050 795.600 ;
        RECT 652.950 793.950 655.050 794.400 ;
        RECT 667.950 793.950 670.050 794.400 ;
        RECT 823.950 795.600 826.050 796.050 ;
        RECT 850.950 795.600 853.050 796.050 ;
        RECT 823.950 794.400 853.050 795.600 ;
        RECT 823.950 793.950 826.050 794.400 ;
        RECT 850.950 793.950 853.050 794.400 ;
        RECT 13.950 792.600 16.050 793.050 ;
        RECT 46.800 792.600 48.900 793.050 ;
        RECT 13.950 791.400 48.900 792.600 ;
        RECT 13.950 790.950 16.050 791.400 ;
        RECT 46.800 790.950 48.900 791.400 ;
        RECT 49.950 792.600 52.050 793.050 ;
        RECT 79.950 792.600 82.050 793.050 ;
        RECT 49.950 791.400 82.050 792.600 ;
        RECT 49.950 790.950 52.050 791.400 ;
        RECT 79.950 790.950 82.050 791.400 ;
        RECT 172.950 792.600 175.050 793.050 ;
        RECT 187.950 792.600 190.050 793.050 ;
        RECT 172.950 791.400 190.050 792.600 ;
        RECT 172.950 790.950 175.050 791.400 ;
        RECT 187.950 790.950 190.050 791.400 ;
        RECT 340.950 792.600 343.050 793.050 ;
        RECT 370.950 792.600 373.050 793.050 ;
        RECT 340.950 791.400 373.050 792.600 ;
        RECT 340.950 790.950 343.050 791.400 ;
        RECT 370.950 790.950 373.050 791.400 ;
        RECT 430.950 792.600 433.050 793.050 ;
        RECT 463.950 792.600 466.050 793.050 ;
        RECT 481.950 792.600 484.050 793.050 ;
        RECT 595.950 792.600 598.050 793.050 ;
        RECT 430.950 791.400 598.050 792.600 ;
        RECT 430.950 790.950 433.050 791.400 ;
        RECT 463.950 790.950 466.050 791.400 ;
        RECT 481.950 790.950 484.050 791.400 ;
        RECT 595.950 790.950 598.050 791.400 ;
        RECT 760.950 792.600 763.050 793.050 ;
        RECT 781.950 792.600 784.050 793.050 ;
        RECT 760.950 791.400 784.050 792.600 ;
        RECT 760.950 790.950 763.050 791.400 ;
        RECT 781.950 790.950 784.050 791.400 ;
        RECT 811.950 792.600 814.050 793.050 ;
        RECT 856.950 792.600 859.050 793.050 ;
        RECT 811.950 791.400 859.050 792.600 ;
        RECT 811.950 790.950 814.050 791.400 ;
        RECT 856.950 790.950 859.050 791.400 ;
        RECT 64.950 789.600 67.050 790.050 ;
        RECT 220.950 789.600 223.050 790.050 ;
        RECT 64.950 788.400 223.050 789.600 ;
        RECT 64.950 787.950 67.050 788.400 ;
        RECT 220.950 787.950 223.050 788.400 ;
        RECT 235.950 789.600 238.050 790.050 ;
        RECT 265.950 789.600 268.050 790.050 ;
        RECT 301.950 789.600 304.050 790.050 ;
        RECT 235.950 788.400 304.050 789.600 ;
        RECT 235.950 787.950 238.050 788.400 ;
        RECT 265.950 787.950 268.050 788.400 ;
        RECT 301.950 787.950 304.050 788.400 ;
        RECT 307.950 789.600 310.050 790.050 ;
        RECT 316.950 789.600 319.050 790.050 ;
        RECT 307.950 788.400 319.050 789.600 ;
        RECT 307.950 787.950 310.050 788.400 ;
        RECT 316.950 787.950 319.050 788.400 ;
        RECT 334.950 789.600 337.050 790.050 ;
        RECT 382.800 789.600 384.900 790.050 ;
        RECT 334.950 788.400 384.900 789.600 ;
        RECT 334.950 787.950 337.050 788.400 ;
        RECT 382.800 787.950 384.900 788.400 ;
        RECT 385.950 789.600 388.050 790.050 ;
        RECT 391.950 789.600 394.050 790.050 ;
        RECT 433.950 789.600 436.050 790.050 ;
        RECT 439.950 789.600 442.050 790.050 ;
        RECT 385.950 788.400 420.600 789.600 ;
        RECT 385.950 787.950 388.050 788.400 ;
        RECT 391.950 787.950 394.050 788.400 ;
        RECT 1.950 786.600 4.050 787.050 ;
        RECT 65.400 786.600 66.600 787.950 ;
        RECT 1.950 785.400 66.600 786.600 ;
        RECT 82.950 786.600 85.050 787.050 ;
        RECT 139.950 786.600 142.050 787.050 ;
        RECT 82.950 785.400 142.050 786.600 ;
        RECT 1.950 784.950 4.050 785.400 ;
        RECT 82.950 784.950 85.050 785.400 ;
        RECT 139.950 784.950 142.050 785.400 ;
        RECT 169.950 786.600 172.050 787.050 ;
        RECT 184.950 786.600 187.050 787.050 ;
        RECT 169.950 785.400 187.050 786.600 ;
        RECT 169.950 784.950 172.050 785.400 ;
        RECT 184.950 784.950 187.050 785.400 ;
        RECT 223.950 786.600 226.050 787.050 ;
        RECT 247.950 786.600 250.050 787.050 ;
        RECT 286.800 786.600 288.900 787.050 ;
        RECT 223.950 785.400 288.900 786.600 ;
        RECT 223.950 784.950 226.050 785.400 ;
        RECT 247.950 784.950 250.050 785.400 ;
        RECT 286.800 784.950 288.900 785.400 ;
        RECT 289.950 786.600 292.050 787.050 ;
        RECT 328.950 786.600 331.050 787.050 ;
        RECT 289.950 785.400 331.050 786.600 ;
        RECT 289.950 784.950 292.050 785.400 ;
        RECT 328.950 784.950 331.050 785.400 ;
        RECT 343.950 786.600 346.050 787.050 ;
        RECT 349.950 786.600 352.050 787.050 ;
        RECT 343.950 785.400 352.050 786.600 ;
        RECT 419.400 786.600 420.600 788.400 ;
        RECT 433.950 788.400 442.050 789.600 ;
        RECT 433.950 787.950 436.050 788.400 ;
        RECT 439.950 787.950 442.050 788.400 ;
        RECT 517.950 789.600 520.050 790.050 ;
        RECT 559.950 789.600 562.050 790.050 ;
        RECT 517.950 788.400 562.050 789.600 ;
        RECT 517.950 787.950 520.050 788.400 ;
        RECT 559.950 787.950 562.050 788.400 ;
        RECT 586.950 789.600 589.050 790.050 ;
        RECT 634.950 789.600 637.050 790.050 ;
        RECT 586.950 788.400 637.050 789.600 ;
        RECT 586.950 787.950 589.050 788.400 ;
        RECT 634.950 787.950 637.050 788.400 ;
        RECT 670.950 789.600 673.050 790.050 ;
        RECT 733.950 789.600 736.050 790.050 ;
        RECT 862.950 789.600 865.050 790.050 ;
        RECT 670.950 788.400 736.050 789.600 ;
        RECT 670.950 787.950 673.050 788.400 ;
        RECT 733.950 787.950 736.050 788.400 ;
        RECT 767.400 788.400 865.050 789.600 ;
        RECT 451.950 786.600 454.050 787.050 ;
        RECT 419.400 785.400 454.050 786.600 ;
        RECT 343.950 784.950 346.050 785.400 ;
        RECT 349.950 784.950 352.050 785.400 ;
        RECT 451.950 784.950 454.050 785.400 ;
        RECT 475.950 786.600 478.050 787.050 ;
        RECT 481.950 786.600 484.050 787.050 ;
        RECT 475.950 785.400 484.050 786.600 ;
        RECT 475.950 784.950 478.050 785.400 ;
        RECT 481.950 784.950 484.050 785.400 ;
        RECT 499.950 786.600 502.050 787.050 ;
        RECT 523.950 786.600 526.050 787.050 ;
        RECT 556.950 786.600 559.050 787.050 ;
        RECT 499.950 785.400 559.050 786.600 ;
        RECT 499.950 784.950 502.050 785.400 ;
        RECT 523.950 784.950 526.050 785.400 ;
        RECT 556.950 784.950 559.050 785.400 ;
        RECT 580.950 786.600 583.050 787.050 ;
        RECT 589.950 786.600 592.050 787.050 ;
        RECT 580.950 785.400 592.050 786.600 ;
        RECT 580.950 784.950 583.050 785.400 ;
        RECT 589.950 784.950 592.050 785.400 ;
        RECT 595.950 786.600 598.050 787.050 ;
        RECT 649.950 786.600 652.050 787.050 ;
        RECT 595.950 785.400 652.050 786.600 ;
        RECT 595.950 784.950 598.050 785.400 ;
        RECT 649.950 784.950 652.050 785.400 ;
        RECT 673.950 786.600 676.050 787.050 ;
        RECT 767.400 786.600 768.600 788.400 ;
        RECT 862.950 787.950 865.050 788.400 ;
        RECT 673.950 785.400 768.600 786.600 ;
        RECT 769.950 786.600 772.050 787.050 ;
        RECT 811.950 786.600 814.050 787.050 ;
        RECT 769.950 785.400 814.050 786.600 ;
        RECT 673.950 784.950 676.050 785.400 ;
        RECT 769.950 784.950 772.050 785.400 ;
        RECT 811.950 784.950 814.050 785.400 ;
        RECT 28.950 783.600 31.050 784.050 ;
        RECT 52.950 783.600 55.050 784.050 ;
        RECT 28.950 782.400 55.050 783.600 ;
        RECT 28.950 781.950 31.050 782.400 ;
        RECT 52.950 781.950 55.050 782.400 ;
        RECT 301.950 783.600 304.050 784.050 ;
        RECT 310.950 783.600 313.050 784.050 ;
        RECT 301.950 782.400 313.050 783.600 ;
        RECT 301.950 781.950 304.050 782.400 ;
        RECT 310.950 781.950 313.050 782.400 ;
        RECT 415.950 783.600 418.050 784.050 ;
        RECT 457.950 783.600 460.050 784.050 ;
        RECT 415.950 782.400 460.050 783.600 ;
        RECT 415.950 781.950 418.050 782.400 ;
        RECT 457.950 781.950 460.050 782.400 ;
        RECT 502.950 783.600 505.050 784.050 ;
        RECT 565.950 783.600 568.050 784.050 ;
        RECT 502.950 782.400 568.050 783.600 ;
        RECT 502.950 781.950 505.050 782.400 ;
        RECT 565.950 781.950 568.050 782.400 ;
        RECT 604.950 783.600 607.050 784.050 ;
        RECT 622.950 783.600 625.050 784.050 ;
        RECT 604.950 782.400 625.050 783.600 ;
        RECT 604.950 781.950 607.050 782.400 ;
        RECT 622.950 781.950 625.050 782.400 ;
        RECT 655.950 783.600 658.050 784.050 ;
        RECT 667.950 783.600 670.050 784.050 ;
        RECT 655.950 782.400 670.050 783.600 ;
        RECT 655.950 781.950 658.050 782.400 ;
        RECT 667.950 781.950 670.050 782.400 ;
        RECT 757.950 783.600 760.050 784.050 ;
        RECT 796.950 783.600 799.050 784.050 ;
        RECT 757.950 782.400 799.050 783.600 ;
        RECT 757.950 781.950 760.050 782.400 ;
        RECT 796.950 781.950 799.050 782.400 ;
        RECT 76.950 780.600 79.050 781.050 ;
        RECT 103.950 780.600 106.050 781.050 ;
        RECT 76.950 779.400 106.050 780.600 ;
        RECT 76.950 778.950 79.050 779.400 ;
        RECT 103.950 778.950 106.050 779.400 ;
        RECT 163.950 780.600 166.050 781.050 ;
        RECT 175.950 780.600 178.050 781.050 ;
        RECT 163.950 779.400 178.050 780.600 ;
        RECT 163.950 778.950 166.050 779.400 ;
        RECT 175.950 778.950 178.050 779.400 ;
        RECT 229.950 780.600 232.050 781.050 ;
        RECT 280.950 780.600 283.050 781.050 ;
        RECT 229.950 779.400 283.050 780.600 ;
        RECT 229.950 778.950 232.050 779.400 ;
        RECT 280.950 778.950 283.050 779.400 ;
        RECT 286.950 780.600 289.050 781.050 ;
        RECT 322.950 780.600 325.050 781.050 ;
        RECT 286.950 779.400 325.050 780.600 ;
        RECT 286.950 778.950 289.050 779.400 ;
        RECT 322.950 778.950 325.050 779.400 ;
        RECT 391.950 780.600 394.050 781.050 ;
        RECT 406.950 780.600 409.050 781.050 ;
        RECT 391.950 779.400 409.050 780.600 ;
        RECT 391.950 778.950 394.050 779.400 ;
        RECT 406.950 778.950 409.050 779.400 ;
        RECT 436.950 780.600 439.050 781.050 ;
        RECT 487.950 780.600 490.050 781.050 ;
        RECT 436.950 779.400 490.050 780.600 ;
        RECT 436.950 778.950 439.050 779.400 ;
        RECT 487.950 778.950 490.050 779.400 ;
        RECT 508.950 780.600 511.050 781.050 ;
        RECT 526.950 780.600 529.050 781.050 ;
        RECT 508.950 779.400 529.050 780.600 ;
        RECT 508.950 778.950 511.050 779.400 ;
        RECT 526.950 778.950 529.050 779.400 ;
        RECT 625.950 780.600 628.050 781.050 ;
        RECT 643.950 780.600 646.050 781.050 ;
        RECT 625.950 779.400 646.050 780.600 ;
        RECT 625.950 778.950 628.050 779.400 ;
        RECT 643.950 778.950 646.050 779.400 ;
        RECT 649.950 780.600 652.050 781.050 ;
        RECT 676.950 780.600 679.050 781.050 ;
        RECT 649.950 779.400 679.050 780.600 ;
        RECT 649.950 778.950 652.050 779.400 ;
        RECT 676.950 778.950 679.050 779.400 ;
        RECT 736.950 780.600 739.050 781.050 ;
        RECT 760.950 780.600 763.050 781.050 ;
        RECT 736.950 779.400 763.050 780.600 ;
        RECT 736.950 778.950 739.050 779.400 ;
        RECT 760.950 778.950 763.050 779.400 ;
        RECT 787.950 780.600 790.050 781.050 ;
        RECT 826.950 780.600 829.050 781.050 ;
        RECT 859.950 780.600 862.050 781.050 ;
        RECT 904.950 780.600 907.050 781.050 ;
        RECT 787.950 779.400 907.050 780.600 ;
        RECT 787.950 778.950 790.050 779.400 ;
        RECT 826.950 778.950 829.050 779.400 ;
        RECT 859.950 778.950 862.050 779.400 ;
        RECT 904.950 778.950 907.050 779.400 ;
        RECT 208.950 777.600 211.050 778.050 ;
        RECT 310.950 777.600 313.050 778.050 ;
        RECT 208.950 776.400 313.050 777.600 ;
        RECT 208.950 775.950 211.050 776.400 ;
        RECT 310.950 775.950 313.050 776.400 ;
        RECT 319.950 777.600 322.050 778.050 ;
        RECT 328.950 777.600 331.050 778.050 ;
        RECT 319.950 776.400 331.050 777.600 ;
        RECT 319.950 775.950 322.050 776.400 ;
        RECT 328.950 775.950 331.050 776.400 ;
        RECT 388.950 777.600 391.050 778.050 ;
        RECT 412.950 777.600 415.050 778.050 ;
        RECT 388.950 776.400 415.050 777.600 ;
        RECT 388.950 775.950 391.050 776.400 ;
        RECT 412.950 775.950 415.050 776.400 ;
        RECT 445.950 777.600 448.050 778.050 ;
        RECT 451.950 777.600 454.050 778.050 ;
        RECT 445.950 776.400 454.050 777.600 ;
        RECT 445.950 775.950 448.050 776.400 ;
        RECT 451.950 775.950 454.050 776.400 ;
        RECT 529.950 777.600 532.050 778.050 ;
        RECT 544.950 777.600 547.050 778.050 ;
        RECT 529.950 776.400 547.050 777.600 ;
        RECT 529.950 775.950 532.050 776.400 ;
        RECT 544.950 775.950 547.050 776.400 ;
        RECT 592.950 777.600 595.050 778.050 ;
        RECT 604.950 777.600 607.050 778.050 ;
        RECT 592.950 776.400 607.050 777.600 ;
        RECT 592.950 775.950 595.050 776.400 ;
        RECT 604.950 775.950 607.050 776.400 ;
        RECT 637.950 777.600 640.050 778.050 ;
        RECT 682.950 777.600 685.050 778.050 ;
        RECT 637.950 776.400 685.050 777.600 ;
        RECT 637.950 775.950 640.050 776.400 ;
        RECT 682.950 775.950 685.050 776.400 ;
        RECT 715.950 777.600 718.050 778.050 ;
        RECT 808.950 777.600 811.050 778.050 ;
        RECT 850.950 777.600 853.050 778.050 ;
        RECT 715.950 776.400 750.600 777.600 ;
        RECT 715.950 775.950 718.050 776.400 ;
        RECT 749.400 775.050 750.600 776.400 ;
        RECT 808.950 776.400 853.050 777.600 ;
        RECT 808.950 775.950 811.050 776.400 ;
        RECT 850.950 775.950 853.050 776.400 ;
        RECT 115.950 774.600 118.050 775.050 ;
        RECT 145.950 774.600 148.050 775.050 ;
        RECT 115.950 773.400 148.050 774.600 ;
        RECT 115.950 772.950 118.050 773.400 ;
        RECT 145.950 772.950 148.050 773.400 ;
        RECT 163.950 774.600 166.050 775.050 ;
        RECT 205.950 774.600 208.050 775.050 ;
        RECT 163.950 773.400 208.050 774.600 ;
        RECT 163.950 772.950 166.050 773.400 ;
        RECT 205.950 772.950 208.050 773.400 ;
        RECT 217.950 774.600 220.050 775.050 ;
        RECT 241.950 774.600 244.050 775.050 ;
        RECT 217.950 773.400 244.050 774.600 ;
        RECT 217.950 772.950 220.050 773.400 ;
        RECT 241.950 772.950 244.050 773.400 ;
        RECT 376.950 774.600 379.050 775.050 ;
        RECT 400.950 774.600 403.050 775.050 ;
        RECT 376.950 773.400 403.050 774.600 ;
        RECT 376.950 772.950 379.050 773.400 ;
        RECT 400.950 772.950 403.050 773.400 ;
        RECT 445.950 774.600 448.050 774.900 ;
        RECT 466.950 774.600 469.050 775.050 ;
        RECT 445.950 773.400 469.050 774.600 ;
        RECT 445.950 772.800 448.050 773.400 ;
        RECT 466.950 772.950 469.050 773.400 ;
        RECT 472.950 774.600 475.050 775.050 ;
        RECT 514.950 774.600 517.050 775.050 ;
        RECT 472.950 773.400 517.050 774.600 ;
        RECT 472.950 772.950 475.050 773.400 ;
        RECT 514.950 772.950 517.050 773.400 ;
        RECT 556.950 774.600 559.050 775.050 ;
        RECT 571.950 774.600 574.050 775.050 ;
        RECT 556.950 773.400 574.050 774.600 ;
        RECT 556.950 772.950 559.050 773.400 ;
        RECT 571.950 772.950 574.050 773.400 ;
        RECT 601.950 774.600 604.050 775.050 ;
        RECT 619.950 774.600 622.050 775.050 ;
        RECT 601.950 773.400 622.050 774.600 ;
        RECT 601.950 772.950 604.050 773.400 ;
        RECT 619.950 772.950 622.050 773.400 ;
        RECT 628.950 774.600 631.050 774.900 ;
        RECT 685.950 774.600 688.050 775.050 ;
        RECT 628.950 773.400 688.050 774.600 ;
        RECT 628.950 772.800 631.050 773.400 ;
        RECT 685.950 772.950 688.050 773.400 ;
        RECT 694.950 774.600 697.050 775.050 ;
        RECT 739.950 774.600 742.050 775.050 ;
        RECT 694.950 773.400 742.050 774.600 ;
        RECT 694.950 772.950 697.050 773.400 ;
        RECT 739.950 772.950 742.050 773.400 ;
        RECT 748.950 774.600 751.050 775.050 ;
        RECT 766.950 774.600 769.050 775.050 ;
        RECT 748.950 773.400 769.050 774.600 ;
        RECT 748.950 772.950 751.050 773.400 ;
        RECT 766.950 772.950 769.050 773.400 ;
        RECT 13.950 771.600 16.050 772.050 ;
        RECT 49.950 771.600 52.050 772.050 ;
        RECT 13.950 770.400 52.050 771.600 ;
        RECT 13.950 769.950 16.050 770.400 ;
        RECT 49.950 769.950 52.050 770.400 ;
        RECT 67.950 771.600 70.050 772.050 ;
        RECT 82.950 771.600 85.050 772.050 ;
        RECT 67.950 770.400 85.050 771.600 ;
        RECT 67.950 769.950 70.050 770.400 ;
        RECT 82.950 769.950 85.050 770.400 ;
        RECT 490.950 771.600 493.050 772.050 ;
        RECT 532.950 771.600 535.050 772.050 ;
        RECT 490.950 770.400 535.050 771.600 ;
        RECT 490.950 769.950 493.050 770.400 ;
        RECT 532.950 769.950 535.050 770.400 ;
        RECT 538.950 771.600 541.050 772.050 ;
        RECT 583.950 771.600 586.050 772.050 ;
        RECT 538.950 770.400 586.050 771.600 ;
        RECT 538.950 769.950 541.050 770.400 ;
        RECT 583.950 769.950 586.050 770.400 ;
        RECT 850.950 771.600 853.050 772.050 ;
        RECT 877.950 771.600 880.050 772.050 ;
        RECT 850.950 770.400 880.050 771.600 ;
        RECT 850.950 769.950 853.050 770.400 ;
        RECT 877.950 769.950 880.050 770.400 ;
        RECT 172.950 768.600 175.050 769.050 ;
        RECT 202.950 768.600 205.050 769.050 ;
        RECT 172.950 767.400 205.050 768.600 ;
        RECT 172.950 766.950 175.050 767.400 ;
        RECT 202.950 766.950 205.050 767.400 ;
        RECT 262.950 768.600 265.050 769.050 ;
        RECT 316.950 768.600 319.050 769.050 ;
        RECT 376.950 768.600 379.050 769.050 ;
        RECT 385.950 768.600 388.050 769.050 ;
        RECT 262.950 767.400 330.600 768.600 ;
        RECT 262.950 766.950 265.050 767.400 ;
        RECT 316.950 766.950 319.050 767.400 ;
        RECT 52.950 765.600 55.050 766.050 ;
        RECT 100.950 765.600 103.050 766.050 ;
        RECT 52.950 764.400 103.050 765.600 ;
        RECT 52.950 763.950 55.050 764.400 ;
        RECT 100.950 763.950 103.050 764.400 ;
        RECT 193.950 765.600 196.050 766.050 ;
        RECT 199.950 765.600 202.050 766.050 ;
        RECT 193.950 764.400 202.050 765.600 ;
        RECT 193.950 763.950 196.050 764.400 ;
        RECT 199.950 763.950 202.050 764.400 ;
        RECT 220.950 765.600 223.050 766.050 ;
        RECT 229.950 765.600 232.050 766.050 ;
        RECT 220.950 764.400 232.050 765.600 ;
        RECT 329.400 765.600 330.600 767.400 ;
        RECT 376.950 767.400 388.050 768.600 ;
        RECT 376.950 766.950 379.050 767.400 ;
        RECT 385.950 766.950 388.050 767.400 ;
        RECT 394.950 768.600 397.050 769.050 ;
        RECT 403.950 768.600 406.050 769.050 ;
        RECT 394.950 767.400 406.050 768.600 ;
        RECT 394.950 766.950 397.050 767.400 ;
        RECT 403.950 766.950 406.050 767.400 ;
        RECT 553.950 768.600 556.050 769.050 ;
        RECT 565.950 768.600 568.050 769.050 ;
        RECT 553.950 767.400 568.050 768.600 ;
        RECT 553.950 766.950 556.050 767.400 ;
        RECT 565.950 766.950 568.050 767.400 ;
        RECT 574.950 768.600 577.050 769.050 ;
        RECT 592.950 768.600 595.050 769.050 ;
        RECT 600.000 768.600 604.050 769.050 ;
        RECT 574.950 767.400 595.050 768.600 ;
        RECT 574.950 766.950 577.050 767.400 ;
        RECT 592.950 766.950 595.050 767.400 ;
        RECT 599.400 766.950 604.050 768.600 ;
        RECT 607.800 768.000 609.900 769.050 ;
        RECT 610.950 768.600 613.050 769.050 ;
        RECT 682.950 768.600 685.050 769.050 ;
        RECT 724.950 768.600 727.050 769.050 ;
        RECT 607.800 766.950 610.050 768.000 ;
        RECT 610.950 767.400 633.600 768.600 ;
        RECT 610.950 766.950 613.050 767.400 ;
        RECT 352.950 765.600 355.050 766.050 ;
        RECT 329.400 764.400 355.050 765.600 ;
        RECT 220.950 763.950 223.050 764.400 ;
        RECT 229.950 763.950 232.050 764.400 ;
        RECT 352.950 763.950 355.050 764.400 ;
        RECT 358.950 765.600 361.050 766.050 ;
        RECT 391.950 765.600 394.050 766.050 ;
        RECT 424.950 765.600 427.050 766.050 ;
        RECT 358.950 764.400 394.050 765.600 ;
        RECT 358.950 763.950 361.050 764.400 ;
        RECT 7.950 762.750 10.050 763.200 ;
        RECT 19.950 762.750 22.050 763.200 ;
        RECT 7.950 762.600 22.050 762.750 ;
        RECT 37.950 762.600 40.050 763.200 ;
        RECT 7.950 761.550 40.050 762.600 ;
        RECT 7.950 761.100 10.050 761.550 ;
        RECT 19.950 761.400 40.050 761.550 ;
        RECT 19.950 761.100 22.050 761.400 ;
        RECT 37.950 761.100 40.050 761.400 ;
        RECT 43.950 762.750 46.050 763.200 ;
        RECT 76.950 762.750 79.050 763.200 ;
        RECT 43.950 761.550 79.050 762.750 ;
        RECT 43.950 761.100 46.050 761.550 ;
        RECT 76.950 761.100 79.050 761.550 ;
        RECT 106.950 762.750 109.050 763.200 ;
        RECT 112.950 762.750 115.050 763.200 ;
        RECT 106.950 761.550 115.050 762.750 ;
        RECT 106.950 761.100 109.050 761.550 ;
        RECT 112.950 761.100 115.050 761.550 ;
        RECT 121.950 762.600 124.050 763.200 ;
        RECT 130.950 762.600 133.050 763.050 ;
        RECT 163.950 762.600 166.050 763.200 ;
        RECT 121.950 761.400 133.050 762.600 ;
        RECT 121.950 761.100 124.050 761.400 ;
        RECT 130.950 760.950 133.050 761.400 ;
        RECT 134.400 761.400 166.050 762.600 ;
        RECT 134.400 759.600 135.600 761.400 ;
        RECT 163.950 761.100 166.050 761.400 ;
        RECT 211.950 762.750 214.050 763.200 ;
        RECT 217.950 762.750 220.050 763.200 ;
        RECT 211.950 761.550 220.050 762.750 ;
        RECT 211.950 761.100 214.050 761.550 ;
        RECT 217.950 761.100 220.050 761.550 ;
        RECT 241.950 762.750 244.050 763.200 ;
        RECT 247.950 762.750 250.050 763.200 ;
        RECT 241.950 762.600 250.050 762.750 ;
        RECT 262.950 762.600 265.050 763.200 ;
        RECT 241.950 761.550 265.050 762.600 ;
        RECT 241.950 761.100 244.050 761.550 ;
        RECT 247.950 761.400 265.050 761.550 ;
        RECT 247.950 761.100 250.050 761.400 ;
        RECT 262.950 761.100 265.050 761.400 ;
        RECT 271.800 762.000 273.900 763.050 ;
        RECT 271.800 760.950 274.050 762.000 ;
        RECT 274.950 761.100 277.050 763.200 ;
        RECT 286.950 762.750 289.050 763.200 ;
        RECT 292.950 762.750 295.050 763.200 ;
        RECT 286.950 761.550 295.050 762.750 ;
        RECT 286.950 761.100 289.050 761.550 ;
        RECT 292.950 761.100 295.050 761.550 ;
        RECT 322.950 762.600 325.050 763.200 ;
        RECT 322.950 761.400 345.600 762.600 ;
        RECT 322.950 761.100 325.050 761.400 ;
        RECT 271.950 759.600 274.050 760.950 ;
        RECT 125.400 758.400 135.600 759.600 ;
        RECT 263.400 759.000 274.050 759.600 ;
        RECT 263.400 758.400 273.450 759.000 ;
        RECT 125.400 756.900 126.600 758.400 ;
        RECT 4.950 756.450 7.050 756.900 ;
        RECT 22.950 756.600 25.050 756.900 ;
        RECT 34.950 756.600 37.050 756.900 ;
        RECT 22.950 756.450 37.050 756.600 ;
        RECT 4.950 755.400 37.050 756.450 ;
        RECT 4.950 755.250 25.050 755.400 ;
        RECT 4.950 754.800 7.050 755.250 ;
        RECT 22.950 754.800 25.050 755.250 ;
        RECT 34.950 754.800 37.050 755.400 ;
        RECT 124.950 754.800 127.050 756.900 ;
        RECT 202.950 756.600 205.050 756.900 ;
        RECT 238.950 756.600 241.050 756.900 ;
        RECT 202.950 755.400 241.050 756.600 ;
        RECT 202.950 754.800 205.050 755.400 ;
        RECT 238.950 754.800 241.050 755.400 ;
        RECT 259.950 756.600 262.050 756.900 ;
        RECT 263.400 756.600 264.600 758.400 ;
        RECT 259.950 755.400 264.600 756.600 ;
        RECT 265.950 756.600 268.050 757.050 ;
        RECT 275.400 756.600 276.600 761.100 ;
        RECT 344.400 757.050 345.600 761.400 ;
        RECT 382.950 761.100 385.050 763.200 ;
        RECT 349.950 759.600 352.050 760.050 ;
        RECT 383.400 759.600 384.600 761.100 ;
        RECT 349.950 758.400 384.600 759.600 ;
        RECT 349.950 757.950 352.050 758.400 ;
        RECT 265.950 755.400 276.600 756.600 ;
        RECT 283.950 756.600 286.050 757.050 ;
        RECT 307.950 756.600 310.050 757.050 ;
        RECT 283.950 755.400 310.050 756.600 ;
        RECT 259.950 754.800 262.050 755.400 ;
        RECT 265.950 754.950 268.050 755.400 ;
        RECT 283.950 754.950 286.050 755.400 ;
        RECT 307.950 754.950 310.050 755.400 ;
        RECT 343.950 754.950 346.050 757.050 ;
        RECT 386.400 756.900 387.600 764.400 ;
        RECT 391.950 763.950 394.050 764.400 ;
        RECT 419.400 764.400 427.050 765.600 ;
        RECT 391.950 762.600 394.050 762.900 ;
        RECT 403.950 762.600 406.050 763.200 ;
        RECT 391.950 761.400 406.050 762.600 ;
        RECT 391.950 760.800 394.050 761.400 ;
        RECT 403.950 761.100 406.050 761.400 ;
        RECT 419.400 759.600 420.600 764.400 ;
        RECT 424.950 763.950 427.050 764.400 ;
        RECT 532.950 765.600 535.050 766.050 ;
        RECT 599.400 765.600 600.600 766.950 ;
        RECT 532.950 764.400 600.600 765.600 ;
        RECT 607.950 765.600 610.050 766.950 ;
        RECT 613.950 765.600 616.050 766.050 ;
        RECT 607.950 765.000 616.050 765.600 ;
        RECT 608.250 764.400 616.050 765.000 ;
        RECT 532.950 763.950 535.050 764.400 ;
        RECT 613.950 763.950 616.050 764.400 ;
        RECT 619.950 765.600 622.050 766.050 ;
        RECT 619.950 764.400 630.600 765.600 ;
        RECT 619.950 763.950 622.050 764.400 ;
        RECT 421.950 762.600 424.050 763.200 ;
        RECT 445.950 762.600 448.050 763.200 ;
        RECT 421.950 761.400 448.050 762.600 ;
        RECT 421.950 761.100 424.050 761.400 ;
        RECT 445.950 761.100 448.050 761.400 ;
        RECT 451.950 761.100 454.050 763.200 ;
        RECT 493.950 762.600 496.050 763.200 ;
        RECT 508.950 762.600 511.050 763.050 ;
        RECT 493.950 761.400 511.050 762.600 ;
        RECT 493.950 761.100 496.050 761.400 ;
        RECT 452.400 759.600 453.600 761.100 ;
        RECT 508.950 760.950 511.050 761.400 ;
        RECT 520.950 762.600 523.050 763.200 ;
        RECT 538.950 762.600 541.050 763.200 ;
        RECT 520.950 761.400 541.050 762.600 ;
        RECT 520.950 761.100 523.050 761.400 ;
        RECT 538.950 761.100 541.050 761.400 ;
        RECT 559.950 761.100 562.050 763.200 ;
        RECT 580.950 762.600 583.050 763.050 ;
        RECT 569.400 761.400 583.050 762.600 ;
        RECT 560.400 759.600 561.600 761.100 ;
        RECT 419.400 758.400 423.600 759.600 ;
        RECT 452.400 758.400 462.600 759.600 ;
        RECT 367.950 756.450 370.050 756.900 ;
        RECT 373.950 756.450 376.050 756.900 ;
        RECT 367.950 755.250 376.050 756.450 ;
        RECT 367.950 754.800 370.050 755.250 ;
        RECT 373.950 754.800 376.050 755.250 ;
        RECT 385.950 756.600 388.050 756.900 ;
        RECT 406.950 756.600 409.050 756.900 ;
        RECT 385.950 755.400 409.050 756.600 ;
        RECT 385.950 754.800 388.050 755.400 ;
        RECT 406.950 754.800 409.050 755.400 ;
        RECT 422.400 754.050 423.600 758.400 ;
        RECT 436.950 756.600 439.050 757.050 ;
        RECT 448.950 756.600 451.050 756.900 ;
        RECT 436.950 755.400 451.050 756.600 ;
        RECT 461.400 756.600 462.600 758.400 ;
        RECT 554.400 758.400 561.600 759.600 ;
        RECT 463.950 756.600 466.050 756.900 ;
        RECT 461.400 755.400 466.050 756.600 ;
        RECT 436.950 754.950 439.050 755.400 ;
        RECT 448.950 754.800 451.050 755.400 ;
        RECT 463.950 754.800 466.050 755.400 ;
        RECT 475.950 756.450 478.050 756.900 ;
        RECT 490.950 756.450 493.050 756.900 ;
        RECT 475.950 755.250 493.050 756.450 ;
        RECT 475.950 754.800 478.050 755.250 ;
        RECT 490.950 754.800 493.050 755.250 ;
        RECT 502.950 756.450 505.050 756.900 ;
        RECT 523.950 756.600 526.050 756.900 ;
        RECT 529.950 756.600 532.050 757.050 ;
        RECT 523.950 756.450 532.050 756.600 ;
        RECT 502.950 755.400 532.050 756.450 ;
        RECT 502.950 755.250 526.050 755.400 ;
        RECT 502.950 754.800 505.050 755.250 ;
        RECT 523.950 754.800 526.050 755.250 ;
        RECT 529.950 754.950 532.050 755.400 ;
        RECT 541.950 756.600 544.050 756.900 ;
        RECT 554.400 756.600 555.600 758.400 ;
        RECT 541.950 755.400 555.600 756.600 ;
        RECT 556.950 756.600 559.050 757.050 ;
        RECT 569.400 756.600 570.600 761.400 ;
        RECT 580.950 760.950 583.050 761.400 ;
        RECT 589.950 762.600 594.000 763.050 ;
        RECT 589.950 760.950 594.600 762.600 ;
        RECT 616.950 761.100 619.050 763.200 ;
        RECT 556.950 755.400 570.600 756.600 ;
        RECT 593.400 756.600 594.600 760.950 ;
        RECT 617.400 757.050 618.600 761.100 ;
        RECT 601.950 756.600 604.050 757.050 ;
        RECT 593.400 755.400 604.050 756.600 ;
        RECT 617.400 755.400 622.050 757.050 ;
        RECT 629.400 756.600 630.600 764.400 ;
        RECT 632.400 762.600 633.600 767.400 ;
        RECT 682.950 767.400 727.050 768.600 ;
        RECT 682.950 766.950 685.050 767.400 ;
        RECT 724.950 766.950 727.050 767.400 ;
        RECT 820.950 768.600 823.050 769.050 ;
        RECT 841.950 768.600 844.050 769.050 ;
        RECT 898.950 768.600 901.050 769.050 ;
        RECT 913.950 768.600 916.050 769.050 ;
        RECT 820.950 767.400 916.050 768.600 ;
        RECT 820.950 766.950 823.050 767.400 ;
        RECT 841.950 766.950 844.050 767.400 ;
        RECT 898.950 766.950 901.050 767.400 ;
        RECT 913.950 766.950 916.050 767.400 ;
        RECT 634.950 765.600 637.050 766.050 ;
        RECT 661.950 765.600 664.050 766.050 ;
        RECT 685.950 765.600 688.050 766.050 ;
        RECT 634.950 764.400 651.600 765.600 ;
        RECT 634.950 763.950 637.050 764.400 ;
        RECT 650.400 762.600 651.600 764.400 ;
        RECT 661.950 764.400 688.050 765.600 ;
        RECT 661.950 763.950 664.050 764.400 ;
        RECT 685.950 763.950 688.050 764.400 ;
        RECT 721.950 765.600 724.050 766.050 ;
        RECT 736.950 765.600 739.050 766.050 ;
        RECT 721.950 764.400 739.050 765.600 ;
        RECT 721.950 763.950 724.050 764.400 ;
        RECT 736.950 763.950 739.050 764.400 ;
        RECT 772.950 765.600 775.050 766.050 ;
        RECT 778.950 765.600 781.050 766.050 ;
        RECT 883.950 765.600 886.050 766.050 ;
        RECT 895.950 765.600 898.050 766.050 ;
        RECT 772.950 764.400 781.050 765.600 ;
        RECT 772.950 763.950 775.050 764.400 ;
        RECT 778.950 763.950 781.050 764.400 ;
        RECT 875.400 764.400 898.050 765.600 ;
        RECT 673.800 762.600 675.900 763.050 ;
        RECT 632.400 761.400 636.600 762.600 ;
        RECT 650.400 761.400 675.900 762.600 ;
        RECT 635.400 759.600 636.600 761.400 ;
        RECT 653.400 759.600 654.600 761.400 ;
        RECT 673.800 760.950 675.900 761.400 ;
        RECT 676.950 762.600 679.050 763.200 ;
        RECT 685.950 762.600 688.050 763.200 ;
        RECT 703.950 762.600 706.050 763.200 ;
        RECT 676.950 761.400 681.600 762.600 ;
        RECT 676.950 761.100 679.050 761.400 ;
        RECT 635.400 758.400 651.600 759.600 ;
        RECT 653.400 758.400 657.600 759.600 ;
        RECT 650.400 757.050 651.600 758.400 ;
        RECT 634.950 756.600 637.050 756.900 ;
        RECT 646.950 756.600 649.050 757.050 ;
        RECT 629.400 755.400 649.050 756.600 ;
        RECT 650.400 755.400 655.050 757.050 ;
        RECT 656.400 756.600 657.600 758.400 ;
        RECT 680.400 757.050 681.600 761.400 ;
        RECT 685.950 761.400 706.050 762.600 ;
        RECT 685.950 761.100 688.050 761.400 ;
        RECT 703.950 761.100 706.050 761.400 ;
        RECT 730.950 761.100 733.050 763.200 ;
        RECT 787.950 762.600 790.050 763.200 ;
        RECT 776.400 761.400 790.050 762.600 ;
        RECT 673.950 756.600 676.050 757.050 ;
        RECT 656.400 755.400 676.050 756.600 ;
        RECT 541.950 754.800 544.050 755.400 ;
        RECT 556.950 754.950 559.050 755.400 ;
        RECT 601.950 754.950 604.050 755.400 ;
        RECT 618.000 754.950 622.050 755.400 ;
        RECT 634.950 754.800 637.050 755.400 ;
        RECT 646.950 754.950 649.050 755.400 ;
        RECT 651.000 754.950 655.050 755.400 ;
        RECT 673.950 754.950 676.050 755.400 ;
        RECT 679.950 754.950 682.050 757.050 ;
        RECT 706.950 756.600 709.050 756.900 ;
        RECT 721.950 756.600 724.050 756.900 ;
        RECT 706.950 755.400 724.050 756.600 ;
        RECT 731.400 756.600 732.600 761.100 ;
        RECT 776.400 756.900 777.600 761.400 ;
        RECT 787.950 761.100 790.050 761.400 ;
        RECT 793.950 762.750 796.050 763.200 ;
        RECT 802.800 762.750 804.900 763.200 ;
        RECT 793.950 761.550 804.900 762.750 ;
        RECT 793.950 761.100 796.050 761.550 ;
        RECT 802.800 761.100 804.900 761.550 ;
        RECT 805.950 762.750 808.050 763.200 ;
        RECT 811.950 762.750 814.050 763.200 ;
        RECT 805.950 761.550 814.050 762.750 ;
        RECT 805.950 761.100 808.050 761.550 ;
        RECT 811.950 761.100 814.050 761.550 ;
        RECT 823.950 760.950 826.050 763.050 ;
        RECT 856.950 762.600 859.050 763.200 ;
        RECT 875.400 762.600 876.600 764.400 ;
        RECT 883.950 763.950 886.050 764.400 ;
        RECT 895.950 763.950 898.050 764.400 ;
        RECT 839.400 761.400 876.600 762.600 ;
        RECT 877.950 762.600 880.050 763.200 ;
        RECT 904.950 762.750 907.050 763.200 ;
        RECT 910.950 762.750 913.050 763.200 ;
        RECT 877.950 761.400 897.600 762.600 ;
        RECT 748.950 756.600 751.050 756.900 ;
        RECT 731.400 755.400 751.050 756.600 ;
        RECT 706.950 754.800 709.050 755.400 ;
        RECT 721.950 754.800 724.050 755.400 ;
        RECT 748.950 754.800 751.050 755.400 ;
        RECT 775.950 754.800 778.050 756.900 ;
        RECT 824.400 756.600 825.600 760.950 ;
        RECT 839.400 759.600 840.600 761.400 ;
        RECT 856.950 761.100 859.050 761.400 ;
        RECT 877.950 761.100 880.050 761.400 ;
        RECT 836.400 758.400 840.600 759.600 ;
        RECT 836.400 756.900 837.600 758.400 ;
        RECT 896.400 756.900 897.600 761.400 ;
        RECT 904.950 761.550 913.050 762.750 ;
        RECT 904.950 761.100 907.050 761.550 ;
        RECT 910.950 761.100 913.050 761.550 ;
        RECT 829.950 756.600 832.050 756.900 ;
        RECT 824.400 755.400 832.050 756.600 ;
        RECT 829.950 754.800 832.050 755.400 ;
        RECT 835.950 754.800 838.050 756.900 ;
        RECT 841.950 756.450 844.050 756.900 ;
        RECT 853.950 756.450 856.050 756.900 ;
        RECT 841.950 755.250 856.050 756.450 ;
        RECT 841.950 754.800 844.050 755.250 ;
        RECT 853.950 754.800 856.050 755.250 ;
        RECT 895.950 754.800 898.050 756.900 ;
        RECT 16.950 753.600 19.050 754.050 ;
        RECT 52.950 753.600 55.050 754.050 ;
        RECT 16.950 752.400 55.050 753.600 ;
        RECT 16.950 751.950 19.050 752.400 ;
        RECT 52.950 751.950 55.050 752.400 ;
        RECT 103.950 753.600 106.050 754.050 ;
        RECT 115.950 753.600 118.050 754.050 ;
        RECT 103.950 752.400 118.050 753.600 ;
        RECT 103.950 751.950 106.050 752.400 ;
        RECT 115.950 751.950 118.050 752.400 ;
        RECT 130.950 753.600 133.050 754.050 ;
        RECT 148.950 753.600 151.050 754.050 ;
        RECT 130.950 752.400 151.050 753.600 ;
        RECT 130.950 751.950 133.050 752.400 ;
        RECT 148.950 751.950 151.050 752.400 ;
        RECT 181.950 753.600 184.050 754.050 ;
        RECT 187.950 753.600 190.050 754.050 ;
        RECT 181.950 752.400 190.050 753.600 ;
        RECT 181.950 751.950 184.050 752.400 ;
        RECT 187.950 751.950 190.050 752.400 ;
        RECT 193.950 753.600 196.050 754.050 ;
        RECT 199.950 753.600 202.050 754.050 ;
        RECT 220.950 753.600 223.050 754.050 ;
        RECT 193.950 752.400 223.050 753.600 ;
        RECT 193.950 751.950 196.050 752.400 ;
        RECT 199.950 751.950 202.050 752.400 ;
        RECT 220.950 751.950 223.050 752.400 ;
        RECT 268.950 753.600 271.050 754.050 ;
        RECT 277.950 753.600 280.050 754.050 ;
        RECT 268.950 752.400 280.050 753.600 ;
        RECT 268.950 751.950 271.050 752.400 ;
        RECT 277.950 751.950 280.050 752.400 ;
        RECT 286.950 753.600 289.050 754.050 ;
        RECT 292.950 753.600 295.050 754.050 ;
        RECT 286.950 752.400 295.050 753.600 ;
        RECT 286.950 751.950 289.050 752.400 ;
        RECT 292.950 751.950 295.050 752.400 ;
        RECT 352.950 753.600 355.050 754.050 ;
        RECT 361.950 753.600 364.050 754.050 ;
        RECT 352.950 752.400 364.050 753.600 ;
        RECT 352.950 751.950 355.050 752.400 ;
        RECT 361.950 751.950 364.050 752.400 ;
        RECT 421.950 751.950 424.050 754.050 ;
        RECT 457.950 753.600 460.050 754.050 ;
        RECT 496.950 753.600 499.050 754.050 ;
        RECT 457.950 752.400 499.050 753.600 ;
        RECT 457.950 751.950 460.050 752.400 ;
        RECT 496.950 751.950 499.050 752.400 ;
        RECT 577.950 753.600 580.050 754.050 ;
        RECT 583.800 753.600 585.900 754.050 ;
        RECT 577.950 752.400 585.900 753.600 ;
        RECT 577.950 751.950 580.050 752.400 ;
        RECT 583.800 751.950 585.900 752.400 ;
        RECT 586.950 753.600 589.050 754.050 ;
        RECT 610.950 753.600 613.050 754.050 ;
        RECT 586.950 752.400 613.050 753.600 ;
        RECT 586.950 751.950 589.050 752.400 ;
        RECT 610.950 751.950 613.050 752.400 ;
        RECT 664.950 753.600 667.050 754.050 ;
        RECT 694.950 753.600 697.050 754.050 ;
        RECT 664.950 752.400 697.050 753.600 ;
        RECT 664.950 751.950 667.050 752.400 ;
        RECT 694.950 751.950 697.050 752.400 ;
        RECT 709.950 753.600 712.050 754.050 ;
        RECT 715.950 753.600 718.050 754.050 ;
        RECT 709.950 752.400 718.050 753.600 ;
        RECT 709.950 751.950 712.050 752.400 ;
        RECT 715.950 751.950 718.050 752.400 ;
        RECT 757.950 753.600 760.050 754.050 ;
        RECT 772.950 753.600 775.050 754.050 ;
        RECT 757.950 752.400 775.050 753.600 ;
        RECT 757.950 751.950 760.050 752.400 ;
        RECT 772.950 751.950 775.050 752.400 ;
        RECT 889.950 753.600 892.050 754.050 ;
        RECT 913.950 753.600 916.050 754.050 ;
        RECT 889.950 752.400 916.050 753.600 ;
        RECT 889.950 751.950 892.050 752.400 ;
        RECT 913.950 751.950 916.050 752.400 ;
        RECT 73.950 750.600 76.050 751.050 ;
        RECT 94.950 750.600 97.050 751.050 ;
        RECT 73.950 749.400 97.050 750.600 ;
        RECT 73.950 748.950 76.050 749.400 ;
        RECT 94.950 748.950 97.050 749.400 ;
        RECT 235.950 750.600 238.050 751.050 ;
        RECT 250.950 750.600 253.050 751.050 ;
        RECT 262.950 750.600 265.050 751.050 ;
        RECT 235.950 749.400 265.050 750.600 ;
        RECT 235.950 748.950 238.050 749.400 ;
        RECT 250.950 748.950 253.050 749.400 ;
        RECT 262.950 748.950 265.050 749.400 ;
        RECT 304.950 750.600 307.050 751.050 ;
        RECT 328.950 750.600 331.050 751.050 ;
        RECT 304.950 749.400 331.050 750.600 ;
        RECT 304.950 748.950 307.050 749.400 ;
        RECT 328.950 748.950 331.050 749.400 ;
        RECT 523.950 750.600 526.050 751.050 ;
        RECT 556.950 750.600 559.050 751.050 ;
        RECT 523.950 749.400 559.050 750.600 ;
        RECT 523.950 748.950 526.050 749.400 ;
        RECT 556.950 748.950 559.050 749.400 ;
        RECT 568.950 750.600 571.050 751.050 ;
        RECT 587.400 750.600 588.600 751.950 ;
        RECT 568.950 749.400 588.600 750.600 ;
        RECT 616.950 750.600 619.050 751.050 ;
        RECT 631.950 750.600 634.050 751.050 ;
        RECT 616.950 749.400 634.050 750.600 ;
        RECT 568.950 748.950 571.050 749.400 ;
        RECT 616.950 748.950 619.050 749.400 ;
        RECT 631.950 748.950 634.050 749.400 ;
        RECT 727.950 750.600 730.050 751.050 ;
        RECT 796.950 750.600 799.050 751.050 ;
        RECT 811.950 750.600 814.050 751.050 ;
        RECT 727.950 749.400 795.600 750.600 ;
        RECT 727.950 748.950 730.050 749.400 ;
        RECT 40.950 747.600 43.050 748.050 ;
        RECT 64.950 747.600 67.050 748.050 ;
        RECT 40.950 746.400 67.050 747.600 ;
        RECT 40.950 745.950 43.050 746.400 ;
        RECT 64.950 745.950 67.050 746.400 ;
        RECT 136.950 747.600 139.050 748.050 ;
        RECT 160.950 747.600 163.050 748.050 ;
        RECT 175.950 747.600 178.050 748.050 ;
        RECT 136.950 746.400 159.600 747.600 ;
        RECT 136.950 745.950 139.050 746.400 ;
        RECT 61.950 744.600 64.050 745.050 ;
        RECT 76.950 744.600 79.050 745.050 ;
        RECT 61.950 743.400 79.050 744.600 ;
        RECT 61.950 742.950 64.050 743.400 ;
        RECT 76.950 742.950 79.050 743.400 ;
        RECT 85.950 744.600 88.050 745.050 ;
        RECT 112.950 744.600 115.050 745.050 ;
        RECT 118.800 744.600 120.900 745.050 ;
        RECT 85.950 743.400 120.900 744.600 ;
        RECT 85.950 742.950 88.050 743.400 ;
        RECT 112.950 742.950 115.050 743.400 ;
        RECT 118.800 742.950 120.900 743.400 ;
        RECT 121.950 744.600 124.050 745.050 ;
        RECT 142.950 744.600 145.050 745.050 ;
        RECT 121.950 743.400 145.050 744.600 ;
        RECT 158.400 744.600 159.600 746.400 ;
        RECT 160.950 746.400 178.050 747.600 ;
        RECT 160.950 745.950 163.050 746.400 ;
        RECT 175.950 745.950 178.050 746.400 ;
        RECT 238.950 747.600 241.050 748.050 ;
        RECT 265.950 747.600 268.050 748.050 ;
        RECT 238.950 746.400 268.050 747.600 ;
        RECT 238.950 745.950 241.050 746.400 ;
        RECT 265.950 745.950 268.050 746.400 ;
        RECT 295.950 747.600 298.050 748.050 ;
        RECT 319.950 747.600 322.050 748.050 ;
        RECT 337.950 747.600 340.050 748.050 ;
        RECT 295.950 746.400 340.050 747.600 ;
        RECT 295.950 745.950 298.050 746.400 ;
        RECT 319.950 745.950 322.050 746.400 ;
        RECT 337.950 745.950 340.050 746.400 ;
        RECT 361.950 747.600 364.050 748.050 ;
        RECT 439.950 747.600 442.050 748.050 ;
        RECT 361.950 746.400 442.050 747.600 ;
        RECT 361.950 745.950 364.050 746.400 ;
        RECT 439.950 745.950 442.050 746.400 ;
        RECT 493.950 747.600 496.050 748.050 ;
        RECT 520.950 747.600 523.050 748.050 ;
        RECT 493.950 746.400 523.050 747.600 ;
        RECT 493.950 745.950 496.050 746.400 ;
        RECT 520.950 745.950 523.050 746.400 ;
        RECT 532.950 747.600 535.050 748.050 ;
        RECT 538.950 747.600 541.050 748.050 ;
        RECT 532.950 746.400 541.050 747.600 ;
        RECT 532.950 745.950 535.050 746.400 ;
        RECT 538.950 745.950 541.050 746.400 ;
        RECT 547.950 747.600 550.050 748.050 ;
        RECT 562.950 747.600 565.050 748.050 ;
        RECT 547.950 746.400 565.050 747.600 ;
        RECT 547.950 745.950 550.050 746.400 ;
        RECT 562.950 745.950 565.050 746.400 ;
        RECT 571.950 747.600 574.050 748.050 ;
        RECT 601.950 747.600 604.050 748.050 ;
        RECT 613.950 747.600 616.050 748.050 ;
        RECT 640.950 747.600 643.050 748.050 ;
        RECT 571.950 746.400 643.050 747.600 ;
        RECT 571.950 745.950 574.050 746.400 ;
        RECT 601.950 745.950 604.050 746.400 ;
        RECT 613.950 745.950 616.050 746.400 ;
        RECT 640.950 745.950 643.050 746.400 ;
        RECT 655.950 747.600 658.050 748.050 ;
        RECT 667.950 747.600 670.050 748.050 ;
        RECT 700.950 747.600 703.050 748.050 ;
        RECT 655.950 746.400 703.050 747.600 ;
        RECT 655.950 745.950 658.050 746.400 ;
        RECT 667.950 745.950 670.050 746.400 ;
        RECT 700.950 745.950 703.050 746.400 ;
        RECT 709.950 747.600 712.050 748.050 ;
        RECT 724.950 747.600 727.050 748.050 ;
        RECT 709.950 746.400 727.050 747.600 ;
        RECT 709.950 745.950 712.050 746.400 ;
        RECT 724.950 745.950 727.050 746.400 ;
        RECT 742.950 747.600 745.050 748.050 ;
        RECT 781.950 747.600 784.050 748.050 ;
        RECT 742.950 746.400 784.050 747.600 ;
        RECT 794.400 747.600 795.600 749.400 ;
        RECT 796.950 749.400 814.050 750.600 ;
        RECT 796.950 748.950 799.050 749.400 ;
        RECT 811.950 748.950 814.050 749.400 ;
        RECT 859.950 750.600 862.050 751.050 ;
        RECT 874.950 750.600 877.050 751.050 ;
        RECT 859.950 749.400 877.050 750.600 ;
        RECT 859.950 748.950 862.050 749.400 ;
        RECT 874.950 748.950 877.050 749.400 ;
        RECT 880.950 750.600 883.050 751.050 ;
        RECT 886.950 750.600 889.050 751.050 ;
        RECT 910.950 750.600 913.050 751.050 ;
        RECT 880.950 749.400 913.050 750.600 ;
        RECT 880.950 748.950 883.050 749.400 ;
        RECT 886.950 748.950 889.050 749.400 ;
        RECT 910.950 748.950 913.050 749.400 ;
        RECT 799.950 747.600 802.050 748.050 ;
        RECT 794.400 746.400 802.050 747.600 ;
        RECT 742.950 745.950 745.050 746.400 ;
        RECT 781.950 745.950 784.050 746.400 ;
        RECT 799.950 745.950 802.050 746.400 ;
        RECT 805.950 747.600 808.050 748.050 ;
        RECT 814.950 747.600 817.050 748.050 ;
        RECT 805.950 746.400 817.050 747.600 ;
        RECT 805.950 745.950 808.050 746.400 ;
        RECT 814.950 745.950 817.050 746.400 ;
        RECT 847.950 747.600 850.050 748.050 ;
        RECT 856.950 747.600 859.050 748.050 ;
        RECT 847.950 746.400 859.050 747.600 ;
        RECT 847.950 745.950 850.050 746.400 ;
        RECT 856.950 745.950 859.050 746.400 ;
        RECT 259.950 744.600 262.050 745.050 ;
        RECT 158.400 743.400 262.050 744.600 ;
        RECT 121.950 742.950 124.050 743.400 ;
        RECT 142.950 742.950 145.050 743.400 ;
        RECT 259.950 742.950 262.050 743.400 ;
        RECT 343.950 744.600 346.050 745.050 ;
        RECT 424.950 744.600 427.050 745.050 ;
        RECT 442.950 744.600 445.050 745.050 ;
        RECT 457.950 744.600 460.050 745.050 ;
        RECT 343.950 743.400 460.050 744.600 ;
        RECT 343.950 742.950 346.050 743.400 ;
        RECT 424.950 742.950 427.050 743.400 ;
        RECT 442.950 742.950 445.050 743.400 ;
        RECT 457.950 742.950 460.050 743.400 ;
        RECT 481.950 744.600 484.050 745.050 ;
        RECT 508.950 744.600 511.050 745.050 ;
        RECT 481.950 743.400 511.050 744.600 ;
        RECT 481.950 742.950 484.050 743.400 ;
        RECT 508.950 742.950 511.050 743.400 ;
        RECT 628.950 744.600 631.050 745.050 ;
        RECT 634.950 744.600 637.050 745.050 ;
        RECT 628.950 743.400 637.050 744.600 ;
        RECT 628.950 742.950 631.050 743.400 ;
        RECT 634.950 742.950 637.050 743.400 ;
        RECT 646.950 744.600 649.050 745.050 ;
        RECT 682.950 744.600 685.050 745.050 ;
        RECT 646.950 743.400 685.050 744.600 ;
        RECT 701.400 744.600 702.600 745.950 ;
        RECT 706.950 744.600 709.050 745.050 ;
        RECT 701.400 743.400 709.050 744.600 ;
        RECT 646.950 742.950 649.050 743.400 ;
        RECT 682.950 742.950 685.050 743.400 ;
        RECT 706.950 742.950 709.050 743.400 ;
        RECT 769.950 744.600 772.050 745.050 ;
        RECT 802.950 744.600 805.050 745.050 ;
        RECT 769.950 743.400 805.050 744.600 ;
        RECT 769.950 742.950 772.050 743.400 ;
        RECT 802.950 742.950 805.050 743.400 ;
        RECT 151.950 741.600 154.050 742.050 ;
        RECT 190.950 741.600 193.050 742.050 ;
        RECT 151.950 740.400 193.050 741.600 ;
        RECT 151.950 739.950 154.050 740.400 ;
        RECT 190.950 739.950 193.050 740.400 ;
        RECT 217.950 741.600 220.050 742.050 ;
        RECT 256.950 741.600 259.050 742.050 ;
        RECT 217.950 740.400 259.050 741.600 ;
        RECT 217.950 739.950 220.050 740.400 ;
        RECT 256.950 739.950 259.050 740.400 ;
        RECT 475.950 741.600 478.050 742.050 ;
        RECT 493.950 741.600 496.050 742.050 ;
        RECT 475.950 740.400 496.050 741.600 ;
        RECT 475.950 739.950 478.050 740.400 ;
        RECT 493.950 739.950 496.050 740.400 ;
        RECT 520.950 741.600 523.050 742.050 ;
        RECT 565.950 741.600 568.050 742.050 ;
        RECT 571.950 741.600 574.050 742.050 ;
        RECT 520.950 740.400 574.050 741.600 ;
        RECT 520.950 739.950 523.050 740.400 ;
        RECT 565.950 739.950 568.050 740.400 ;
        RECT 571.950 739.950 574.050 740.400 ;
        RECT 619.950 741.600 622.050 742.050 ;
        RECT 643.950 741.600 646.050 742.050 ;
        RECT 619.950 740.400 646.050 741.600 ;
        RECT 619.950 739.950 622.050 740.400 ;
        RECT 643.950 739.950 646.050 740.400 ;
        RECT 691.950 741.600 694.050 742.050 ;
        RECT 709.950 741.600 712.050 742.050 ;
        RECT 691.950 740.400 712.050 741.600 ;
        RECT 691.950 739.950 694.050 740.400 ;
        RECT 709.950 739.950 712.050 740.400 ;
        RECT 715.950 741.600 718.050 742.050 ;
        RECT 748.950 741.600 751.050 742.050 ;
        RECT 715.950 740.400 751.050 741.600 ;
        RECT 715.950 739.950 718.050 740.400 ;
        RECT 748.950 739.950 751.050 740.400 ;
        RECT 805.950 741.600 808.050 742.050 ;
        RECT 838.950 741.600 841.050 742.050 ;
        RECT 805.950 740.400 841.050 741.600 ;
        RECT 805.950 739.950 808.050 740.400 ;
        RECT 838.950 739.950 841.050 740.400 ;
        RECT 196.950 738.600 199.050 739.050 ;
        RECT 247.950 738.600 250.050 739.050 ;
        RECT 196.950 737.400 250.050 738.600 ;
        RECT 196.950 736.950 199.050 737.400 ;
        RECT 247.950 736.950 250.050 737.400 ;
        RECT 358.950 738.600 361.050 739.050 ;
        RECT 370.950 738.600 373.050 739.050 ;
        RECT 376.800 738.600 378.900 739.050 ;
        RECT 358.950 737.400 378.900 738.600 ;
        RECT 358.950 736.950 361.050 737.400 ;
        RECT 370.950 736.950 373.050 737.400 ;
        RECT 376.800 736.950 378.900 737.400 ;
        RECT 379.950 738.600 382.050 739.050 ;
        RECT 388.950 738.600 391.050 739.050 ;
        RECT 379.950 737.400 391.050 738.600 ;
        RECT 379.950 736.950 382.050 737.400 ;
        RECT 388.950 736.950 391.050 737.400 ;
        RECT 469.950 738.600 472.050 739.050 ;
        RECT 508.950 738.600 511.050 739.050 ;
        RECT 469.950 737.400 511.050 738.600 ;
        RECT 469.950 736.950 472.050 737.400 ;
        RECT 508.950 736.950 511.050 737.400 ;
        RECT 517.950 738.600 520.050 739.050 ;
        RECT 568.950 738.600 571.050 739.050 ;
        RECT 517.950 737.400 571.050 738.600 ;
        RECT 517.950 736.950 520.050 737.400 ;
        RECT 568.950 736.950 571.050 737.400 ;
        RECT 589.950 738.600 592.050 739.050 ;
        RECT 598.950 738.600 601.050 739.050 ;
        RECT 589.950 737.400 601.050 738.600 ;
        RECT 589.950 736.950 592.050 737.400 ;
        RECT 598.950 736.950 601.050 737.400 ;
        RECT 607.950 738.600 610.050 739.050 ;
        RECT 616.950 738.600 619.050 739.050 ;
        RECT 607.950 737.400 619.050 738.600 ;
        RECT 607.950 736.950 610.050 737.400 ;
        RECT 616.950 736.950 619.050 737.400 ;
        RECT 628.950 738.600 631.050 739.050 ;
        RECT 694.950 738.600 697.050 739.050 ;
        RECT 628.950 737.400 697.050 738.600 ;
        RECT 628.950 736.950 631.050 737.400 ;
        RECT 694.950 736.950 697.050 737.400 ;
        RECT 754.950 738.600 757.050 739.050 ;
        RECT 766.950 738.600 769.050 739.050 ;
        RECT 754.950 737.400 769.050 738.600 ;
        RECT 754.950 736.950 757.050 737.400 ;
        RECT 766.950 736.950 769.050 737.400 ;
        RECT 901.950 738.600 904.050 739.050 ;
        RECT 901.950 737.400 918.600 738.600 ;
        RECT 901.950 736.950 904.050 737.400 ;
        RECT 917.400 736.050 918.600 737.400 ;
        RECT 58.950 735.600 61.050 736.050 ;
        RECT 73.950 735.600 76.050 736.050 ;
        RECT 58.950 734.400 76.050 735.600 ;
        RECT 58.950 733.950 61.050 734.400 ;
        RECT 73.950 733.950 76.050 734.400 ;
        RECT 232.950 735.600 235.050 736.050 ;
        RECT 253.950 735.600 256.050 736.050 ;
        RECT 271.950 735.600 274.050 736.050 ;
        RECT 232.950 734.400 274.050 735.600 ;
        RECT 232.950 733.950 235.050 734.400 ;
        RECT 253.950 733.950 256.050 734.400 ;
        RECT 271.950 733.950 274.050 734.400 ;
        RECT 310.950 735.600 313.050 736.050 ;
        RECT 322.950 735.600 325.050 736.050 ;
        RECT 310.950 734.400 325.050 735.600 ;
        RECT 310.950 733.950 313.050 734.400 ;
        RECT 322.950 733.950 325.050 734.400 ;
        RECT 352.950 735.600 355.050 736.050 ;
        RECT 364.950 735.600 367.050 736.050 ;
        RECT 352.950 734.400 367.050 735.600 ;
        RECT 352.950 733.950 355.050 734.400 ;
        RECT 364.950 733.950 367.050 734.400 ;
        RECT 391.950 735.600 394.050 736.050 ;
        RECT 418.950 735.600 421.050 736.050 ;
        RECT 391.950 734.400 421.050 735.600 ;
        RECT 391.950 733.950 394.050 734.400 ;
        RECT 418.950 733.950 421.050 734.400 ;
        RECT 424.950 735.600 427.050 736.050 ;
        RECT 448.950 735.600 451.050 736.050 ;
        RECT 457.950 735.600 460.050 736.050 ;
        RECT 424.950 734.400 460.050 735.600 ;
        RECT 424.950 733.950 427.050 734.400 ;
        RECT 448.950 733.950 451.050 734.400 ;
        RECT 457.950 733.950 460.050 734.400 ;
        RECT 514.950 735.600 517.050 736.050 ;
        RECT 586.950 735.600 589.050 736.050 ;
        RECT 514.950 734.400 589.050 735.600 ;
        RECT 514.950 733.950 517.050 734.400 ;
        RECT 586.950 733.950 589.050 734.400 ;
        RECT 625.950 735.600 628.050 736.050 ;
        RECT 658.950 735.600 661.050 736.050 ;
        RECT 625.950 734.400 661.050 735.600 ;
        RECT 625.950 733.950 628.050 734.400 ;
        RECT 658.950 733.950 661.050 734.400 ;
        RECT 682.950 735.600 685.050 736.050 ;
        RECT 697.950 735.600 700.050 736.050 ;
        RECT 682.950 734.400 700.050 735.600 ;
        RECT 682.950 733.950 685.050 734.400 ;
        RECT 697.950 733.950 700.050 734.400 ;
        RECT 739.950 735.600 742.050 736.050 ;
        RECT 799.950 735.600 802.050 736.050 ;
        RECT 739.950 734.400 802.050 735.600 ;
        RECT 739.950 733.950 742.050 734.400 ;
        RECT 799.950 733.950 802.050 734.400 ;
        RECT 844.950 735.600 847.050 736.050 ;
        RECT 856.950 735.600 859.050 735.900 ;
        RECT 844.950 734.400 859.050 735.600 ;
        RECT 917.400 734.400 922.050 736.050 ;
        RECT 844.950 733.950 847.050 734.400 ;
        RECT 856.950 733.800 859.050 734.400 ;
        RECT 918.000 733.950 922.050 734.400 ;
        RECT 25.950 732.600 28.050 733.050 ;
        RECT 34.950 732.600 37.050 733.050 ;
        RECT 82.950 732.600 85.050 733.050 ;
        RECT 103.950 732.600 106.050 733.050 ;
        RECT 151.950 732.600 154.050 733.050 ;
        RECT 25.950 731.400 106.050 732.600 ;
        RECT 25.950 730.950 28.050 731.400 ;
        RECT 34.950 730.950 37.050 731.400 ;
        RECT 82.950 730.950 85.050 731.400 ;
        RECT 103.950 730.950 106.050 731.400 ;
        RECT 146.400 731.400 154.050 732.600 ;
        RECT 16.950 729.600 19.050 730.200 ;
        RECT 40.950 729.600 43.050 730.200 ;
        RECT 46.950 729.600 49.050 730.050 ;
        RECT 16.950 728.400 24.600 729.600 ;
        RECT 16.950 728.100 19.050 728.400 ;
        RECT 23.400 724.050 24.600 728.400 ;
        RECT 40.950 728.400 49.050 729.600 ;
        RECT 40.950 728.100 43.050 728.400 ;
        RECT 46.950 727.950 49.050 728.400 ;
        RECT 55.950 729.750 58.050 730.200 ;
        RECT 70.950 729.750 73.050 730.200 ;
        RECT 55.950 728.550 73.050 729.750 ;
        RECT 88.950 729.600 91.050 730.200 ;
        RECT 55.950 728.100 58.050 728.550 ;
        RECT 70.950 728.100 73.050 728.550 ;
        RECT 86.400 728.400 91.050 729.600 ;
        RECT 86.400 726.600 87.600 728.400 ;
        RECT 88.950 728.100 91.050 728.400 ;
        RECT 109.950 729.600 112.050 730.200 ;
        RECT 127.950 729.600 130.050 730.200 ;
        RECT 109.950 728.400 130.050 729.600 ;
        RECT 109.950 728.100 112.050 728.400 ;
        RECT 127.950 728.100 130.050 728.400 ;
        RECT 146.400 726.600 147.600 731.400 ;
        RECT 151.950 730.950 154.050 731.400 ;
        RECT 349.950 730.950 352.050 733.050 ;
        RECT 388.950 732.600 391.050 733.050 ;
        RECT 553.950 732.600 556.050 733.050 ;
        RECT 388.950 731.400 402.600 732.600 ;
        RECT 388.950 730.950 391.050 731.400 ;
        RECT 163.950 729.750 166.050 730.200 ;
        RECT 166.950 729.750 169.050 730.050 ;
        RECT 169.950 729.750 172.050 730.200 ;
        RECT 163.950 728.550 172.050 729.750 ;
        RECT 163.950 728.100 166.050 728.550 ;
        RECT 166.950 727.950 169.050 728.550 ;
        RECT 169.950 728.100 172.050 728.550 ;
        RECT 178.950 729.600 181.050 730.050 ;
        RECT 196.950 729.600 199.050 730.050 ;
        RECT 178.950 728.400 199.050 729.600 ;
        RECT 178.950 727.950 181.050 728.400 ;
        RECT 196.950 727.950 199.050 728.400 ;
        RECT 202.950 729.750 205.050 730.200 ;
        RECT 211.950 729.750 214.050 730.200 ;
        RECT 202.950 728.550 214.050 729.750 ;
        RECT 202.950 728.100 205.050 728.550 ;
        RECT 211.950 728.100 214.050 728.550 ;
        RECT 238.950 729.600 241.050 730.050 ;
        RECT 247.950 729.600 250.050 730.200 ;
        RECT 238.950 728.400 250.050 729.600 ;
        RECT 238.950 727.950 241.050 728.400 ;
        RECT 247.950 728.100 250.050 728.400 ;
        RECT 271.950 728.100 274.050 730.200 ;
        RECT 331.950 729.600 334.050 730.200 ;
        RECT 340.950 729.600 343.050 730.050 ;
        RECT 331.950 728.400 343.050 729.600 ;
        RECT 331.950 728.100 334.050 728.400 ;
        RECT 77.400 725.400 87.600 726.600 ;
        RECT 131.400 725.400 147.600 726.600 ;
        RECT 272.400 726.600 273.600 728.100 ;
        RECT 340.950 727.950 343.050 728.400 ;
        RECT 272.400 725.400 294.600 726.600 ;
        RECT 22.950 721.950 25.050 724.050 ;
        RECT 46.950 723.450 49.050 723.900 ;
        RECT 58.950 723.450 61.050 723.900 ;
        RECT 46.950 722.250 61.050 723.450 ;
        RECT 46.950 721.800 49.050 722.250 ;
        RECT 58.950 721.800 61.050 722.250 ;
        RECT 64.950 723.600 67.050 723.900 ;
        RECT 77.400 723.600 78.600 725.400 ;
        RECT 97.950 723.600 100.050 724.050 ;
        RECT 121.950 723.600 124.050 724.050 ;
        RECT 131.400 723.900 132.600 725.400 ;
        RECT 146.400 723.900 147.600 725.400 ;
        RECT 64.950 723.000 84.600 723.600 ;
        RECT 64.950 722.400 85.050 723.000 ;
        RECT 64.950 721.800 67.050 722.400 ;
        RECT 19.950 720.600 22.050 721.050 ;
        RECT 25.950 720.600 28.050 721.050 ;
        RECT 19.950 719.400 28.050 720.600 ;
        RECT 19.950 718.950 22.050 719.400 ;
        RECT 25.950 718.950 28.050 719.400 ;
        RECT 82.950 718.950 85.050 722.400 ;
        RECT 97.950 722.400 124.050 723.600 ;
        RECT 97.950 721.950 100.050 722.400 ;
        RECT 121.950 721.950 124.050 722.400 ;
        RECT 130.950 721.800 133.050 723.900 ;
        RECT 145.950 721.800 148.050 723.900 ;
        RECT 151.950 723.600 154.050 723.900 ;
        RECT 172.950 723.600 175.050 723.900 ;
        RECT 151.950 722.400 175.050 723.600 ;
        RECT 151.950 721.800 154.050 722.400 ;
        RECT 172.950 721.800 175.050 722.400 ;
        RECT 229.950 723.600 232.050 723.900 ;
        RECT 256.950 723.600 259.050 724.050 ;
        RECT 277.950 723.600 280.050 723.900 ;
        RECT 229.950 723.450 280.050 723.600 ;
        RECT 286.950 723.450 289.050 723.900 ;
        RECT 229.950 722.400 289.050 723.450 ;
        RECT 293.400 723.600 294.600 725.400 ;
        RECT 295.950 723.600 298.050 723.900 ;
        RECT 293.400 722.400 298.050 723.600 ;
        RECT 229.950 721.800 232.050 722.400 ;
        RECT 256.950 721.950 259.050 722.400 ;
        RECT 277.950 722.250 289.050 722.400 ;
        RECT 277.950 721.800 280.050 722.250 ;
        RECT 286.950 721.800 289.050 722.250 ;
        RECT 295.950 721.800 298.050 722.400 ;
        RECT 310.950 723.600 313.050 723.900 ;
        RECT 328.950 723.600 331.050 723.900 ;
        RECT 310.950 722.400 331.050 723.600 ;
        RECT 310.950 721.800 313.050 722.400 ;
        RECT 328.950 721.800 331.050 722.400 ;
        RECT 334.950 723.450 337.050 723.900 ;
        RECT 343.950 723.450 346.050 723.900 ;
        RECT 334.950 722.250 346.050 723.450 ;
        RECT 350.400 723.600 351.600 730.950 ;
        RECT 361.950 723.600 364.050 724.050 ;
        RECT 401.400 723.900 402.600 731.400 ;
        RECT 553.950 731.400 573.600 732.600 ;
        RECT 553.950 730.950 556.050 731.400 ;
        RECT 412.950 729.600 415.050 730.050 ;
        RECT 424.950 729.600 427.050 730.200 ;
        RECT 412.950 728.400 427.050 729.600 ;
        RECT 412.950 727.950 415.050 728.400 ;
        RECT 424.950 728.100 427.050 728.400 ;
        RECT 430.950 728.100 433.050 730.200 ;
        RECT 454.950 729.600 457.050 730.200 ;
        RECT 472.950 729.600 475.050 730.200 ;
        RECT 484.950 729.600 487.050 730.050 ;
        RECT 454.950 728.400 468.600 729.600 ;
        RECT 454.950 728.100 457.050 728.400 ;
        RECT 431.400 726.600 432.600 728.100 ;
        RECT 431.400 725.400 450.600 726.600 ;
        RECT 350.400 722.400 364.050 723.600 ;
        RECT 334.950 721.800 337.050 722.250 ;
        RECT 343.950 721.800 346.050 722.250 ;
        RECT 361.950 721.950 364.050 722.400 ;
        RECT 400.950 721.800 403.050 723.900 ;
        RECT 406.950 723.450 409.050 723.900 ;
        RECT 412.950 723.450 415.050 723.900 ;
        RECT 406.950 722.250 415.050 723.450 ;
        RECT 406.950 721.800 409.050 722.250 ;
        RECT 412.950 721.800 415.050 722.250 ;
        RECT 418.950 723.450 421.050 724.050 ;
        RECT 427.950 723.450 430.050 723.900 ;
        RECT 418.950 722.250 430.050 723.450 ;
        RECT 449.400 723.600 450.600 725.400 ;
        RECT 449.400 722.400 453.600 723.600 ;
        RECT 418.950 721.950 421.050 722.250 ;
        RECT 427.950 721.800 430.050 722.250 ;
        RECT 452.400 721.050 453.600 722.400 ;
        RECT 199.950 720.600 202.050 721.050 ;
        RECT 217.950 720.600 220.050 721.050 ;
        RECT 289.950 720.600 292.050 721.050 ;
        RECT 199.950 719.400 292.050 720.600 ;
        RECT 199.950 718.950 202.050 719.400 ;
        RECT 217.950 718.950 220.050 719.400 ;
        RECT 289.950 718.950 292.050 719.400 ;
        RECT 355.950 720.600 358.050 721.050 ;
        RECT 391.950 720.600 394.050 721.050 ;
        RECT 355.950 719.400 394.050 720.600 ;
        RECT 355.950 718.950 358.050 719.400 ;
        RECT 391.950 718.950 394.050 719.400 ;
        RECT 427.950 720.600 430.050 721.050 ;
        RECT 445.950 720.600 448.050 721.050 ;
        RECT 427.950 719.400 448.050 720.600 ;
        RECT 452.400 719.400 457.050 721.050 ;
        RECT 467.400 720.600 468.600 728.400 ;
        RECT 472.950 728.400 487.050 729.600 ;
        RECT 472.950 728.100 475.050 728.400 ;
        RECT 484.950 727.950 487.050 728.400 ;
        RECT 532.950 729.600 535.050 730.200 ;
        RECT 541.950 729.600 544.050 730.050 ;
        RECT 532.950 728.400 544.050 729.600 ;
        RECT 532.950 728.100 535.050 728.400 ;
        RECT 541.950 727.950 544.050 728.400 ;
        RECT 547.950 729.600 550.050 730.050 ;
        RECT 556.950 729.600 559.050 730.200 ;
        RECT 547.950 728.400 559.050 729.600 ;
        RECT 547.950 727.950 550.050 728.400 ;
        RECT 556.950 728.100 559.050 728.400 ;
        RECT 562.950 727.950 565.050 730.050 ;
        RECT 478.950 723.450 481.050 723.900 ;
        RECT 493.950 723.450 496.050 723.900 ;
        RECT 478.950 722.250 496.050 723.450 ;
        RECT 478.950 721.800 481.050 722.250 ;
        RECT 493.950 721.800 496.050 722.250 ;
        RECT 475.950 720.600 478.050 721.050 ;
        RECT 467.400 719.400 478.050 720.600 ;
        RECT 563.400 720.600 564.600 727.950 ;
        RECT 572.400 723.900 573.600 731.400 ;
        RECT 595.950 730.950 598.050 733.050 ;
        RECT 604.950 732.600 607.050 733.050 ;
        RECT 628.950 732.600 631.050 733.050 ;
        RECT 604.950 731.400 631.050 732.600 ;
        RECT 604.950 730.950 607.050 731.400 ;
        RECT 574.950 729.600 577.050 730.200 ;
        RECT 574.950 728.400 582.600 729.600 ;
        RECT 574.950 728.100 577.050 728.400 ;
        RECT 581.400 724.050 582.600 728.400 ;
        RECT 571.950 721.800 574.050 723.900 ;
        RECT 580.950 721.950 583.050 724.050 ;
        RECT 596.400 723.900 597.600 730.950 ;
        RECT 598.950 729.600 601.050 730.200 ;
        RECT 610.950 729.750 613.050 730.200 ;
        RECT 619.950 729.750 622.050 730.200 ;
        RECT 598.950 728.400 609.600 729.600 ;
        RECT 598.950 728.100 601.050 728.400 ;
        RECT 608.400 726.600 609.600 728.400 ;
        RECT 610.950 728.550 622.050 729.750 ;
        RECT 610.950 728.100 613.050 728.550 ;
        RECT 619.950 728.100 622.050 728.550 ;
        RECT 608.400 725.400 624.600 726.600 ;
        RECT 595.950 721.800 598.050 723.900 ;
        RECT 601.950 723.600 604.050 723.900 ;
        RECT 610.950 723.600 613.050 724.050 ;
        RECT 623.400 723.900 624.600 725.400 ;
        RECT 601.950 722.400 613.050 723.600 ;
        RECT 601.950 721.800 604.050 722.400 ;
        RECT 610.950 721.950 613.050 722.400 ;
        RECT 622.950 721.800 625.050 723.900 ;
        RECT 626.400 721.050 627.600 731.400 ;
        RECT 628.950 730.950 631.050 731.400 ;
        RECT 670.950 732.600 673.050 733.050 ;
        RECT 676.950 732.600 679.050 733.050 ;
        RECT 670.950 731.400 679.050 732.600 ;
        RECT 670.950 730.950 673.050 731.400 ;
        RECT 676.950 730.950 679.050 731.400 ;
        RECT 709.950 732.600 712.050 733.050 ;
        RECT 727.950 732.600 730.050 733.050 ;
        RECT 709.950 731.400 730.050 732.600 ;
        RECT 709.950 730.950 712.050 731.400 ;
        RECT 727.950 730.950 730.050 731.400 ;
        RECT 775.950 732.600 778.050 733.050 ;
        RECT 784.950 732.600 787.050 733.050 ;
        RECT 790.950 732.600 793.050 733.050 ;
        RECT 775.950 731.400 793.050 732.600 ;
        RECT 775.950 730.950 778.050 731.400 ;
        RECT 784.950 730.950 787.050 731.400 ;
        RECT 790.950 730.950 793.050 731.400 ;
        RECT 628.950 727.800 631.050 729.900 ;
        RECT 664.950 728.100 667.050 730.200 ;
        RECT 629.400 724.050 630.600 727.800 ;
        RECT 631.950 726.600 634.050 727.050 ;
        RECT 665.400 726.600 666.600 728.100 ;
        RECT 673.950 727.950 676.050 730.050 ;
        RECT 682.950 728.100 685.050 730.200 ;
        RECT 688.950 729.600 691.050 730.200 ;
        RECT 706.950 729.600 709.050 730.200 ;
        RECT 712.950 729.600 715.050 730.200 ;
        RECT 688.950 728.400 709.050 729.600 ;
        RECT 688.950 728.100 691.050 728.400 ;
        RECT 706.950 728.100 709.050 728.400 ;
        RECT 710.400 728.400 715.050 729.600 ;
        RECT 631.950 725.400 666.600 726.600 ;
        RECT 631.950 724.950 634.050 725.400 ;
        RECT 628.950 721.950 631.050 724.050 ;
        RECT 646.950 723.600 649.050 723.900 ;
        RECT 661.950 723.600 664.050 723.900 ;
        RECT 667.950 723.600 670.050 724.050 ;
        RECT 646.950 722.400 670.050 723.600 ;
        RECT 646.950 721.800 649.050 722.400 ;
        RECT 661.950 721.800 664.050 722.400 ;
        RECT 667.950 721.950 670.050 722.400 ;
        RECT 568.950 720.600 571.050 721.050 ;
        RECT 563.400 719.400 571.050 720.600 ;
        RECT 427.950 718.950 430.050 719.400 ;
        RECT 445.950 718.950 448.050 719.400 ;
        RECT 453.000 718.950 457.050 719.400 ;
        RECT 475.950 718.950 478.050 719.400 ;
        RECT 568.950 718.950 571.050 719.400 ;
        RECT 616.950 720.600 619.050 721.050 ;
        RECT 625.950 720.600 628.050 721.050 ;
        RECT 616.950 719.400 628.050 720.600 ;
        RECT 674.400 720.600 675.600 727.950 ;
        RECT 683.400 726.600 684.600 728.100 ;
        RECT 680.400 726.000 684.600 726.600 ;
        RECT 679.950 725.400 684.600 726.000 ;
        RECT 700.950 726.600 703.050 726.900 ;
        RECT 710.400 726.600 711.600 728.400 ;
        RECT 712.950 728.100 715.050 728.400 ;
        RECT 739.950 729.600 742.050 730.050 ;
        RECT 748.950 729.600 751.050 730.200 ;
        RECT 754.950 729.600 757.050 730.200 ;
        RECT 739.950 728.400 751.050 729.600 ;
        RECT 739.950 727.950 742.050 728.400 ;
        RECT 748.950 728.100 751.050 728.400 ;
        RECT 752.400 728.400 757.050 729.600 ;
        RECT 752.400 726.600 753.600 728.400 ;
        RECT 754.950 728.100 757.050 728.400 ;
        RECT 760.950 727.950 763.050 730.050 ;
        RECT 769.950 729.600 772.050 730.050 ;
        RECT 778.950 729.600 781.050 730.200 ;
        RECT 769.950 728.400 781.050 729.600 ;
        RECT 769.950 727.950 772.050 728.400 ;
        RECT 778.950 728.100 781.050 728.400 ;
        RECT 787.950 727.950 790.050 730.050 ;
        RECT 817.950 729.600 820.050 733.050 ;
        RECT 835.950 732.600 838.050 733.050 ;
        RECT 841.950 732.600 844.050 733.050 ;
        RECT 835.950 731.400 844.050 732.600 ;
        RECT 835.950 730.950 838.050 731.400 ;
        RECT 841.950 730.950 844.050 731.400 ;
        RECT 862.950 732.600 865.050 733.050 ;
        RECT 862.950 731.400 870.600 732.600 ;
        RECT 862.950 730.950 865.050 731.400 ;
        RECT 826.950 729.600 829.050 730.200 ;
        RECT 817.950 729.000 829.050 729.600 ;
        RECT 818.400 728.400 829.050 729.000 ;
        RECT 826.950 728.100 829.050 728.400 ;
        RECT 832.950 727.950 835.050 730.050 ;
        RECT 700.950 725.400 711.600 726.600 ;
        RECT 749.400 725.400 753.600 726.600 ;
        RECT 679.950 721.950 682.050 725.400 ;
        RECT 700.950 724.800 703.050 725.400 ;
        RECT 715.950 723.600 718.050 723.900 ;
        RECT 733.950 723.600 736.050 723.900 ;
        RECT 715.950 722.400 736.050 723.600 ;
        RECT 715.950 721.800 718.050 722.400 ;
        RECT 733.950 721.800 736.050 722.400 ;
        RECT 749.400 721.050 750.600 725.400 ;
        RECT 761.400 724.050 762.600 727.950 ;
        RECT 760.950 721.950 763.050 724.050 ;
        RECT 766.950 723.450 769.050 723.900 ;
        RECT 775.950 723.450 778.050 723.900 ;
        RECT 788.400 723.600 789.600 727.950 ;
        RECT 833.400 724.050 834.600 727.950 ;
        RECT 838.950 726.600 841.050 730.050 ;
        RECT 865.950 728.100 868.050 730.200 ;
        RECT 866.400 726.600 867.600 728.100 ;
        RECT 838.950 726.000 846.600 726.600 ;
        RECT 863.400 726.000 867.600 726.600 ;
        RECT 839.400 725.400 846.600 726.000 ;
        RECT 766.950 722.250 778.050 723.450 ;
        RECT 785.400 723.000 789.600 723.600 ;
        RECT 766.950 721.800 769.050 722.250 ;
        RECT 775.950 721.800 778.050 722.250 ;
        RECT 784.950 722.400 789.600 723.000 ;
        RECT 790.950 723.450 793.050 723.900 ;
        RECT 796.950 723.450 799.050 723.900 ;
        RECT 682.950 720.600 685.050 721.050 ;
        RECT 674.400 719.400 685.050 720.600 ;
        RECT 616.950 718.950 619.050 719.400 ;
        RECT 625.950 718.950 628.050 719.400 ;
        RECT 682.950 718.950 685.050 719.400 ;
        RECT 748.950 718.950 751.050 721.050 ;
        RECT 784.950 718.950 787.050 722.400 ;
        RECT 790.950 722.250 799.050 723.450 ;
        RECT 790.950 721.800 793.050 722.250 ;
        RECT 796.950 721.800 799.050 722.250 ;
        RECT 811.950 723.450 814.050 723.900 ;
        RECT 823.950 723.450 826.050 723.900 ;
        RECT 811.950 722.250 826.050 723.450 ;
        RECT 811.950 721.800 814.050 722.250 ;
        RECT 823.950 721.800 826.050 722.250 ;
        RECT 832.950 721.950 835.050 724.050 ;
        RECT 845.400 723.900 846.600 725.400 ;
        RECT 862.950 725.400 867.600 726.000 ;
        RECT 869.400 726.600 870.600 731.400 ;
        RECT 871.950 729.600 874.050 730.200 ;
        RECT 913.950 729.600 916.050 730.050 ;
        RECT 871.950 728.400 916.050 729.600 ;
        RECT 871.950 728.100 874.050 728.400 ;
        RECT 913.950 727.950 916.050 728.400 ;
        RECT 869.400 725.400 876.600 726.600 ;
        RECT 844.950 721.800 847.050 723.900 ;
        RECT 862.950 721.950 865.050 725.400 ;
        RECT 875.400 723.900 876.600 725.400 ;
        RECT 874.950 721.800 877.050 723.900 ;
        RECT 37.950 717.600 40.050 718.050 ;
        RECT 49.950 717.600 52.050 718.050 ;
        RECT 37.950 716.400 52.050 717.600 ;
        RECT 37.950 715.950 40.050 716.400 ;
        RECT 49.950 715.950 52.050 716.400 ;
        RECT 106.950 717.600 109.050 718.050 ;
        RECT 130.950 717.600 133.050 718.050 ;
        RECT 106.950 716.400 133.050 717.600 ;
        RECT 106.950 715.950 109.050 716.400 ;
        RECT 130.950 715.950 133.050 716.400 ;
        RECT 187.950 717.600 190.050 718.050 ;
        RECT 208.950 717.600 211.050 718.050 ;
        RECT 187.950 716.400 211.050 717.600 ;
        RECT 187.950 715.950 190.050 716.400 ;
        RECT 208.950 715.950 211.050 716.400 ;
        RECT 244.950 717.600 247.050 718.050 ;
        RECT 280.950 717.600 283.050 718.050 ;
        RECT 244.950 716.400 283.050 717.600 ;
        RECT 244.950 715.950 247.050 716.400 ;
        RECT 280.950 715.950 283.050 716.400 ;
        RECT 298.950 717.600 301.050 718.050 ;
        RECT 316.950 717.600 319.050 718.050 ;
        RECT 298.950 716.400 319.050 717.600 ;
        RECT 298.950 715.950 301.050 716.400 ;
        RECT 316.950 715.950 319.050 716.400 ;
        RECT 481.950 717.600 484.050 718.050 ;
        RECT 511.950 717.600 514.050 718.050 ;
        RECT 481.950 716.400 514.050 717.600 ;
        RECT 481.950 715.950 484.050 716.400 ;
        RECT 511.950 715.950 514.050 716.400 ;
        RECT 517.950 717.600 520.050 718.050 ;
        RECT 541.950 717.600 544.050 718.050 ;
        RECT 517.950 716.400 544.050 717.600 ;
        RECT 517.950 715.950 520.050 716.400 ;
        RECT 541.950 715.950 544.050 716.400 ;
        RECT 547.950 717.600 550.050 718.050 ;
        RECT 577.950 717.600 580.050 718.050 ;
        RECT 547.950 716.400 580.050 717.600 ;
        RECT 547.950 715.950 550.050 716.400 ;
        RECT 577.950 715.950 580.050 716.400 ;
        RECT 610.950 717.600 613.050 718.050 ;
        RECT 649.950 717.600 652.050 718.050 ;
        RECT 610.950 716.400 652.050 717.600 ;
        RECT 610.950 715.950 613.050 716.400 ;
        RECT 649.950 715.950 652.050 716.400 ;
        RECT 667.950 717.600 670.050 718.050 ;
        RECT 685.950 717.600 688.050 718.050 ;
        RECT 667.950 716.400 688.050 717.600 ;
        RECT 667.950 715.950 670.050 716.400 ;
        RECT 685.950 715.950 688.050 716.400 ;
        RECT 700.950 717.600 703.050 718.050 ;
        RECT 730.950 717.600 733.050 718.050 ;
        RECT 700.950 716.400 733.050 717.600 ;
        RECT 700.950 715.950 703.050 716.400 ;
        RECT 730.950 715.950 733.050 716.400 ;
        RECT 769.950 717.600 772.050 718.050 ;
        RECT 802.950 717.600 805.050 718.050 ;
        RECT 769.950 716.400 805.050 717.600 ;
        RECT 769.950 715.950 772.050 716.400 ;
        RECT 802.950 715.950 805.050 716.400 ;
        RECT 844.950 717.600 847.050 718.050 ;
        RECT 868.950 717.600 871.050 718.050 ;
        RECT 844.950 716.400 871.050 717.600 ;
        RECT 844.950 715.950 847.050 716.400 ;
        RECT 868.950 715.950 871.050 716.400 ;
        RECT 163.950 714.600 166.050 715.050 ;
        RECT 232.950 714.600 235.050 715.050 ;
        RECT 238.950 714.600 241.050 715.050 ;
        RECT 163.950 713.400 241.050 714.600 ;
        RECT 163.950 712.950 166.050 713.400 ;
        RECT 232.950 712.950 235.050 713.400 ;
        RECT 238.950 712.950 241.050 713.400 ;
        RECT 319.950 714.600 322.050 715.050 ;
        RECT 379.950 714.600 382.050 715.050 ;
        RECT 319.950 713.400 382.050 714.600 ;
        RECT 319.950 712.950 322.050 713.400 ;
        RECT 379.950 712.950 382.050 713.400 ;
        RECT 493.950 714.600 496.050 715.050 ;
        RECT 502.950 714.600 505.050 715.050 ;
        RECT 493.950 713.400 505.050 714.600 ;
        RECT 493.950 712.950 496.050 713.400 ;
        RECT 502.950 712.950 505.050 713.400 ;
        RECT 592.950 714.600 595.050 715.050 ;
        RECT 655.950 714.600 658.050 715.050 ;
        RECT 661.950 714.600 664.050 715.050 ;
        RECT 678.000 714.600 682.050 715.050 ;
        RECT 592.950 713.400 664.050 714.600 ;
        RECT 592.950 712.950 595.050 713.400 ;
        RECT 655.950 712.950 658.050 713.400 ;
        RECT 661.950 712.950 664.050 713.400 ;
        RECT 677.400 712.950 682.050 714.600 ;
        RECT 697.950 714.600 700.050 715.050 ;
        RECT 733.950 714.600 736.050 715.050 ;
        RECT 907.950 714.600 910.050 715.050 ;
        RECT 697.950 713.400 726.600 714.600 ;
        RECT 697.950 712.950 700.050 713.400 ;
        RECT 13.950 711.600 16.050 712.050 ;
        RECT 28.950 711.600 31.050 712.050 ;
        RECT 31.950 711.600 34.050 712.050 ;
        RECT 79.950 711.600 82.050 712.050 ;
        RECT 109.950 711.600 112.050 712.050 ;
        RECT 13.950 710.400 112.050 711.600 ;
        RECT 13.950 709.950 16.050 710.400 ;
        RECT 28.950 709.950 31.050 710.400 ;
        RECT 31.950 709.950 34.050 710.400 ;
        RECT 79.950 709.950 82.050 710.400 ;
        RECT 109.950 709.950 112.050 710.400 ;
        RECT 202.950 711.600 205.050 712.050 ;
        RECT 298.950 711.600 301.050 712.050 ;
        RECT 337.950 711.600 340.050 712.050 ;
        RECT 358.950 711.600 361.050 712.050 ;
        RECT 202.950 710.400 340.050 711.600 ;
        RECT 202.950 709.950 205.050 710.400 ;
        RECT 298.950 709.950 301.050 710.400 ;
        RECT 337.950 709.950 340.050 710.400 ;
        RECT 341.400 710.400 361.050 711.600 ;
        RECT 49.950 708.600 52.050 709.050 ;
        RECT 85.950 708.600 88.050 709.050 ;
        RECT 49.950 707.400 88.050 708.600 ;
        RECT 49.950 706.950 52.050 707.400 ;
        RECT 85.950 706.950 88.050 707.400 ;
        RECT 112.950 708.600 115.050 709.050 ;
        RECT 157.950 708.600 160.050 709.050 ;
        RECT 202.950 708.600 205.050 708.900 ;
        RECT 112.950 707.400 160.050 708.600 ;
        RECT 112.950 706.950 115.050 707.400 ;
        RECT 157.950 706.950 160.050 707.400 ;
        RECT 188.400 707.400 205.050 708.600 ;
        RECT 115.950 705.600 118.050 706.050 ;
        RECT 178.950 705.600 181.050 706.050 ;
        RECT 188.400 705.600 189.600 707.400 ;
        RECT 202.950 706.800 205.050 707.400 ;
        RECT 208.950 708.600 211.050 709.050 ;
        RECT 268.950 708.600 271.050 709.050 ;
        RECT 208.950 707.400 271.050 708.600 ;
        RECT 208.950 706.950 211.050 707.400 ;
        RECT 268.950 706.950 271.050 707.400 ;
        RECT 316.950 708.600 319.050 709.050 ;
        RECT 341.400 708.600 342.600 710.400 ;
        RECT 358.950 709.950 361.050 710.400 ;
        RECT 433.950 711.600 436.050 712.050 ;
        RECT 535.950 711.600 538.050 712.050 ;
        RECT 634.950 711.600 637.050 712.050 ;
        RECT 433.950 710.400 538.050 711.600 ;
        RECT 433.950 709.950 436.050 710.400 ;
        RECT 535.950 709.950 538.050 710.400 ;
        RECT 587.400 710.400 637.050 711.600 ;
        RECT 316.950 707.400 342.600 708.600 ;
        RECT 364.950 708.600 367.050 709.050 ;
        RECT 451.950 708.600 454.050 709.050 ;
        RECT 499.950 708.600 502.050 709.050 ;
        RECT 364.950 707.400 502.050 708.600 ;
        RECT 316.950 706.950 319.050 707.400 ;
        RECT 364.950 706.950 367.050 707.400 ;
        RECT 451.950 706.950 454.050 707.400 ;
        RECT 499.950 706.950 502.050 707.400 ;
        RECT 565.950 708.600 568.050 709.050 ;
        RECT 587.400 708.600 588.600 710.400 ;
        RECT 634.950 709.950 637.050 710.400 ;
        RECT 640.950 711.600 643.050 712.050 ;
        RECT 677.400 711.600 678.600 712.950 ;
        RECT 640.950 710.400 678.600 711.600 ;
        RECT 725.400 711.600 726.600 713.400 ;
        RECT 733.950 713.400 910.050 714.600 ;
        RECT 733.950 712.950 736.050 713.400 ;
        RECT 907.950 712.950 910.050 713.400 ;
        RECT 775.950 711.600 778.050 712.050 ;
        RECT 725.400 710.400 778.050 711.600 ;
        RECT 640.950 709.950 643.050 710.400 ;
        RECT 775.950 709.950 778.050 710.400 ;
        RECT 781.950 711.600 784.050 712.050 ;
        RECT 787.950 711.600 790.050 712.050 ;
        RECT 805.950 711.600 808.050 712.050 ;
        RECT 781.950 710.400 808.050 711.600 ;
        RECT 781.950 709.950 784.050 710.400 ;
        RECT 787.950 709.950 790.050 710.400 ;
        RECT 805.950 709.950 808.050 710.400 ;
        RECT 565.950 707.400 588.600 708.600 ;
        RECT 589.950 708.600 592.050 709.050 ;
        RECT 607.950 708.600 610.050 709.050 ;
        RECT 589.950 707.400 610.050 708.600 ;
        RECT 565.950 706.950 568.050 707.400 ;
        RECT 589.950 706.950 592.050 707.400 ;
        RECT 607.950 706.950 610.050 707.400 ;
        RECT 628.950 708.600 631.050 709.050 ;
        RECT 673.800 708.600 675.900 709.050 ;
        RECT 628.950 707.400 675.900 708.600 ;
        RECT 628.950 706.950 631.050 707.400 ;
        RECT 673.800 706.950 675.900 707.400 ;
        RECT 703.950 708.600 706.050 709.050 ;
        RECT 751.950 708.600 754.050 709.050 ;
        RECT 703.950 707.400 754.050 708.600 ;
        RECT 703.950 706.950 706.050 707.400 ;
        RECT 751.950 706.950 754.050 707.400 ;
        RECT 115.950 704.400 189.600 705.600 ;
        RECT 193.950 705.600 196.050 706.050 ;
        RECT 271.950 705.600 274.050 706.050 ;
        RECT 313.950 705.600 316.050 706.050 ;
        RECT 352.950 705.600 355.050 706.050 ;
        RECT 193.950 704.400 316.050 705.600 ;
        RECT 115.950 703.950 118.050 704.400 ;
        RECT 178.950 703.950 181.050 704.400 ;
        RECT 193.950 703.950 196.050 704.400 ;
        RECT 271.950 703.950 274.050 704.400 ;
        RECT 313.950 703.950 316.050 704.400 ;
        RECT 326.400 704.400 355.050 705.600 ;
        RECT 70.950 702.600 73.050 703.050 ;
        RECT 91.950 702.600 94.050 703.050 ;
        RECT 70.950 701.400 94.050 702.600 ;
        RECT 70.950 700.950 73.050 701.400 ;
        RECT 91.950 700.950 94.050 701.400 ;
        RECT 223.950 702.600 226.050 703.050 ;
        RECT 241.950 702.600 244.050 703.050 ;
        RECT 250.950 702.600 253.050 703.050 ;
        RECT 223.950 701.400 253.050 702.600 ;
        RECT 223.950 700.950 226.050 701.400 ;
        RECT 241.950 700.950 244.050 701.400 ;
        RECT 250.950 700.950 253.050 701.400 ;
        RECT 289.950 702.600 292.050 703.050 ;
        RECT 326.400 702.600 327.600 704.400 ;
        RECT 352.950 703.950 355.050 704.400 ;
        RECT 361.950 705.600 364.050 706.050 ;
        RECT 436.950 705.600 439.050 706.050 ;
        RECT 361.950 704.400 439.050 705.600 ;
        RECT 361.950 703.950 364.050 704.400 ;
        RECT 436.950 703.950 439.050 704.400 ;
        RECT 454.950 705.600 457.050 706.050 ;
        RECT 490.950 705.600 493.050 706.050 ;
        RECT 454.950 704.400 493.050 705.600 ;
        RECT 454.950 703.950 457.050 704.400 ;
        RECT 490.950 703.950 493.050 704.400 ;
        RECT 541.950 705.600 544.050 706.050 ;
        RECT 553.950 705.600 556.050 706.050 ;
        RECT 541.950 704.400 556.050 705.600 ;
        RECT 541.950 703.950 544.050 704.400 ;
        RECT 553.950 703.950 556.050 704.400 ;
        RECT 598.950 705.600 601.050 706.050 ;
        RECT 631.950 705.600 634.050 706.050 ;
        RECT 598.950 704.400 634.050 705.600 ;
        RECT 598.950 703.950 601.050 704.400 ;
        RECT 631.950 703.950 634.050 704.400 ;
        RECT 652.950 705.600 655.050 706.050 ;
        RECT 706.800 705.600 708.900 706.050 ;
        RECT 652.950 704.400 708.900 705.600 ;
        RECT 652.950 703.950 655.050 704.400 ;
        RECT 706.800 703.950 708.900 704.400 ;
        RECT 709.950 705.600 712.050 706.050 ;
        RECT 781.950 705.600 784.050 706.050 ;
        RECT 709.950 704.400 784.050 705.600 ;
        RECT 709.950 703.950 712.050 704.400 ;
        RECT 781.950 703.950 784.050 704.400 ;
        RECT 787.950 705.600 790.050 706.050 ;
        RECT 820.950 705.600 823.050 706.050 ;
        RECT 832.950 705.600 835.050 706.050 ;
        RECT 787.950 704.400 835.050 705.600 ;
        RECT 787.950 703.950 790.050 704.400 ;
        RECT 820.950 703.950 823.050 704.400 ;
        RECT 832.950 703.950 835.050 704.400 ;
        RECT 289.950 701.400 327.600 702.600 ;
        RECT 328.950 702.600 331.050 703.050 ;
        RECT 532.950 702.600 535.050 703.050 ;
        RECT 547.950 702.600 550.050 703.050 ;
        RECT 553.950 702.600 556.050 702.900 ;
        RECT 328.950 701.400 441.600 702.600 ;
        RECT 289.950 700.950 292.050 701.400 ;
        RECT 328.950 700.950 331.050 701.400 ;
        RECT 1.950 699.600 4.050 700.050 ;
        RECT 115.950 699.600 118.050 700.050 ;
        RECT 1.950 698.400 118.050 699.600 ;
        RECT 1.950 697.950 4.050 698.400 ;
        RECT 115.950 697.950 118.050 698.400 ;
        RECT 181.950 699.600 184.050 700.050 ;
        RECT 193.950 699.600 196.050 700.050 ;
        RECT 181.950 698.400 196.050 699.600 ;
        RECT 181.950 697.950 184.050 698.400 ;
        RECT 193.950 697.950 196.050 698.400 ;
        RECT 259.950 699.600 262.050 700.050 ;
        RECT 349.950 699.600 352.050 700.050 ;
        RECT 259.950 698.400 352.050 699.600 ;
        RECT 259.950 697.950 262.050 698.400 ;
        RECT 349.950 697.950 352.050 698.400 ;
        RECT 358.950 699.600 361.050 700.050 ;
        RECT 403.950 699.600 406.050 700.050 ;
        RECT 358.950 698.400 406.050 699.600 ;
        RECT 440.400 699.600 441.600 701.400 ;
        RECT 532.950 701.400 556.050 702.600 ;
        RECT 532.950 700.950 535.050 701.400 ;
        RECT 547.950 700.950 550.050 701.400 ;
        RECT 553.950 700.800 556.050 701.400 ;
        RECT 586.950 702.600 589.050 703.050 ;
        RECT 649.950 702.600 652.050 703.050 ;
        RECT 586.950 701.400 652.050 702.600 ;
        RECT 586.950 700.950 589.050 701.400 ;
        RECT 649.950 700.950 652.050 701.400 ;
        RECT 691.950 702.600 694.050 703.050 ;
        RECT 721.950 702.600 724.050 703.050 ;
        RECT 691.950 701.400 724.050 702.600 ;
        RECT 691.950 700.950 694.050 701.400 ;
        RECT 721.950 700.950 724.050 701.400 ;
        RECT 730.950 702.600 733.050 703.050 ;
        RECT 847.950 702.600 850.050 703.050 ;
        RECT 730.950 701.400 850.050 702.600 ;
        RECT 730.950 700.950 733.050 701.400 ;
        RECT 847.950 700.950 850.050 701.400 ;
        RECT 460.950 699.600 463.050 700.050 ;
        RECT 440.400 698.400 463.050 699.600 ;
        RECT 358.950 697.950 361.050 698.400 ;
        RECT 403.950 697.950 406.050 698.400 ;
        RECT 460.950 697.950 463.050 698.400 ;
        RECT 490.950 699.600 493.050 700.050 ;
        RECT 598.950 699.600 601.050 700.050 ;
        RECT 490.950 698.400 601.050 699.600 ;
        RECT 490.950 697.950 493.050 698.400 ;
        RECT 598.950 697.950 601.050 698.400 ;
        RECT 673.950 699.600 676.050 700.050 ;
        RECT 691.950 699.600 694.050 699.900 ;
        RECT 673.950 698.400 694.050 699.600 ;
        RECT 673.950 697.950 676.050 698.400 ;
        RECT 691.950 697.800 694.050 698.400 ;
        RECT 802.950 699.600 805.050 700.050 ;
        RECT 844.950 699.600 847.050 700.050 ;
        RECT 802.950 698.400 847.050 699.600 ;
        RECT 802.950 697.950 805.050 698.400 ;
        RECT 844.950 697.950 847.050 698.400 ;
        RECT 883.950 699.600 886.050 700.050 ;
        RECT 913.950 699.600 916.050 700.050 ;
        RECT 883.950 698.400 916.050 699.600 ;
        RECT 883.950 697.950 886.050 698.400 ;
        RECT 913.950 697.950 916.050 698.400 ;
        RECT 130.950 696.600 133.050 697.050 ;
        RECT 172.950 696.600 175.050 697.050 ;
        RECT 130.950 695.400 175.050 696.600 ;
        RECT 130.950 694.950 133.050 695.400 ;
        RECT 172.950 694.950 175.050 695.400 ;
        RECT 208.950 696.600 211.050 697.050 ;
        RECT 238.950 696.600 241.050 697.050 ;
        RECT 409.950 696.600 412.050 697.050 ;
        RECT 208.950 695.400 412.050 696.600 ;
        RECT 208.950 694.950 211.050 695.400 ;
        RECT 238.950 694.950 241.050 695.400 ;
        RECT 409.950 694.950 412.050 695.400 ;
        RECT 430.950 696.600 433.050 697.050 ;
        RECT 439.950 696.600 442.050 697.050 ;
        RECT 430.950 695.400 442.050 696.600 ;
        RECT 430.950 694.950 433.050 695.400 ;
        RECT 439.950 694.950 442.050 695.400 ;
        RECT 487.950 696.600 490.050 697.050 ;
        RECT 532.800 696.600 534.900 697.050 ;
        RECT 487.950 695.400 534.900 696.600 ;
        RECT 487.950 694.950 490.050 695.400 ;
        RECT 532.800 694.950 534.900 695.400 ;
        RECT 535.950 696.600 538.050 697.050 ;
        RECT 649.950 696.600 652.050 697.050 ;
        RECT 697.950 696.600 700.050 697.050 ;
        RECT 535.950 695.400 627.600 696.600 ;
        RECT 535.950 694.950 538.050 695.400 ;
        RECT 73.950 693.600 76.050 694.050 ;
        RECT 145.950 693.600 148.050 694.050 ;
        RECT 73.950 692.400 148.050 693.600 ;
        RECT 73.950 691.950 76.050 692.400 ;
        RECT 145.950 691.950 148.050 692.400 ;
        RECT 256.950 693.600 259.050 694.050 ;
        RECT 283.800 693.600 285.900 694.050 ;
        RECT 256.950 692.400 285.900 693.600 ;
        RECT 256.950 691.950 259.050 692.400 ;
        RECT 283.800 691.950 285.900 692.400 ;
        RECT 286.950 693.600 289.050 694.050 ;
        RECT 343.950 693.600 346.050 694.050 ;
        RECT 364.950 693.600 367.050 694.050 ;
        RECT 286.950 692.400 327.600 693.600 ;
        RECT 286.950 691.950 289.050 692.400 ;
        RECT 10.950 690.600 13.050 691.050 ;
        RECT 34.950 690.600 37.050 691.050 ;
        RECT 10.950 689.400 37.050 690.600 ;
        RECT 10.950 688.950 13.050 689.400 ;
        RECT 34.950 688.950 37.050 689.400 ;
        RECT 154.950 690.600 157.050 691.050 ;
        RECT 160.950 690.600 163.050 691.050 ;
        RECT 154.950 689.400 163.050 690.600 ;
        RECT 326.400 690.600 327.600 692.400 ;
        RECT 343.950 692.400 367.050 693.600 ;
        RECT 343.950 691.950 346.050 692.400 ;
        RECT 364.950 691.950 367.050 692.400 ;
        RECT 571.950 693.600 574.050 694.050 ;
        RECT 622.950 693.600 625.050 694.050 ;
        RECT 571.950 692.400 625.050 693.600 ;
        RECT 626.400 693.600 627.600 695.400 ;
        RECT 649.950 695.400 700.050 696.600 ;
        RECT 649.950 694.950 652.050 695.400 ;
        RECT 697.950 694.950 700.050 695.400 ;
        RECT 760.950 696.600 763.050 697.050 ;
        RECT 772.950 696.600 775.050 697.050 ;
        RECT 760.950 695.400 775.050 696.600 ;
        RECT 760.950 694.950 763.050 695.400 ;
        RECT 772.950 694.950 775.050 695.400 ;
        RECT 781.950 696.600 784.050 697.050 ;
        RECT 829.950 696.600 832.050 697.050 ;
        RECT 781.950 695.400 832.050 696.600 ;
        RECT 781.950 694.950 784.050 695.400 ;
        RECT 829.950 694.950 832.050 695.400 ;
        RECT 856.950 696.600 859.050 697.050 ;
        RECT 874.950 696.600 877.050 697.050 ;
        RECT 856.950 695.400 877.050 696.600 ;
        RECT 856.950 694.950 859.050 695.400 ;
        RECT 874.950 694.950 877.050 695.400 ;
        RECT 640.950 693.600 643.050 694.050 ;
        RECT 626.400 692.400 643.050 693.600 ;
        RECT 571.950 691.950 574.050 692.400 ;
        RECT 622.950 691.950 625.050 692.400 ;
        RECT 640.950 691.950 643.050 692.400 ;
        RECT 679.950 693.600 682.050 694.050 ;
        RECT 694.950 693.600 697.050 694.050 ;
        RECT 679.950 692.400 697.050 693.600 ;
        RECT 679.950 691.950 682.050 692.400 ;
        RECT 694.950 691.950 697.050 692.400 ;
        RECT 826.950 693.600 829.050 694.050 ;
        RECT 835.950 693.600 838.050 694.050 ;
        RECT 826.950 692.400 838.050 693.600 ;
        RECT 826.950 691.950 829.050 692.400 ;
        RECT 835.950 691.950 838.050 692.400 ;
        RECT 847.950 693.600 850.050 694.050 ;
        RECT 886.950 693.600 889.050 694.050 ;
        RECT 847.950 692.400 889.050 693.600 ;
        RECT 847.950 691.950 850.050 692.400 ;
        RECT 886.950 691.950 889.050 692.400 ;
        RECT 355.950 690.600 358.050 691.050 ;
        RECT 326.400 689.400 358.050 690.600 ;
        RECT 154.950 688.950 157.050 689.400 ;
        RECT 160.950 688.950 163.050 689.400 ;
        RECT 355.950 688.950 358.050 689.400 ;
        RECT 379.950 690.600 382.050 691.050 ;
        RECT 391.950 690.600 394.050 691.050 ;
        RECT 379.950 689.400 394.050 690.600 ;
        RECT 379.950 688.950 382.050 689.400 ;
        RECT 391.950 688.950 394.050 689.400 ;
        RECT 397.950 690.600 400.050 691.050 ;
        RECT 439.950 690.600 442.050 691.050 ;
        RECT 397.950 689.400 442.050 690.600 ;
        RECT 397.950 688.950 400.050 689.400 ;
        RECT 439.950 688.950 442.050 689.400 ;
        RECT 463.950 690.600 466.050 691.050 ;
        RECT 523.950 690.600 526.050 691.050 ;
        RECT 463.950 689.400 526.050 690.600 ;
        RECT 463.950 688.950 466.050 689.400 ;
        RECT 523.950 688.950 526.050 689.400 ;
        RECT 580.950 690.600 583.050 691.050 ;
        RECT 667.800 690.600 669.900 691.050 ;
        RECT 580.950 689.400 669.900 690.600 ;
        RECT 580.950 688.950 583.050 689.400 ;
        RECT 667.800 688.950 669.900 689.400 ;
        RECT 670.950 690.600 673.050 691.050 ;
        RECT 685.950 690.600 688.050 691.050 ;
        RECT 670.950 689.400 688.050 690.600 ;
        RECT 670.950 688.950 673.050 689.400 ;
        RECT 685.950 688.950 688.050 689.400 ;
        RECT 709.950 690.600 712.050 690.900 ;
        RECT 721.950 690.600 724.050 691.050 ;
        RECT 709.950 689.400 724.050 690.600 ;
        RECT 709.950 688.800 712.050 689.400 ;
        RECT 721.950 688.950 724.050 689.400 ;
        RECT 745.950 690.600 748.050 691.050 ;
        RECT 802.950 690.600 805.050 691.050 ;
        RECT 745.950 689.400 805.050 690.600 ;
        RECT 745.950 688.950 748.050 689.400 ;
        RECT 802.950 688.950 805.050 689.400 ;
        RECT 811.950 690.600 814.050 691.050 ;
        RECT 832.950 690.600 835.050 691.050 ;
        RECT 811.950 689.400 835.050 690.600 ;
        RECT 811.950 688.950 814.050 689.400 ;
        RECT 832.950 688.950 835.050 689.400 ;
        RECT 109.950 687.600 112.050 688.050 ;
        RECT 169.950 687.600 172.050 688.050 ;
        RECT 181.950 687.600 184.050 688.050 ;
        RECT 109.950 686.400 162.600 687.600 ;
        RECT 109.950 685.950 112.050 686.400 ;
        RECT 4.950 684.750 7.050 685.200 ;
        RECT 10.950 684.750 13.050 685.200 ;
        RECT 4.950 683.550 13.050 684.750 ;
        RECT 4.950 683.100 7.050 683.550 ;
        RECT 10.950 683.100 13.050 683.550 ;
        RECT 16.950 684.750 19.050 685.200 ;
        RECT 22.800 684.750 24.900 685.200 ;
        RECT 16.950 683.550 24.900 684.750 ;
        RECT 16.950 683.100 19.050 683.550 ;
        RECT 22.800 683.100 24.900 683.550 ;
        RECT 25.950 682.950 28.050 685.050 ;
        RECT 43.950 684.600 46.050 685.050 ;
        RECT 58.950 684.600 61.050 685.050 ;
        RECT 43.950 683.400 61.050 684.600 ;
        RECT 43.950 682.950 46.050 683.400 ;
        RECT 58.950 682.950 61.050 683.400 ;
        RECT 64.950 684.600 67.050 685.200 ;
        RECT 76.950 684.600 79.050 685.200 ;
        RECT 64.950 683.400 79.050 684.600 ;
        RECT 64.950 683.100 67.050 683.400 ;
        RECT 76.950 683.100 79.050 683.400 ;
        RECT 82.950 684.600 85.050 685.200 ;
        RECT 100.950 684.600 103.050 685.200 ;
        RECT 82.950 683.400 103.050 684.600 ;
        RECT 82.950 683.100 85.050 683.400 ;
        RECT 100.950 683.100 103.050 683.400 ;
        RECT 106.950 683.100 109.050 685.200 ;
        RECT 115.950 684.600 118.050 685.050 ;
        RECT 121.950 684.600 124.050 685.050 ;
        RECT 115.950 683.400 124.050 684.600 ;
        RECT 26.400 678.600 27.600 682.950 ;
        RECT 77.400 681.600 78.600 683.100 ;
        RECT 107.400 681.600 108.600 683.100 ;
        RECT 115.950 682.950 118.050 683.400 ;
        RECT 121.950 682.950 124.050 683.400 ;
        RECT 154.950 684.600 159.000 685.050 ;
        RECT 161.400 684.600 162.600 686.400 ;
        RECT 169.950 686.400 184.050 687.600 ;
        RECT 169.950 685.950 172.050 686.400 ;
        RECT 181.950 685.950 184.050 686.400 ;
        RECT 322.950 687.600 325.050 688.050 ;
        RECT 331.950 687.600 334.050 688.050 ;
        RECT 322.950 686.400 334.050 687.600 ;
        RECT 322.950 685.950 325.050 686.400 ;
        RECT 331.950 685.950 334.050 686.400 ;
        RECT 442.950 687.600 445.050 688.050 ;
        RECT 451.950 687.600 454.050 688.050 ;
        RECT 442.950 686.400 454.050 687.600 ;
        RECT 442.950 685.950 445.050 686.400 ;
        RECT 451.950 685.950 454.050 686.400 ;
        RECT 694.950 687.600 697.050 688.050 ;
        RECT 706.950 687.600 709.050 688.050 ;
        RECT 694.950 686.400 709.050 687.600 ;
        RECT 694.950 685.950 697.050 686.400 ;
        RECT 706.950 685.950 709.050 686.400 ;
        RECT 733.950 687.600 736.050 688.050 ;
        RECT 742.950 687.600 745.050 688.050 ;
        RECT 733.950 686.400 745.050 687.600 ;
        RECT 733.950 685.950 736.050 686.400 ;
        RECT 742.950 685.950 745.050 686.400 ;
        RECT 766.950 687.600 769.050 688.050 ;
        RECT 796.950 687.600 799.050 688.050 ;
        RECT 766.950 686.400 799.050 687.600 ;
        RECT 766.950 685.950 769.050 686.400 ;
        RECT 796.950 685.950 799.050 686.400 ;
        RECT 814.950 685.950 817.050 688.050 ;
        RECT 856.950 685.950 859.050 688.050 ;
        RECT 919.950 687.600 924.000 688.050 ;
        RECT 919.950 685.950 924.600 687.600 ;
        RECT 187.950 684.750 190.050 685.200 ;
        RECT 196.950 684.750 199.050 685.200 ;
        RECT 154.950 682.950 159.600 684.600 ;
        RECT 161.400 683.400 183.600 684.600 ;
        RECT 77.400 680.400 108.600 681.600 ;
        RECT 158.400 681.600 159.600 682.950 ;
        RECT 158.400 680.400 180.600 681.600 ;
        RECT 31.950 678.600 34.050 678.900 ;
        RECT 26.400 677.400 34.050 678.600 ;
        RECT 31.950 676.800 34.050 677.400 ;
        RECT 46.950 678.600 49.050 679.050 ;
        RECT 55.950 678.600 58.050 678.900 ;
        RECT 46.950 677.400 58.050 678.600 ;
        RECT 46.950 676.950 49.050 677.400 ;
        RECT 55.950 676.800 58.050 677.400 ;
        RECT 79.950 678.600 82.050 678.900 ;
        RECT 103.950 678.600 106.050 678.900 ;
        RECT 79.950 677.400 106.050 678.600 ;
        RECT 79.950 676.800 82.050 677.400 ;
        RECT 103.950 676.800 106.050 677.400 ;
        RECT 88.950 675.600 91.050 676.050 ;
        RECT 94.950 675.600 97.050 676.050 ;
        RECT 88.950 674.400 97.050 675.600 ;
        RECT 107.400 675.600 108.600 680.400 ;
        RECT 118.950 678.600 121.050 679.050 ;
        RECT 154.950 678.600 157.050 679.050 ;
        RECT 179.400 678.900 180.600 680.400 ;
        RECT 118.950 677.400 157.050 678.600 ;
        RECT 118.950 676.950 121.050 677.400 ;
        RECT 154.950 676.950 157.050 677.400 ;
        RECT 163.950 678.450 166.050 678.900 ;
        RECT 175.800 678.450 177.900 678.900 ;
        RECT 163.950 677.250 177.900 678.450 ;
        RECT 163.950 676.800 166.050 677.250 ;
        RECT 175.800 676.800 177.900 677.250 ;
        RECT 178.950 676.800 181.050 678.900 ;
        RECT 182.400 678.600 183.600 683.400 ;
        RECT 187.950 683.550 199.050 684.750 ;
        RECT 187.950 683.100 190.050 683.550 ;
        RECT 196.950 683.100 199.050 683.550 ;
        RECT 226.950 683.100 229.050 685.200 ;
        RECT 232.950 684.600 235.050 685.200 ;
        RECT 250.950 684.600 253.050 685.200 ;
        RECT 256.950 684.600 259.050 685.200 ;
        RECT 232.950 683.400 253.050 684.600 ;
        RECT 232.950 683.100 235.050 683.400 ;
        RECT 250.950 683.100 253.050 683.400 ;
        RECT 254.400 683.400 259.050 684.600 ;
        RECT 227.400 681.600 228.600 683.100 ;
        RECT 254.400 681.600 255.600 683.400 ;
        RECT 256.950 683.100 259.050 683.400 ;
        RECT 274.950 683.100 277.050 685.200 ;
        RECT 280.950 684.600 283.050 685.050 ;
        RECT 292.950 684.750 295.050 685.200 ;
        RECT 307.950 684.750 310.050 685.200 ;
        RECT 292.950 684.600 310.050 684.750 ;
        RECT 280.950 683.550 310.050 684.600 ;
        RECT 280.950 683.400 295.050 683.550 ;
        RECT 221.400 681.000 228.600 681.600 ;
        RECT 220.950 680.400 228.600 681.000 ;
        RECT 230.400 680.400 255.600 681.600 ;
        RECT 184.950 678.600 187.050 678.900 ;
        RECT 182.400 677.400 187.050 678.600 ;
        RECT 184.950 676.800 187.050 677.400 ;
        RECT 196.950 678.600 199.050 679.050 ;
        RECT 205.950 678.600 208.050 678.900 ;
        RECT 196.950 677.400 208.050 678.600 ;
        RECT 196.950 676.950 199.050 677.400 ;
        RECT 205.950 676.800 208.050 677.400 ;
        RECT 220.950 676.950 223.050 680.400 ;
        RECT 230.400 678.900 231.600 680.400 ;
        RECT 229.950 676.800 232.050 678.900 ;
        RECT 265.950 678.600 268.050 679.050 ;
        RECT 271.950 678.600 274.050 678.900 ;
        RECT 265.950 677.400 274.050 678.600 ;
        RECT 265.950 676.950 268.050 677.400 ;
        RECT 271.950 676.800 274.050 677.400 ;
        RECT 133.950 675.600 136.050 676.050 ;
        RECT 107.400 674.400 136.050 675.600 ;
        RECT 88.950 673.950 91.050 674.400 ;
        RECT 94.950 673.950 97.050 674.400 ;
        RECT 133.950 673.950 136.050 674.400 ;
        RECT 259.950 675.600 262.050 676.050 ;
        RECT 275.400 675.600 276.600 683.100 ;
        RECT 280.950 682.950 283.050 683.400 ;
        RECT 292.950 683.100 295.050 683.400 ;
        RECT 307.950 683.100 310.050 683.550 ;
        RECT 319.950 683.100 322.050 685.200 ;
        RECT 352.950 684.750 355.050 685.200 ;
        RECT 421.950 684.750 424.050 685.200 ;
        RECT 352.950 684.600 424.050 684.750 ;
        RECT 433.950 684.600 436.050 685.050 ;
        RECT 463.950 684.600 466.050 685.050 ;
        RECT 352.950 683.550 436.050 684.600 ;
        RECT 352.950 683.100 355.050 683.550 ;
        RECT 421.950 683.400 436.050 683.550 ;
        RECT 421.950 683.100 424.050 683.400 ;
        RECT 283.950 678.600 286.050 679.050 ;
        RECT 316.950 678.600 319.050 678.900 ;
        RECT 283.950 677.400 319.050 678.600 ;
        RECT 320.400 678.600 321.600 683.100 ;
        RECT 433.950 682.950 436.050 683.400 ;
        RECT 458.400 683.400 466.050 684.600 ;
        RECT 367.950 681.600 370.050 682.050 ;
        RECT 458.400 681.600 459.600 683.400 ;
        RECT 463.950 682.950 466.050 683.400 ;
        RECT 472.950 684.600 475.050 685.050 ;
        RECT 484.950 684.600 487.050 685.050 ;
        RECT 472.950 683.400 487.050 684.600 ;
        RECT 472.950 682.950 475.050 683.400 ;
        RECT 484.950 682.950 487.050 683.400 ;
        RECT 496.950 684.600 499.050 685.050 ;
        RECT 541.950 684.600 544.050 685.050 ;
        RECT 496.950 683.400 544.050 684.600 ;
        RECT 496.950 682.950 499.050 683.400 ;
        RECT 541.950 682.950 544.050 683.400 ;
        RECT 559.950 684.750 562.050 685.200 ;
        RECT 571.950 684.750 574.050 685.200 ;
        RECT 559.950 683.550 574.050 684.750 ;
        RECT 559.950 683.100 562.050 683.550 ;
        RECT 571.950 683.100 574.050 683.550 ;
        RECT 601.950 684.600 604.050 685.200 ;
        RECT 616.950 684.600 619.050 685.200 ;
        RECT 624.000 684.600 628.050 685.050 ;
        RECT 601.950 683.400 619.050 684.600 ;
        RECT 601.950 683.100 604.050 683.400 ;
        RECT 616.950 683.100 619.050 683.400 ;
        RECT 623.400 682.950 628.050 684.600 ;
        RECT 637.950 684.750 640.050 685.200 ;
        RECT 643.950 684.750 646.050 685.200 ;
        RECT 637.950 683.550 646.050 684.750 ;
        RECT 637.950 683.100 640.050 683.550 ;
        RECT 643.950 683.100 646.050 683.550 ;
        RECT 667.950 684.600 670.050 685.200 ;
        RECT 685.950 684.600 688.050 685.050 ;
        RECT 757.950 684.750 760.050 684.900 ;
        RECT 766.950 684.750 769.050 685.200 ;
        RECT 667.950 683.400 684.600 684.600 ;
        RECT 667.950 683.100 670.050 683.400 ;
        RECT 367.950 680.400 405.600 681.600 ;
        RECT 367.950 679.950 370.050 680.400 ;
        RECT 325.950 678.600 328.050 679.050 ;
        RECT 320.400 677.400 328.050 678.600 ;
        RECT 404.400 678.600 405.600 680.400 ;
        RECT 449.400 680.400 459.600 681.600 ;
        RECT 424.950 678.600 427.050 678.900 ;
        RECT 436.950 678.600 439.050 678.900 ;
        RECT 404.400 677.400 439.050 678.600 ;
        RECT 283.950 676.950 286.050 677.400 ;
        RECT 316.950 676.800 319.050 677.400 ;
        RECT 325.950 676.950 328.050 677.400 ;
        RECT 424.950 676.800 427.050 677.400 ;
        RECT 436.950 676.800 439.050 677.400 ;
        RECT 442.950 678.600 445.050 678.900 ;
        RECT 449.400 678.600 450.600 680.400 ;
        RECT 442.950 677.400 450.600 678.600 ;
        RECT 451.950 678.450 454.050 678.900 ;
        RECT 460.950 678.450 463.050 678.900 ;
        RECT 442.950 676.800 445.050 677.400 ;
        RECT 451.950 677.250 463.050 678.450 ;
        RECT 451.950 676.800 454.050 677.250 ;
        RECT 460.950 676.800 463.050 677.250 ;
        RECT 565.950 678.600 568.050 679.050 ;
        RECT 574.950 678.600 577.050 679.050 ;
        RECT 565.950 677.400 577.050 678.600 ;
        RECT 565.950 676.950 568.050 677.400 ;
        RECT 574.950 676.950 577.050 677.400 ;
        RECT 623.400 676.050 624.600 682.950 ;
        RECT 683.400 681.600 684.600 683.400 ;
        RECT 685.950 683.400 753.600 684.600 ;
        RECT 685.950 682.950 688.050 683.400 ;
        RECT 752.400 682.050 753.600 683.400 ;
        RECT 757.950 683.550 769.050 684.750 ;
        RECT 757.950 682.800 760.050 683.550 ;
        RECT 766.950 683.100 769.050 683.550 ;
        RECT 772.950 683.100 775.050 685.200 ;
        RECT 790.950 683.100 793.050 685.200 ;
        RECT 804.000 684.600 808.050 685.050 ;
        RECT 683.400 681.000 687.600 681.600 ;
        RECT 683.400 680.400 688.050 681.000 ;
        RECT 752.400 680.400 757.050 682.050 ;
        RECT 685.950 676.950 688.050 680.400 ;
        RECT 753.000 679.950 757.050 680.400 ;
        RECT 773.400 679.050 774.600 683.100 ;
        RECT 791.400 679.050 792.600 683.100 ;
        RECT 803.400 682.950 808.050 684.600 ;
        RECT 803.400 679.050 804.600 682.950 ;
        RECT 703.950 678.450 706.050 678.900 ;
        RECT 742.950 678.450 745.050 678.900 ;
        RECT 703.950 677.250 745.050 678.450 ;
        RECT 773.400 677.400 778.050 679.050 ;
        RECT 703.950 676.800 706.050 677.250 ;
        RECT 742.950 676.800 745.050 677.250 ;
        RECT 774.000 676.950 778.050 677.400 ;
        RECT 787.950 677.400 792.600 679.050 ;
        RECT 787.950 676.950 792.000 677.400 ;
        RECT 802.950 676.950 805.050 679.050 ;
        RECT 815.400 678.600 816.600 685.950 ;
        RECT 817.950 684.600 820.050 685.200 ;
        RECT 823.950 684.600 826.050 685.050 ;
        RECT 817.950 683.400 826.050 684.600 ;
        RECT 817.950 683.100 820.050 683.400 ;
        RECT 823.950 682.950 826.050 683.400 ;
        RECT 841.950 684.600 844.050 685.200 ;
        RECT 841.950 683.400 846.600 684.600 ;
        RECT 841.950 683.100 844.050 683.400 ;
        RECT 845.400 679.050 846.600 683.400 ;
        RECT 820.950 678.600 823.050 679.050 ;
        RECT 815.400 677.400 823.050 678.600 ;
        RECT 820.950 676.950 823.050 677.400 ;
        RECT 844.950 676.950 847.050 679.050 ;
        RECT 857.400 676.050 858.600 685.950 ;
        RECT 883.950 681.600 886.050 685.050 ;
        RECT 889.950 684.600 892.050 685.200 ;
        RECT 910.950 684.750 913.050 685.200 ;
        RECT 919.950 684.750 922.050 684.900 ;
        RECT 889.950 683.400 909.600 684.600 ;
        RECT 889.950 683.100 892.050 683.400 ;
        RECT 883.950 681.000 888.600 681.600 ;
        RECT 884.400 680.400 888.600 681.000 ;
        RECT 887.400 678.900 888.600 680.400 ;
        RECT 908.400 678.900 909.600 683.400 ;
        RECT 910.950 683.550 922.050 684.750 ;
        RECT 910.950 683.100 913.050 683.550 ;
        RECT 919.950 682.800 922.050 683.550 ;
        RECT 923.400 681.600 924.600 685.950 ;
        RECT 917.400 681.000 924.600 681.600 ;
        RECT 916.950 680.400 924.600 681.000 ;
        RECT 886.950 676.800 889.050 678.900 ;
        RECT 907.950 676.800 910.050 678.900 ;
        RECT 916.950 676.950 919.050 680.400 ;
        RECT 259.950 674.400 276.600 675.600 ;
        RECT 283.950 675.600 286.050 675.900 ;
        RECT 328.950 675.600 331.050 676.050 ;
        RECT 283.950 674.400 331.050 675.600 ;
        RECT 259.950 673.950 262.050 674.400 ;
        RECT 283.950 673.800 286.050 674.400 ;
        RECT 328.950 673.950 331.050 674.400 ;
        RECT 352.950 675.600 355.050 676.050 ;
        RECT 421.950 675.600 424.050 676.050 ;
        RECT 352.950 674.400 424.050 675.600 ;
        RECT 352.950 673.950 355.050 674.400 ;
        RECT 421.950 673.950 424.050 674.400 ;
        RECT 469.950 675.600 472.050 676.050 ;
        RECT 475.950 675.600 478.050 676.050 ;
        RECT 469.950 674.400 478.050 675.600 ;
        RECT 469.950 673.950 472.050 674.400 ;
        RECT 475.950 673.950 478.050 674.400 ;
        RECT 598.950 675.600 601.050 676.050 ;
        RECT 619.800 675.600 621.900 676.050 ;
        RECT 598.950 674.400 621.900 675.600 ;
        RECT 598.950 673.950 601.050 674.400 ;
        RECT 619.800 673.950 621.900 674.400 ;
        RECT 622.950 673.950 625.050 676.050 ;
        RECT 688.950 675.600 691.050 676.050 ;
        RECT 697.950 675.600 700.050 676.050 ;
        RECT 688.950 674.400 700.050 675.600 ;
        RECT 688.950 673.950 691.050 674.400 ;
        RECT 697.950 673.950 700.050 674.400 ;
        RECT 748.950 675.600 751.050 676.050 ;
        RECT 757.950 675.600 760.050 676.050 ;
        RECT 748.950 674.400 760.050 675.600 ;
        RECT 748.950 673.950 751.050 674.400 ;
        RECT 757.950 673.950 760.050 674.400 ;
        RECT 808.950 675.600 811.050 676.050 ;
        RECT 829.950 675.600 832.050 676.050 ;
        RECT 808.950 674.400 832.050 675.600 ;
        RECT 808.950 673.950 811.050 674.400 ;
        RECT 829.950 673.950 832.050 674.400 ;
        RECT 856.950 673.950 859.050 676.050 ;
        RECT 25.950 672.600 28.050 673.050 ;
        RECT 43.950 672.600 46.050 673.050 ;
        RECT 25.950 671.400 46.050 672.600 ;
        RECT 25.950 670.950 28.050 671.400 ;
        RECT 43.950 670.950 46.050 671.400 ;
        RECT 121.950 672.600 124.050 673.050 ;
        RECT 127.950 672.600 130.050 673.050 ;
        RECT 121.950 671.400 130.050 672.600 ;
        RECT 121.950 670.950 124.050 671.400 ;
        RECT 127.950 670.950 130.050 671.400 ;
        RECT 157.950 672.600 160.050 673.050 ;
        RECT 184.950 672.600 187.050 673.050 ;
        RECT 157.950 671.400 187.050 672.600 ;
        RECT 157.950 670.950 160.050 671.400 ;
        RECT 184.950 670.950 187.050 671.400 ;
        RECT 220.950 672.600 223.050 673.050 ;
        RECT 253.950 672.600 256.050 673.050 ;
        RECT 220.950 671.400 256.050 672.600 ;
        RECT 220.950 670.950 223.050 671.400 ;
        RECT 253.950 670.950 256.050 671.400 ;
        RECT 262.950 672.600 265.050 673.050 ;
        RECT 277.950 672.600 280.050 673.050 ;
        RECT 286.950 672.600 289.050 673.050 ;
        RECT 262.950 671.400 289.050 672.600 ;
        RECT 262.950 670.950 265.050 671.400 ;
        RECT 277.950 670.950 280.050 671.400 ;
        RECT 286.950 670.950 289.050 671.400 ;
        RECT 310.950 672.600 313.050 673.050 ;
        RECT 325.800 672.600 327.900 673.050 ;
        RECT 310.950 671.400 327.900 672.600 ;
        RECT 310.950 670.950 313.050 671.400 ;
        RECT 325.800 670.950 327.900 671.400 ;
        RECT 328.950 672.600 331.050 672.900 ;
        RECT 343.950 672.600 346.050 673.050 ;
        RECT 328.950 671.400 346.050 672.600 ;
        RECT 328.950 670.800 331.050 671.400 ;
        RECT 343.950 670.950 346.050 671.400 ;
        RECT 436.950 672.600 439.050 673.050 ;
        RECT 496.950 672.600 499.050 673.050 ;
        RECT 532.950 672.600 535.050 673.050 ;
        RECT 436.950 671.400 535.050 672.600 ;
        RECT 436.950 670.950 439.050 671.400 ;
        RECT 496.950 670.950 499.050 671.400 ;
        RECT 532.950 670.950 535.050 671.400 ;
        RECT 541.950 672.600 544.050 673.050 ;
        RECT 577.950 672.600 580.050 673.050 ;
        RECT 541.950 671.400 580.050 672.600 ;
        RECT 541.950 670.950 544.050 671.400 ;
        RECT 577.950 670.950 580.050 671.400 ;
        RECT 631.950 672.600 634.050 673.050 ;
        RECT 643.800 672.600 645.900 673.050 ;
        RECT 631.950 671.400 645.900 672.600 ;
        RECT 631.950 670.950 634.050 671.400 ;
        RECT 643.800 670.950 645.900 671.400 ;
        RECT 646.950 672.600 649.050 673.050 ;
        RECT 685.950 672.600 688.050 673.050 ;
        RECT 646.950 671.400 688.050 672.600 ;
        RECT 646.950 670.950 649.050 671.400 ;
        RECT 685.950 670.950 688.050 671.400 ;
        RECT 691.950 672.600 694.050 673.050 ;
        RECT 700.950 672.600 703.050 673.050 ;
        RECT 691.950 671.400 703.050 672.600 ;
        RECT 691.950 670.950 694.050 671.400 ;
        RECT 700.950 670.950 703.050 671.400 ;
        RECT 715.950 672.600 718.050 673.050 ;
        RECT 763.950 672.600 766.050 673.050 ;
        RECT 787.950 672.600 790.050 673.050 ;
        RECT 715.950 671.400 790.050 672.600 ;
        RECT 715.950 670.950 718.050 671.400 ;
        RECT 763.950 670.950 766.050 671.400 ;
        RECT 787.950 670.950 790.050 671.400 ;
        RECT 805.950 672.600 808.050 673.050 ;
        RECT 820.950 672.600 823.050 673.050 ;
        RECT 805.950 671.400 823.050 672.600 ;
        RECT 805.950 670.950 808.050 671.400 ;
        RECT 820.950 670.950 823.050 671.400 ;
        RECT 883.950 672.600 886.050 673.050 ;
        RECT 913.950 672.600 916.050 673.050 ;
        RECT 883.950 671.400 916.050 672.600 ;
        RECT 883.950 670.950 886.050 671.400 ;
        RECT 913.950 670.950 916.050 671.400 ;
        RECT 13.950 669.600 16.050 670.050 ;
        RECT 61.950 669.600 64.050 670.050 ;
        RECT 79.950 669.600 82.050 670.050 ;
        RECT 13.950 668.400 82.050 669.600 ;
        RECT 13.950 667.950 16.050 668.400 ;
        RECT 61.950 667.950 64.050 668.400 ;
        RECT 79.950 667.950 82.050 668.400 ;
        RECT 85.950 669.600 88.050 670.050 ;
        RECT 115.950 669.600 118.050 670.050 ;
        RECT 85.950 668.400 118.050 669.600 ;
        RECT 85.950 667.950 88.050 668.400 ;
        RECT 115.950 667.950 118.050 668.400 ;
        RECT 172.950 669.600 175.050 670.050 ;
        RECT 217.950 669.600 220.050 670.050 ;
        RECT 172.950 668.400 220.050 669.600 ;
        RECT 172.950 667.950 175.050 668.400 ;
        RECT 217.950 667.950 220.050 668.400 ;
        RECT 322.950 669.600 325.050 670.050 ;
        RECT 367.950 669.600 370.050 670.050 ;
        RECT 322.950 668.400 370.050 669.600 ;
        RECT 322.950 667.950 325.050 668.400 ;
        RECT 367.950 667.950 370.050 668.400 ;
        RECT 430.950 669.600 433.050 670.050 ;
        RECT 589.950 669.600 592.050 670.050 ;
        RECT 430.950 668.400 592.050 669.600 ;
        RECT 430.950 667.950 433.050 668.400 ;
        RECT 589.950 667.950 592.050 668.400 ;
        RECT 673.950 669.600 676.050 670.050 ;
        RECT 712.950 669.600 715.050 670.050 ;
        RECT 673.950 668.400 715.050 669.600 ;
        RECT 673.950 667.950 676.050 668.400 ;
        RECT 712.950 667.950 715.050 668.400 ;
        RECT 721.950 669.600 724.050 670.050 ;
        RECT 799.950 669.600 802.050 670.050 ;
        RECT 826.950 669.600 829.050 670.050 ;
        RECT 835.950 669.600 838.050 670.050 ;
        RECT 721.950 668.400 838.050 669.600 ;
        RECT 721.950 667.950 724.050 668.400 ;
        RECT 799.950 667.950 802.050 668.400 ;
        RECT 826.950 667.950 829.050 668.400 ;
        RECT 835.950 667.950 838.050 668.400 ;
        RECT 898.950 669.600 901.050 670.050 ;
        RECT 913.950 669.600 916.050 669.900 ;
        RECT 898.950 668.400 916.050 669.600 ;
        RECT 898.950 667.950 901.050 668.400 ;
        RECT 913.950 667.800 916.050 668.400 ;
        RECT 175.950 666.600 178.050 667.050 ;
        RECT 196.800 666.600 198.900 667.050 ;
        RECT 175.950 665.400 198.900 666.600 ;
        RECT 175.950 664.950 178.050 665.400 ;
        RECT 196.800 664.950 198.900 665.400 ;
        RECT 199.950 666.600 202.050 667.050 ;
        RECT 211.950 666.600 214.050 667.050 ;
        RECT 199.950 665.400 214.050 666.600 ;
        RECT 199.950 664.950 202.050 665.400 ;
        RECT 211.950 664.950 214.050 665.400 ;
        RECT 370.950 666.600 373.050 667.050 ;
        RECT 397.950 666.600 400.050 667.050 ;
        RECT 370.950 665.400 400.050 666.600 ;
        RECT 370.950 664.950 373.050 665.400 ;
        RECT 397.950 664.950 400.050 665.400 ;
        RECT 403.950 666.600 406.050 667.050 ;
        RECT 418.950 666.600 421.050 667.050 ;
        RECT 403.950 665.400 421.050 666.600 ;
        RECT 403.950 664.950 406.050 665.400 ;
        RECT 418.950 664.950 421.050 665.400 ;
        RECT 439.950 666.600 442.050 667.050 ;
        RECT 454.950 666.600 457.050 667.050 ;
        RECT 439.950 665.400 457.050 666.600 ;
        RECT 439.950 664.950 442.050 665.400 ;
        RECT 454.950 664.950 457.050 665.400 ;
        RECT 535.950 666.600 538.050 667.050 ;
        RECT 556.950 666.600 559.050 667.050 ;
        RECT 535.950 665.400 559.050 666.600 ;
        RECT 535.950 664.950 538.050 665.400 ;
        RECT 556.950 664.950 559.050 665.400 ;
        RECT 676.950 666.600 679.050 667.050 ;
        RECT 688.950 666.600 691.050 667.050 ;
        RECT 676.950 665.400 691.050 666.600 ;
        RECT 676.950 664.950 679.050 665.400 ;
        RECT 688.950 664.950 691.050 665.400 ;
        RECT 694.950 666.600 697.050 667.050 ;
        RECT 736.950 666.600 739.050 667.050 ;
        RECT 694.950 665.400 739.050 666.600 ;
        RECT 694.950 664.950 697.050 665.400 ;
        RECT 736.950 664.950 739.050 665.400 ;
        RECT 763.950 666.600 766.050 667.050 ;
        RECT 769.950 666.600 772.050 667.050 ;
        RECT 763.950 665.400 772.050 666.600 ;
        RECT 763.950 664.950 766.050 665.400 ;
        RECT 769.950 664.950 772.050 665.400 ;
        RECT 781.950 666.600 784.050 667.050 ;
        RECT 808.950 666.600 811.050 667.050 ;
        RECT 781.950 665.400 811.050 666.600 ;
        RECT 781.950 664.950 784.050 665.400 ;
        RECT 808.950 664.950 811.050 665.400 ;
        RECT 856.950 666.600 859.050 667.050 ;
        RECT 871.950 666.600 874.050 667.050 ;
        RECT 856.950 665.400 874.050 666.600 ;
        RECT 856.950 664.950 859.050 665.400 ;
        RECT 871.950 664.950 874.050 665.400 ;
        RECT 145.950 663.600 148.050 664.050 ;
        RECT 166.800 663.600 168.900 664.050 ;
        RECT 145.950 662.400 168.900 663.600 ;
        RECT 145.950 661.950 148.050 662.400 ;
        RECT 166.800 661.950 168.900 662.400 ;
        RECT 169.950 663.600 172.050 664.050 ;
        RECT 247.950 663.600 250.050 664.050 ;
        RECT 169.950 662.400 250.050 663.600 ;
        RECT 169.950 661.950 172.050 662.400 ;
        RECT 247.950 661.950 250.050 662.400 ;
        RECT 277.950 663.600 280.050 664.050 ;
        RECT 295.950 663.600 298.050 664.050 ;
        RECT 277.950 662.400 298.050 663.600 ;
        RECT 277.950 661.950 280.050 662.400 ;
        RECT 295.950 661.950 298.050 662.400 ;
        RECT 343.950 663.600 346.050 664.050 ;
        RECT 364.950 663.600 367.050 664.050 ;
        RECT 343.950 662.400 367.050 663.600 ;
        RECT 343.950 661.950 346.050 662.400 ;
        RECT 364.950 661.950 367.050 662.400 ;
        RECT 373.950 663.600 376.050 664.050 ;
        RECT 379.950 663.600 382.050 664.050 ;
        RECT 373.950 662.400 382.050 663.600 ;
        RECT 373.950 661.950 376.050 662.400 ;
        RECT 379.950 661.950 382.050 662.400 ;
        RECT 409.950 663.600 412.050 664.050 ;
        RECT 457.950 663.600 460.050 664.050 ;
        RECT 481.950 663.600 484.050 664.050 ;
        RECT 409.950 662.400 484.050 663.600 ;
        RECT 409.950 661.950 412.050 662.400 ;
        RECT 457.950 661.950 460.050 662.400 ;
        RECT 481.950 661.950 484.050 662.400 ;
        RECT 493.950 663.600 496.050 664.050 ;
        RECT 595.950 663.600 598.050 664.050 ;
        RECT 493.950 662.400 598.050 663.600 ;
        RECT 493.950 661.950 496.050 662.400 ;
        RECT 595.950 661.950 598.050 662.400 ;
        RECT 607.950 663.600 610.050 664.050 ;
        RECT 634.950 663.600 637.050 664.050 ;
        RECT 607.950 662.400 637.050 663.600 ;
        RECT 607.950 661.950 610.050 662.400 ;
        RECT 634.950 661.950 637.050 662.400 ;
        RECT 670.950 663.600 673.050 664.050 ;
        RECT 691.950 663.600 694.050 664.050 ;
        RECT 670.950 662.400 694.050 663.600 ;
        RECT 670.950 661.950 673.050 662.400 ;
        RECT 691.950 661.950 694.050 662.400 ;
        RECT 697.950 663.600 700.050 664.050 ;
        RECT 709.950 663.600 712.050 664.050 ;
        RECT 697.950 662.400 712.050 663.600 ;
        RECT 697.950 661.950 700.050 662.400 ;
        RECT 709.950 661.950 712.050 662.400 ;
        RECT 838.950 663.600 841.050 664.050 ;
        RECT 844.950 663.600 847.050 664.050 ;
        RECT 838.950 662.400 847.050 663.600 ;
        RECT 838.950 661.950 841.050 662.400 ;
        RECT 844.950 661.950 847.050 662.400 ;
        RECT 892.950 663.600 895.050 664.050 ;
        RECT 901.950 663.600 904.050 664.050 ;
        RECT 916.950 663.600 919.050 664.050 ;
        RECT 892.950 662.400 919.050 663.600 ;
        RECT 892.950 661.950 895.050 662.400 ;
        RECT 901.950 661.950 904.050 662.400 ;
        RECT 916.950 661.950 919.050 662.400 ;
        RECT 91.950 660.600 94.050 661.050 ;
        RECT 97.950 660.600 100.050 661.050 ;
        RECT 130.950 660.600 133.050 661.050 ;
        RECT 91.950 659.400 133.050 660.600 ;
        RECT 91.950 658.950 94.050 659.400 ;
        RECT 97.950 658.950 100.050 659.400 ;
        RECT 130.950 658.950 133.050 659.400 ;
        RECT 142.950 660.600 145.050 661.050 ;
        RECT 148.950 660.600 151.050 661.050 ;
        RECT 250.950 660.600 253.050 661.050 ;
        RECT 142.950 659.400 253.050 660.600 ;
        RECT 142.950 658.950 145.050 659.400 ;
        RECT 148.950 658.950 151.050 659.400 ;
        RECT 250.950 658.950 253.050 659.400 ;
        RECT 280.950 660.600 283.050 661.050 ;
        RECT 319.950 660.600 322.050 661.050 ;
        RECT 280.950 659.400 322.050 660.600 ;
        RECT 280.950 658.950 283.050 659.400 ;
        RECT 319.950 658.950 322.050 659.400 ;
        RECT 361.950 660.600 364.050 661.050 ;
        RECT 394.950 660.600 397.050 661.050 ;
        RECT 361.950 659.400 397.050 660.600 ;
        RECT 361.950 658.950 364.050 659.400 ;
        RECT 394.950 658.950 397.050 659.400 ;
        RECT 400.950 660.600 403.050 661.050 ;
        RECT 406.950 660.600 409.050 661.050 ;
        RECT 415.950 660.600 418.050 661.050 ;
        RECT 400.950 659.400 418.050 660.600 ;
        RECT 400.950 658.950 403.050 659.400 ;
        RECT 406.950 658.950 409.050 659.400 ;
        RECT 415.950 658.950 418.050 659.400 ;
        RECT 511.950 660.600 514.050 661.050 ;
        RECT 538.950 660.600 541.050 661.050 ;
        RECT 511.950 659.400 541.050 660.600 ;
        RECT 511.950 658.950 514.050 659.400 ;
        RECT 538.950 658.950 541.050 659.400 ;
        RECT 556.950 660.600 559.050 661.050 ;
        RECT 592.950 660.600 595.050 661.050 ;
        RECT 556.950 659.400 595.050 660.600 ;
        RECT 556.950 658.950 559.050 659.400 ;
        RECT 592.950 658.950 595.050 659.400 ;
        RECT 667.950 660.600 670.050 661.050 ;
        RECT 694.950 660.600 697.050 661.050 ;
        RECT 667.950 659.400 697.050 660.600 ;
        RECT 667.950 658.950 670.050 659.400 ;
        RECT 694.950 658.950 697.050 659.400 ;
        RECT 709.950 660.600 712.050 660.900 ;
        RECT 715.950 660.600 718.050 661.050 ;
        RECT 709.950 659.400 718.050 660.600 ;
        RECT 709.950 658.800 712.050 659.400 ;
        RECT 715.950 658.950 718.050 659.400 ;
        RECT 856.950 660.600 859.050 661.050 ;
        RECT 865.950 660.600 868.050 661.050 ;
        RECT 856.950 659.400 868.050 660.600 ;
        RECT 856.950 658.950 859.050 659.400 ;
        RECT 865.950 658.950 868.050 659.400 ;
        RECT 34.950 657.600 37.050 658.050 ;
        RECT 55.950 657.600 58.050 658.050 ;
        RECT 34.950 656.400 58.050 657.600 ;
        RECT 34.950 655.950 37.050 656.400 ;
        RECT 55.950 655.950 58.050 656.400 ;
        RECT 127.950 657.600 130.050 658.050 ;
        RECT 223.950 657.600 226.050 658.050 ;
        RECT 127.950 656.400 226.050 657.600 ;
        RECT 127.950 655.950 130.050 656.400 ;
        RECT 223.950 655.950 226.050 656.400 ;
        RECT 235.950 657.600 238.050 658.050 ;
        RECT 271.950 657.600 274.050 658.050 ;
        RECT 235.950 656.400 274.050 657.600 ;
        RECT 235.950 655.950 238.050 656.400 ;
        RECT 271.950 655.950 274.050 656.400 ;
        RECT 367.950 657.600 370.050 658.050 ;
        RECT 409.950 657.600 412.050 658.050 ;
        RECT 367.950 656.400 412.050 657.600 ;
        RECT 367.950 655.950 370.050 656.400 ;
        RECT 409.950 655.950 412.050 656.400 ;
        RECT 418.950 657.600 421.050 658.050 ;
        RECT 436.950 657.600 439.050 658.050 ;
        RECT 418.950 656.400 439.050 657.600 ;
        RECT 418.950 655.950 421.050 656.400 ;
        RECT 436.950 655.950 439.050 656.400 ;
        RECT 493.950 657.600 496.050 658.050 ;
        RECT 499.950 657.600 502.050 658.050 ;
        RECT 493.950 656.400 502.050 657.600 ;
        RECT 493.950 655.950 496.050 656.400 ;
        RECT 499.950 655.950 502.050 656.400 ;
        RECT 517.950 657.600 520.050 658.050 ;
        RECT 529.950 657.600 532.050 658.050 ;
        RECT 517.950 656.400 532.050 657.600 ;
        RECT 517.950 655.950 520.050 656.400 ;
        RECT 529.950 655.950 532.050 656.400 ;
        RECT 643.950 657.600 646.050 658.050 ;
        RECT 676.800 657.600 678.900 658.050 ;
        RECT 643.950 656.400 678.900 657.600 ;
        RECT 643.950 655.950 646.050 656.400 ;
        RECT 676.800 655.950 678.900 656.400 ;
        RECT 679.950 657.600 682.050 658.050 ;
        RECT 721.950 657.600 724.050 658.050 ;
        RECT 679.950 656.400 724.050 657.600 ;
        RECT 679.950 655.950 682.050 656.400 ;
        RECT 721.950 655.950 724.050 656.400 ;
        RECT 757.950 657.600 760.050 658.050 ;
        RECT 766.950 657.600 769.050 658.050 ;
        RECT 757.950 656.400 769.050 657.600 ;
        RECT 757.950 655.950 760.050 656.400 ;
        RECT 766.950 655.950 769.050 656.400 ;
        RECT 790.950 657.600 793.050 658.050 ;
        RECT 844.950 657.600 847.050 658.050 ;
        RECT 790.950 656.400 847.050 657.600 ;
        RECT 790.950 655.950 793.050 656.400 ;
        RECT 844.950 655.950 847.050 656.400 ;
        RECT 889.950 657.600 892.050 658.050 ;
        RECT 910.950 657.600 913.050 658.050 ;
        RECT 889.950 656.400 913.050 657.600 ;
        RECT 889.950 655.950 892.050 656.400 ;
        RECT 910.950 655.950 913.050 656.400 ;
        RECT 37.950 652.950 40.050 655.050 ;
        RECT 43.950 654.600 46.050 655.050 ;
        RECT 67.950 654.600 70.050 655.050 ;
        RECT 43.950 653.400 70.050 654.600 ;
        RECT 43.950 652.950 46.050 653.400 ;
        RECT 67.950 652.950 70.050 653.400 ;
        RECT 109.950 654.600 112.050 655.050 ;
        RECT 118.950 654.600 121.050 655.050 ;
        RECT 109.950 653.400 121.050 654.600 ;
        RECT 109.950 652.950 112.050 653.400 ;
        RECT 118.950 652.950 121.050 653.400 ;
        RECT 163.950 654.600 166.050 655.050 ;
        RECT 172.950 654.600 175.050 655.050 ;
        RECT 163.950 653.400 175.050 654.600 ;
        RECT 163.950 652.950 166.050 653.400 ;
        RECT 172.950 652.950 175.050 653.400 ;
        RECT 178.950 654.600 181.050 655.050 ;
        RECT 199.950 654.600 202.050 655.050 ;
        RECT 178.950 653.400 202.050 654.600 ;
        RECT 178.950 652.950 181.050 653.400 ;
        RECT 199.950 652.950 202.050 653.400 ;
        RECT 298.950 654.600 303.000 655.050 ;
        RECT 364.950 654.600 367.050 655.050 ;
        RECT 403.950 654.600 406.050 655.050 ;
        RECT 298.950 652.950 303.600 654.600 ;
        RECT 364.950 653.400 406.050 654.600 ;
        RECT 364.950 652.950 367.050 653.400 ;
        RECT 403.950 652.950 406.050 653.400 ;
        RECT 592.950 654.600 595.050 655.050 ;
        RECT 610.950 654.600 613.050 655.050 ;
        RECT 592.950 653.400 613.050 654.600 ;
        RECT 592.950 652.950 595.050 653.400 ;
        RECT 610.950 652.950 613.050 653.400 ;
        RECT 658.950 654.600 661.050 655.050 ;
        RECT 682.950 654.600 685.050 655.050 ;
        RECT 658.950 653.400 685.050 654.600 ;
        RECT 658.950 652.950 661.050 653.400 ;
        RECT 682.950 652.950 685.050 653.400 ;
        RECT 688.950 654.600 691.050 655.050 ;
        RECT 703.950 654.600 706.050 655.050 ;
        RECT 688.950 653.400 706.050 654.600 ;
        RECT 688.950 652.950 691.050 653.400 ;
        RECT 703.950 652.950 706.050 653.400 ;
        RECT 748.950 654.600 751.050 655.050 ;
        RECT 754.950 654.600 757.050 655.050 ;
        RECT 748.950 653.400 757.050 654.600 ;
        RECT 748.950 652.950 751.050 653.400 ;
        RECT 754.950 652.950 757.050 653.400 ;
        RECT 760.950 652.950 763.050 655.050 ;
        RECT 847.950 654.600 850.050 655.050 ;
        RECT 859.950 654.600 862.050 655.050 ;
        RECT 886.950 654.600 889.050 655.050 ;
        RECT 847.950 653.400 858.600 654.600 ;
        RECT 847.950 652.950 850.050 653.400 ;
        RECT 7.950 651.750 10.050 652.200 ;
        RECT 13.950 651.750 16.050 652.200 ;
        RECT 7.950 650.550 16.050 651.750 ;
        RECT 7.950 650.100 10.050 650.550 ;
        RECT 13.950 650.100 16.050 650.550 ;
        RECT 22.950 651.600 25.050 652.050 ;
        RECT 22.950 650.400 33.600 651.600 ;
        RECT 22.950 649.950 25.050 650.400 ;
        RECT 16.950 645.600 19.050 645.900 ;
        RECT 25.950 645.600 28.050 646.050 ;
        RECT 32.400 645.900 33.600 650.400 ;
        RECT 38.400 648.600 39.600 652.950 ;
        RECT 40.950 651.750 43.050 652.200 ;
        RECT 46.800 651.750 48.900 652.200 ;
        RECT 40.950 650.550 48.900 651.750 ;
        RECT 40.950 650.100 43.050 650.550 ;
        RECT 46.800 650.100 48.900 650.550 ;
        RECT 49.950 648.600 52.050 652.050 ;
        RECT 79.950 651.600 82.050 652.200 ;
        RECT 71.400 650.400 82.050 651.600 ;
        RECT 38.400 647.400 48.600 648.600 ;
        RECT 49.950 648.000 57.600 648.600 ;
        RECT 50.400 647.400 57.600 648.000 ;
        RECT 16.950 644.400 28.050 645.600 ;
        RECT 16.950 643.800 19.050 644.400 ;
        RECT 25.950 643.950 28.050 644.400 ;
        RECT 31.950 643.800 34.050 645.900 ;
        RECT 47.400 645.600 48.600 647.400 ;
        RECT 52.950 645.600 55.050 645.900 ;
        RECT 47.400 644.400 55.050 645.600 ;
        RECT 56.400 645.600 57.600 647.400 ;
        RECT 71.400 646.050 72.600 650.400 ;
        RECT 79.950 650.100 82.050 650.400 ;
        RECT 100.950 650.100 103.050 652.200 ;
        RECT 175.950 651.600 178.050 652.200 ;
        RECT 175.950 650.400 180.600 651.600 ;
        RECT 175.950 650.100 178.050 650.400 ;
        RECT 101.400 646.050 102.600 650.100 ;
        RECT 179.400 646.050 180.600 650.400 ;
        RECT 265.950 650.100 268.050 652.200 ;
        RECT 280.950 651.600 283.050 652.050 ;
        RECT 275.400 650.400 283.050 651.600 ;
        RECT 302.400 651.600 303.600 652.950 ;
        RECT 352.950 651.600 355.050 652.050 ;
        RECT 302.400 650.400 355.050 651.600 ;
        RECT 190.950 648.600 193.050 649.050 ;
        RECT 208.800 648.600 210.900 649.050 ;
        RECT 190.950 647.400 210.900 648.600 ;
        RECT 190.950 646.950 193.050 647.400 ;
        RECT 208.800 646.950 210.900 647.400 ;
        RECT 64.950 645.600 67.050 646.050 ;
        RECT 56.400 644.400 67.050 645.600 ;
        RECT 52.950 643.800 55.050 644.400 ;
        RECT 64.950 643.950 67.050 644.400 ;
        RECT 70.950 643.950 73.050 646.050 ;
        RECT 101.400 644.400 106.050 646.050 ;
        RECT 102.000 643.950 106.050 644.400 ;
        RECT 121.950 645.450 124.050 645.900 ;
        RECT 151.950 645.450 154.050 645.900 ;
        RECT 121.950 644.250 154.050 645.450 ;
        RECT 121.950 643.800 124.050 644.250 ;
        RECT 151.950 643.800 154.050 644.250 ;
        RECT 157.950 645.450 160.050 645.900 ;
        RECT 163.950 645.450 166.050 645.900 ;
        RECT 157.950 644.250 166.050 645.450 ;
        RECT 179.400 644.400 184.050 646.050 ;
        RECT 211.950 645.600 214.050 649.050 ;
        RECT 244.950 645.600 247.050 646.050 ;
        RECT 211.950 645.000 247.050 645.600 ;
        RECT 212.400 644.400 247.050 645.000 ;
        RECT 157.950 643.800 160.050 644.250 ;
        RECT 163.950 643.800 166.050 644.250 ;
        RECT 180.000 643.950 184.050 644.400 ;
        RECT 244.950 643.950 247.050 644.400 ;
        RECT 256.950 645.600 259.050 646.050 ;
        RECT 266.400 645.600 267.600 650.100 ;
        RECT 275.400 645.900 276.600 650.400 ;
        RECT 280.950 649.950 283.050 650.400 ;
        RECT 352.950 649.950 355.050 650.400 ;
        RECT 361.950 649.950 364.050 652.050 ;
        RECT 412.950 651.600 415.050 652.200 ;
        RECT 404.400 650.400 415.050 651.600 ;
        RECT 362.400 646.050 363.600 649.950 ;
        RECT 404.400 646.050 405.600 650.400 ;
        RECT 412.950 650.100 415.050 650.400 ;
        RECT 418.950 651.600 423.000 652.050 ;
        RECT 433.950 651.600 436.050 652.050 ;
        RECT 439.950 651.600 442.050 652.050 ;
        RECT 505.950 651.600 508.050 652.200 ;
        RECT 418.950 649.950 423.600 651.600 ;
        RECT 433.950 650.400 442.050 651.600 ;
        RECT 433.950 649.950 436.050 650.400 ;
        RECT 439.950 649.950 442.050 650.400 ;
        RECT 446.400 650.400 508.050 651.600 ;
        RECT 422.400 646.050 423.600 649.950 ;
        RECT 446.400 646.050 447.600 650.400 ;
        RECT 505.950 650.100 508.050 650.400 ;
        RECT 511.950 651.600 514.050 652.200 ;
        RECT 523.950 651.600 526.050 652.200 ;
        RECT 534.000 651.600 538.050 652.050 ;
        RECT 511.950 650.400 526.050 651.600 ;
        RECT 511.950 650.100 514.050 650.400 ;
        RECT 523.950 650.100 526.050 650.400 ;
        RECT 533.400 649.950 538.050 651.600 ;
        RECT 553.950 650.100 556.050 652.200 ;
        RECT 559.950 650.400 562.050 652.500 ;
        RECT 256.950 644.400 267.600 645.600 ;
        RECT 256.950 643.950 259.050 644.400 ;
        RECT 274.950 643.800 277.050 645.900 ;
        RECT 361.950 643.950 364.050 646.050 ;
        RECT 403.950 643.950 406.050 646.050 ;
        RECT 421.950 643.950 424.050 646.050 ;
        RECT 445.950 643.950 448.050 646.050 ;
        RECT 533.400 645.900 534.600 649.950 ;
        RECT 554.400 646.050 555.600 650.100 ;
        RECT 532.950 643.800 535.050 645.900 ;
        RECT 554.400 644.400 559.050 646.050 ;
        RECT 555.000 643.950 559.050 644.400 ;
        RECT 58.950 642.600 61.050 643.050 ;
        RECT 82.950 642.600 85.050 643.050 ;
        RECT 91.950 642.600 94.050 643.050 ;
        RECT 58.950 641.400 94.050 642.600 ;
        RECT 58.950 640.950 61.050 641.400 ;
        RECT 82.950 640.950 85.050 641.400 ;
        RECT 91.950 640.950 94.050 641.400 ;
        RECT 115.950 642.600 118.050 643.050 ;
        RECT 139.950 642.600 142.050 643.050 ;
        RECT 196.950 642.600 199.050 643.050 ;
        RECT 232.950 642.600 235.050 643.050 ;
        RECT 115.950 641.400 150.600 642.600 ;
        RECT 115.950 640.950 118.050 641.400 ;
        RECT 139.950 640.950 142.050 641.400 ;
        RECT 67.950 639.600 70.050 640.050 ;
        RECT 76.950 639.600 79.050 640.050 ;
        RECT 67.950 638.400 79.050 639.600 ;
        RECT 149.400 639.600 150.600 641.400 ;
        RECT 196.950 641.400 235.050 642.600 ;
        RECT 196.950 640.950 199.050 641.400 ;
        RECT 232.950 640.950 235.050 641.400 ;
        RECT 295.950 642.600 298.050 643.050 ;
        RECT 310.950 642.600 313.050 643.050 ;
        RECT 295.950 641.400 313.050 642.600 ;
        RECT 295.950 640.950 298.050 641.400 ;
        RECT 310.950 640.950 313.050 641.400 ;
        RECT 397.950 642.600 400.050 643.050 ;
        RECT 418.950 642.600 421.050 643.050 ;
        RECT 397.950 641.400 421.050 642.600 ;
        RECT 397.950 640.950 400.050 641.400 ;
        RECT 418.950 640.950 421.050 641.400 ;
        RECT 535.950 642.600 538.050 643.050 ;
        RECT 560.400 642.600 561.600 650.400 ;
        RECT 574.950 649.950 577.050 652.050 ;
        RECT 607.950 650.100 610.050 652.200 ;
        RECT 613.950 650.100 616.050 652.200 ;
        RECT 694.950 650.100 697.050 652.200 ;
        RECT 700.950 650.100 703.050 652.200 ;
        RECT 718.950 651.600 721.050 652.200 ;
        RECT 704.400 650.400 721.050 651.600 ;
        RECT 575.400 646.050 576.600 649.950 ;
        RECT 608.400 648.600 609.600 650.100 ;
        RECT 596.400 647.400 609.600 648.600 ;
        RECT 574.950 643.950 577.050 646.050 ;
        RECT 580.950 645.600 583.050 646.050 ;
        RECT 596.400 645.600 597.600 647.400 ;
        RECT 580.950 644.400 597.600 645.600 ;
        RECT 598.950 645.450 601.050 645.900 ;
        RECT 604.950 645.450 607.050 645.900 ;
        RECT 580.950 643.950 583.050 644.400 ;
        RECT 598.950 644.250 607.050 645.450 ;
        RECT 614.400 645.600 615.600 650.100 ;
        RECT 619.950 645.600 622.050 646.050 ;
        RECT 614.400 644.400 622.050 645.600 ;
        RECT 598.950 643.800 601.050 644.250 ;
        RECT 604.950 643.800 607.050 644.250 ;
        RECT 619.950 643.950 622.050 644.400 ;
        RECT 628.950 645.600 631.050 646.050 ;
        RECT 682.800 645.600 684.900 646.050 ;
        RECT 628.950 644.400 684.900 645.600 ;
        RECT 628.950 643.950 631.050 644.400 ;
        RECT 682.800 643.950 684.900 644.400 ;
        RECT 685.950 645.600 688.050 646.050 ;
        RECT 691.950 645.600 694.050 646.050 ;
        RECT 685.950 644.400 694.050 645.600 ;
        RECT 685.950 643.950 688.050 644.400 ;
        RECT 691.950 643.950 694.050 644.400 ;
        RECT 695.400 643.050 696.600 650.100 ;
        RECT 701.400 643.050 702.600 650.100 ;
        RECT 704.400 645.900 705.600 650.400 ;
        RECT 718.950 650.100 721.050 650.400 ;
        RECT 724.950 651.750 727.050 652.200 ;
        RECT 733.950 651.750 736.050 652.200 ;
        RECT 724.950 651.600 736.050 651.750 ;
        RECT 745.950 651.600 748.050 652.050 ;
        RECT 724.950 650.550 748.050 651.600 ;
        RECT 724.950 650.100 727.050 650.550 ;
        RECT 733.950 650.400 748.050 650.550 ;
        RECT 733.950 650.100 736.050 650.400 ;
        RECT 745.950 649.950 748.050 650.400 ;
        RECT 761.400 648.600 762.600 652.950 ;
        RECT 763.950 650.100 766.050 652.200 ;
        RECT 772.950 651.600 775.050 652.050 ;
        RECT 781.950 651.600 784.050 652.200 ;
        RECT 772.950 650.400 784.050 651.600 ;
        RECT 752.400 648.000 762.600 648.600 ;
        RECT 751.950 647.400 762.600 648.000 ;
        RECT 703.950 643.800 706.050 645.900 ;
        RECT 721.950 645.600 724.050 645.900 ;
        RECT 739.950 645.600 742.050 645.900 ;
        RECT 721.950 644.400 742.050 645.600 ;
        RECT 721.950 643.800 724.050 644.400 ;
        RECT 739.950 643.800 742.050 644.400 ;
        RECT 751.950 643.950 754.050 647.400 ;
        RECT 764.400 643.050 765.600 650.100 ;
        RECT 772.950 649.950 775.050 650.400 ;
        RECT 781.950 650.100 784.050 650.400 ;
        RECT 799.950 651.600 802.050 652.200 ;
        RECT 811.950 651.600 814.050 652.200 ;
        RECT 799.950 650.400 814.050 651.600 ;
        RECT 799.950 650.100 802.050 650.400 ;
        RECT 811.950 650.100 814.050 650.400 ;
        RECT 817.950 650.100 820.050 652.200 ;
        RECT 790.950 645.600 793.050 646.050 ;
        RECT 796.950 645.600 799.050 645.900 ;
        RECT 790.950 644.400 799.050 645.600 ;
        RECT 790.950 643.950 793.050 644.400 ;
        RECT 796.950 643.800 799.050 644.400 ;
        RECT 818.400 643.050 819.600 650.100 ;
        RECT 823.950 649.950 826.050 652.050 ;
        RECT 820.950 645.600 823.050 645.900 ;
        RECT 824.400 645.600 825.600 649.950 ;
        RECT 857.400 646.050 858.600 653.400 ;
        RECT 859.950 653.400 889.050 654.600 ;
        RECT 859.950 652.950 862.050 653.400 ;
        RECT 865.950 651.600 868.050 652.200 ;
        RECT 880.950 651.600 883.050 652.050 ;
        RECT 865.950 650.400 883.050 651.600 ;
        RECT 865.950 650.100 868.050 650.400 ;
        RECT 880.950 649.950 883.050 650.400 ;
        RECT 884.400 646.050 885.600 653.400 ;
        RECT 886.950 652.950 889.050 653.400 ;
        RECT 895.950 649.950 898.050 652.050 ;
        RECT 896.400 646.050 897.600 649.950 ;
        RECT 820.950 644.400 825.600 645.600 ;
        RECT 829.950 645.450 832.050 645.900 ;
        RECT 835.950 645.450 838.050 645.900 ;
        RECT 820.950 643.800 823.050 644.400 ;
        RECT 829.950 644.250 838.050 645.450 ;
        RECT 829.950 643.800 832.050 644.250 ;
        RECT 835.950 643.800 838.050 644.250 ;
        RECT 856.950 643.950 859.050 646.050 ;
        RECT 883.950 643.950 886.050 646.050 ;
        RECT 895.950 643.950 898.050 646.050 ;
        RECT 535.950 641.400 561.600 642.600 ;
        RECT 535.950 640.950 538.050 641.400 ;
        RECT 694.950 640.950 697.050 643.050 ;
        RECT 700.950 640.950 703.050 643.050 ;
        RECT 763.950 640.950 766.050 643.050 ;
        RECT 787.950 642.600 790.050 643.050 ;
        RECT 770.400 641.400 790.050 642.600 ;
        RECT 818.400 642.750 822.000 643.050 ;
        RECT 818.400 641.400 823.050 642.750 ;
        RECT 172.950 639.600 175.050 640.050 ;
        RECT 149.400 638.400 175.050 639.600 ;
        RECT 67.950 637.950 70.050 638.400 ;
        RECT 76.950 637.950 79.050 638.400 ;
        RECT 172.950 637.950 175.050 638.400 ;
        RECT 250.950 639.600 253.050 640.050 ;
        RECT 259.950 639.600 262.050 640.050 ;
        RECT 250.950 638.400 262.050 639.600 ;
        RECT 250.950 637.950 253.050 638.400 ;
        RECT 259.950 637.950 262.050 638.400 ;
        RECT 373.950 639.600 376.050 640.050 ;
        RECT 409.950 639.600 412.050 640.050 ;
        RECT 373.950 638.400 412.050 639.600 ;
        RECT 373.950 637.950 376.050 638.400 ;
        RECT 409.950 637.950 412.050 638.400 ;
        RECT 451.950 639.600 454.050 640.050 ;
        RECT 490.950 639.600 493.050 640.050 ;
        RECT 451.950 638.400 493.050 639.600 ;
        RECT 451.950 637.950 454.050 638.400 ;
        RECT 490.950 637.950 493.050 638.400 ;
        RECT 541.950 639.600 544.050 640.050 ;
        RECT 550.800 639.600 552.900 640.050 ;
        RECT 541.950 638.400 552.900 639.600 ;
        RECT 541.950 637.950 544.050 638.400 ;
        RECT 550.800 637.950 552.900 638.400 ;
        RECT 553.950 639.600 556.050 640.050 ;
        RECT 586.950 639.600 589.050 640.050 ;
        RECT 553.950 638.400 589.050 639.600 ;
        RECT 553.950 637.950 556.050 638.400 ;
        RECT 586.950 637.950 589.050 638.400 ;
        RECT 595.950 639.600 598.050 640.050 ;
        RECT 613.950 639.600 616.050 640.050 ;
        RECT 595.950 638.400 616.050 639.600 ;
        RECT 595.950 637.950 598.050 638.400 ;
        RECT 613.950 637.950 616.050 638.400 ;
        RECT 727.950 639.600 730.050 640.050 ;
        RECT 733.950 639.600 736.050 640.050 ;
        RECT 742.950 639.600 745.050 640.050 ;
        RECT 727.950 638.400 745.050 639.600 ;
        RECT 727.950 637.950 730.050 638.400 ;
        RECT 733.950 637.950 736.050 638.400 ;
        RECT 742.950 637.950 745.050 638.400 ;
        RECT 757.950 639.600 760.050 640.050 ;
        RECT 770.400 639.600 771.600 641.400 ;
        RECT 787.950 640.950 790.050 641.400 ;
        RECT 819.000 640.950 823.050 641.400 ;
        RECT 841.950 642.600 844.050 643.050 ;
        RECT 844.950 642.600 847.050 643.050 ;
        RECT 862.950 642.600 865.050 643.050 ;
        RECT 841.950 641.400 865.050 642.600 ;
        RECT 841.950 640.950 844.050 641.400 ;
        RECT 844.950 640.950 847.050 641.400 ;
        RECT 862.950 640.950 865.050 641.400 ;
        RECT 880.950 642.600 883.050 643.050 ;
        RECT 886.950 642.600 889.050 643.050 ;
        RECT 880.950 641.400 889.050 642.600 ;
        RECT 880.950 640.950 883.050 641.400 ;
        RECT 886.950 640.950 889.050 641.400 ;
        RECT 820.950 640.650 823.050 640.950 ;
        RECT 757.950 638.400 771.600 639.600 ;
        RECT 757.950 637.950 760.050 638.400 ;
        RECT 88.950 636.600 91.050 637.050 ;
        RECT 106.950 636.600 109.050 637.050 ;
        RECT 88.950 635.400 109.050 636.600 ;
        RECT 88.950 634.950 91.050 635.400 ;
        RECT 106.950 634.950 109.050 635.400 ;
        RECT 112.950 636.600 115.050 637.050 ;
        RECT 160.950 636.600 163.050 637.050 ;
        RECT 112.950 635.400 163.050 636.600 ;
        RECT 112.950 634.950 115.050 635.400 ;
        RECT 160.950 634.950 163.050 635.400 ;
        RECT 184.950 636.600 187.050 637.050 ;
        RECT 220.950 636.600 223.050 637.050 ;
        RECT 184.950 635.400 223.050 636.600 ;
        RECT 184.950 634.950 187.050 635.400 ;
        RECT 220.950 634.950 223.050 635.400 ;
        RECT 253.950 636.600 256.050 637.050 ;
        RECT 259.950 636.600 262.050 636.900 ;
        RECT 283.950 636.600 286.050 637.050 ;
        RECT 253.950 635.400 286.050 636.600 ;
        RECT 253.950 634.950 256.050 635.400 ;
        RECT 259.950 634.800 262.050 635.400 ;
        RECT 283.950 634.950 286.050 635.400 ;
        RECT 313.950 636.600 316.050 637.050 ;
        RECT 328.950 636.600 331.050 637.050 ;
        RECT 313.950 635.400 331.050 636.600 ;
        RECT 313.950 634.950 316.050 635.400 ;
        RECT 328.950 634.950 331.050 635.400 ;
        RECT 478.950 636.600 481.050 637.050 ;
        RECT 517.950 636.600 520.050 637.050 ;
        RECT 478.950 635.400 520.050 636.600 ;
        RECT 478.950 634.950 481.050 635.400 ;
        RECT 517.950 634.950 520.050 635.400 ;
        RECT 637.950 636.600 640.050 637.050 ;
        RECT 670.950 636.600 673.050 637.050 ;
        RECT 637.950 635.400 673.050 636.600 ;
        RECT 637.950 634.950 640.050 635.400 ;
        RECT 670.950 634.950 673.050 635.400 ;
        RECT 754.950 636.600 757.050 637.050 ;
        RECT 772.950 636.600 775.050 637.050 ;
        RECT 754.950 635.400 775.050 636.600 ;
        RECT 754.950 634.950 757.050 635.400 ;
        RECT 772.950 634.950 775.050 635.400 ;
        RECT 796.950 636.600 799.050 637.050 ;
        RECT 832.950 636.600 835.050 637.050 ;
        RECT 796.950 635.400 835.050 636.600 ;
        RECT 796.950 634.950 799.050 635.400 ;
        RECT 832.950 634.950 835.050 635.400 ;
        RECT 892.950 636.600 895.050 637.050 ;
        RECT 904.950 636.600 907.050 637.050 ;
        RECT 892.950 635.400 907.050 636.600 ;
        RECT 892.950 634.950 895.050 635.400 ;
        RECT 904.950 634.950 907.050 635.400 ;
        RECT 169.950 633.600 172.050 634.050 ;
        RECT 238.800 633.600 240.900 634.050 ;
        RECT 169.950 632.400 240.900 633.600 ;
        RECT 169.950 631.950 172.050 632.400 ;
        RECT 238.800 631.950 240.900 632.400 ;
        RECT 241.950 633.600 244.050 634.050 ;
        RECT 298.950 633.600 301.050 634.050 ;
        RECT 241.950 632.400 301.050 633.600 ;
        RECT 241.950 631.950 244.050 632.400 ;
        RECT 298.950 631.950 301.050 632.400 ;
        RECT 355.950 633.600 358.050 634.050 ;
        RECT 397.950 633.600 400.050 634.050 ;
        RECT 355.950 632.400 400.050 633.600 ;
        RECT 355.950 631.950 358.050 632.400 ;
        RECT 397.950 631.950 400.050 632.400 ;
        RECT 403.950 633.600 406.050 634.050 ;
        RECT 676.950 633.600 679.050 634.050 ;
        RECT 718.950 633.600 721.050 634.050 ;
        RECT 403.950 632.400 417.600 633.600 ;
        RECT 403.950 631.950 406.050 632.400 ;
        RECT 97.950 630.600 100.050 631.050 ;
        RECT 115.950 630.600 118.050 631.050 ;
        RECT 97.950 629.400 118.050 630.600 ;
        RECT 97.950 628.950 100.050 629.400 ;
        RECT 115.950 628.950 118.050 629.400 ;
        RECT 178.950 630.600 181.050 631.050 ;
        RECT 193.950 630.600 196.050 631.050 ;
        RECT 178.950 629.400 196.050 630.600 ;
        RECT 178.950 628.950 181.050 629.400 ;
        RECT 193.950 628.950 196.050 629.400 ;
        RECT 238.950 630.600 241.050 630.900 ;
        RECT 295.950 630.600 298.050 631.050 ;
        RECT 238.950 629.400 298.050 630.600 ;
        RECT 416.400 630.600 417.600 632.400 ;
        RECT 676.950 632.400 721.050 633.600 ;
        RECT 676.950 631.950 679.050 632.400 ;
        RECT 718.950 631.950 721.050 632.400 ;
        RECT 724.950 633.600 727.050 634.050 ;
        RECT 748.950 633.600 751.050 634.050 ;
        RECT 724.950 632.400 751.050 633.600 ;
        RECT 724.950 631.950 727.050 632.400 ;
        RECT 748.950 631.950 751.050 632.400 ;
        RECT 775.950 633.600 778.050 634.050 ;
        RECT 847.950 633.600 850.050 634.050 ;
        RECT 775.950 632.400 850.050 633.600 ;
        RECT 775.950 631.950 778.050 632.400 ;
        RECT 847.950 631.950 850.050 632.400 ;
        RECT 442.950 630.600 445.050 631.050 ;
        RECT 416.400 629.400 445.050 630.600 ;
        RECT 238.950 628.800 241.050 629.400 ;
        RECT 295.950 628.950 298.050 629.400 ;
        RECT 442.950 628.950 445.050 629.400 ;
        RECT 487.950 630.600 490.050 631.050 ;
        RECT 535.950 630.600 538.050 631.050 ;
        RECT 487.950 629.400 538.050 630.600 ;
        RECT 487.950 628.950 490.050 629.400 ;
        RECT 535.950 628.950 538.050 629.400 ;
        RECT 619.950 630.600 622.050 631.050 ;
        RECT 805.950 630.600 808.050 631.050 ;
        RECT 619.950 629.400 808.050 630.600 ;
        RECT 619.950 628.950 622.050 629.400 ;
        RECT 805.950 628.950 808.050 629.400 ;
        RECT 118.950 627.600 121.050 628.050 ;
        RECT 136.950 627.600 139.050 628.050 ;
        RECT 118.950 626.400 139.050 627.600 ;
        RECT 118.950 625.950 121.050 626.400 ;
        RECT 136.950 625.950 139.050 626.400 ;
        RECT 166.950 627.600 169.050 628.050 ;
        RECT 199.950 627.600 202.050 628.050 ;
        RECT 166.950 626.400 202.050 627.600 ;
        RECT 166.950 625.950 169.050 626.400 ;
        RECT 199.950 625.950 202.050 626.400 ;
        RECT 235.950 627.600 238.050 628.050 ;
        RECT 379.950 627.600 382.050 628.050 ;
        RECT 430.950 627.600 433.050 628.050 ;
        RECT 235.950 626.400 382.050 627.600 ;
        RECT 235.950 625.950 238.050 626.400 ;
        RECT 379.950 625.950 382.050 626.400 ;
        RECT 407.400 626.400 433.050 627.600 ;
        RECT 407.400 625.050 408.600 626.400 ;
        RECT 430.950 625.950 433.050 626.400 ;
        RECT 544.950 627.600 547.050 628.050 ;
        RECT 628.950 627.600 631.050 628.050 ;
        RECT 544.950 626.400 631.050 627.600 ;
        RECT 544.950 625.950 547.050 626.400 ;
        RECT 628.950 625.950 631.050 626.400 ;
        RECT 718.950 627.600 721.050 628.050 ;
        RECT 757.950 627.600 760.050 628.050 ;
        RECT 718.950 626.400 760.050 627.600 ;
        RECT 718.950 625.950 721.050 626.400 ;
        RECT 757.950 625.950 760.050 626.400 ;
        RECT 826.950 627.600 829.050 628.050 ;
        RECT 835.950 627.600 838.050 628.050 ;
        RECT 826.950 626.400 838.050 627.600 ;
        RECT 826.950 625.950 829.050 626.400 ;
        RECT 835.950 625.950 838.050 626.400 ;
        RECT 229.950 624.600 232.050 625.050 ;
        RECT 385.950 624.600 388.050 625.050 ;
        RECT 406.950 624.600 409.050 625.050 ;
        RECT 229.950 623.400 339.600 624.600 ;
        RECT 229.950 622.950 232.050 623.400 ;
        RECT 338.400 622.050 339.600 623.400 ;
        RECT 385.950 623.400 409.050 624.600 ;
        RECT 385.950 622.950 388.050 623.400 ;
        RECT 406.950 622.950 409.050 623.400 ;
        RECT 433.950 624.600 436.050 625.050 ;
        RECT 451.950 624.600 454.050 625.050 ;
        RECT 556.950 624.600 559.050 625.050 ;
        RECT 433.950 623.400 454.050 624.600 ;
        RECT 433.950 622.950 436.050 623.400 ;
        RECT 451.950 622.950 454.050 623.400 ;
        RECT 467.400 623.400 559.050 624.600 ;
        RECT 103.950 621.600 106.050 622.050 ;
        RECT 133.950 621.600 136.050 622.050 ;
        RECT 163.950 621.600 166.050 622.050 ;
        RECT 181.950 621.600 184.050 622.050 ;
        RECT 103.950 620.400 184.050 621.600 ;
        RECT 103.950 619.950 106.050 620.400 ;
        RECT 133.950 619.950 136.050 620.400 ;
        RECT 163.950 619.950 166.050 620.400 ;
        RECT 181.950 619.950 184.050 620.400 ;
        RECT 337.950 621.600 340.050 622.050 ;
        RECT 364.950 621.600 367.050 622.050 ;
        RECT 467.400 621.600 468.600 623.400 ;
        RECT 556.950 622.950 559.050 623.400 ;
        RECT 568.950 624.600 571.050 625.050 ;
        RECT 601.950 624.600 604.050 625.050 ;
        RECT 568.950 623.400 604.050 624.600 ;
        RECT 568.950 622.950 571.050 623.400 ;
        RECT 601.950 622.950 604.050 623.400 ;
        RECT 634.950 624.600 637.050 625.050 ;
        RECT 709.950 624.600 712.050 625.050 ;
        RECT 634.950 623.400 712.050 624.600 ;
        RECT 634.950 622.950 637.050 623.400 ;
        RECT 709.950 622.950 712.050 623.400 ;
        RECT 718.950 624.600 721.050 624.900 ;
        RECT 739.950 624.600 742.050 625.050 ;
        RECT 883.950 624.600 886.050 625.050 ;
        RECT 718.950 623.400 742.050 624.600 ;
        RECT 718.950 622.800 721.050 623.400 ;
        RECT 739.950 622.950 742.050 623.400 ;
        RECT 854.400 623.400 886.050 624.600 ;
        RECT 337.950 620.400 468.600 621.600 ;
        RECT 538.950 621.600 541.050 622.050 ;
        RECT 547.950 621.600 550.050 622.050 ;
        RECT 538.950 620.400 550.050 621.600 ;
        RECT 337.950 619.950 340.050 620.400 ;
        RECT 364.950 619.950 367.050 620.400 ;
        RECT 538.950 619.950 541.050 620.400 ;
        RECT 547.950 619.950 550.050 620.400 ;
        RECT 694.950 621.600 697.050 622.050 ;
        RECT 760.950 621.600 763.050 622.050 ;
        RECT 694.950 620.400 763.050 621.600 ;
        RECT 694.950 619.950 697.050 620.400 ;
        RECT 760.950 619.950 763.050 620.400 ;
        RECT 808.950 621.600 811.050 622.050 ;
        RECT 814.950 621.600 817.050 622.050 ;
        RECT 808.950 620.400 817.050 621.600 ;
        RECT 808.950 619.950 811.050 620.400 ;
        RECT 814.950 619.950 817.050 620.400 ;
        RECT 829.950 621.600 832.050 622.050 ;
        RECT 854.400 621.600 855.600 623.400 ;
        RECT 883.950 622.950 886.050 623.400 ;
        RECT 829.950 620.400 855.600 621.600 ;
        RECT 829.950 619.950 832.050 620.400 ;
        RECT 247.950 618.600 250.050 619.050 ;
        RECT 307.950 618.600 310.050 619.050 ;
        RECT 316.950 618.600 319.050 619.050 ;
        RECT 247.950 617.400 319.050 618.600 ;
        RECT 247.950 616.950 250.050 617.400 ;
        RECT 307.950 616.950 310.050 617.400 ;
        RECT 316.950 616.950 319.050 617.400 ;
        RECT 325.950 618.600 328.050 619.050 ;
        RECT 337.950 618.600 340.050 618.900 ;
        RECT 394.950 618.600 397.050 619.050 ;
        RECT 487.950 618.600 490.050 619.050 ;
        RECT 325.950 617.400 354.600 618.600 ;
        RECT 325.950 616.950 328.050 617.400 ;
        RECT 337.950 616.800 340.050 617.400 ;
        RECT 160.950 615.600 163.050 616.050 ;
        RECT 187.950 615.600 190.050 616.050 ;
        RECT 205.950 615.600 208.050 616.050 ;
        RECT 160.950 614.400 208.050 615.600 ;
        RECT 160.950 613.950 163.050 614.400 ;
        RECT 187.950 613.950 190.050 614.400 ;
        RECT 205.950 613.950 208.050 614.400 ;
        RECT 214.950 615.600 217.050 616.050 ;
        RECT 256.950 615.600 259.050 616.050 ;
        RECT 214.950 614.400 259.050 615.600 ;
        RECT 353.400 615.600 354.600 617.400 ;
        RECT 394.950 617.400 490.050 618.600 ;
        RECT 394.950 616.950 397.050 617.400 ;
        RECT 487.950 616.950 490.050 617.400 ;
        RECT 526.950 618.600 529.050 619.050 ;
        RECT 550.950 618.600 553.050 619.050 ;
        RECT 571.950 618.600 574.050 619.050 ;
        RECT 610.950 618.600 613.050 619.050 ;
        RECT 526.950 617.400 613.050 618.600 ;
        RECT 526.950 616.950 529.050 617.400 ;
        RECT 550.950 616.950 553.050 617.400 ;
        RECT 571.950 616.950 574.050 617.400 ;
        RECT 610.950 616.950 613.050 617.400 ;
        RECT 625.950 618.600 628.050 619.050 ;
        RECT 634.950 618.600 637.050 619.050 ;
        RECT 625.950 617.400 637.050 618.600 ;
        RECT 625.950 616.950 628.050 617.400 ;
        RECT 634.950 616.950 637.050 617.400 ;
        RECT 646.950 618.600 649.050 619.050 ;
        RECT 667.950 618.600 670.050 619.050 ;
        RECT 682.950 618.600 685.050 619.050 ;
        RECT 646.950 617.400 685.050 618.600 ;
        RECT 646.950 616.950 649.050 617.400 ;
        RECT 667.950 616.950 670.050 617.400 ;
        RECT 682.950 616.950 685.050 617.400 ;
        RECT 694.950 618.600 697.050 618.900 ;
        RECT 700.950 618.600 703.050 619.050 ;
        RECT 694.950 617.400 703.050 618.600 ;
        RECT 694.950 616.800 697.050 617.400 ;
        RECT 700.950 616.950 703.050 617.400 ;
        RECT 739.950 618.600 742.050 619.050 ;
        RECT 751.950 618.600 754.050 619.050 ;
        RECT 739.950 617.400 754.050 618.600 ;
        RECT 739.950 616.950 742.050 617.400 ;
        RECT 751.950 616.950 754.050 617.400 ;
        RECT 781.950 618.600 784.050 619.050 ;
        RECT 802.950 618.600 805.050 619.050 ;
        RECT 781.950 617.400 805.050 618.600 ;
        RECT 781.950 616.950 784.050 617.400 ;
        RECT 802.950 616.950 805.050 617.400 ;
        RECT 862.950 618.600 865.050 619.050 ;
        RECT 868.950 618.600 871.050 619.050 ;
        RECT 892.950 618.600 895.050 619.050 ;
        RECT 904.950 618.600 907.050 619.050 ;
        RECT 862.950 617.400 907.050 618.600 ;
        RECT 862.950 616.950 865.050 617.400 ;
        RECT 868.950 616.950 871.050 617.400 ;
        RECT 892.950 616.950 895.050 617.400 ;
        RECT 904.950 616.950 907.050 617.400 ;
        RECT 370.950 615.600 373.050 616.050 ;
        RECT 353.400 614.400 373.050 615.600 ;
        RECT 214.950 613.950 217.050 614.400 ;
        RECT 256.950 613.950 259.050 614.400 ;
        RECT 370.950 613.950 373.050 614.400 ;
        RECT 403.950 615.600 406.050 616.050 ;
        RECT 424.950 615.600 427.050 616.050 ;
        RECT 403.950 614.400 427.050 615.600 ;
        RECT 403.950 613.950 406.050 614.400 ;
        RECT 424.950 613.950 427.050 614.400 ;
        RECT 496.950 615.600 499.050 616.050 ;
        RECT 523.950 615.600 526.050 616.050 ;
        RECT 496.950 614.400 526.050 615.600 ;
        RECT 496.950 613.950 499.050 614.400 ;
        RECT 523.950 613.950 526.050 614.400 ;
        RECT 652.950 615.600 655.050 616.050 ;
        RECT 697.950 615.600 700.050 616.050 ;
        RECT 652.950 614.400 700.050 615.600 ;
        RECT 652.950 613.950 655.050 614.400 ;
        RECT 697.950 613.950 700.050 614.400 ;
        RECT 820.950 615.600 823.050 616.050 ;
        RECT 868.950 615.600 871.050 615.900 ;
        RECT 820.950 614.400 871.050 615.600 ;
        RECT 820.950 613.950 823.050 614.400 ;
        RECT 868.950 613.800 871.050 614.400 ;
        RECT 16.950 612.600 19.050 613.050 ;
        RECT 46.950 612.600 49.050 613.050 ;
        RECT 58.950 612.600 61.050 613.050 ;
        RECT 16.950 611.400 61.050 612.600 ;
        RECT 16.950 610.950 19.050 611.400 ;
        RECT 46.950 610.950 49.050 611.400 ;
        RECT 58.950 610.950 61.050 611.400 ;
        RECT 73.950 612.600 76.050 613.050 ;
        RECT 112.950 612.600 115.050 613.050 ;
        RECT 73.950 611.400 115.050 612.600 ;
        RECT 73.950 610.950 76.050 611.400 ;
        RECT 112.950 610.950 115.050 611.400 ;
        RECT 268.950 612.600 271.050 613.050 ;
        RECT 343.950 612.600 346.050 613.050 ;
        RECT 268.950 611.400 346.050 612.600 ;
        RECT 268.950 610.950 271.050 611.400 ;
        RECT 37.950 609.600 40.050 610.050 ;
        RECT 32.400 608.400 40.050 609.600 ;
        RECT 22.950 606.750 25.050 607.200 ;
        RECT 28.950 606.750 31.050 607.200 ;
        RECT 22.950 605.550 31.050 606.750 ;
        RECT 22.950 605.100 25.050 605.550 ;
        RECT 28.950 605.100 31.050 605.550 ;
        RECT 32.400 601.050 33.600 608.400 ;
        RECT 37.950 607.950 40.050 608.400 ;
        RECT 199.950 609.600 202.050 610.050 ;
        RECT 214.950 609.600 217.050 610.050 ;
        RECT 259.950 609.600 262.050 610.050 ;
        RECT 199.950 608.400 217.050 609.600 ;
        RECT 199.950 607.950 202.050 608.400 ;
        RECT 214.950 607.950 217.050 608.400 ;
        RECT 242.400 608.400 262.050 609.600 ;
        RECT 34.950 606.600 37.050 607.200 ;
        RECT 49.950 606.600 52.050 607.050 ;
        RECT 73.950 606.750 76.050 607.200 ;
        RECT 79.950 606.750 82.050 607.200 ;
        RECT 73.950 606.600 82.050 606.750 ;
        RECT 34.950 605.550 82.050 606.600 ;
        RECT 34.950 605.400 76.050 605.550 ;
        RECT 34.950 605.100 37.050 605.400 ;
        RECT 49.950 604.950 52.050 605.400 ;
        RECT 73.950 605.100 76.050 605.400 ;
        RECT 79.950 605.100 82.050 605.550 ;
        RECT 85.950 606.600 88.050 607.200 ;
        RECT 100.950 606.600 103.050 607.200 ;
        RECT 85.950 605.400 103.050 606.600 ;
        RECT 85.950 605.100 88.050 605.400 ;
        RECT 100.950 605.100 103.050 605.400 ;
        RECT 178.950 606.750 181.050 607.200 ;
        RECT 190.950 606.750 193.050 607.200 ;
        RECT 178.950 605.550 193.050 606.750 ;
        RECT 178.950 605.100 181.050 605.550 ;
        RECT 190.950 605.100 193.050 605.550 ;
        RECT 211.950 606.600 214.050 607.050 ;
        RECT 220.950 606.600 223.050 607.200 ;
        RECT 211.950 605.400 223.050 606.600 ;
        RECT 211.950 604.950 214.050 605.400 ;
        RECT 220.950 605.100 223.050 605.400 ;
        RECT 115.950 603.600 118.050 604.050 ;
        RECT 142.950 603.600 145.050 603.900 ;
        RECT 115.950 602.400 145.050 603.600 ;
        RECT 115.950 601.950 118.050 602.400 ;
        RECT 142.950 601.800 145.050 602.400 ;
        RECT 7.950 600.600 10.050 601.050 ;
        RECT 13.950 600.600 16.050 600.900 ;
        RECT 7.950 599.400 16.050 600.600 ;
        RECT 7.950 598.950 10.050 599.400 ;
        RECT 13.950 598.800 16.050 599.400 ;
        RECT 31.950 598.950 34.050 601.050 ;
        RECT 82.950 600.600 85.050 600.900 ;
        RECT 77.400 600.000 85.050 600.600 ;
        RECT 76.950 599.400 85.050 600.000 ;
        RECT 19.950 597.600 22.050 598.050 ;
        RECT 37.950 597.600 40.050 598.050 ;
        RECT 19.950 596.400 40.050 597.600 ;
        RECT 19.950 595.950 22.050 596.400 ;
        RECT 37.950 595.950 40.050 596.400 ;
        RECT 76.950 595.950 79.050 599.400 ;
        RECT 82.950 598.800 85.050 599.400 ;
        RECT 193.950 600.600 196.050 601.050 ;
        RECT 223.950 600.600 226.050 600.900 ;
        RECT 193.950 599.400 226.050 600.600 ;
        RECT 193.950 598.950 196.050 599.400 ;
        RECT 223.950 598.800 226.050 599.400 ;
        RECT 232.950 600.600 235.050 601.050 ;
        RECT 242.400 600.600 243.600 608.400 ;
        RECT 259.950 607.950 262.050 608.400 ;
        RECT 280.950 609.600 283.050 610.050 ;
        RECT 286.950 609.600 289.050 610.200 ;
        RECT 280.950 608.400 289.050 609.600 ;
        RECT 280.950 607.950 283.050 608.400 ;
        RECT 286.950 608.100 289.050 608.400 ;
        RECT 244.950 606.600 247.050 607.200 ;
        RECT 271.950 606.600 274.050 607.200 ;
        RECT 286.950 606.600 289.050 607.050 ;
        RECT 244.950 605.400 274.050 606.600 ;
        RECT 244.950 605.100 247.050 605.400 ;
        RECT 271.950 605.100 274.050 605.400 ;
        RECT 275.400 605.400 289.050 606.600 ;
        RECT 275.400 603.600 276.600 605.400 ;
        RECT 286.950 604.950 289.050 605.400 ;
        RECT 290.400 603.600 291.600 611.400 ;
        RECT 343.950 610.950 346.050 611.400 ;
        RECT 349.950 612.600 352.050 613.050 ;
        RECT 400.950 612.600 403.050 612.900 ;
        RECT 349.950 611.400 403.050 612.600 ;
        RECT 349.950 610.950 352.050 611.400 ;
        RECT 400.950 610.800 403.050 611.400 ;
        RECT 427.950 612.600 430.050 613.050 ;
        RECT 493.950 612.600 496.050 613.050 ;
        RECT 499.950 612.600 502.050 613.050 ;
        RECT 427.950 611.400 502.050 612.600 ;
        RECT 427.950 610.950 430.050 611.400 ;
        RECT 493.950 610.950 496.050 611.400 ;
        RECT 499.950 610.950 502.050 611.400 ;
        RECT 562.950 612.600 565.050 613.050 ;
        RECT 586.950 612.600 589.050 613.050 ;
        RECT 595.950 612.600 598.050 613.050 ;
        RECT 562.950 611.400 598.050 612.600 ;
        RECT 562.950 610.950 565.050 611.400 ;
        RECT 586.950 610.950 589.050 611.400 ;
        RECT 595.950 610.950 598.050 611.400 ;
        RECT 601.950 612.600 604.050 613.050 ;
        RECT 616.950 612.600 619.050 613.050 ;
        RECT 601.950 611.400 619.050 612.600 ;
        RECT 601.950 610.950 604.050 611.400 ;
        RECT 616.950 610.950 619.050 611.400 ;
        RECT 655.950 612.600 658.050 613.050 ;
        RECT 661.950 612.600 664.050 613.050 ;
        RECT 655.950 611.400 664.050 612.600 ;
        RECT 655.950 610.950 658.050 611.400 ;
        RECT 661.950 610.950 664.050 611.400 ;
        RECT 745.950 612.600 748.050 613.050 ;
        RECT 760.950 612.600 763.050 613.050 ;
        RECT 745.950 611.400 763.050 612.600 ;
        RECT 745.950 610.950 748.050 611.400 ;
        RECT 760.950 610.950 763.050 611.400 ;
        RECT 841.950 612.600 844.050 613.050 ;
        RECT 862.950 612.600 865.050 613.050 ;
        RECT 841.950 611.400 865.050 612.600 ;
        RECT 869.400 612.600 870.600 613.800 ;
        RECT 913.950 612.600 916.050 613.050 ;
        RECT 869.400 611.400 916.050 612.600 ;
        RECT 841.950 610.950 844.050 611.400 ;
        RECT 862.950 610.950 865.050 611.400 ;
        RECT 913.950 610.950 916.050 611.400 ;
        RECT 319.950 609.600 322.050 610.050 ;
        RECT 331.950 609.600 334.050 610.050 ;
        RECT 319.950 608.400 334.050 609.600 ;
        RECT 319.950 607.950 322.050 608.400 ;
        RECT 331.950 607.950 334.050 608.400 ;
        RECT 370.950 609.600 373.050 610.050 ;
        RECT 391.950 609.600 394.050 610.050 ;
        RECT 397.950 609.600 400.050 610.050 ;
        RECT 421.950 609.600 424.050 610.050 ;
        RECT 370.950 608.400 400.050 609.600 ;
        RECT 370.950 607.950 373.050 608.400 ;
        RECT 391.950 607.950 394.050 608.400 ;
        RECT 397.950 607.950 400.050 608.400 ;
        RECT 410.400 608.400 424.050 609.600 ;
        RECT 295.950 606.750 298.050 607.200 ;
        RECT 307.950 606.750 310.050 607.200 ;
        RECT 295.950 605.550 310.050 606.750 ;
        RECT 295.950 605.100 298.050 605.550 ;
        RECT 307.950 605.100 310.050 605.550 ;
        RECT 322.950 606.600 325.050 607.200 ;
        RECT 331.950 606.600 334.050 606.900 ;
        RECT 349.950 606.600 352.050 607.200 ;
        RECT 322.950 605.400 352.050 606.600 ;
        RECT 322.950 605.100 325.050 605.400 ;
        RECT 331.950 604.800 334.050 605.400 ;
        RECT 349.950 605.100 352.050 605.400 ;
        RECT 394.950 603.600 397.050 607.050 ;
        RECT 269.400 602.400 276.600 603.600 ;
        RECT 284.400 602.400 291.600 603.600 ;
        RECT 380.400 603.000 397.050 603.600 ;
        RECT 410.400 603.600 411.600 608.400 ;
        RECT 421.950 607.950 424.050 608.400 ;
        RECT 502.950 607.950 505.050 610.050 ;
        RECT 607.950 609.600 610.050 610.050 ;
        RECT 628.800 609.600 630.900 610.050 ;
        RECT 607.950 608.400 630.900 609.600 ;
        RECT 607.950 607.950 610.050 608.400 ;
        RECT 628.800 607.950 630.900 608.400 ;
        RECT 631.950 609.600 634.050 610.050 ;
        RECT 766.950 609.600 769.050 610.050 ;
        RECT 772.950 609.600 775.050 610.050 ;
        RECT 631.950 608.400 642.600 609.600 ;
        RECT 631.950 607.950 634.050 608.400 ;
        RECT 412.950 606.600 415.050 607.200 ;
        RECT 427.950 606.600 430.050 607.200 ;
        RECT 439.950 606.600 442.050 607.050 ;
        RECT 412.950 605.400 442.050 606.600 ;
        RECT 475.950 605.400 478.050 607.500 ;
        RECT 484.950 605.400 487.050 607.500 ;
        RECT 412.950 605.100 415.050 605.400 ;
        RECT 427.950 605.100 430.050 605.400 ;
        RECT 439.950 604.950 442.050 605.400 ;
        RECT 380.400 602.400 396.600 603.000 ;
        RECT 410.400 602.400 426.600 603.600 ;
        RECT 269.400 600.900 270.600 602.400 ;
        RECT 284.400 600.900 285.600 602.400 ;
        RECT 232.950 599.400 243.600 600.600 ;
        RECT 232.950 598.950 235.050 599.400 ;
        RECT 268.950 598.800 271.050 600.900 ;
        RECT 283.950 598.800 286.050 600.900 ;
        RECT 313.950 600.600 316.050 601.050 ;
        RECT 352.950 600.600 355.050 601.050 ;
        RECT 380.400 600.600 381.600 602.400 ;
        RECT 425.400 600.900 426.600 602.400 ;
        RECT 476.400 601.050 477.600 605.400 ;
        RECT 485.400 603.600 486.600 605.400 ;
        RECT 493.950 603.600 496.050 604.050 ;
        RECT 485.400 602.400 496.050 603.600 ;
        RECT 493.950 601.950 496.050 602.400 ;
        RECT 313.950 599.400 381.600 600.600 ;
        RECT 385.950 600.450 388.050 600.900 ;
        RECT 403.950 600.450 406.050 600.900 ;
        RECT 313.950 598.950 316.050 599.400 ;
        RECT 352.950 598.950 355.050 599.400 ;
        RECT 385.950 599.250 406.050 600.450 ;
        RECT 385.950 598.800 388.050 599.250 ;
        RECT 403.950 598.800 406.050 599.250 ;
        RECT 409.950 600.600 412.050 600.900 ;
        RECT 409.950 600.000 417.600 600.600 ;
        RECT 409.950 599.400 418.050 600.000 ;
        RECT 409.950 598.800 412.050 599.400 ;
        RECT 106.950 597.600 109.050 598.050 ;
        RECT 151.950 597.600 154.050 598.050 ;
        RECT 265.950 597.600 268.050 598.050 ;
        RECT 106.950 596.400 154.050 597.600 ;
        RECT 106.950 595.950 109.050 596.400 ;
        RECT 151.950 595.950 154.050 596.400 ;
        RECT 257.400 596.400 268.050 597.600 ;
        RECT 70.950 594.600 73.050 595.050 ;
        RECT 100.950 594.600 103.050 595.050 ;
        RECT 70.950 593.400 103.050 594.600 ;
        RECT 70.950 592.950 73.050 593.400 ;
        RECT 100.950 592.950 103.050 593.400 ;
        RECT 187.950 594.600 190.050 595.050 ;
        RECT 208.950 594.600 211.050 595.050 ;
        RECT 187.950 593.400 211.050 594.600 ;
        RECT 187.950 592.950 190.050 593.400 ;
        RECT 208.950 592.950 211.050 593.400 ;
        RECT 217.950 594.600 220.050 595.050 ;
        RECT 235.950 594.600 238.050 595.050 ;
        RECT 217.950 593.400 238.050 594.600 ;
        RECT 217.950 592.950 220.050 593.400 ;
        RECT 235.950 592.950 238.050 593.400 ;
        RECT 241.950 594.600 244.050 595.050 ;
        RECT 257.400 594.600 258.600 596.400 ;
        RECT 265.950 595.950 268.050 596.400 ;
        RECT 415.950 595.950 418.050 599.400 ;
        RECT 424.950 598.800 427.050 600.900 ;
        RECT 430.950 600.600 433.050 601.050 ;
        RECT 436.950 600.600 439.050 601.050 ;
        RECT 445.950 600.600 448.050 600.900 ;
        RECT 430.950 599.400 448.050 600.600 ;
        RECT 430.950 598.950 433.050 599.400 ;
        RECT 436.950 598.950 439.050 599.400 ;
        RECT 445.950 598.800 448.050 599.400 ;
        RECT 472.950 599.400 477.600 601.050 ;
        RECT 503.400 600.900 504.600 607.950 ;
        RECT 505.950 605.100 508.050 607.200 ;
        RECT 526.950 606.600 529.050 607.050 ;
        RECT 532.950 606.600 535.050 607.500 ;
        RECT 526.950 605.400 535.050 606.600 ;
        RECT 541.950 606.600 544.050 607.500 ;
        RECT 553.950 606.600 556.050 607.050 ;
        RECT 541.950 605.400 556.050 606.600 ;
        RECT 506.400 601.050 507.600 605.100 ;
        RECT 526.950 604.950 529.050 605.400 ;
        RECT 542.400 601.050 543.600 605.400 ;
        RECT 553.950 604.950 556.050 605.400 ;
        RECT 574.950 606.750 577.050 607.200 ;
        RECT 580.950 606.750 583.050 607.200 ;
        RECT 574.950 605.550 583.050 606.750 ;
        RECT 574.950 605.100 577.050 605.550 ;
        RECT 580.950 605.100 583.050 605.550 ;
        RECT 592.950 604.950 595.050 607.050 ;
        RECT 610.950 604.950 613.050 607.050 ;
        RECT 619.950 604.950 622.050 607.050 ;
        RECT 628.950 606.750 631.050 607.200 ;
        RECT 637.950 606.750 640.050 607.200 ;
        RECT 628.950 605.550 640.050 606.750 ;
        RECT 628.950 605.100 631.050 605.550 ;
        RECT 637.950 605.100 640.050 605.550 ;
        RECT 472.950 598.950 477.000 599.400 ;
        RECT 502.950 598.800 505.050 600.900 ;
        RECT 506.400 599.400 511.050 601.050 ;
        RECT 507.000 598.950 511.050 599.400 ;
        RECT 514.950 600.150 517.050 600.600 ;
        RECT 523.950 600.150 526.050 600.600 ;
        RECT 514.950 598.950 526.050 600.150 ;
        RECT 542.400 599.400 547.050 601.050 ;
        RECT 543.000 598.950 547.050 599.400 ;
        RECT 559.950 600.600 562.050 600.900 ;
        RECT 574.950 600.600 577.050 601.050 ;
        RECT 559.950 599.400 577.050 600.600 ;
        RECT 514.950 598.500 517.050 598.950 ;
        RECT 523.950 598.500 526.050 598.950 ;
        RECT 559.950 598.800 562.050 599.400 ;
        RECT 574.950 598.950 577.050 599.400 ;
        RECT 577.950 597.600 580.050 598.050 ;
        RECT 593.400 597.600 594.600 604.950 ;
        RECT 604.950 600.600 607.050 600.900 ;
        RECT 611.400 600.600 612.600 604.950 ;
        RECT 620.400 601.050 621.600 604.950 ;
        RECT 604.950 599.400 612.600 600.600 ;
        RECT 604.950 598.800 607.050 599.400 ;
        RECT 619.950 598.950 622.050 601.050 ;
        RECT 631.950 600.600 634.050 600.900 ;
        RECT 641.400 600.600 642.600 608.400 ;
        RECT 766.950 608.400 775.050 609.600 ;
        RECT 766.950 607.950 769.050 608.400 ;
        RECT 772.950 607.950 775.050 608.400 ;
        RECT 805.950 609.600 808.050 610.050 ;
        RECT 829.950 609.600 832.050 610.050 ;
        RECT 805.950 608.400 832.050 609.600 ;
        RECT 805.950 607.950 808.050 608.400 ;
        RECT 829.950 607.950 832.050 608.400 ;
        RECT 893.400 608.400 912.600 609.600 ;
        RECT 658.950 604.950 661.050 607.050 ;
        RECT 688.950 606.600 691.050 607.200 ;
        RECT 703.950 606.600 706.050 607.200 ;
        RECT 688.950 605.400 706.050 606.600 ;
        RECT 688.950 605.100 691.050 605.400 ;
        RECT 703.950 605.100 706.050 605.400 ;
        RECT 712.950 606.600 715.050 607.050 ;
        RECT 724.950 606.600 727.050 607.200 ;
        RECT 733.950 606.600 736.050 607.050 ;
        RECT 787.950 606.600 790.050 607.200 ;
        RECT 841.950 606.600 844.050 607.050 ;
        RECT 712.950 605.400 727.050 606.600 ;
        RECT 712.950 604.950 715.050 605.400 ;
        RECT 724.950 605.100 727.050 605.400 ;
        RECT 728.400 605.400 736.050 606.600 ;
        RECT 659.400 601.050 660.600 604.950 ;
        RECT 728.400 603.600 729.600 605.400 ;
        RECT 733.950 604.950 736.050 605.400 ;
        RECT 785.400 605.400 790.050 606.600 ;
        RECT 809.400 606.000 844.050 606.600 ;
        RECT 725.400 602.400 729.600 603.600 ;
        RECT 631.950 599.400 642.600 600.600 ;
        RECT 646.950 600.450 649.050 600.900 ;
        RECT 652.950 600.450 655.050 600.900 ;
        RECT 631.950 598.800 634.050 599.400 ;
        RECT 646.950 599.250 655.050 600.450 ;
        RECT 646.950 598.800 649.050 599.250 ;
        RECT 652.950 598.800 655.050 599.250 ;
        RECT 658.950 598.950 661.050 601.050 ;
        RECT 685.950 600.600 688.050 600.900 ;
        RECT 691.950 600.600 694.050 601.050 ;
        RECT 685.950 599.400 694.050 600.600 ;
        RECT 685.950 598.800 688.050 599.400 ;
        RECT 691.950 598.950 694.050 599.400 ;
        RECT 706.950 600.450 709.050 600.900 ;
        RECT 712.950 600.450 715.050 600.900 ;
        RECT 706.950 599.250 715.050 600.450 ;
        RECT 706.950 598.800 709.050 599.250 ;
        RECT 712.950 598.800 715.050 599.250 ;
        RECT 725.400 598.050 726.600 602.400 ;
        RECT 785.400 601.050 786.600 605.400 ;
        RECT 787.950 605.100 790.050 605.400 ;
        RECT 808.950 605.400 844.050 606.000 ;
        RECT 808.950 601.800 811.050 605.400 ;
        RECT 841.950 604.950 844.050 605.400 ;
        RECT 859.950 604.950 862.050 607.050 ;
        RECT 868.950 606.600 871.050 607.200 ;
        RECT 886.950 606.600 889.050 607.050 ;
        RECT 893.400 606.600 894.600 608.400 ;
        RECT 911.400 607.050 912.600 608.400 ;
        RECT 919.950 607.950 922.050 610.050 ;
        RECT 868.950 605.400 873.600 606.600 ;
        RECT 868.950 605.100 871.050 605.400 ;
        RECT 860.400 601.050 861.600 604.950 ;
        RECT 872.400 601.050 873.600 605.400 ;
        RECT 886.950 605.400 894.600 606.600 ;
        RECT 895.950 606.600 900.000 607.050 ;
        RECT 886.950 604.950 889.050 605.400 ;
        RECT 895.950 604.950 900.600 606.600 ;
        RECT 763.950 600.450 766.050 600.900 ;
        RECT 769.950 600.450 772.050 600.900 ;
        RECT 763.950 599.250 772.050 600.450 ;
        RECT 763.950 598.800 766.050 599.250 ;
        RECT 769.950 598.800 772.050 599.250 ;
        RECT 784.950 598.950 787.050 601.050 ;
        RECT 859.950 598.950 862.050 601.050 ;
        RECT 871.950 598.950 874.050 601.050 ;
        RECT 880.950 600.600 883.050 601.050 ;
        RECT 887.400 600.600 888.600 604.950 ;
        RECT 880.950 599.400 888.600 600.600 ;
        RECT 899.400 600.600 900.600 604.950 ;
        RECT 901.950 603.600 904.050 607.050 ;
        RECT 910.950 604.950 913.050 607.050 ;
        RECT 901.950 603.000 909.600 603.600 ;
        RECT 902.400 602.400 909.600 603.000 ;
        RECT 908.400 600.900 909.600 602.400 ;
        RECT 899.400 600.000 906.600 600.600 ;
        RECT 899.400 599.400 907.050 600.000 ;
        RECT 880.950 598.950 883.050 599.400 ;
        RECT 577.950 596.400 594.600 597.600 ;
        RECT 598.950 597.600 601.050 598.050 ;
        RECT 613.950 597.600 616.050 598.050 ;
        RECT 598.950 596.400 616.050 597.600 ;
        RECT 577.950 595.950 580.050 596.400 ;
        RECT 598.950 595.950 601.050 596.400 ;
        RECT 613.950 595.950 616.050 596.400 ;
        RECT 694.950 597.600 697.050 598.050 ;
        RECT 700.950 597.600 703.050 598.050 ;
        RECT 694.950 596.400 703.050 597.600 ;
        RECT 694.950 595.950 697.050 596.400 ;
        RECT 700.950 595.950 703.050 596.400 ;
        RECT 724.950 595.950 727.050 598.050 ;
        RECT 904.950 595.950 907.050 599.400 ;
        RECT 907.950 598.800 910.050 600.900 ;
        RECT 920.400 600.600 921.600 607.950 ;
        RECT 920.400 599.400 924.600 600.600 ;
        RECT 241.950 593.400 258.600 594.600 ;
        RECT 268.950 594.600 271.050 595.050 ;
        RECT 274.950 594.600 277.050 595.050 ;
        RECT 268.950 593.400 277.050 594.600 ;
        RECT 241.950 592.950 244.050 593.400 ;
        RECT 268.950 592.950 271.050 593.400 ;
        RECT 274.950 592.950 277.050 593.400 ;
        RECT 295.950 594.600 298.050 595.050 ;
        RECT 313.950 594.600 316.050 595.050 ;
        RECT 295.950 593.400 316.050 594.600 ;
        RECT 295.950 592.950 298.050 593.400 ;
        RECT 313.950 592.950 316.050 593.400 ;
        RECT 319.950 594.600 322.050 595.050 ;
        RECT 430.950 594.600 433.050 595.050 ;
        RECT 319.950 593.400 433.050 594.600 ;
        RECT 319.950 592.950 322.050 593.400 ;
        RECT 430.950 592.950 433.050 593.400 ;
        RECT 493.950 594.600 496.050 595.050 ;
        RECT 511.950 594.600 514.050 595.050 ;
        RECT 544.950 594.600 547.050 595.050 ;
        RECT 682.950 594.600 685.050 594.900 ;
        RECT 493.950 593.400 685.050 594.600 ;
        RECT 493.950 592.950 496.050 593.400 ;
        RECT 511.950 592.950 514.050 593.400 ;
        RECT 544.950 592.950 547.050 593.400 ;
        RECT 682.950 592.800 685.050 593.400 ;
        RECT 688.950 594.600 691.050 595.050 ;
        RECT 727.950 594.600 730.050 595.050 ;
        RECT 688.950 593.400 730.050 594.600 ;
        RECT 688.950 592.950 691.050 593.400 ;
        RECT 727.950 592.950 730.050 593.400 ;
        RECT 766.950 594.600 769.050 595.050 ;
        RECT 790.950 594.600 793.050 595.050 ;
        RECT 766.950 593.400 793.050 594.600 ;
        RECT 766.950 592.950 769.050 593.400 ;
        RECT 790.950 592.950 793.050 593.400 ;
        RECT 865.950 594.600 868.050 595.050 ;
        RECT 880.950 594.600 883.050 595.050 ;
        RECT 865.950 593.400 883.050 594.600 ;
        RECT 865.950 592.950 868.050 593.400 ;
        RECT 880.950 592.950 883.050 593.400 ;
        RECT 889.950 594.600 892.050 595.050 ;
        RECT 919.950 594.600 922.050 595.050 ;
        RECT 889.950 593.400 922.050 594.600 ;
        RECT 889.950 592.950 892.050 593.400 ;
        RECT 919.950 592.950 922.050 593.400 ;
        RECT 1.950 591.600 4.050 592.050 ;
        RECT 61.950 591.600 64.050 592.050 ;
        RECT 1.950 590.400 64.050 591.600 ;
        RECT 1.950 589.950 4.050 590.400 ;
        RECT 61.950 589.950 64.050 590.400 ;
        RECT 73.950 591.600 76.050 592.050 ;
        RECT 103.950 591.600 106.050 592.050 ;
        RECT 73.950 590.400 106.050 591.600 ;
        RECT 73.950 589.950 76.050 590.400 ;
        RECT 103.950 589.950 106.050 590.400 ;
        RECT 121.950 591.600 124.050 592.050 ;
        RECT 130.950 591.600 133.050 592.050 ;
        RECT 121.950 590.400 133.050 591.600 ;
        RECT 121.950 589.950 124.050 590.400 ;
        RECT 130.950 589.950 133.050 590.400 ;
        RECT 148.950 591.600 151.050 592.050 ;
        RECT 178.950 591.600 181.050 592.050 ;
        RECT 148.950 590.400 181.050 591.600 ;
        RECT 148.950 589.950 151.050 590.400 ;
        RECT 178.950 589.950 181.050 590.400 ;
        RECT 184.950 591.600 187.050 592.050 ;
        RECT 211.950 591.600 214.050 592.050 ;
        RECT 184.950 590.400 214.050 591.600 ;
        RECT 184.950 589.950 187.050 590.400 ;
        RECT 211.950 589.950 214.050 590.400 ;
        RECT 238.950 591.600 241.050 592.050 ;
        RECT 265.950 591.600 268.050 592.050 ;
        RECT 238.950 590.400 268.050 591.600 ;
        RECT 238.950 589.950 241.050 590.400 ;
        RECT 265.950 589.950 268.050 590.400 ;
        RECT 277.950 591.600 280.050 592.050 ;
        RECT 304.950 591.600 307.050 592.050 ;
        RECT 523.950 591.600 526.050 592.050 ;
        RECT 277.950 590.400 307.050 591.600 ;
        RECT 515.400 591.000 526.050 591.600 ;
        RECT 277.950 589.950 280.050 590.400 ;
        RECT 304.950 589.950 307.050 590.400 ;
        RECT 514.950 590.400 526.050 591.000 ;
        RECT 16.950 588.600 19.050 589.050 ;
        RECT 49.950 588.600 52.050 589.050 ;
        RECT 16.950 587.400 52.050 588.600 ;
        RECT 16.950 586.950 19.050 587.400 ;
        RECT 49.950 586.950 52.050 587.400 ;
        RECT 100.950 588.600 103.050 589.050 ;
        RECT 127.950 588.600 130.050 589.050 ;
        RECT 262.950 588.600 265.050 589.050 ;
        RECT 100.950 587.400 130.050 588.600 ;
        RECT 100.950 586.950 103.050 587.400 ;
        RECT 127.950 586.950 130.050 587.400 ;
        RECT 134.400 587.400 265.050 588.600 ;
        RECT 22.950 585.600 25.050 586.050 ;
        RECT 40.950 585.600 43.050 586.050 ;
        RECT 112.950 585.600 115.050 586.050 ;
        RECT 134.400 585.600 135.600 587.400 ;
        RECT 262.950 586.950 265.050 587.400 ;
        RECT 334.950 588.600 337.050 589.050 ;
        RECT 493.950 588.600 496.050 589.050 ;
        RECT 508.950 588.600 511.050 589.050 ;
        RECT 334.950 587.400 399.600 588.600 ;
        RECT 334.950 586.950 337.050 587.400 ;
        RECT 398.400 586.050 399.600 587.400 ;
        RECT 493.950 587.400 511.050 588.600 ;
        RECT 493.950 586.950 496.050 587.400 ;
        RECT 508.950 586.950 511.050 587.400 ;
        RECT 514.950 586.950 517.050 590.400 ;
        RECT 523.950 589.950 526.050 590.400 ;
        RECT 574.950 591.600 577.050 592.050 ;
        RECT 661.950 591.600 664.050 592.050 ;
        RECT 574.950 590.400 664.050 591.600 ;
        RECT 574.950 589.950 577.050 590.400 ;
        RECT 661.950 589.950 664.050 590.400 ;
        RECT 697.950 591.600 700.050 592.050 ;
        RECT 718.950 591.600 721.050 592.050 ;
        RECT 697.950 590.400 721.050 591.600 ;
        RECT 697.950 589.950 700.050 590.400 ;
        RECT 718.950 589.950 721.050 590.400 ;
        RECT 730.950 591.600 733.050 592.050 ;
        RECT 763.950 591.600 766.050 592.050 ;
        RECT 730.950 590.400 766.050 591.600 ;
        RECT 730.950 589.950 733.050 590.400 ;
        RECT 763.950 589.950 766.050 590.400 ;
        RECT 923.400 589.050 924.600 599.400 ;
        RECT 526.950 588.600 529.050 589.050 ;
        RECT 583.950 588.600 586.050 589.050 ;
        RECT 526.950 587.400 586.050 588.600 ;
        RECT 526.950 586.950 529.050 587.400 ;
        RECT 583.950 586.950 586.050 587.400 ;
        RECT 589.950 588.600 592.050 589.050 ;
        RECT 631.950 588.600 634.050 589.050 ;
        RECT 589.950 587.400 634.050 588.600 ;
        RECT 589.950 586.950 592.050 587.400 ;
        RECT 631.950 586.950 634.050 587.400 ;
        RECT 736.950 588.600 739.050 589.050 ;
        RECT 751.950 588.600 754.050 589.050 ;
        RECT 736.950 587.400 754.050 588.600 ;
        RECT 736.950 586.950 739.050 587.400 ;
        RECT 751.950 586.950 754.050 587.400 ;
        RECT 781.950 588.600 784.050 589.050 ;
        RECT 787.950 588.600 790.050 589.050 ;
        RECT 781.950 587.400 790.050 588.600 ;
        RECT 781.950 586.950 784.050 587.400 ;
        RECT 787.950 586.950 790.050 587.400 ;
        RECT 907.950 588.600 910.050 589.050 ;
        RECT 913.950 588.600 916.050 589.050 ;
        RECT 907.950 587.400 916.050 588.600 ;
        RECT 907.950 586.950 910.050 587.400 ;
        RECT 913.950 586.950 916.050 587.400 ;
        RECT 919.950 587.400 924.600 589.050 ;
        RECT 919.950 586.950 924.000 587.400 ;
        RECT 22.950 584.400 135.600 585.600 ;
        RECT 154.950 585.600 157.050 586.050 ;
        RECT 166.950 585.600 169.050 586.050 ;
        RECT 154.950 584.400 169.050 585.600 ;
        RECT 22.950 583.950 25.050 584.400 ;
        RECT 40.950 583.950 43.050 584.400 ;
        RECT 112.950 583.950 115.050 584.400 ;
        RECT 154.950 583.950 157.050 584.400 ;
        RECT 166.950 583.950 169.050 584.400 ;
        RECT 175.950 585.600 178.050 586.050 ;
        RECT 190.950 585.600 193.050 586.050 ;
        RECT 175.950 584.400 193.050 585.600 ;
        RECT 175.950 583.950 178.050 584.400 ;
        RECT 190.950 583.950 193.050 584.400 ;
        RECT 238.950 585.600 241.050 586.050 ;
        RECT 244.950 585.600 247.050 586.050 ;
        RECT 253.950 585.600 256.050 586.050 ;
        RECT 238.950 584.400 256.050 585.600 ;
        RECT 238.950 583.950 241.050 584.400 ;
        RECT 244.950 583.950 247.050 584.400 ;
        RECT 253.950 583.950 256.050 584.400 ;
        RECT 379.950 585.600 382.050 586.050 ;
        RECT 391.950 585.600 394.050 586.050 ;
        RECT 379.950 584.400 394.050 585.600 ;
        RECT 379.950 583.950 382.050 584.400 ;
        RECT 391.950 583.950 394.050 584.400 ;
        RECT 397.950 585.600 400.050 586.050 ;
        RECT 439.950 585.600 442.050 586.050 ;
        RECT 397.950 584.400 442.050 585.600 ;
        RECT 397.950 583.950 400.050 584.400 ;
        RECT 439.950 583.950 442.050 584.400 ;
        RECT 466.950 585.600 469.050 586.050 ;
        RECT 478.950 585.600 481.050 586.050 ;
        RECT 466.950 584.400 481.050 585.600 ;
        RECT 466.950 583.950 469.050 584.400 ;
        RECT 478.950 583.950 481.050 584.400 ;
        RECT 511.950 585.600 514.050 586.050 ;
        RECT 517.950 585.600 520.050 586.050 ;
        RECT 511.950 584.400 520.050 585.600 ;
        RECT 511.950 583.950 514.050 584.400 ;
        RECT 517.950 583.950 520.050 584.400 ;
        RECT 541.950 585.600 544.050 586.050 ;
        RECT 550.950 585.600 553.050 586.050 ;
        RECT 541.950 584.400 553.050 585.600 ;
        RECT 541.950 583.950 544.050 584.400 ;
        RECT 550.950 583.950 553.050 584.400 ;
        RECT 625.950 585.600 628.050 586.050 ;
        RECT 631.950 585.600 634.050 585.900 ;
        RECT 625.950 584.400 634.050 585.600 ;
        RECT 625.950 583.950 628.050 584.400 ;
        RECT 631.950 583.800 634.050 584.400 ;
        RECT 664.950 585.600 667.050 586.050 ;
        RECT 737.400 585.600 738.600 586.950 ;
        RECT 664.950 584.400 738.600 585.600 ;
        RECT 763.950 585.600 766.050 586.050 ;
        RECT 790.950 585.600 793.050 586.050 ;
        RECT 763.950 584.400 793.050 585.600 ;
        RECT 664.950 583.950 667.050 584.400 ;
        RECT 763.950 583.950 766.050 584.400 ;
        RECT 790.950 583.950 793.050 584.400 ;
        RECT 55.950 582.600 58.050 583.050 ;
        RECT 76.950 582.600 79.050 583.050 ;
        RECT 124.950 582.600 127.050 583.050 ;
        RECT 55.950 581.400 127.050 582.600 ;
        RECT 55.950 580.950 58.050 581.400 ;
        RECT 76.950 580.950 79.050 581.400 ;
        RECT 124.950 580.950 127.050 581.400 ;
        RECT 214.950 582.600 217.050 583.050 ;
        RECT 229.950 582.600 232.050 583.050 ;
        RECT 214.950 581.400 232.050 582.600 ;
        RECT 214.950 580.950 217.050 581.400 ;
        RECT 229.950 580.950 232.050 581.400 ;
        RECT 262.950 582.600 265.050 583.050 ;
        RECT 283.950 582.600 286.050 583.050 ;
        RECT 262.950 581.400 286.050 582.600 ;
        RECT 262.950 580.950 265.050 581.400 ;
        RECT 283.950 580.950 286.050 581.400 ;
        RECT 325.950 582.600 328.050 583.050 ;
        RECT 340.950 582.600 343.050 583.050 ;
        RECT 325.950 581.400 343.050 582.600 ;
        RECT 325.950 580.950 328.050 581.400 ;
        RECT 340.950 580.950 343.050 581.400 ;
        RECT 412.950 582.600 415.050 583.050 ;
        RECT 436.950 582.600 439.050 583.050 ;
        RECT 412.950 581.400 439.050 582.600 ;
        RECT 412.950 580.950 415.050 581.400 ;
        RECT 436.950 580.950 439.050 581.400 ;
        RECT 481.950 582.600 484.050 583.050 ;
        RECT 520.950 582.600 523.050 583.050 ;
        RECT 481.950 581.400 523.050 582.600 ;
        RECT 481.950 580.950 484.050 581.400 ;
        RECT 520.950 580.950 523.050 581.400 ;
        RECT 691.950 582.600 694.050 583.050 ;
        RECT 733.950 582.600 736.050 583.050 ;
        RECT 691.950 581.400 736.050 582.600 ;
        RECT 691.950 580.950 694.050 581.400 ;
        RECT 733.950 580.950 736.050 581.400 ;
        RECT 760.950 582.600 763.050 583.050 ;
        RECT 793.950 582.600 796.050 583.050 ;
        RECT 760.950 581.400 796.050 582.600 ;
        RECT 760.950 580.950 763.050 581.400 ;
        RECT 793.950 580.950 796.050 581.400 ;
        RECT 844.950 582.600 847.050 583.050 ;
        RECT 868.950 582.600 871.050 583.050 ;
        RECT 844.950 581.400 871.050 582.600 ;
        RECT 844.950 580.950 847.050 581.400 ;
        RECT 868.950 580.950 871.050 581.400 ;
        RECT 901.950 582.600 904.050 583.050 ;
        RECT 910.950 582.600 913.050 583.050 ;
        RECT 901.950 581.400 913.050 582.600 ;
        RECT 901.950 580.950 904.050 581.400 ;
        RECT 910.950 580.950 913.050 581.400 ;
        RECT 133.950 579.600 136.050 580.050 ;
        RECT 172.950 579.600 175.050 580.050 ;
        RECT 133.950 578.400 175.050 579.600 ;
        RECT 133.950 577.950 136.050 578.400 ;
        RECT 172.950 577.950 175.050 578.400 ;
        RECT 190.950 579.600 193.050 580.050 ;
        RECT 226.950 579.600 229.050 580.050 ;
        RECT 190.950 578.400 229.050 579.600 ;
        RECT 190.950 577.950 193.050 578.400 ;
        RECT 226.950 577.950 229.050 578.400 ;
        RECT 244.950 579.600 247.050 580.050 ;
        RECT 253.950 579.600 256.050 580.050 ;
        RECT 244.950 578.400 256.050 579.600 ;
        RECT 244.950 577.950 247.050 578.400 ;
        RECT 253.950 577.950 256.050 578.400 ;
        RECT 259.950 579.600 262.050 580.050 ;
        RECT 277.950 579.600 280.050 580.050 ;
        RECT 259.950 578.400 280.050 579.600 ;
        RECT 259.950 577.950 262.050 578.400 ;
        RECT 277.950 577.950 280.050 578.400 ;
        RECT 286.950 579.600 289.050 580.050 ;
        RECT 301.950 579.600 304.050 580.050 ;
        RECT 286.950 578.400 304.050 579.600 ;
        RECT 286.950 577.950 289.050 578.400 ;
        RECT 301.950 577.950 304.050 578.400 ;
        RECT 382.950 579.600 385.050 580.050 ;
        RECT 391.950 579.600 394.050 579.900 ;
        RECT 382.950 578.400 394.050 579.600 ;
        RECT 382.950 577.950 385.050 578.400 ;
        RECT 391.950 577.800 394.050 578.400 ;
        RECT 403.950 579.600 406.050 580.050 ;
        RECT 418.950 579.600 421.050 580.050 ;
        RECT 454.950 579.600 457.050 580.050 ;
        RECT 403.950 578.400 457.050 579.600 ;
        RECT 403.950 577.950 406.050 578.400 ;
        RECT 418.950 577.950 421.050 578.400 ;
        RECT 454.950 577.950 457.050 578.400 ;
        RECT 460.950 579.600 463.050 580.050 ;
        RECT 469.950 579.600 472.050 580.050 ;
        RECT 460.950 578.400 472.050 579.600 ;
        RECT 460.950 577.950 463.050 578.400 ;
        RECT 469.950 577.950 472.050 578.400 ;
        RECT 478.950 579.600 481.050 580.050 ;
        RECT 580.950 579.600 583.050 580.050 ;
        RECT 610.950 579.600 613.050 580.050 ;
        RECT 478.950 578.400 531.600 579.600 ;
        RECT 478.950 577.950 481.050 578.400 ;
        RECT 7.950 576.600 10.050 577.050 ;
        RECT 37.950 576.600 40.050 577.050 ;
        RECT 61.950 576.600 64.050 577.050 ;
        RECT 7.950 575.400 64.050 576.600 ;
        RECT 7.950 574.950 10.050 575.400 ;
        RECT 37.950 574.950 40.050 575.400 ;
        RECT 61.950 574.950 64.050 575.400 ;
        RECT 88.950 576.600 91.050 577.050 ;
        RECT 94.950 576.600 97.050 577.050 ;
        RECT 121.950 576.600 124.050 577.050 ;
        RECT 88.950 575.400 124.050 576.600 ;
        RECT 88.950 574.950 91.050 575.400 ;
        RECT 94.950 574.950 97.050 575.400 ;
        RECT 121.950 574.950 124.050 575.400 ;
        RECT 256.950 574.950 259.050 577.050 ;
        RECT 331.950 576.600 334.050 577.050 ;
        RECT 337.950 576.600 340.050 577.050 ;
        RECT 331.950 575.400 340.050 576.600 ;
        RECT 331.950 574.950 334.050 575.400 ;
        RECT 337.950 574.950 340.050 575.400 ;
        RECT 370.950 576.600 373.050 577.050 ;
        RECT 376.950 576.600 379.050 577.050 ;
        RECT 370.950 575.400 379.050 576.600 ;
        RECT 370.950 574.950 373.050 575.400 ;
        RECT 376.950 574.950 379.050 575.400 ;
        RECT 406.950 576.600 409.050 577.050 ;
        RECT 418.950 576.600 421.050 576.900 ;
        RECT 433.950 576.600 436.050 577.050 ;
        RECT 406.950 575.400 436.050 576.600 ;
        RECT 406.950 574.950 409.050 575.400 ;
        RECT 28.950 571.950 31.050 574.050 ;
        RECT 43.950 573.600 46.050 574.050 ;
        RECT 52.950 573.600 55.050 574.050 ;
        RECT 43.950 572.400 55.050 573.600 ;
        RECT 43.950 571.950 46.050 572.400 ;
        RECT 52.950 571.950 55.050 572.400 ;
        RECT 85.950 573.600 88.050 574.200 ;
        RECT 85.950 572.400 90.600 573.600 ;
        RECT 85.950 572.100 88.050 572.400 ;
        RECT 7.950 567.450 10.050 567.900 ;
        RECT 13.950 567.450 16.050 567.900 ;
        RECT 7.950 566.250 16.050 567.450 ;
        RECT 29.400 567.600 30.600 571.950 ;
        RECT 89.400 568.050 90.600 572.400 ;
        RECT 97.950 571.950 100.050 574.050 ;
        RECT 108.000 573.600 112.050 574.050 ;
        RECT 136.950 573.600 139.050 574.050 ;
        RECT 107.400 571.950 112.050 573.600 ;
        RECT 128.400 572.400 139.050 573.600 ;
        RECT 37.950 567.600 40.050 567.900 ;
        RECT 29.400 566.400 40.050 567.600 ;
        RECT 7.950 565.800 10.050 566.250 ;
        RECT 13.950 565.800 16.050 566.250 ;
        RECT 37.950 565.800 40.050 566.400 ;
        RECT 58.950 567.600 61.050 567.900 ;
        RECT 76.950 567.600 79.050 567.900 ;
        RECT 58.950 567.450 79.050 567.600 ;
        RECT 82.950 567.450 85.050 567.900 ;
        RECT 58.950 566.400 85.050 567.450 ;
        RECT 89.400 566.400 94.050 568.050 ;
        RECT 98.400 567.600 99.600 571.950 ;
        RECT 107.400 567.900 108.600 571.950 ;
        RECT 128.400 568.050 129.600 572.400 ;
        RECT 136.950 571.950 139.050 572.400 ;
        RECT 142.950 573.600 145.050 574.200 ;
        RECT 163.950 573.600 166.050 574.200 ;
        RECT 142.950 572.400 166.050 573.600 ;
        RECT 142.950 572.100 145.050 572.400 ;
        RECT 163.950 572.100 166.050 572.400 ;
        RECT 169.950 573.600 172.050 574.200 ;
        RECT 169.950 572.400 195.600 573.600 ;
        RECT 169.950 572.100 172.050 572.400 ;
        RECT 100.950 567.600 103.050 567.900 ;
        RECT 98.400 566.400 103.050 567.600 ;
        RECT 58.950 565.800 61.050 566.400 ;
        RECT 76.950 566.250 85.050 566.400 ;
        RECT 76.950 565.800 79.050 566.250 ;
        RECT 82.950 565.800 85.050 566.250 ;
        RECT 90.000 565.950 94.050 566.400 ;
        RECT 100.950 565.800 103.050 566.400 ;
        RECT 106.950 565.800 109.050 567.900 ;
        RECT 112.950 567.450 115.050 567.900 ;
        RECT 118.950 567.450 121.050 567.900 ;
        RECT 112.950 566.250 121.050 567.450 ;
        RECT 112.950 565.800 115.050 566.250 ;
        RECT 118.950 565.800 121.050 566.250 ;
        RECT 127.950 565.950 130.050 568.050 ;
        RECT 133.950 567.450 136.050 567.900 ;
        RECT 139.950 567.600 142.050 567.900 ;
        RECT 157.950 567.600 160.050 568.050 ;
        RECT 194.400 567.900 195.600 572.400 ;
        RECT 196.950 572.100 199.050 574.200 ;
        RECT 223.950 573.600 226.050 573.900 ;
        RECT 232.950 573.600 235.050 574.050 ;
        RECT 244.950 573.600 247.050 574.050 ;
        RECT 223.950 572.400 235.050 573.600 ;
        RECT 197.400 568.050 198.600 572.100 ;
        RECT 223.950 571.800 226.050 572.400 ;
        RECT 232.950 571.950 235.050 572.400 ;
        RECT 236.400 572.400 247.050 573.600 ;
        RECT 202.950 570.600 205.050 570.900 ;
        RECT 236.400 570.600 237.600 572.400 ;
        RECT 244.950 571.950 247.050 572.400 ;
        RECT 250.950 573.600 255.000 574.050 ;
        RECT 250.950 571.950 255.600 573.600 ;
        RECT 202.950 569.400 237.600 570.600 ;
        RECT 202.950 568.800 205.050 569.400 ;
        RECT 139.950 567.450 160.050 567.600 ;
        RECT 133.950 566.400 160.050 567.450 ;
        RECT 133.950 566.250 142.050 566.400 ;
        RECT 133.950 565.800 136.050 566.250 ;
        RECT 139.950 565.800 142.050 566.250 ;
        RECT 157.950 565.950 160.050 566.400 ;
        RECT 181.950 567.450 184.050 567.900 ;
        RECT 187.950 567.450 190.050 567.900 ;
        RECT 181.950 566.250 190.050 567.450 ;
        RECT 181.950 565.800 184.050 566.250 ;
        RECT 187.950 565.800 190.050 566.250 ;
        RECT 193.950 565.800 196.050 567.900 ;
        RECT 197.400 566.400 202.050 568.050 ;
        RECT 198.000 565.950 202.050 566.400 ;
        RECT 214.950 567.450 217.050 567.900 ;
        RECT 226.950 567.450 229.050 567.900 ;
        RECT 214.950 566.250 229.050 567.450 ;
        RECT 214.950 565.800 217.050 566.250 ;
        RECT 226.950 565.800 229.050 566.250 ;
        RECT 235.950 567.450 238.050 567.900 ;
        RECT 250.950 567.450 253.050 567.900 ;
        RECT 235.950 566.250 253.050 567.450 ;
        RECT 235.950 565.800 238.050 566.250 ;
        RECT 250.950 565.800 253.050 566.250 ;
        RECT 55.950 564.600 58.050 565.050 ;
        RECT 106.950 564.600 109.050 565.050 ;
        RECT 55.950 563.400 109.050 564.600 ;
        RECT 55.950 562.950 58.050 563.400 ;
        RECT 106.950 562.950 109.050 563.400 ;
        RECT 166.950 564.600 169.050 565.050 ;
        RECT 175.950 564.600 178.050 565.050 ;
        RECT 254.400 564.750 255.600 571.950 ;
        RECT 257.400 570.600 258.600 574.950 ;
        RECT 418.950 574.800 421.050 575.400 ;
        RECT 433.950 574.950 436.050 575.400 ;
        RECT 448.950 576.600 451.050 577.050 ;
        RECT 457.950 576.600 460.050 577.050 ;
        RECT 448.950 575.400 460.050 576.600 ;
        RECT 448.950 574.950 451.050 575.400 ;
        RECT 457.950 574.950 460.050 575.400 ;
        RECT 496.950 576.600 499.050 577.050 ;
        RECT 523.950 576.600 526.050 577.050 ;
        RECT 496.950 575.400 526.050 576.600 ;
        RECT 496.950 574.950 499.050 575.400 ;
        RECT 523.950 574.950 526.050 575.400 ;
        RECT 265.950 570.600 268.050 574.050 ;
        RECT 283.950 571.950 286.050 574.050 ;
        RECT 289.950 573.750 292.050 573.900 ;
        RECT 295.950 573.750 298.050 574.200 ;
        RECT 289.950 573.600 298.050 573.750 ;
        RECT 328.950 573.600 331.050 574.050 ;
        RECT 289.950 572.550 331.050 573.600 ;
        RECT 257.400 569.400 261.600 570.600 ;
        RECT 265.950 570.000 270.600 570.600 ;
        RECT 266.400 569.400 270.600 570.000 ;
        RECT 256.950 565.800 259.050 567.900 ;
        RECT 260.400 567.600 261.600 569.400 ;
        RECT 265.950 567.600 268.050 568.050 ;
        RECT 260.400 566.400 268.050 567.600 ;
        RECT 269.400 567.600 270.600 569.400 ;
        RECT 274.950 567.600 277.050 567.900 ;
        RECT 269.400 566.400 277.050 567.600 ;
        RECT 284.400 567.600 285.600 571.950 ;
        RECT 289.950 571.800 292.050 572.550 ;
        RECT 295.950 572.400 331.050 572.550 ;
        RECT 295.950 572.100 298.050 572.400 ;
        RECT 328.950 571.950 331.050 572.400 ;
        RECT 334.950 570.600 337.050 574.050 ;
        RECT 349.800 571.950 351.900 574.050 ;
        RECT 352.950 573.600 355.050 574.200 ;
        RECT 352.950 572.400 366.600 573.600 ;
        RECT 352.950 572.100 355.050 572.400 ;
        RECT 332.400 570.000 337.050 570.600 ;
        RECT 332.400 569.400 336.600 570.000 ;
        RECT 332.400 567.900 333.600 569.400 ;
        RECT 350.250 568.050 351.450 571.950 ;
        RECT 298.950 567.600 301.050 567.900 ;
        RECT 284.400 567.450 301.050 567.600 ;
        RECT 328.800 567.450 330.900 567.900 ;
        RECT 284.400 566.400 330.900 567.450 ;
        RECT 265.950 565.950 268.050 566.400 ;
        RECT 274.950 565.800 277.050 566.400 ;
        RECT 298.950 566.250 330.900 566.400 ;
        RECT 298.950 565.800 301.050 566.250 ;
        RECT 328.800 565.800 330.900 566.250 ;
        RECT 331.950 565.800 334.050 567.900 ;
        RECT 340.950 567.600 343.050 568.050 ;
        RECT 346.800 567.600 348.900 567.900 ;
        RECT 340.950 566.400 348.900 567.600 ;
        RECT 340.950 565.950 343.050 566.400 ;
        RECT 346.800 565.800 348.900 566.400 ;
        RECT 349.950 565.950 352.050 568.050 ;
        RECT 166.950 563.400 178.050 564.600 ;
        RECT 166.950 562.950 169.050 563.400 ;
        RECT 175.950 562.950 178.050 563.400 ;
        RECT 253.950 562.650 256.050 564.750 ;
        RECT 257.400 564.600 258.600 565.800 ;
        RECT 365.400 565.050 366.600 572.400 ;
        RECT 367.950 571.950 370.050 574.050 ;
        RECT 388.950 573.600 391.050 574.200 ;
        RECT 394.950 573.600 397.050 574.050 ;
        RECT 388.950 572.400 397.050 573.600 ;
        RECT 388.950 572.100 391.050 572.400 ;
        RECT 394.950 571.950 397.050 572.400 ;
        RECT 403.950 571.950 406.050 574.050 ;
        RECT 427.950 572.100 430.050 574.200 ;
        RECT 442.950 573.600 445.050 574.050 ;
        RECT 463.950 573.600 466.050 574.050 ;
        RECT 442.950 572.400 466.050 573.600 ;
        RECT 368.400 567.600 369.600 571.950 ;
        RECT 404.400 568.050 405.600 571.950 ;
        RECT 373.950 567.600 376.050 568.050 ;
        RECT 368.400 566.400 376.050 567.600 ;
        RECT 373.950 565.950 376.050 566.400 ;
        RECT 403.950 565.950 406.050 568.050 ;
        RECT 418.950 567.450 421.050 568.050 ;
        RECT 424.950 567.450 427.050 567.900 ;
        RECT 418.950 566.250 427.050 567.450 ;
        RECT 418.950 565.950 421.050 566.250 ;
        RECT 424.950 565.800 427.050 566.250 ;
        RECT 428.400 565.050 429.600 572.100 ;
        RECT 442.950 571.950 445.050 572.400 ;
        RECT 463.950 571.950 466.050 572.400 ;
        RECT 481.950 570.600 484.050 574.050 ;
        RECT 514.950 573.600 517.050 574.050 ;
        RECT 437.400 570.000 484.050 570.600 ;
        RECT 506.400 572.400 517.050 573.600 ;
        RECT 437.400 569.400 483.600 570.000 ;
        RECT 437.400 565.050 438.600 569.400 ;
        RECT 506.400 568.050 507.600 572.400 ;
        RECT 514.950 571.950 517.050 572.400 ;
        RECT 526.950 573.600 529.050 574.200 ;
        RECT 530.400 573.600 531.600 578.400 ;
        RECT 580.950 578.400 613.050 579.600 ;
        RECT 580.950 577.950 583.050 578.400 ;
        RECT 610.950 577.950 613.050 578.400 ;
        RECT 751.950 579.600 754.050 580.050 ;
        RECT 784.950 579.600 787.050 580.050 ;
        RECT 751.950 578.400 787.050 579.600 ;
        RECT 751.950 577.950 754.050 578.400 ;
        RECT 784.950 577.950 787.050 578.400 ;
        RECT 811.950 579.600 814.050 580.050 ;
        RECT 820.950 579.600 823.050 580.050 ;
        RECT 811.950 578.400 823.050 579.600 ;
        RECT 811.950 577.950 814.050 578.400 ;
        RECT 820.950 577.950 823.050 578.400 ;
        RECT 829.950 579.600 832.050 580.050 ;
        RECT 838.950 579.600 841.050 580.050 ;
        RECT 829.950 578.400 841.050 579.600 ;
        RECT 829.950 577.950 832.050 578.400 ;
        RECT 838.950 577.950 841.050 578.400 ;
        RECT 865.950 579.600 868.050 580.050 ;
        RECT 874.950 579.600 877.050 580.050 ;
        RECT 865.950 578.400 877.050 579.600 ;
        RECT 865.950 577.950 868.050 578.400 ;
        RECT 874.950 577.950 877.050 578.400 ;
        RECT 883.950 579.600 886.050 580.050 ;
        RECT 889.950 579.600 892.050 580.050 ;
        RECT 883.950 578.400 892.050 579.600 ;
        RECT 883.950 577.950 886.050 578.400 ;
        RECT 889.950 577.950 892.050 578.400 ;
        RECT 547.950 576.600 550.050 577.050 ;
        RECT 559.950 576.600 562.050 577.050 ;
        RECT 547.950 575.400 562.050 576.600 ;
        RECT 547.950 574.950 550.050 575.400 ;
        RECT 559.950 574.950 562.050 575.400 ;
        RECT 526.950 572.400 531.600 573.600 ;
        RECT 550.950 573.600 553.050 574.200 ;
        RECT 562.800 573.600 564.900 574.050 ;
        RECT 550.950 572.400 564.900 573.600 ;
        RECT 526.950 572.100 529.050 572.400 ;
        RECT 550.950 572.100 553.050 572.400 ;
        RECT 562.800 571.950 564.900 572.400 ;
        RECT 571.950 571.950 574.050 574.050 ;
        RECT 577.950 571.950 580.050 574.050 ;
        RECT 589.950 573.600 592.050 574.200 ;
        RECT 584.400 572.400 592.050 573.600 ;
        RECT 601.950 574.050 604.050 574.500 ;
        RECT 616.950 574.050 619.050 577.050 ;
        RECT 790.950 576.600 793.050 577.050 ;
        RECT 823.950 576.600 826.050 577.050 ;
        RECT 847.950 576.600 850.050 577.050 ;
        RECT 790.950 575.400 826.050 576.600 ;
        RECT 790.950 574.950 793.050 575.400 ;
        RECT 823.950 574.950 826.050 575.400 ;
        RECT 842.400 575.400 850.050 576.600 ;
        RECT 622.950 574.050 625.050 574.500 ;
        RECT 601.950 572.850 625.050 574.050 ;
        RECT 601.950 572.400 604.050 572.850 ;
        RECT 617.400 572.400 618.600 572.850 ;
        RECT 622.950 572.400 625.050 572.850 ;
        RECT 439.950 567.450 442.050 567.900 ;
        RECT 445.950 567.450 448.050 567.900 ;
        RECT 439.950 566.250 448.050 567.450 ;
        RECT 439.950 565.800 442.050 566.250 ;
        RECT 445.950 565.800 448.050 566.250 ;
        RECT 451.950 567.600 454.050 567.900 ;
        RECT 475.950 567.600 478.050 567.900 ;
        RECT 451.950 566.400 478.050 567.600 ;
        RECT 451.950 565.800 454.050 566.400 ;
        RECT 475.950 565.800 478.050 566.400 ;
        RECT 496.950 567.600 499.050 568.050 ;
        RECT 496.950 566.400 504.900 567.600 ;
        RECT 496.950 565.950 499.050 566.400 ;
        RECT 502.800 565.500 504.900 566.400 ;
        RECT 505.950 565.950 508.050 568.050 ;
        RECT 568.950 567.600 571.050 567.900 ;
        RECT 572.400 567.600 573.600 571.950 ;
        RECT 578.400 568.050 579.600 571.950 ;
        RECT 584.400 568.050 585.600 572.400 ;
        RECT 589.950 572.100 592.050 572.400 ;
        RECT 511.950 567.150 514.050 567.600 ;
        RECT 517.950 567.150 520.050 567.600 ;
        RECT 511.950 565.950 520.050 567.150 ;
        RECT 511.950 565.500 514.050 565.950 ;
        RECT 517.950 565.500 520.050 565.950 ;
        RECT 568.950 566.400 573.600 567.600 ;
        RECT 568.950 565.800 571.050 566.400 ;
        RECT 577.950 565.950 580.050 568.050 ;
        RECT 583.950 565.950 586.050 568.050 ;
        RECT 592.950 567.600 595.050 567.900 ;
        RECT 598.950 567.600 601.050 571.050 ;
        RECT 637.950 570.600 640.050 574.050 ;
        RECT 661.950 573.750 664.050 574.200 ;
        RECT 673.950 573.750 676.050 574.200 ;
        RECT 661.950 572.550 676.050 573.750 ;
        RECT 661.950 572.100 664.050 572.550 ;
        RECT 673.950 572.100 676.050 572.550 ;
        RECT 682.950 571.950 685.050 574.050 ;
        RECT 763.950 572.100 766.050 574.200 ;
        RECT 805.950 573.600 808.050 574.050 ;
        RECT 817.950 573.750 820.050 574.200 ;
        RECT 826.950 573.750 829.050 574.200 ;
        RECT 805.950 572.400 816.600 573.600 ;
        RECT 592.950 567.000 601.050 567.600 ;
        RECT 629.400 570.000 640.050 570.600 ;
        RECT 629.400 569.400 639.600 570.000 ;
        RECT 592.950 566.400 600.600 567.000 ;
        RECT 592.950 565.800 595.050 566.400 ;
        RECT 629.400 565.050 630.600 569.400 ;
        RECT 631.950 567.150 634.050 568.050 ;
        RECT 683.400 567.600 684.600 571.950 ;
        RECT 764.400 570.600 765.600 572.100 ;
        RECT 805.950 571.950 808.050 572.400 ;
        RECT 755.400 569.400 765.600 570.600 ;
        RECT 815.400 570.600 816.600 572.400 ;
        RECT 817.950 572.550 829.050 573.750 ;
        RECT 817.950 572.100 820.050 572.550 ;
        RECT 826.950 572.100 829.050 572.550 ;
        RECT 815.400 570.000 837.600 570.600 ;
        RECT 815.400 569.400 838.050 570.000 ;
        RECT 685.950 567.600 688.050 567.900 ;
        RECT 640.950 567.150 643.050 567.600 ;
        RECT 631.950 565.950 643.050 567.150 ;
        RECT 683.400 566.400 688.050 567.600 ;
        RECT 640.950 565.500 643.050 565.950 ;
        RECT 685.950 565.800 688.050 566.400 ;
        RECT 739.950 567.600 742.050 567.900 ;
        RECT 755.400 567.600 756.600 569.400 ;
        RECT 739.950 566.400 756.600 567.600 ;
        RECT 757.950 567.600 760.050 568.050 ;
        RECT 787.950 567.600 790.050 568.050 ;
        RECT 757.950 566.400 790.050 567.600 ;
        RECT 739.950 565.800 742.050 566.400 ;
        RECT 757.950 565.950 760.050 566.400 ;
        RECT 787.950 565.950 790.050 566.400 ;
        RECT 835.950 565.950 838.050 569.400 ;
        RECT 842.400 567.900 843.600 575.400 ;
        RECT 847.950 574.950 850.050 575.400 ;
        RECT 904.950 576.600 907.050 577.050 ;
        RECT 913.950 576.600 916.050 577.050 ;
        RECT 904.950 575.400 916.050 576.600 ;
        RECT 904.950 574.950 907.050 575.400 ;
        RECT 913.950 574.950 916.050 575.400 ;
        RECT 859.950 573.600 862.050 574.050 ;
        RECT 883.950 573.600 886.050 574.200 ;
        RECT 859.950 572.400 867.600 573.600 ;
        RECT 859.950 571.950 862.050 572.400 ;
        RECT 841.950 565.800 844.050 567.900 ;
        RECT 866.400 565.050 867.600 572.400 ;
        RECT 869.400 572.400 886.050 573.600 ;
        RECT 869.400 567.900 870.600 572.400 ;
        RECT 883.950 572.100 886.050 572.400 ;
        RECT 892.950 573.600 895.050 574.050 ;
        RECT 898.950 573.600 901.050 574.050 ;
        RECT 892.950 572.400 901.050 573.600 ;
        RECT 892.950 571.950 895.050 572.400 ;
        RECT 898.950 571.950 901.050 572.400 ;
        RECT 907.950 571.950 910.050 574.050 ;
        RECT 908.400 568.050 909.600 571.950 ;
        RECT 868.950 565.800 871.050 567.900 ;
        RECT 907.950 565.950 910.050 568.050 ;
        RECT 286.950 564.600 289.050 565.050 ;
        RECT 257.400 563.400 289.050 564.600 ;
        RECT 286.950 562.950 289.050 563.400 ;
        RECT 304.950 564.600 307.050 565.050 ;
        RECT 313.950 564.600 316.050 565.050 ;
        RECT 322.950 564.600 325.050 565.050 ;
        RECT 304.950 563.400 325.050 564.600 ;
        RECT 304.950 562.950 307.050 563.400 ;
        RECT 313.950 562.950 316.050 563.400 ;
        RECT 322.950 562.950 325.050 563.400 ;
        RECT 331.950 564.600 334.050 564.750 ;
        RECT 355.950 564.600 358.050 565.050 ;
        RECT 331.950 563.400 358.050 564.600 ;
        RECT 365.400 563.400 370.050 565.050 ;
        RECT 331.950 562.650 334.050 563.400 ;
        RECT 355.950 562.950 358.050 563.400 ;
        RECT 366.000 562.950 370.050 563.400 ;
        RECT 382.950 564.600 385.050 565.050 ;
        RECT 397.950 564.600 400.050 565.050 ;
        RECT 382.950 563.400 400.050 564.600 ;
        RECT 382.950 562.950 385.050 563.400 ;
        RECT 397.950 562.950 400.050 563.400 ;
        RECT 427.950 562.950 430.050 565.050 ;
        RECT 433.950 563.400 438.600 565.050 ;
        RECT 463.950 564.600 466.050 565.050 ;
        RECT 481.950 564.600 484.050 565.050 ;
        RECT 463.950 563.400 484.050 564.600 ;
        RECT 433.950 562.950 438.000 563.400 ;
        RECT 463.950 562.950 466.050 563.400 ;
        RECT 481.950 562.950 484.050 563.400 ;
        RECT 520.950 564.600 523.050 565.050 ;
        RECT 547.950 564.600 550.050 565.050 ;
        RECT 520.950 563.400 550.050 564.600 ;
        RECT 629.400 564.900 633.000 565.050 ;
        RECT 629.400 563.400 634.050 564.900 ;
        RECT 520.950 562.950 523.050 563.400 ;
        RECT 547.950 562.950 550.050 563.400 ;
        RECT 630.000 562.950 634.050 563.400 ;
        RECT 658.950 564.600 661.050 565.050 ;
        RECT 667.950 564.600 670.050 565.050 ;
        RECT 658.950 563.400 670.050 564.600 ;
        RECT 658.950 562.950 661.050 563.400 ;
        RECT 667.950 562.950 670.050 563.400 ;
        RECT 739.950 564.600 742.050 564.750 ;
        RECT 796.950 564.600 799.050 565.050 ;
        RECT 739.950 563.400 799.050 564.600 ;
        RECT 631.950 562.800 634.050 562.950 ;
        RECT 739.950 562.650 742.050 563.400 ;
        RECT 796.950 562.950 799.050 563.400 ;
        RECT 865.950 562.950 868.050 565.050 ;
        RECT 25.950 561.600 28.050 562.050 ;
        RECT 46.950 561.600 49.050 562.050 ;
        RECT 124.950 561.600 127.050 562.050 ;
        RECT 202.950 561.600 205.050 562.050 ;
        RECT 25.950 560.400 205.050 561.600 ;
        RECT 25.950 559.950 28.050 560.400 ;
        RECT 46.950 559.950 49.050 560.400 ;
        RECT 124.950 559.950 127.050 560.400 ;
        RECT 202.950 559.950 205.050 560.400 ;
        RECT 208.950 561.600 211.050 562.050 ;
        RECT 229.950 561.600 232.050 562.050 ;
        RECT 208.950 560.400 232.050 561.600 ;
        RECT 208.950 559.950 211.050 560.400 ;
        RECT 229.950 559.950 232.050 560.400 ;
        RECT 250.950 561.600 253.050 562.050 ;
        RECT 262.950 561.600 265.050 561.900 ;
        RECT 250.950 560.400 265.050 561.600 ;
        RECT 250.950 559.950 253.050 560.400 ;
        RECT 262.950 559.800 265.050 560.400 ;
        RECT 268.950 561.600 271.050 562.050 ;
        RECT 274.950 561.600 277.050 562.050 ;
        RECT 268.950 560.400 277.050 561.600 ;
        RECT 268.950 559.950 271.050 560.400 ;
        RECT 274.950 559.950 277.050 560.400 ;
        RECT 343.950 561.600 346.050 562.050 ;
        RECT 349.950 561.600 352.050 562.050 ;
        RECT 343.950 560.400 352.050 561.600 ;
        RECT 343.950 559.950 346.050 560.400 ;
        RECT 349.950 559.950 352.050 560.400 ;
        RECT 358.950 561.600 361.050 562.050 ;
        RECT 385.950 561.600 388.050 562.050 ;
        RECT 358.950 560.400 388.050 561.600 ;
        RECT 358.950 559.950 361.050 560.400 ;
        RECT 385.950 559.950 388.050 560.400 ;
        RECT 475.950 561.600 478.050 562.050 ;
        RECT 496.950 561.600 499.050 562.050 ;
        RECT 475.950 560.400 499.050 561.600 ;
        RECT 475.950 559.950 478.050 560.400 ;
        RECT 496.950 559.950 499.050 560.400 ;
        RECT 535.950 561.600 538.050 562.050 ;
        RECT 562.950 561.600 565.050 562.050 ;
        RECT 535.950 560.400 565.050 561.600 ;
        RECT 535.950 559.950 538.050 560.400 ;
        RECT 562.950 559.950 565.050 560.400 ;
        RECT 673.950 561.600 676.050 562.050 ;
        RECT 697.950 561.600 700.050 562.050 ;
        RECT 673.950 560.400 700.050 561.600 ;
        RECT 673.950 559.950 676.050 560.400 ;
        RECT 697.950 559.950 700.050 560.400 ;
        RECT 751.950 561.600 754.050 562.050 ;
        RECT 769.950 561.600 772.050 562.050 ;
        RECT 751.950 560.400 772.050 561.600 ;
        RECT 751.950 559.950 754.050 560.400 ;
        RECT 769.950 559.950 772.050 560.400 ;
        RECT 811.950 561.600 814.050 562.050 ;
        RECT 826.950 561.600 829.050 562.050 ;
        RECT 847.950 561.600 850.050 562.050 ;
        RECT 811.950 560.400 850.050 561.600 ;
        RECT 811.950 559.950 814.050 560.400 ;
        RECT 826.950 559.950 829.050 560.400 ;
        RECT 847.950 559.950 850.050 560.400 ;
        RECT 877.950 561.600 880.050 562.050 ;
        RECT 886.950 561.600 889.050 562.050 ;
        RECT 877.950 560.400 889.050 561.600 ;
        RECT 877.950 559.950 880.050 560.400 ;
        RECT 886.950 559.950 889.050 560.400 ;
        RECT 88.950 558.600 91.050 559.050 ;
        RECT 100.950 558.600 103.050 559.050 ;
        RECT 133.950 558.600 136.050 559.050 ;
        RECT 88.950 557.400 136.050 558.600 ;
        RECT 88.950 556.950 91.050 557.400 ;
        RECT 100.950 556.950 103.050 557.400 ;
        RECT 133.950 556.950 136.050 557.400 ;
        RECT 154.950 558.600 157.050 559.050 ;
        RECT 172.950 558.600 175.050 559.050 ;
        RECT 154.950 557.400 175.050 558.600 ;
        RECT 154.950 556.950 157.050 557.400 ;
        RECT 172.950 556.950 175.050 557.400 ;
        RECT 265.950 558.600 268.050 559.050 ;
        RECT 313.800 558.600 315.900 559.050 ;
        RECT 265.950 557.400 315.900 558.600 ;
        RECT 265.950 556.950 268.050 557.400 ;
        RECT 313.800 556.950 315.900 557.400 ;
        RECT 316.950 558.600 319.050 559.050 ;
        RECT 346.950 558.600 349.050 559.050 ;
        RECT 316.950 557.400 349.050 558.600 ;
        RECT 316.950 556.950 319.050 557.400 ;
        RECT 346.950 556.950 349.050 557.400 ;
        RECT 613.950 558.600 616.050 559.050 ;
        RECT 634.950 558.600 637.050 559.050 ;
        RECT 613.950 557.400 637.050 558.600 ;
        RECT 613.950 556.950 616.050 557.400 ;
        RECT 634.950 556.950 637.050 557.400 ;
        RECT 661.950 558.600 664.050 559.050 ;
        RECT 667.950 558.600 670.050 559.050 ;
        RECT 661.950 557.400 670.050 558.600 ;
        RECT 661.950 556.950 664.050 557.400 ;
        RECT 667.950 556.950 670.050 557.400 ;
        RECT 682.950 558.600 685.050 559.050 ;
        RECT 694.950 558.600 697.050 559.050 ;
        RECT 682.950 557.400 697.050 558.600 ;
        RECT 682.950 556.950 685.050 557.400 ;
        RECT 694.950 556.950 697.050 557.400 ;
        RECT 772.950 558.600 775.050 559.050 ;
        RECT 820.950 558.600 823.050 559.050 ;
        RECT 772.950 557.400 823.050 558.600 ;
        RECT 772.950 556.950 775.050 557.400 ;
        RECT 820.950 556.950 823.050 557.400 ;
        RECT 241.950 555.600 244.050 556.050 ;
        RECT 268.950 555.600 271.050 556.050 ;
        RECT 241.950 554.400 271.050 555.600 ;
        RECT 241.950 553.950 244.050 554.400 ;
        RECT 268.950 553.950 271.050 554.400 ;
        RECT 274.950 555.600 277.050 556.050 ;
        RECT 292.950 555.600 295.050 556.050 ;
        RECT 319.950 555.600 322.050 556.050 ;
        RECT 349.950 555.600 352.050 556.050 ;
        RECT 274.950 554.400 303.600 555.600 ;
        RECT 274.950 553.950 277.050 554.400 ;
        RECT 292.950 553.950 295.050 554.400 ;
        RECT 148.950 552.600 151.050 553.050 ;
        RECT 229.950 552.600 232.050 553.050 ;
        RECT 271.950 552.600 274.050 553.050 ;
        RECT 148.950 551.400 274.050 552.600 ;
        RECT 302.400 552.600 303.600 554.400 ;
        RECT 319.950 554.400 352.050 555.600 ;
        RECT 319.950 553.950 322.050 554.400 ;
        RECT 349.950 553.950 352.050 554.400 ;
        RECT 379.950 555.600 382.050 556.050 ;
        RECT 418.950 555.600 421.050 556.050 ;
        RECT 379.950 554.400 421.050 555.600 ;
        RECT 379.950 553.950 382.050 554.400 ;
        RECT 418.950 553.950 421.050 554.400 ;
        RECT 448.950 555.600 451.050 556.050 ;
        RECT 478.950 555.600 481.050 556.050 ;
        RECT 448.950 554.400 481.050 555.600 ;
        RECT 448.950 553.950 451.050 554.400 ;
        RECT 478.950 553.950 481.050 554.400 ;
        RECT 553.950 555.600 556.050 556.050 ;
        RECT 601.950 555.600 604.050 556.050 ;
        RECT 553.950 554.400 604.050 555.600 ;
        RECT 553.950 553.950 556.050 554.400 ;
        RECT 601.950 553.950 604.050 554.400 ;
        RECT 697.950 555.600 700.050 556.050 ;
        RECT 760.950 555.600 763.050 556.050 ;
        RECT 697.950 554.400 763.050 555.600 ;
        RECT 697.950 553.950 700.050 554.400 ;
        RECT 760.950 553.950 763.050 554.400 ;
        RECT 361.950 552.600 364.050 553.050 ;
        RECT 433.950 552.600 436.050 553.050 ;
        RECT 302.400 551.400 436.050 552.600 ;
        RECT 148.950 550.950 151.050 551.400 ;
        RECT 229.950 550.950 232.050 551.400 ;
        RECT 271.950 550.950 274.050 551.400 ;
        RECT 361.950 550.950 364.050 551.400 ;
        RECT 433.950 550.950 436.050 551.400 ;
        RECT 454.950 552.600 457.050 553.050 ;
        RECT 502.950 552.600 505.050 553.050 ;
        RECT 454.950 551.400 505.050 552.600 ;
        RECT 454.950 550.950 457.050 551.400 ;
        RECT 502.950 550.950 505.050 551.400 ;
        RECT 583.950 552.600 586.050 553.050 ;
        RECT 607.950 552.600 610.050 553.050 ;
        RECT 583.950 551.400 610.050 552.600 ;
        RECT 583.950 550.950 586.050 551.400 ;
        RECT 607.950 550.950 610.050 551.400 ;
        RECT 754.950 552.600 757.050 553.050 ;
        RECT 772.950 552.600 775.050 553.050 ;
        RECT 754.950 551.400 775.050 552.600 ;
        RECT 754.950 550.950 757.050 551.400 ;
        RECT 772.950 550.950 775.050 551.400 ;
        RECT 901.950 552.600 904.050 553.050 ;
        RECT 916.950 552.600 919.050 553.050 ;
        RECT 901.950 551.400 919.050 552.600 ;
        RECT 901.950 550.950 904.050 551.400 ;
        RECT 916.950 550.950 919.050 551.400 ;
        RECT 103.950 549.600 106.050 550.050 ;
        RECT 130.950 549.600 133.050 550.050 ;
        RECT 103.950 548.400 133.050 549.600 ;
        RECT 103.950 547.950 106.050 548.400 ;
        RECT 130.950 547.950 133.050 548.400 ;
        RECT 247.950 549.600 250.050 550.050 ;
        RECT 256.950 549.600 259.050 550.050 ;
        RECT 247.950 548.400 259.050 549.600 ;
        RECT 247.950 547.950 250.050 548.400 ;
        RECT 256.950 547.950 259.050 548.400 ;
        RECT 280.950 549.600 283.050 550.050 ;
        RECT 322.950 549.600 325.050 550.050 ;
        RECT 364.950 549.600 367.050 550.050 ;
        RECT 280.950 548.400 321.600 549.600 ;
        RECT 280.950 547.950 283.050 548.400 ;
        RECT 187.950 546.600 190.050 547.050 ;
        RECT 247.950 546.600 250.050 546.900 ;
        RECT 295.950 546.600 298.050 547.050 ;
        RECT 187.950 545.400 246.600 546.600 ;
        RECT 187.950 544.950 190.050 545.400 ;
        RECT 1.950 543.600 4.050 544.050 ;
        RECT 49.950 543.600 52.050 544.050 ;
        RECT 64.950 543.600 67.050 544.050 ;
        RECT 1.950 542.400 67.050 543.600 ;
        RECT 245.400 543.600 246.600 545.400 ;
        RECT 247.950 545.400 298.050 546.600 ;
        RECT 320.400 546.600 321.600 548.400 ;
        RECT 322.950 548.400 367.050 549.600 ;
        RECT 322.950 547.950 325.050 548.400 ;
        RECT 364.950 547.950 367.050 548.400 ;
        RECT 436.950 549.600 439.050 550.050 ;
        RECT 490.950 549.600 493.050 550.050 ;
        RECT 436.950 548.400 493.050 549.600 ;
        RECT 436.950 547.950 439.050 548.400 ;
        RECT 490.950 547.950 493.050 548.400 ;
        RECT 496.950 549.600 499.050 550.050 ;
        RECT 622.950 549.600 625.050 550.050 ;
        RECT 652.950 549.600 655.050 550.050 ;
        RECT 751.950 549.600 754.050 550.050 ;
        RECT 496.950 548.400 534.600 549.600 ;
        RECT 496.950 547.950 499.050 548.400 ;
        RECT 352.800 546.600 354.900 547.050 ;
        RECT 320.400 545.400 354.900 546.600 ;
        RECT 247.950 544.800 250.050 545.400 ;
        RECT 295.950 544.950 298.050 545.400 ;
        RECT 352.800 544.950 354.900 545.400 ;
        RECT 355.950 546.600 358.050 547.050 ;
        RECT 394.950 546.600 397.050 547.050 ;
        RECT 355.950 545.400 397.050 546.600 ;
        RECT 355.950 544.950 358.050 545.400 ;
        RECT 394.950 544.950 397.050 545.400 ;
        RECT 409.950 546.600 412.050 547.050 ;
        RECT 457.950 546.600 460.050 547.050 ;
        RECT 409.950 545.400 460.050 546.600 ;
        RECT 409.950 544.950 412.050 545.400 ;
        RECT 457.950 544.950 460.050 545.400 ;
        RECT 475.950 546.600 478.050 547.050 ;
        RECT 487.950 546.600 490.050 547.050 ;
        RECT 475.950 545.400 490.050 546.600 ;
        RECT 533.400 546.600 534.600 548.400 ;
        RECT 622.950 548.400 754.050 549.600 ;
        RECT 622.950 547.950 625.050 548.400 ;
        RECT 652.950 547.950 655.050 548.400 ;
        RECT 751.950 547.950 754.050 548.400 ;
        RECT 787.950 549.600 790.050 550.050 ;
        RECT 838.950 549.600 841.050 550.050 ;
        RECT 787.950 548.400 841.050 549.600 ;
        RECT 787.950 547.950 790.050 548.400 ;
        RECT 838.950 547.950 841.050 548.400 ;
        RECT 880.950 549.600 883.050 550.050 ;
        RECT 913.950 549.600 916.050 550.050 ;
        RECT 880.950 548.400 916.050 549.600 ;
        RECT 880.950 547.950 883.050 548.400 ;
        RECT 913.950 547.950 916.050 548.400 ;
        RECT 583.950 546.600 586.050 547.050 ;
        RECT 533.400 545.400 586.050 546.600 ;
        RECT 475.950 544.950 478.050 545.400 ;
        RECT 487.950 544.950 490.050 545.400 ;
        RECT 583.950 544.950 586.050 545.400 ;
        RECT 649.950 546.600 652.050 547.050 ;
        RECT 673.950 546.600 676.050 547.050 ;
        RECT 649.950 545.400 676.050 546.600 ;
        RECT 649.950 544.950 652.050 545.400 ;
        RECT 673.950 544.950 676.050 545.400 ;
        RECT 679.950 546.600 682.050 547.050 ;
        RECT 715.950 546.600 718.050 547.050 ;
        RECT 679.950 545.400 718.050 546.600 ;
        RECT 679.950 544.950 682.050 545.400 ;
        RECT 715.950 544.950 718.050 545.400 ;
        RECT 904.950 546.600 907.050 547.050 ;
        RECT 916.950 546.600 919.050 547.050 ;
        RECT 904.950 545.400 919.050 546.600 ;
        RECT 904.950 544.950 907.050 545.400 ;
        RECT 916.950 544.950 919.050 545.400 ;
        RECT 259.950 543.600 262.050 544.050 ;
        RECT 245.400 542.400 262.050 543.600 ;
        RECT 1.950 541.950 4.050 542.400 ;
        RECT 49.950 541.950 52.050 542.400 ;
        RECT 64.950 541.950 67.050 542.400 ;
        RECT 259.950 541.950 262.050 542.400 ;
        RECT 292.950 543.600 295.050 544.050 ;
        RECT 370.950 543.600 373.050 544.050 ;
        RECT 292.950 542.400 373.050 543.600 ;
        RECT 292.950 541.950 295.050 542.400 ;
        RECT 370.950 541.950 373.050 542.400 ;
        RECT 430.950 543.600 433.050 544.050 ;
        RECT 499.950 543.600 502.050 544.050 ;
        RECT 430.950 542.400 502.050 543.600 ;
        RECT 430.950 541.950 433.050 542.400 ;
        RECT 499.950 541.950 502.050 542.400 ;
        RECT 529.950 543.600 532.050 544.050 ;
        RECT 541.950 543.600 544.050 544.050 ;
        RECT 637.950 543.600 640.050 544.050 ;
        RECT 529.950 542.400 640.050 543.600 ;
        RECT 529.950 541.950 532.050 542.400 ;
        RECT 541.950 541.950 544.050 542.400 ;
        RECT 637.950 541.950 640.050 542.400 ;
        RECT 751.950 543.600 754.050 544.050 ;
        RECT 781.950 543.600 784.050 544.050 ;
        RECT 787.950 543.600 790.050 544.050 ;
        RECT 751.950 542.400 790.050 543.600 ;
        RECT 751.950 541.950 754.050 542.400 ;
        RECT 781.950 541.950 784.050 542.400 ;
        RECT 787.950 541.950 790.050 542.400 ;
        RECT 859.950 543.600 862.050 544.050 ;
        RECT 877.950 543.600 880.050 544.050 ;
        RECT 859.950 542.400 880.050 543.600 ;
        RECT 859.950 541.950 862.050 542.400 ;
        RECT 877.950 541.950 880.050 542.400 ;
        RECT 28.950 540.600 31.050 541.050 ;
        RECT 112.950 540.600 115.050 541.050 ;
        RECT 28.950 539.400 115.050 540.600 ;
        RECT 28.950 538.950 31.050 539.400 ;
        RECT 112.950 538.950 115.050 539.400 ;
        RECT 142.950 540.600 145.050 541.050 ;
        RECT 160.950 540.600 163.050 541.050 ;
        RECT 142.950 539.400 163.050 540.600 ;
        RECT 142.950 538.950 145.050 539.400 ;
        RECT 160.950 538.950 163.050 539.400 ;
        RECT 175.950 540.600 178.050 541.050 ;
        RECT 184.950 540.600 187.050 541.050 ;
        RECT 175.950 539.400 187.050 540.600 ;
        RECT 175.950 538.950 178.050 539.400 ;
        RECT 184.950 538.950 187.050 539.400 ;
        RECT 232.950 540.600 235.050 541.050 ;
        RECT 241.950 540.600 244.050 541.050 ;
        RECT 232.950 539.400 244.050 540.600 ;
        RECT 232.950 538.950 235.050 539.400 ;
        RECT 241.950 538.950 244.050 539.400 ;
        RECT 262.950 540.600 265.050 541.050 ;
        RECT 283.950 540.600 286.050 541.050 ;
        RECT 262.950 539.400 286.050 540.600 ;
        RECT 262.950 538.950 265.050 539.400 ;
        RECT 283.950 538.950 286.050 539.400 ;
        RECT 364.950 540.600 367.050 541.050 ;
        RECT 373.950 540.600 376.050 541.050 ;
        RECT 364.950 539.400 376.050 540.600 ;
        RECT 364.950 538.950 367.050 539.400 ;
        RECT 373.950 538.950 376.050 539.400 ;
        RECT 397.950 540.600 400.050 541.050 ;
        RECT 475.800 540.600 477.900 541.050 ;
        RECT 397.950 539.400 477.900 540.600 ;
        RECT 397.950 538.950 400.050 539.400 ;
        RECT 475.800 538.950 477.900 539.400 ;
        RECT 478.950 540.600 481.050 541.050 ;
        RECT 484.950 540.600 487.050 541.050 ;
        RECT 478.950 539.400 487.050 540.600 ;
        RECT 478.950 538.950 481.050 539.400 ;
        RECT 484.950 538.950 487.050 539.400 ;
        RECT 547.950 540.600 550.050 541.050 ;
        RECT 676.950 540.600 679.050 541.050 ;
        RECT 547.950 539.400 679.050 540.600 ;
        RECT 547.950 538.950 550.050 539.400 ;
        RECT 676.950 538.950 679.050 539.400 ;
        RECT 694.950 540.600 697.050 541.050 ;
        RECT 718.950 540.600 721.050 541.050 ;
        RECT 694.950 539.400 721.050 540.600 ;
        RECT 694.950 538.950 697.050 539.400 ;
        RECT 718.950 538.950 721.050 539.400 ;
        RECT 832.950 540.600 835.050 541.050 ;
        RECT 856.950 540.600 859.050 541.050 ;
        RECT 832.950 539.400 859.050 540.600 ;
        RECT 832.950 538.950 835.050 539.400 ;
        RECT 856.950 538.950 859.050 539.400 ;
        RECT 889.950 540.600 892.050 541.050 ;
        RECT 913.950 540.600 916.050 541.050 ;
        RECT 889.950 539.400 916.050 540.600 ;
        RECT 889.950 538.950 892.050 539.400 ;
        RECT 913.950 538.950 916.050 539.400 ;
        RECT 40.950 537.600 43.050 538.050 ;
        RECT 52.950 537.600 55.050 538.050 ;
        RECT 40.950 536.400 55.050 537.600 ;
        RECT 40.950 535.950 43.050 536.400 ;
        RECT 52.950 535.950 55.050 536.400 ;
        RECT 205.950 537.600 208.050 538.050 ;
        RECT 232.950 537.600 235.050 537.900 ;
        RECT 205.950 536.400 235.050 537.600 ;
        RECT 205.950 535.950 208.050 536.400 ;
        RECT 232.950 535.800 235.050 536.400 ;
        RECT 259.950 537.600 262.050 538.050 ;
        RECT 286.950 537.600 289.050 538.050 ;
        RECT 259.950 536.400 289.050 537.600 ;
        RECT 259.950 535.950 262.050 536.400 ;
        RECT 286.950 535.950 289.050 536.400 ;
        RECT 328.950 537.600 331.050 538.050 ;
        RECT 340.950 537.600 343.050 538.050 ;
        RECT 355.950 537.600 358.050 538.050 ;
        RECT 328.950 536.400 358.050 537.600 ;
        RECT 328.950 535.950 331.050 536.400 ;
        RECT 340.950 535.950 343.050 536.400 ;
        RECT 355.950 535.950 358.050 536.400 ;
        RECT 427.950 537.600 430.050 538.050 ;
        RECT 451.950 537.600 454.050 538.050 ;
        RECT 427.950 536.400 454.050 537.600 ;
        RECT 427.950 535.950 430.050 536.400 ;
        RECT 451.950 535.950 454.050 536.400 ;
        RECT 625.950 537.600 628.050 538.050 ;
        RECT 655.950 537.600 658.050 538.050 ;
        RECT 625.950 536.400 658.050 537.600 ;
        RECT 625.950 535.950 628.050 536.400 ;
        RECT 655.950 535.950 658.050 536.400 ;
        RECT 835.950 537.600 838.050 538.050 ;
        RECT 868.950 537.600 871.050 538.050 ;
        RECT 835.950 536.400 871.050 537.600 ;
        RECT 835.950 535.950 838.050 536.400 ;
        RECT 868.950 535.950 871.050 536.400 ;
        RECT 100.950 534.600 103.050 535.050 ;
        RECT 92.400 533.400 103.050 534.600 ;
        RECT 92.400 532.050 93.600 533.400 ;
        RECT 100.950 532.950 103.050 533.400 ;
        RECT 115.950 534.600 118.050 535.050 ;
        RECT 142.950 534.600 145.050 535.050 ;
        RECT 115.950 533.400 145.050 534.600 ;
        RECT 115.950 532.950 118.050 533.400 ;
        RECT 142.950 532.950 145.050 533.400 ;
        RECT 151.950 534.600 154.050 535.050 ;
        RECT 166.950 534.600 169.050 535.050 ;
        RECT 151.950 533.400 169.050 534.600 ;
        RECT 151.950 532.950 154.050 533.400 ;
        RECT 166.950 532.950 169.050 533.400 ;
        RECT 178.950 534.600 181.050 535.050 ;
        RECT 187.950 534.600 190.050 535.050 ;
        RECT 178.950 533.400 190.050 534.600 ;
        RECT 178.950 532.950 181.050 533.400 ;
        RECT 187.950 532.950 190.050 533.400 ;
        RECT 193.950 534.600 196.050 535.050 ;
        RECT 199.950 534.600 202.050 535.050 ;
        RECT 235.950 534.600 238.050 535.050 ;
        RECT 277.950 534.600 280.050 535.050 ;
        RECT 193.950 533.400 238.050 534.600 ;
        RECT 193.950 532.950 196.050 533.400 ;
        RECT 199.950 532.950 202.050 533.400 ;
        RECT 235.950 532.950 238.050 533.400 ;
        RECT 263.400 533.400 280.050 534.600 ;
        RECT 79.950 531.600 82.050 532.050 ;
        RECT 91.950 531.600 94.050 532.050 ;
        RECT 79.950 530.400 94.050 531.600 ;
        RECT 79.950 529.950 82.050 530.400 ;
        RECT 91.950 529.950 94.050 530.400 ;
        RECT 256.950 531.600 259.050 532.050 ;
        RECT 263.400 531.600 264.600 533.400 ;
        RECT 277.950 532.950 280.050 533.400 ;
        RECT 460.950 534.600 463.050 535.050 ;
        RECT 472.950 534.600 475.050 535.050 ;
        RECT 460.950 533.400 475.050 534.600 ;
        RECT 460.950 532.950 463.050 533.400 ;
        RECT 472.950 532.950 475.050 533.400 ;
        RECT 481.950 534.600 484.050 535.050 ;
        RECT 535.950 534.600 538.050 535.050 ;
        RECT 481.950 533.400 538.050 534.600 ;
        RECT 481.950 532.950 484.050 533.400 ;
        RECT 535.950 532.950 538.050 533.400 ;
        RECT 670.950 534.600 673.050 535.050 ;
        RECT 679.950 534.600 682.050 535.050 ;
        RECT 670.950 533.400 682.050 534.600 ;
        RECT 670.950 532.950 673.050 533.400 ;
        RECT 679.950 532.950 682.050 533.400 ;
        RECT 703.950 534.600 706.050 535.050 ;
        RECT 733.950 534.600 736.050 535.050 ;
        RECT 703.950 533.400 736.050 534.600 ;
        RECT 703.950 532.950 706.050 533.400 ;
        RECT 733.950 532.950 736.050 533.400 ;
        RECT 766.950 534.600 769.050 535.050 ;
        RECT 793.950 534.600 796.050 535.050 ;
        RECT 766.950 533.400 796.050 534.600 ;
        RECT 766.950 532.950 769.050 533.400 ;
        RECT 793.950 532.950 796.050 533.400 ;
        RECT 883.950 534.600 886.050 535.050 ;
        RECT 910.950 534.600 913.050 535.050 ;
        RECT 883.950 533.400 913.050 534.600 ;
        RECT 883.950 532.950 886.050 533.400 ;
        RECT 910.950 532.950 913.050 533.400 ;
        RECT 256.950 530.400 264.600 531.600 ;
        RECT 385.950 531.600 388.050 532.050 ;
        RECT 412.950 531.600 415.050 532.050 ;
        RECT 430.950 531.600 433.050 532.050 ;
        RECT 385.950 530.400 433.050 531.600 ;
        RECT 256.950 529.950 259.050 530.400 ;
        RECT 385.950 529.950 388.050 530.400 ;
        RECT 412.950 529.950 415.050 530.400 ;
        RECT 430.950 529.950 433.050 530.400 ;
        RECT 553.950 531.600 556.050 532.050 ;
        RECT 559.950 531.600 562.050 532.050 ;
        RECT 553.950 530.400 562.050 531.600 ;
        RECT 553.950 529.950 556.050 530.400 ;
        RECT 559.950 529.950 562.050 530.400 ;
        RECT 580.950 531.600 583.050 532.050 ;
        RECT 610.950 531.600 613.050 532.050 ;
        RECT 903.000 531.600 907.050 532.050 ;
        RECT 580.950 530.400 613.050 531.600 ;
        RECT 580.950 529.950 583.050 530.400 ;
        RECT 610.950 529.950 613.050 530.400 ;
        RECT 902.400 529.950 907.050 531.600 ;
        RECT 19.950 528.600 22.050 528.900 ;
        RECT 34.950 528.600 37.050 529.050 ;
        RECT 19.950 527.400 37.050 528.600 ;
        RECT 19.950 526.800 22.050 527.400 ;
        RECT 34.950 526.950 37.050 527.400 ;
        RECT 64.950 528.750 67.050 529.200 ;
        RECT 73.950 528.750 76.050 529.200 ;
        RECT 64.950 527.550 76.050 528.750 ;
        RECT 94.950 528.600 97.050 529.200 ;
        RECT 64.950 527.100 67.050 527.550 ;
        RECT 73.950 527.100 76.050 527.550 ;
        RECT 80.400 527.400 97.050 528.600 ;
        RECT 80.400 525.600 81.600 527.400 ;
        RECT 94.950 527.100 97.050 527.400 ;
        RECT 100.950 526.950 103.050 529.050 ;
        RECT 109.950 527.100 112.050 529.200 ;
        RECT 124.950 528.750 127.050 529.200 ;
        RECT 136.950 528.750 139.050 529.200 ;
        RECT 124.950 527.550 139.050 528.750 ;
        RECT 124.950 527.100 127.050 527.550 ;
        RECT 136.950 527.100 139.050 527.550 ;
        RECT 77.400 524.400 81.600 525.600 ;
        RECT 7.950 522.300 10.050 522.750 ;
        RECT 10.950 522.300 13.050 523.050 ;
        RECT 13.950 522.300 16.050 522.750 ;
        RECT 7.950 521.100 16.050 522.300 ;
        RECT 7.950 520.650 10.050 521.100 ;
        RECT 10.950 520.950 13.050 521.100 ;
        RECT 13.950 520.650 16.050 521.100 ;
        RECT 52.950 522.600 55.050 522.900 ;
        RECT 64.950 522.600 67.050 523.050 ;
        RECT 77.400 522.900 78.600 524.400 ;
        RECT 101.400 523.050 102.600 526.950 ;
        RECT 110.400 525.600 111.600 527.100 ;
        RECT 148.950 526.950 151.050 529.050 ;
        RECT 187.950 528.600 190.050 529.200 ;
        RECT 208.950 528.600 211.050 529.200 ;
        RECT 187.950 527.400 211.050 528.600 ;
        RECT 187.950 527.100 190.050 527.400 ;
        RECT 208.950 527.100 211.050 527.400 ;
        RECT 214.950 527.100 217.050 529.200 ;
        RECT 235.950 528.600 238.050 529.200 ;
        RECT 250.950 528.600 253.050 529.200 ;
        RECT 235.950 527.400 253.050 528.600 ;
        RECT 235.950 527.100 238.050 527.400 ;
        RECT 250.950 527.100 253.050 527.400 ;
        RECT 265.950 527.100 268.050 529.200 ;
        RECT 110.400 524.400 132.600 525.600 ;
        RECT 131.400 523.050 132.600 524.400 ;
        RECT 52.950 521.400 67.050 522.600 ;
        RECT 52.950 520.800 55.050 521.400 ;
        RECT 64.950 520.950 67.050 521.400 ;
        RECT 76.950 520.800 79.050 522.900 ;
        RECT 100.950 520.950 103.050 523.050 ;
        RECT 118.950 522.600 121.050 522.900 ;
        RECT 124.950 522.600 127.050 523.050 ;
        RECT 118.950 521.400 127.050 522.600 ;
        RECT 131.400 521.400 136.050 523.050 ;
        RECT 118.950 520.800 121.050 521.400 ;
        RECT 124.950 520.950 127.050 521.400 ;
        RECT 132.000 520.950 136.050 521.400 ;
        RECT 139.950 522.600 142.050 522.900 ;
        RECT 149.400 522.600 150.600 526.950 ;
        RECT 139.950 521.400 150.600 522.600 ;
        RECT 215.400 523.050 216.600 527.100 ;
        RECT 259.950 525.600 262.050 526.050 ;
        RECT 233.400 524.400 262.050 525.600 ;
        RECT 215.400 521.400 220.050 523.050 ;
        RECT 233.400 522.900 234.600 524.400 ;
        RECT 259.950 523.950 262.050 524.400 ;
        RECT 139.950 520.800 142.050 521.400 ;
        RECT 216.000 520.950 220.050 521.400 ;
        RECT 232.950 520.800 235.050 522.900 ;
        RECT 247.950 522.600 250.050 522.900 ;
        RECT 266.400 522.600 267.600 527.100 ;
        RECT 283.950 525.600 286.050 529.050 ;
        RECT 304.950 528.600 307.050 529.050 ;
        RECT 334.950 528.600 337.050 529.200 ;
        RECT 304.950 527.400 337.050 528.600 ;
        RECT 304.950 526.950 307.050 527.400 ;
        RECT 334.950 527.100 337.050 527.400 ;
        RECT 343.950 526.950 346.050 529.050 ;
        RECT 352.950 528.600 355.050 529.050 ;
        RECT 352.950 527.400 360.600 528.600 ;
        RECT 352.950 526.950 355.050 527.400 ;
        RECT 283.950 525.000 297.600 525.600 ;
        RECT 284.400 524.400 297.600 525.000 ;
        RECT 247.950 521.400 267.600 522.600 ;
        RECT 274.950 522.600 277.050 522.900 ;
        RECT 292.950 522.600 295.050 522.900 ;
        RECT 274.950 521.400 295.050 522.600 ;
        RECT 296.400 522.600 297.600 524.400 ;
        RECT 344.400 523.050 345.600 526.950 ;
        RECT 319.950 522.600 322.050 523.050 ;
        RECT 296.400 521.400 322.050 522.600 ;
        RECT 247.950 520.800 250.050 521.400 ;
        RECT 274.950 520.800 277.050 521.400 ;
        RECT 292.950 520.800 295.050 521.400 ;
        RECT 319.950 520.950 322.050 521.400 ;
        RECT 343.950 520.950 346.050 523.050 ;
        RECT 359.400 522.900 360.600 527.400 ;
        RECT 361.950 525.600 364.050 529.050 ;
        RECT 382.950 526.950 385.050 529.050 ;
        RECT 361.950 525.000 372.600 525.600 ;
        RECT 362.400 524.400 373.050 525.000 ;
        RECT 358.950 520.800 361.050 522.900 ;
        RECT 370.950 520.950 373.050 524.400 ;
        RECT 383.400 522.600 384.600 526.950 ;
        RECT 385.950 525.600 388.050 526.050 ;
        RECT 424.950 525.600 427.050 526.050 ;
        RECT 385.950 524.400 427.050 525.600 ;
        RECT 427.950 525.600 430.050 529.050 ;
        RECT 442.950 528.750 445.050 529.200 ;
        RECT 448.950 528.750 451.050 529.200 ;
        RECT 442.950 527.550 451.050 528.750 ;
        RECT 442.950 527.100 445.050 527.550 ;
        RECT 448.950 527.100 451.050 527.550 ;
        RECT 466.950 527.100 469.050 529.200 ;
        RECT 427.950 525.000 435.600 525.600 ;
        RECT 428.400 524.400 435.600 525.000 ;
        RECT 385.950 523.950 388.050 524.400 ;
        RECT 424.950 523.950 427.050 524.400 ;
        RECT 388.950 522.600 391.050 523.050 ;
        RECT 434.400 522.900 435.600 524.400 ;
        RECT 383.400 521.400 391.050 522.600 ;
        RECT 388.950 520.950 391.050 521.400 ;
        RECT 433.950 520.800 436.050 522.900 ;
        RECT 467.400 522.600 468.600 527.100 ;
        RECT 472.950 525.600 475.050 529.050 ;
        RECT 478.950 527.100 481.050 529.200 ;
        RECT 472.950 525.000 477.600 525.600 ;
        RECT 473.400 524.400 478.050 525.000 ;
        RECT 472.800 522.600 474.900 523.050 ;
        RECT 467.400 521.400 474.900 522.600 ;
        RECT 472.800 520.950 474.900 521.400 ;
        RECT 475.950 520.950 478.050 524.400 ;
        RECT 479.400 520.050 480.600 527.100 ;
        RECT 487.950 526.950 490.050 529.050 ;
        RECT 499.950 527.100 502.050 529.200 ;
        RECT 514.950 528.750 517.050 529.200 ;
        RECT 523.950 528.750 526.050 529.200 ;
        RECT 514.950 527.550 526.050 528.750 ;
        RECT 514.950 527.100 517.050 527.550 ;
        RECT 523.950 527.100 526.050 527.550 ;
        RECT 529.950 528.600 532.050 529.200 ;
        RECT 544.950 528.600 547.050 529.200 ;
        RECT 529.950 527.400 547.050 528.600 ;
        RECT 529.950 527.100 532.050 527.400 ;
        RECT 544.950 527.100 547.050 527.400 ;
        RECT 562.950 528.600 565.050 529.200 ;
        RECT 568.950 528.600 571.050 529.050 ;
        RECT 562.950 527.400 571.050 528.600 ;
        RECT 562.950 527.100 565.050 527.400 ;
        RECT 488.400 523.050 489.600 526.950 ;
        RECT 500.400 525.600 501.600 527.100 ;
        RECT 568.950 526.950 571.050 527.400 ;
        RECT 589.950 525.600 592.050 529.050 ;
        RECT 634.950 528.600 637.050 529.050 ;
        RECT 655.950 528.600 658.050 529.200 ;
        RECT 673.950 528.600 676.050 529.200 ;
        RECT 634.950 527.400 676.050 528.600 ;
        RECT 634.950 526.950 637.050 527.400 ;
        RECT 655.950 527.100 658.050 527.400 ;
        RECT 673.950 527.100 676.050 527.400 ;
        RECT 682.950 526.950 685.050 529.050 ;
        RECT 700.950 526.950 703.050 529.050 ;
        RECT 712.950 528.600 715.050 529.500 ;
        RECT 748.950 528.600 751.050 529.500 ;
        RECT 712.950 527.400 751.050 528.600 ;
        RECT 601.950 525.600 604.050 526.050 ;
        RECT 494.400 525.000 501.600 525.600 ;
        RECT 493.950 524.400 501.600 525.000 ;
        RECT 518.400 524.400 594.600 525.600 ;
        RECT 487.950 520.950 490.050 523.050 ;
        RECT 493.950 520.950 496.050 524.400 ;
        RECT 508.950 522.600 511.050 523.050 ;
        RECT 518.400 522.600 519.600 524.400 ;
        RECT 508.950 521.400 519.600 522.600 ;
        RECT 520.950 522.450 523.050 522.900 ;
        RECT 535.950 522.450 538.050 522.900 ;
        RECT 508.950 520.950 511.050 521.400 ;
        RECT 520.950 521.250 538.050 522.450 ;
        RECT 520.950 520.800 523.050 521.250 ;
        RECT 535.950 520.800 538.050 521.250 ;
        RECT 547.950 522.450 550.050 522.900 ;
        RECT 553.950 522.600 556.050 522.900 ;
        RECT 565.950 522.600 568.050 523.050 ;
        RECT 593.400 522.600 594.600 524.400 ;
        RECT 601.950 524.400 654.600 525.600 ;
        RECT 601.950 523.950 604.050 524.400 ;
        RECT 653.400 522.600 654.600 524.400 ;
        RECT 658.950 522.600 661.050 523.050 ;
        RECT 553.950 522.450 568.050 522.600 ;
        RECT 547.950 521.400 568.050 522.450 ;
        RECT 547.950 521.250 556.050 521.400 ;
        RECT 547.950 520.800 550.050 521.250 ;
        RECT 553.950 520.800 556.050 521.250 ;
        RECT 565.950 520.950 568.050 521.400 ;
        RECT 592.950 520.500 595.050 522.600 ;
        RECT 653.400 521.400 661.050 522.600 ;
        RECT 658.950 520.950 661.050 521.400 ;
        RECT 670.950 522.600 673.050 523.050 ;
        RECT 683.400 522.600 684.600 526.950 ;
        RECT 670.950 521.400 684.600 522.600 ;
        RECT 701.400 522.600 702.600 526.950 ;
        RECT 754.950 525.600 757.050 529.050 ;
        RECT 772.950 526.950 775.050 529.050 ;
        RECT 778.950 528.600 781.050 529.050 ;
        RECT 778.950 527.400 789.600 528.600 ;
        RECT 778.950 526.950 781.050 527.400 ;
        RECT 754.950 525.000 759.600 525.600 ;
        RECT 755.400 524.400 759.600 525.000 ;
        RECT 751.800 522.600 753.900 523.050 ;
        RECT 758.400 522.600 759.600 524.400 ;
        RECT 773.400 523.050 774.600 526.950 ;
        RECT 788.400 523.050 789.600 527.400 ;
        RECT 808.950 525.600 811.050 529.050 ;
        RECT 829.950 528.600 832.050 529.050 ;
        RECT 829.950 527.400 837.600 528.600 ;
        RECT 829.950 526.950 832.050 527.400 ;
        RECT 808.950 525.000 831.600 525.600 ;
        RECT 809.400 524.400 832.050 525.000 ;
        RECT 701.400 521.400 753.900 522.600 ;
        RECT 670.950 520.950 673.050 521.400 ;
        RECT 751.800 520.950 753.900 521.400 ;
        RECT 757.950 520.500 760.050 522.600 ;
        RECT 772.950 520.950 775.050 523.050 ;
        RECT 787.950 520.950 790.050 523.050 ;
        RECT 829.950 520.950 832.050 524.400 ;
        RECT 836.400 522.900 837.600 527.400 ;
        RECT 859.950 527.100 862.050 529.200 ;
        RECT 865.950 528.600 868.050 529.200 ;
        RECT 871.950 528.600 874.050 529.050 ;
        RECT 865.950 527.400 874.050 528.600 ;
        RECT 865.950 527.100 868.050 527.400 ;
        RECT 835.950 520.800 838.050 522.900 ;
        RECT 22.950 519.600 25.050 520.050 ;
        RECT 34.950 519.600 37.050 520.050 ;
        RECT 97.950 519.600 100.050 520.050 ;
        RECT 22.950 518.400 100.050 519.600 ;
        RECT 22.950 517.950 25.050 518.400 ;
        RECT 34.950 517.950 37.050 518.400 ;
        RECT 97.950 517.950 100.050 518.400 ;
        RECT 127.950 519.600 130.050 520.050 ;
        RECT 145.950 519.600 148.050 520.050 ;
        RECT 154.950 519.600 157.050 520.050 ;
        RECT 127.950 518.400 157.050 519.600 ;
        RECT 127.950 517.950 130.050 518.400 ;
        RECT 145.950 517.950 148.050 518.400 ;
        RECT 154.950 517.950 157.050 518.400 ;
        RECT 256.950 519.600 259.050 520.050 ;
        RECT 265.950 519.600 268.050 520.050 ;
        RECT 256.950 518.400 268.050 519.600 ;
        RECT 256.950 517.950 259.050 518.400 ;
        RECT 265.950 517.950 268.050 518.400 ;
        RECT 307.950 519.600 310.050 520.050 ;
        RECT 316.950 519.600 319.050 520.050 ;
        RECT 307.950 518.400 319.050 519.600 ;
        RECT 307.950 517.950 310.050 518.400 ;
        RECT 316.950 517.950 319.050 518.400 ;
        RECT 376.950 519.600 379.050 520.050 ;
        RECT 445.950 519.600 448.050 520.050 ;
        RECT 376.950 518.400 448.050 519.600 ;
        RECT 376.950 517.950 379.050 518.400 ;
        RECT 445.950 517.950 448.050 518.400 ;
        RECT 478.950 517.950 481.050 520.050 ;
        RECT 490.950 519.600 493.050 520.050 ;
        RECT 496.950 519.600 499.050 520.050 ;
        RECT 490.950 518.400 499.050 519.600 ;
        RECT 490.950 517.950 493.050 518.400 ;
        RECT 496.950 517.950 499.050 518.400 ;
        RECT 604.950 519.600 607.050 520.050 ;
        RECT 610.950 519.600 613.050 520.050 ;
        RECT 604.950 518.400 613.050 519.600 ;
        RECT 604.950 517.950 607.050 518.400 ;
        RECT 610.950 517.950 613.050 518.400 ;
        RECT 661.950 519.600 664.050 520.050 ;
        RECT 679.950 519.600 682.050 520.050 ;
        RECT 661.950 518.400 682.050 519.600 ;
        RECT 661.950 517.950 664.050 518.400 ;
        RECT 679.950 517.950 682.050 518.400 ;
        RECT 694.950 519.600 697.050 520.050 ;
        RECT 703.950 519.600 706.050 520.050 ;
        RECT 694.950 518.400 706.050 519.600 ;
        RECT 694.950 517.950 697.050 518.400 ;
        RECT 703.950 517.950 706.050 518.400 ;
        RECT 823.950 519.600 826.050 520.050 ;
        RECT 838.950 519.600 841.050 520.050 ;
        RECT 823.950 518.400 841.050 519.600 ;
        RECT 823.950 517.950 826.050 518.400 ;
        RECT 838.950 517.950 841.050 518.400 ;
        RECT 4.950 516.600 7.050 517.050 ;
        RECT 88.950 516.600 91.050 517.050 ;
        RECT 4.950 515.400 91.050 516.600 ;
        RECT 4.950 514.950 7.050 515.400 ;
        RECT 88.950 514.950 91.050 515.400 ;
        RECT 130.950 516.600 133.050 517.050 ;
        RECT 136.950 516.600 139.050 517.050 ;
        RECT 130.950 515.400 139.050 516.600 ;
        RECT 130.950 514.950 133.050 515.400 ;
        RECT 136.950 514.950 139.050 515.400 ;
        RECT 163.950 516.600 166.050 517.050 ;
        RECT 190.950 516.600 193.050 517.050 ;
        RECT 211.950 516.600 214.050 517.050 ;
        RECT 163.950 515.400 214.050 516.600 ;
        RECT 163.950 514.950 166.050 515.400 ;
        RECT 190.950 514.950 193.050 515.400 ;
        RECT 211.950 514.950 214.050 515.400 ;
        RECT 217.950 516.600 220.050 517.050 ;
        RECT 247.950 516.600 250.050 517.050 ;
        RECT 217.950 515.400 250.050 516.600 ;
        RECT 217.950 514.950 220.050 515.400 ;
        RECT 247.950 514.950 250.050 515.400 ;
        RECT 259.950 516.600 262.050 517.050 ;
        RECT 268.950 516.600 271.050 517.050 ;
        RECT 259.950 515.400 271.050 516.600 ;
        RECT 259.950 514.950 262.050 515.400 ;
        RECT 268.950 514.950 271.050 515.400 ;
        RECT 274.950 516.600 277.050 517.050 ;
        RECT 280.950 516.600 283.050 517.050 ;
        RECT 274.950 515.400 283.050 516.600 ;
        RECT 274.950 514.950 277.050 515.400 ;
        RECT 280.950 514.950 283.050 515.400 ;
        RECT 319.950 516.600 322.050 517.050 ;
        RECT 337.950 516.600 340.050 517.050 ;
        RECT 385.950 516.600 388.050 517.050 ;
        RECT 319.950 515.400 388.050 516.600 ;
        RECT 319.950 514.950 322.050 515.400 ;
        RECT 337.950 514.950 340.050 515.400 ;
        RECT 385.950 514.950 388.050 515.400 ;
        RECT 421.950 516.600 424.050 517.050 ;
        RECT 448.950 516.600 451.050 517.050 ;
        RECT 421.950 515.400 451.050 516.600 ;
        RECT 421.950 514.950 424.050 515.400 ;
        RECT 448.950 514.950 451.050 515.400 ;
        RECT 472.950 516.600 475.050 517.050 ;
        RECT 481.950 516.600 484.050 517.050 ;
        RECT 472.950 515.400 484.050 516.600 ;
        RECT 472.950 514.950 475.050 515.400 ;
        RECT 481.950 514.950 484.050 515.400 ;
        RECT 535.950 516.600 538.050 517.050 ;
        RECT 559.950 516.600 562.050 517.050 ;
        RECT 535.950 515.400 562.050 516.600 ;
        RECT 535.950 514.950 538.050 515.400 ;
        RECT 559.950 514.950 562.050 515.400 ;
        RECT 664.950 516.600 667.050 517.050 ;
        RECT 718.950 516.600 721.050 517.050 ;
        RECT 664.950 515.400 721.050 516.600 ;
        RECT 860.400 516.600 861.600 527.100 ;
        RECT 871.950 526.950 874.050 527.400 ;
        RECT 880.950 526.950 883.050 529.050 ;
        RECT 892.950 528.600 895.050 529.050 ;
        RECT 898.950 528.600 901.050 529.050 ;
        RECT 892.950 527.400 901.050 528.600 ;
        RECT 892.950 526.950 895.050 527.400 ;
        RECT 898.950 526.950 901.050 527.400 ;
        RECT 881.400 523.050 882.600 526.950 ;
        RECT 902.400 525.600 903.600 529.950 ;
        RECT 916.950 528.600 919.050 529.050 ;
        RECT 896.400 524.400 903.600 525.600 ;
        RECT 911.400 527.400 919.050 528.600 ;
        RECT 862.950 522.450 865.050 522.900 ;
        RECT 868.950 522.450 871.050 522.900 ;
        RECT 862.950 521.250 871.050 522.450 ;
        RECT 862.950 520.800 865.050 521.250 ;
        RECT 868.950 520.800 871.050 521.250 ;
        RECT 880.950 520.950 883.050 523.050 ;
        RECT 896.400 522.600 897.600 524.400 ;
        RECT 911.400 522.900 912.600 527.400 ;
        RECT 916.950 526.950 919.050 527.400 ;
        RECT 890.400 522.000 897.600 522.600 ;
        RECT 889.950 521.400 897.600 522.000 ;
        RECT 889.950 517.950 892.050 521.400 ;
        RECT 910.950 520.800 913.050 522.900 ;
        RECT 886.950 516.600 889.050 517.050 ;
        RECT 860.400 515.400 889.050 516.600 ;
        RECT 664.950 514.950 667.050 515.400 ;
        RECT 718.950 514.950 721.050 515.400 ;
        RECT 886.950 514.950 889.050 515.400 ;
        RECT 94.950 513.600 97.050 514.050 ;
        RECT 103.800 513.600 105.900 514.050 ;
        RECT 94.950 512.400 105.900 513.600 ;
        RECT 94.950 511.950 97.050 512.400 ;
        RECT 103.800 511.950 105.900 512.400 ;
        RECT 106.950 513.600 109.050 514.050 ;
        RECT 133.950 513.600 136.050 514.050 ;
        RECT 106.950 512.400 136.050 513.600 ;
        RECT 106.950 511.950 109.050 512.400 ;
        RECT 133.950 511.950 136.050 512.400 ;
        RECT 289.950 513.600 292.050 514.050 ;
        RECT 304.950 513.600 307.050 514.050 ;
        RECT 289.950 512.400 307.050 513.600 ;
        RECT 289.950 511.950 292.050 512.400 ;
        RECT 304.950 511.950 307.050 512.400 ;
        RECT 340.950 513.600 343.050 514.050 ;
        RECT 394.950 513.600 397.050 514.050 ;
        RECT 340.950 512.400 397.050 513.600 ;
        RECT 340.950 511.950 343.050 512.400 ;
        RECT 394.950 511.950 397.050 512.400 ;
        RECT 415.950 513.600 418.050 514.050 ;
        RECT 469.950 513.600 472.050 514.050 ;
        RECT 415.950 512.400 472.050 513.600 ;
        RECT 415.950 511.950 418.050 512.400 ;
        RECT 469.950 511.950 472.050 512.400 ;
        RECT 487.950 513.600 490.050 514.050 ;
        RECT 514.950 513.600 517.050 514.050 ;
        RECT 487.950 512.400 517.050 513.600 ;
        RECT 487.950 511.950 490.050 512.400 ;
        RECT 514.950 511.950 517.050 512.400 ;
        RECT 574.950 513.600 577.050 514.050 ;
        RECT 607.950 513.600 610.050 514.050 ;
        RECT 574.950 512.400 610.050 513.600 ;
        RECT 574.950 511.950 577.050 512.400 ;
        RECT 607.950 511.950 610.050 512.400 ;
        RECT 817.950 513.600 820.050 514.050 ;
        RECT 856.950 513.600 859.050 514.050 ;
        RECT 817.950 512.400 859.050 513.600 ;
        RECT 817.950 511.950 820.050 512.400 ;
        RECT 856.950 511.950 859.050 512.400 ;
        RECT 865.950 513.600 868.050 514.050 ;
        RECT 874.950 513.600 877.050 514.050 ;
        RECT 865.950 512.400 877.050 513.600 ;
        RECT 865.950 511.950 868.050 512.400 ;
        RECT 874.950 511.950 877.050 512.400 ;
        RECT 16.950 510.600 19.050 511.050 ;
        RECT 112.950 510.600 115.050 511.050 ;
        RECT 16.950 509.400 115.050 510.600 ;
        RECT 16.950 508.950 19.050 509.400 ;
        RECT 112.950 508.950 115.050 509.400 ;
        RECT 127.950 510.600 130.050 511.050 ;
        RECT 151.950 510.600 154.050 511.050 ;
        RECT 127.950 509.400 154.050 510.600 ;
        RECT 127.950 508.950 130.050 509.400 ;
        RECT 151.950 508.950 154.050 509.400 ;
        RECT 172.950 510.600 175.050 511.050 ;
        RECT 205.950 510.600 208.050 511.050 ;
        RECT 172.950 509.400 208.050 510.600 ;
        RECT 172.950 508.950 175.050 509.400 ;
        RECT 205.950 508.950 208.050 509.400 ;
        RECT 220.950 510.600 223.050 511.050 ;
        RECT 301.950 510.600 304.050 511.050 ;
        RECT 220.950 509.400 304.050 510.600 ;
        RECT 220.950 508.950 223.050 509.400 ;
        RECT 301.950 508.950 304.050 509.400 ;
        RECT 310.950 510.600 313.050 511.050 ;
        RECT 331.950 510.600 334.050 511.050 ;
        RECT 310.950 509.400 334.050 510.600 ;
        RECT 310.950 508.950 313.050 509.400 ;
        RECT 331.950 508.950 334.050 509.400 ;
        RECT 337.950 510.600 340.050 511.050 ;
        RECT 376.950 510.600 379.050 511.050 ;
        RECT 337.950 509.400 379.050 510.600 ;
        RECT 337.950 508.950 340.050 509.400 ;
        RECT 376.950 508.950 379.050 509.400 ;
        RECT 439.950 510.600 442.050 511.050 ;
        RECT 466.950 510.600 469.050 511.050 ;
        RECT 478.950 510.600 481.050 511.050 ;
        RECT 520.950 510.600 523.050 511.050 ;
        RECT 439.950 509.400 523.050 510.600 ;
        RECT 439.950 508.950 442.050 509.400 ;
        RECT 466.950 508.950 469.050 509.400 ;
        RECT 478.950 508.950 481.050 509.400 ;
        RECT 520.950 508.950 523.050 509.400 ;
        RECT 586.950 510.600 589.050 511.050 ;
        RECT 661.950 510.600 664.050 511.050 ;
        RECT 586.950 509.400 664.050 510.600 ;
        RECT 586.950 508.950 589.050 509.400 ;
        RECT 661.950 508.950 664.050 509.400 ;
        RECT 676.950 510.600 679.050 511.050 ;
        RECT 721.950 510.600 724.050 511.050 ;
        RECT 676.950 509.400 724.050 510.600 ;
        RECT 676.950 508.950 679.050 509.400 ;
        RECT 721.950 508.950 724.050 509.400 ;
        RECT 760.950 510.600 763.050 511.050 ;
        RECT 769.950 510.600 772.050 511.050 ;
        RECT 760.950 509.400 772.050 510.600 ;
        RECT 760.950 508.950 763.050 509.400 ;
        RECT 769.950 508.950 772.050 509.400 ;
        RECT 787.950 510.600 790.050 511.050 ;
        RECT 814.950 510.600 817.050 511.050 ;
        RECT 787.950 509.400 817.050 510.600 ;
        RECT 787.950 508.950 790.050 509.400 ;
        RECT 814.950 508.950 817.050 509.400 ;
        RECT 826.950 510.600 829.050 511.050 ;
        RECT 832.950 510.600 835.050 511.050 ;
        RECT 826.950 509.400 835.050 510.600 ;
        RECT 826.950 508.950 829.050 509.400 ;
        RECT 832.950 508.950 835.050 509.400 ;
        RECT 229.950 507.600 232.050 508.050 ;
        RECT 241.950 507.600 244.050 508.050 ;
        RECT 229.950 506.400 244.050 507.600 ;
        RECT 229.950 505.950 232.050 506.400 ;
        RECT 241.950 505.950 244.050 506.400 ;
        RECT 283.950 507.600 286.050 508.050 ;
        RECT 298.950 507.600 301.050 508.050 ;
        RECT 283.950 506.400 301.050 507.600 ;
        RECT 283.950 505.950 286.050 506.400 ;
        RECT 298.950 505.950 301.050 506.400 ;
        RECT 346.950 507.600 349.050 508.050 ;
        RECT 355.800 507.600 357.900 508.050 ;
        RECT 346.950 506.400 357.900 507.600 ;
        RECT 346.950 505.950 349.050 506.400 ;
        RECT 355.800 505.950 357.900 506.400 ;
        RECT 358.950 507.600 361.050 508.050 ;
        RECT 364.950 507.600 367.050 508.050 ;
        RECT 358.950 506.400 367.050 507.600 ;
        RECT 358.950 505.950 361.050 506.400 ;
        RECT 364.950 505.950 367.050 506.400 ;
        RECT 382.950 507.600 385.050 508.050 ;
        RECT 409.950 507.600 412.050 508.050 ;
        RECT 382.950 506.400 412.050 507.600 ;
        RECT 382.950 505.950 385.050 506.400 ;
        RECT 409.950 505.950 412.050 506.400 ;
        RECT 433.950 507.600 436.050 508.050 ;
        RECT 451.950 507.600 454.050 508.050 ;
        RECT 433.950 506.400 454.050 507.600 ;
        RECT 433.950 505.950 436.050 506.400 ;
        RECT 451.950 505.950 454.050 506.400 ;
        RECT 487.950 507.600 490.050 508.050 ;
        RECT 493.950 507.600 496.050 508.050 ;
        RECT 487.950 506.400 496.050 507.600 ;
        RECT 487.950 505.950 490.050 506.400 ;
        RECT 493.950 505.950 496.050 506.400 ;
        RECT 631.950 507.600 634.050 508.050 ;
        RECT 685.950 507.600 688.050 508.050 ;
        RECT 631.950 506.400 688.050 507.600 ;
        RECT 631.950 505.950 634.050 506.400 ;
        RECT 685.950 505.950 688.050 506.400 ;
        RECT 787.950 507.600 790.050 507.900 ;
        RECT 799.950 507.600 802.050 508.050 ;
        RECT 817.950 507.600 820.050 508.050 ;
        RECT 787.950 506.400 820.050 507.600 ;
        RECT 787.950 505.800 790.050 506.400 ;
        RECT 799.950 505.950 802.050 506.400 ;
        RECT 817.950 505.950 820.050 506.400 ;
        RECT 856.950 507.600 859.050 508.050 ;
        RECT 862.950 507.600 865.050 508.050 ;
        RECT 856.950 506.400 865.050 507.600 ;
        RECT 856.950 505.950 859.050 506.400 ;
        RECT 862.950 505.950 865.050 506.400 ;
        RECT 877.950 507.600 880.050 508.050 ;
        RECT 901.950 507.600 904.050 508.050 ;
        RECT 877.950 506.400 904.050 507.600 ;
        RECT 877.950 505.950 880.050 506.400 ;
        RECT 901.950 505.950 904.050 506.400 ;
        RECT 55.950 504.600 58.050 505.050 ;
        RECT 79.950 504.600 82.050 505.050 ;
        RECT 55.950 503.400 82.050 504.600 ;
        RECT 55.950 502.950 58.050 503.400 ;
        RECT 79.950 502.950 82.050 503.400 ;
        RECT 112.950 504.600 115.050 505.050 ;
        RECT 148.950 504.600 151.050 505.050 ;
        RECT 112.950 503.400 151.050 504.600 ;
        RECT 112.950 502.950 115.050 503.400 ;
        RECT 148.950 502.950 151.050 503.400 ;
        RECT 154.950 504.600 157.050 505.050 ;
        RECT 166.950 504.600 169.050 505.050 ;
        RECT 154.950 503.400 169.050 504.600 ;
        RECT 154.950 502.950 157.050 503.400 ;
        RECT 166.950 502.950 169.050 503.400 ;
        RECT 172.950 504.600 175.050 505.050 ;
        RECT 184.950 504.600 187.050 505.050 ;
        RECT 280.950 504.600 283.050 505.050 ;
        RECT 172.950 503.400 283.050 504.600 ;
        RECT 172.950 502.950 175.050 503.400 ;
        RECT 184.950 502.950 187.050 503.400 ;
        RECT 280.950 502.950 283.050 503.400 ;
        RECT 301.950 504.600 304.050 505.050 ;
        RECT 337.950 504.600 340.050 505.050 ;
        RECT 301.950 503.400 340.050 504.600 ;
        RECT 301.950 502.950 304.050 503.400 ;
        RECT 337.950 502.950 340.050 503.400 ;
        RECT 367.950 504.600 370.050 505.050 ;
        RECT 379.950 504.600 382.050 505.050 ;
        RECT 367.950 503.400 382.050 504.600 ;
        RECT 367.950 502.950 370.050 503.400 ;
        RECT 379.950 502.950 382.050 503.400 ;
        RECT 406.950 504.600 409.050 505.050 ;
        RECT 415.950 504.600 418.050 505.050 ;
        RECT 406.950 503.400 418.050 504.600 ;
        RECT 406.950 502.950 409.050 503.400 ;
        RECT 415.950 502.950 418.050 503.400 ;
        RECT 424.950 504.600 427.050 505.050 ;
        RECT 598.950 504.600 601.050 505.050 ;
        RECT 424.950 503.400 492.600 504.600 ;
        RECT 424.950 502.950 427.050 503.400 ;
        RECT 61.950 501.600 64.050 502.050 ;
        RECT 70.950 501.600 73.050 502.050 ;
        RECT 61.950 500.400 73.050 501.600 ;
        RECT 61.950 499.950 64.050 500.400 ;
        RECT 70.950 499.950 73.050 500.400 ;
        RECT 91.950 501.600 94.050 502.050 ;
        RECT 106.950 501.600 109.050 502.050 ;
        RECT 91.950 500.400 109.050 501.600 ;
        RECT 91.950 499.950 94.050 500.400 ;
        RECT 106.950 499.950 109.050 500.400 ;
        RECT 187.950 501.600 190.050 502.050 ;
        RECT 232.950 501.600 235.050 502.050 ;
        RECT 187.950 500.400 235.050 501.600 ;
        RECT 187.950 499.950 190.050 500.400 ;
        RECT 232.950 499.950 235.050 500.400 ;
        RECT 241.950 501.600 244.050 502.050 ;
        RECT 262.950 501.600 265.050 502.050 ;
        RECT 241.950 500.400 265.050 501.600 ;
        RECT 241.950 499.950 244.050 500.400 ;
        RECT 262.950 499.950 265.050 500.400 ;
        RECT 301.950 501.600 304.050 501.900 ;
        RECT 328.950 501.600 331.050 502.050 ;
        RECT 340.950 501.600 343.050 502.050 ;
        RECT 301.950 500.400 343.050 501.600 ;
        RECT 301.950 499.800 304.050 500.400 ;
        RECT 328.950 499.950 331.050 500.400 ;
        RECT 340.950 499.950 343.050 500.400 ;
        RECT 349.950 501.600 352.050 502.050 ;
        RECT 373.950 501.600 376.050 502.050 ;
        RECT 349.950 500.400 376.050 501.600 ;
        RECT 349.950 499.950 352.050 500.400 ;
        RECT 373.950 499.950 376.050 500.400 ;
        RECT 382.950 501.600 385.050 501.900 ;
        RECT 388.950 501.600 391.050 502.050 ;
        RECT 400.950 501.600 403.050 502.050 ;
        RECT 382.950 500.400 403.050 501.600 ;
        RECT 382.950 499.800 385.050 500.400 ;
        RECT 388.950 499.950 391.050 500.400 ;
        RECT 400.950 499.950 403.050 500.400 ;
        RECT 436.950 501.600 439.050 502.050 ;
        RECT 445.950 501.600 448.050 502.050 ;
        RECT 460.950 501.600 463.050 502.050 ;
        RECT 436.950 500.400 463.050 501.600 ;
        RECT 436.950 499.950 439.050 500.400 ;
        RECT 445.950 499.950 448.050 500.400 ;
        RECT 460.950 499.950 463.050 500.400 ;
        RECT 469.950 501.600 472.050 502.050 ;
        RECT 481.950 501.600 484.050 502.050 ;
        RECT 469.950 500.400 484.050 501.600 ;
        RECT 491.400 501.600 492.600 503.400 ;
        RECT 581.400 503.400 601.050 504.600 ;
        RECT 581.400 502.050 582.600 503.400 ;
        RECT 598.950 502.950 601.050 503.400 ;
        RECT 715.950 504.600 718.050 505.050 ;
        RECT 733.950 504.600 736.050 505.050 ;
        RECT 715.950 503.400 736.050 504.600 ;
        RECT 715.950 502.950 718.050 503.400 ;
        RECT 733.950 502.950 736.050 503.400 ;
        RECT 754.950 504.600 757.050 505.050 ;
        RECT 769.950 504.600 772.050 505.050 ;
        RECT 754.950 503.400 772.050 504.600 ;
        RECT 754.950 502.950 757.050 503.400 ;
        RECT 769.950 502.950 772.050 503.400 ;
        RECT 835.950 504.600 838.050 505.050 ;
        RECT 844.950 504.600 847.050 505.050 ;
        RECT 835.950 503.400 847.050 504.600 ;
        RECT 835.950 502.950 838.050 503.400 ;
        RECT 844.950 502.950 847.050 503.400 ;
        RECT 508.950 501.600 511.050 502.050 ;
        RECT 491.400 500.400 511.050 501.600 ;
        RECT 469.950 499.950 472.050 500.400 ;
        RECT 481.950 499.950 484.050 500.400 ;
        RECT 508.950 499.950 511.050 500.400 ;
        RECT 568.950 501.600 571.050 502.050 ;
        RECT 580.950 501.600 583.050 502.050 ;
        RECT 568.950 500.400 583.050 501.600 ;
        RECT 568.950 499.950 571.050 500.400 ;
        RECT 580.950 499.950 583.050 500.400 ;
        RECT 661.950 501.600 664.050 502.050 ;
        RECT 670.950 501.600 673.050 502.050 ;
        RECT 709.950 501.600 712.050 502.050 ;
        RECT 661.950 500.400 712.050 501.600 ;
        RECT 661.950 499.950 664.050 500.400 ;
        RECT 670.950 499.950 673.050 500.400 ;
        RECT 709.950 499.950 712.050 500.400 ;
        RECT 781.950 501.600 784.050 502.050 ;
        RECT 796.950 501.600 799.050 502.050 ;
        RECT 781.950 500.400 799.050 501.600 ;
        RECT 781.950 499.950 784.050 500.400 ;
        RECT 796.950 499.950 799.050 500.400 ;
        RECT 841.950 501.600 844.050 502.050 ;
        RECT 856.950 501.600 859.050 502.050 ;
        RECT 841.950 500.400 859.050 501.600 ;
        RECT 841.950 499.950 844.050 500.400 ;
        RECT 856.950 499.950 859.050 500.400 ;
        RECT 874.950 501.600 877.050 502.050 ;
        RECT 880.950 501.600 883.050 502.050 ;
        RECT 874.950 500.400 883.050 501.600 ;
        RECT 874.950 499.950 877.050 500.400 ;
        RECT 880.950 499.950 883.050 500.400 ;
        RECT 907.950 501.600 910.050 502.050 ;
        RECT 916.950 501.600 919.050 502.050 ;
        RECT 907.950 500.400 919.050 501.600 ;
        RECT 907.950 499.950 910.050 500.400 ;
        RECT 916.950 499.950 919.050 500.400 ;
        RECT 823.950 499.050 826.050 499.200 ;
        RECT 28.950 498.600 31.050 499.050 ;
        RECT 34.950 498.600 37.050 499.050 ;
        RECT 28.950 497.400 37.050 498.600 ;
        RECT 28.950 496.950 31.050 497.400 ;
        RECT 34.950 496.950 37.050 497.400 ;
        RECT 166.950 498.600 169.050 499.050 ;
        RECT 172.950 498.600 175.050 499.050 ;
        RECT 166.950 497.400 175.050 498.600 ;
        RECT 166.950 496.950 169.050 497.400 ;
        RECT 172.950 496.950 175.050 497.400 ;
        RECT 247.950 498.600 250.050 499.050 ;
        RECT 256.950 498.600 259.050 499.050 ;
        RECT 247.950 497.400 259.050 498.600 ;
        RECT 247.950 496.950 250.050 497.400 ;
        RECT 256.950 496.950 259.050 497.400 ;
        RECT 268.950 498.600 271.050 499.050 ;
        RECT 307.950 498.600 312.000 499.050 ;
        RECT 322.950 498.600 325.050 499.050 ;
        RECT 268.950 497.400 285.600 498.600 ;
        RECT 268.950 496.950 271.050 497.400 ;
        RECT 4.950 495.600 7.050 496.050 ;
        RECT 10.950 495.600 13.050 496.200 ;
        RECT 22.950 495.600 25.050 496.050 ;
        RECT 4.950 494.400 13.050 495.600 ;
        RECT 4.950 493.950 7.050 494.400 ;
        RECT 10.950 494.100 13.050 494.400 ;
        RECT 14.400 494.400 25.050 495.600 ;
        RECT 14.400 489.900 15.600 494.400 ;
        RECT 22.950 493.950 25.050 494.400 ;
        RECT 40.950 495.600 43.050 496.200 ;
        RECT 55.950 495.600 58.050 496.200 ;
        RECT 40.950 494.400 58.050 495.600 ;
        RECT 40.950 494.100 43.050 494.400 ;
        RECT 55.950 494.100 58.050 494.400 ;
        RECT 85.950 495.600 88.050 496.200 ;
        RECT 106.950 495.600 109.050 496.200 ;
        RECT 115.950 495.750 118.050 496.200 ;
        RECT 121.950 495.750 124.050 496.200 ;
        RECT 85.950 494.400 114.600 495.600 ;
        RECT 85.950 494.100 88.050 494.400 ;
        RECT 106.950 494.100 109.050 494.400 ;
        RECT 67.950 492.600 70.050 493.050 ;
        RECT 53.400 491.400 70.050 492.600 ;
        RECT 113.400 492.600 114.600 494.400 ;
        RECT 115.950 494.550 124.050 495.750 ;
        RECT 115.950 494.100 118.050 494.550 ;
        RECT 121.950 494.100 124.050 494.550 ;
        RECT 133.950 495.600 136.050 496.050 ;
        RECT 133.950 494.400 153.600 495.600 ;
        RECT 133.950 493.950 136.050 494.400 ;
        RECT 113.400 491.400 117.600 492.600 ;
        RECT 53.400 489.900 54.600 491.400 ;
        RECT 67.950 490.950 70.050 491.400 ;
        RECT 13.950 487.800 16.050 489.900 ;
        RECT 43.950 489.600 46.050 489.900 ;
        RECT 52.950 489.600 55.050 489.900 ;
        RECT 43.950 488.400 55.050 489.600 ;
        RECT 43.950 487.800 46.050 488.400 ;
        RECT 52.950 487.800 55.050 488.400 ;
        RECT 58.950 489.600 61.050 489.900 ;
        RECT 82.950 489.600 85.050 489.900 ;
        RECT 58.950 488.400 85.050 489.600 ;
        RECT 58.950 487.800 61.050 488.400 ;
        RECT 82.950 487.800 85.050 488.400 ;
        RECT 91.950 489.450 94.050 489.900 ;
        RECT 103.950 489.450 106.050 489.900 ;
        RECT 91.950 488.250 106.050 489.450 ;
        RECT 116.400 489.600 117.600 491.400 ;
        RECT 130.950 489.600 133.050 489.900 ;
        RECT 145.950 489.600 148.050 489.900 ;
        RECT 116.400 488.400 148.050 489.600 ;
        RECT 152.400 489.600 153.600 494.400 ;
        RECT 175.950 492.600 178.050 496.050 ;
        RECT 193.950 495.600 196.050 496.200 ;
        RECT 202.950 495.600 205.050 496.050 ;
        RECT 214.950 495.600 217.050 496.200 ;
        RECT 193.950 494.400 205.050 495.600 ;
        RECT 193.950 494.100 196.050 494.400 ;
        RECT 202.950 493.950 205.050 494.400 ;
        RECT 206.400 494.400 217.050 495.600 ;
        RECT 206.400 492.600 207.600 494.400 ;
        RECT 214.950 494.100 217.050 494.400 ;
        RECT 220.950 494.100 223.050 496.200 ;
        RECT 226.950 495.600 229.050 496.050 ;
        RECT 247.950 495.600 250.050 495.900 ;
        RECT 226.950 494.400 250.050 495.600 ;
        RECT 175.950 492.000 183.600 492.600 ;
        RECT 176.400 491.400 184.050 492.000 ;
        RECT 169.950 489.600 172.050 489.900 ;
        RECT 152.400 488.400 172.050 489.600 ;
        RECT 91.950 487.800 94.050 488.250 ;
        RECT 103.950 487.800 106.050 488.250 ;
        RECT 130.950 487.800 133.050 488.400 ;
        RECT 145.950 487.800 148.050 488.400 ;
        RECT 169.950 487.800 172.050 488.400 ;
        RECT 181.950 487.950 184.050 491.400 ;
        RECT 197.400 491.400 207.600 492.600 ;
        RECT 221.400 492.600 222.600 494.100 ;
        RECT 226.950 493.950 229.050 494.400 ;
        RECT 247.950 493.800 250.050 494.400 ;
        RECT 265.950 493.950 268.050 496.050 ;
        RECT 274.950 493.950 277.050 496.050 ;
        RECT 284.400 495.600 285.600 497.400 ;
        RECT 307.950 496.950 312.600 498.600 ;
        RECT 322.950 497.400 336.600 498.600 ;
        RECT 322.950 496.950 325.050 497.400 ;
        RECT 286.950 495.600 289.050 496.200 ;
        RECT 284.400 494.400 289.050 495.600 ;
        RECT 286.950 494.100 289.050 494.400 ;
        RECT 292.950 495.750 295.050 496.200 ;
        RECT 301.950 495.750 304.050 496.200 ;
        RECT 292.950 494.550 304.050 495.750 ;
        RECT 292.950 494.100 295.050 494.550 ;
        RECT 301.950 494.100 304.050 494.550 ;
        RECT 221.400 491.400 240.600 492.600 ;
        RECT 197.400 489.900 198.600 491.400 ;
        RECT 196.950 487.800 199.050 489.900 ;
        RECT 223.950 489.600 226.050 489.900 ;
        RECT 235.950 489.600 238.050 489.900 ;
        RECT 223.950 488.400 238.050 489.600 ;
        RECT 239.400 489.600 240.600 491.400 ;
        RECT 266.400 490.050 267.600 493.950 ;
        RECT 275.400 490.050 276.600 493.950 ;
        RECT 311.400 490.050 312.600 496.950 ;
        RECT 319.950 495.600 322.050 496.200 ;
        RECT 319.950 494.400 327.600 495.600 ;
        RECT 319.950 494.100 322.050 494.400 ;
        RECT 326.400 490.050 327.600 494.400 ;
        RECT 335.400 490.050 336.600 497.400 ;
        RECT 403.950 496.950 406.050 499.050 ;
        RECT 412.950 498.600 415.050 499.050 ;
        RECT 421.950 498.600 424.050 499.050 ;
        RECT 412.950 497.400 424.050 498.600 ;
        RECT 412.950 496.950 415.050 497.400 ;
        RECT 421.950 496.950 424.050 497.400 ;
        RECT 355.950 495.600 358.050 495.900 ;
        RECT 364.950 495.600 367.050 496.200 ;
        RECT 355.950 494.400 367.050 495.600 ;
        RECT 355.950 493.800 358.050 494.400 ;
        RECT 364.950 494.100 367.050 494.400 ;
        RECT 370.950 493.950 373.050 496.050 ;
        RECT 371.400 490.050 372.600 493.950 ;
        RECT 382.950 492.600 385.050 496.050 ;
        RECT 388.950 495.600 391.050 496.200 ;
        RECT 388.950 494.400 402.600 495.600 ;
        RECT 388.950 494.100 391.050 494.400 ;
        RECT 382.950 492.000 387.600 492.600 ;
        RECT 383.400 491.400 387.600 492.000 ;
        RECT 250.950 489.600 253.050 490.050 ;
        RECT 239.400 488.400 253.050 489.600 ;
        RECT 223.950 487.800 226.050 488.400 ;
        RECT 235.950 487.800 238.050 488.400 ;
        RECT 250.950 487.950 253.050 488.400 ;
        RECT 265.950 487.950 268.050 490.050 ;
        RECT 274.950 487.950 277.050 490.050 ;
        RECT 283.950 489.600 286.050 489.900 ;
        RECT 298.950 489.600 301.050 489.900 ;
        RECT 283.950 488.400 301.050 489.600 ;
        RECT 283.950 487.800 286.050 488.400 ;
        RECT 298.950 487.800 301.050 488.400 ;
        RECT 310.950 487.950 313.050 490.050 ;
        RECT 325.950 487.950 328.050 490.050 ;
        RECT 334.950 487.950 337.050 490.050 ;
        RECT 370.950 487.950 373.050 490.050 ;
        RECT 386.400 489.900 387.600 491.400 ;
        RECT 401.400 490.050 402.600 494.400 ;
        RECT 385.950 487.800 388.050 489.900 ;
        RECT 400.950 487.950 403.050 490.050 ;
        RECT 404.400 489.600 405.600 496.950 ;
        RECT 409.950 495.600 412.050 496.050 ;
        RECT 424.950 495.600 427.050 496.200 ;
        RECT 430.950 495.600 433.050 499.050 ;
        RECT 463.950 498.600 466.050 499.050 ;
        RECT 478.950 498.600 481.050 499.050 ;
        RECT 463.950 497.400 481.050 498.600 ;
        RECT 463.950 496.950 466.050 497.400 ;
        RECT 478.950 496.950 481.050 497.400 ;
        RECT 514.950 498.600 517.050 499.050 ;
        RECT 523.950 498.600 526.050 499.050 ;
        RECT 532.950 498.600 535.050 499.050 ;
        RECT 514.950 497.400 535.050 498.600 ;
        RECT 514.950 496.950 517.050 497.400 ;
        RECT 523.950 496.950 526.050 497.400 ;
        RECT 532.950 496.950 535.050 497.400 ;
        RECT 541.950 498.600 544.050 499.050 ;
        RECT 553.950 498.600 556.050 499.050 ;
        RECT 541.950 497.400 556.050 498.600 ;
        RECT 541.950 496.950 544.050 497.400 ;
        RECT 553.950 496.950 556.050 497.400 ;
        RECT 559.950 498.600 562.050 499.050 ;
        RECT 589.950 498.600 592.050 499.050 ;
        RECT 559.950 497.400 592.050 498.600 ;
        RECT 559.950 496.950 562.050 497.400 ;
        RECT 589.950 496.950 592.050 497.400 ;
        RECT 613.950 498.600 616.050 499.050 ;
        RECT 625.950 498.600 628.050 499.050 ;
        RECT 613.950 497.400 628.050 498.600 ;
        RECT 613.950 496.950 616.050 497.400 ;
        RECT 625.950 496.950 628.050 497.400 ;
        RECT 655.950 498.600 658.050 499.050 ;
        RECT 667.950 498.600 670.050 499.050 ;
        RECT 682.950 498.600 685.050 499.050 ;
        RECT 655.950 497.400 685.050 498.600 ;
        RECT 655.950 496.950 658.050 497.400 ;
        RECT 667.950 496.950 670.050 497.400 ;
        RECT 682.950 496.950 685.050 497.400 ;
        RECT 691.950 498.600 694.050 499.050 ;
        RECT 724.950 498.600 727.050 499.050 ;
        RECT 691.950 497.400 727.050 498.600 ;
        RECT 691.950 496.950 694.050 497.400 ;
        RECT 724.950 496.950 727.050 497.400 ;
        RECT 730.950 498.600 733.050 499.050 ;
        RECT 736.950 498.600 739.050 499.050 ;
        RECT 730.950 497.400 739.050 498.600 ;
        RECT 730.950 496.950 733.050 497.400 ;
        RECT 736.950 496.950 739.050 497.400 ;
        RECT 823.950 498.600 828.000 499.050 ;
        RECT 862.950 498.600 865.050 499.050 ;
        RECT 883.950 498.600 886.050 499.050 ;
        RECT 823.950 497.100 828.600 498.600 ;
        RECT 825.000 496.950 828.600 497.100 ;
        RECT 862.950 497.400 886.050 498.600 ;
        RECT 862.950 496.950 865.050 497.400 ;
        RECT 883.950 496.950 886.050 497.400 ;
        RECT 889.800 496.950 891.900 499.050 ;
        RECT 892.950 496.950 895.050 499.050 ;
        RECT 904.950 498.600 909.000 499.050 ;
        RECT 904.950 496.950 909.600 498.600 ;
        RECT 409.950 494.400 420.600 495.600 ;
        RECT 409.950 493.950 412.050 494.400 ;
        RECT 419.400 492.600 420.600 494.400 ;
        RECT 424.950 495.000 433.050 495.600 ;
        RECT 445.950 495.600 448.050 496.200 ;
        RECT 493.950 495.600 496.050 496.200 ;
        RECT 511.950 495.600 514.050 496.200 ;
        RECT 424.950 494.400 432.600 495.000 ;
        RECT 445.950 494.400 471.600 495.600 ;
        RECT 424.950 494.100 427.050 494.400 ;
        RECT 445.950 494.100 448.050 494.400 ;
        RECT 419.400 491.400 423.600 492.600 ;
        RECT 409.950 489.600 412.050 490.050 ;
        RECT 422.400 489.900 423.600 491.400 ;
        RECT 470.400 489.900 471.600 494.400 ;
        RECT 493.950 494.400 514.050 495.600 ;
        RECT 493.950 494.100 496.050 494.400 ;
        RECT 511.950 494.100 514.050 494.400 ;
        RECT 520.950 495.600 523.050 496.050 ;
        RECT 574.950 495.600 577.050 496.200 ;
        RECT 520.950 494.400 552.600 495.600 ;
        RECT 404.400 488.400 412.050 489.600 ;
        RECT 409.950 487.950 412.050 488.400 ;
        RECT 421.950 487.800 424.050 489.900 ;
        RECT 427.950 489.600 430.050 489.900 ;
        RECT 442.950 489.600 445.050 489.900 ;
        RECT 427.950 488.400 445.050 489.600 ;
        RECT 427.950 487.800 430.050 488.400 ;
        RECT 442.950 487.800 445.050 488.400 ;
        RECT 469.950 487.800 472.050 489.900 ;
        RECT 481.950 489.450 484.050 489.900 ;
        RECT 490.950 489.450 493.050 489.900 ;
        RECT 481.950 488.250 493.050 489.450 ;
        RECT 481.950 487.800 484.050 488.250 ;
        RECT 490.950 487.800 493.050 488.250 ;
        RECT 494.400 487.050 495.600 494.100 ;
        RECT 520.950 493.950 523.050 494.400 ;
        RECT 514.950 489.450 517.050 489.900 ;
        RECT 523.950 489.450 526.050 489.900 ;
        RECT 514.950 488.250 526.050 489.450 ;
        RECT 514.950 487.800 517.050 488.250 ;
        RECT 523.950 487.800 526.050 488.250 ;
        RECT 535.950 489.600 538.050 489.900 ;
        RECT 541.950 489.600 544.050 490.050 ;
        RECT 551.400 489.900 552.600 494.400 ;
        RECT 560.400 494.400 577.050 495.600 ;
        RECT 535.950 488.400 544.050 489.600 ;
        RECT 535.950 487.800 538.050 488.400 ;
        RECT 541.950 487.950 544.050 488.400 ;
        RECT 550.950 487.800 553.050 489.900 ;
        RECT 106.950 486.600 109.050 487.050 ;
        RECT 124.950 486.600 127.050 487.050 ;
        RECT 106.950 485.400 127.050 486.600 ;
        RECT 106.950 484.950 109.050 485.400 ;
        RECT 124.950 484.950 127.050 485.400 ;
        RECT 193.950 484.950 199.050 487.050 ;
        RECT 301.950 486.600 304.050 487.050 ;
        RECT 307.950 486.600 310.050 487.050 ;
        RECT 301.950 485.400 310.050 486.600 ;
        RECT 301.950 484.950 304.050 485.400 ;
        RECT 307.950 484.950 310.050 485.400 ;
        RECT 319.950 486.600 322.050 487.050 ;
        RECT 328.950 486.600 331.050 487.050 ;
        RECT 319.950 485.400 331.050 486.600 ;
        RECT 319.950 484.950 322.050 485.400 ;
        RECT 328.950 484.950 331.050 485.400 ;
        RECT 385.950 486.600 388.050 486.750 ;
        RECT 391.950 486.600 394.050 487.050 ;
        RECT 385.950 485.400 394.050 486.600 ;
        RECT 385.950 484.650 388.050 485.400 ;
        RECT 391.950 484.950 394.050 485.400 ;
        RECT 415.950 486.600 418.050 487.050 ;
        RECT 427.950 486.600 430.050 487.050 ;
        RECT 415.950 485.400 430.050 486.600 ;
        RECT 415.950 484.950 418.050 485.400 ;
        RECT 427.950 484.950 430.050 485.400 ;
        RECT 433.950 486.600 436.050 487.050 ;
        RECT 484.950 486.600 487.050 487.050 ;
        RECT 433.950 485.400 487.050 486.600 ;
        RECT 433.950 484.950 436.050 485.400 ;
        RECT 484.950 484.950 487.050 485.400 ;
        RECT 493.950 484.950 496.050 487.050 ;
        RECT 547.950 486.600 550.050 487.050 ;
        RECT 560.400 486.600 561.600 494.400 ;
        RECT 574.950 494.100 577.050 494.400 ;
        RECT 604.950 495.600 607.050 496.200 ;
        RECT 622.950 495.600 625.050 496.200 ;
        RECT 604.950 494.400 625.050 495.600 ;
        RECT 604.950 494.100 607.050 494.400 ;
        RECT 622.950 494.100 625.050 494.400 ;
        RECT 628.950 495.600 631.050 496.200 ;
        RECT 634.800 495.600 636.900 496.050 ;
        RECT 628.950 494.400 636.900 495.600 ;
        RECT 628.950 494.100 631.050 494.400 ;
        RECT 634.800 493.950 636.900 494.400 ;
        RECT 637.950 495.750 640.050 496.200 ;
        RECT 643.950 495.750 646.050 496.200 ;
        RECT 637.950 494.550 646.050 495.750 ;
        RECT 637.950 494.100 640.050 494.550 ;
        RECT 643.950 494.100 646.050 494.550 ;
        RECT 652.950 493.950 655.050 496.050 ;
        RECT 670.950 495.600 673.050 496.200 ;
        RECT 670.950 494.400 675.600 495.600 ;
        RECT 670.950 494.100 673.050 494.400 ;
        RECT 653.400 490.050 654.600 493.950 ;
        RECT 565.950 489.450 568.050 489.900 ;
        RECT 577.950 489.450 580.050 489.900 ;
        RECT 565.950 488.250 580.050 489.450 ;
        RECT 565.950 487.800 568.050 488.250 ;
        RECT 577.950 487.800 580.050 488.250 ;
        RECT 583.950 489.450 586.050 489.900 ;
        RECT 589.950 489.600 592.050 489.900 ;
        RECT 601.950 489.600 604.050 489.900 ;
        RECT 589.950 489.450 604.050 489.600 ;
        RECT 583.950 488.400 604.050 489.450 ;
        RECT 583.950 488.250 592.050 488.400 ;
        RECT 583.950 487.800 586.050 488.250 ;
        RECT 589.950 487.800 592.050 488.250 ;
        RECT 601.950 487.800 604.050 488.400 ;
        RECT 616.950 489.450 619.050 489.900 ;
        RECT 625.950 489.450 628.050 489.900 ;
        RECT 616.950 488.250 628.050 489.450 ;
        RECT 616.950 487.800 619.050 488.250 ;
        RECT 625.950 487.800 628.050 488.250 ;
        RECT 637.950 489.600 640.050 490.050 ;
        RECT 646.950 489.600 649.050 490.050 ;
        RECT 637.950 488.400 649.050 489.600 ;
        RECT 637.950 487.950 640.050 488.400 ;
        RECT 646.950 487.950 649.050 488.400 ;
        RECT 652.950 487.950 655.050 490.050 ;
        RECT 674.400 489.600 675.600 494.400 ;
        RECT 685.950 494.100 688.050 496.200 ;
        RECT 721.950 495.600 724.050 496.050 ;
        RECT 745.950 495.600 748.050 496.050 ;
        RECT 796.950 495.600 799.050 496.200 ;
        RECT 721.950 494.400 748.050 495.600 ;
        RECT 682.950 489.600 685.050 490.050 ;
        RECT 674.400 488.400 685.050 489.600 ;
        RECT 682.950 487.950 685.050 488.400 ;
        RECT 547.950 485.400 561.600 486.600 ;
        RECT 577.950 486.600 580.050 487.050 ;
        RECT 595.950 486.600 598.050 487.050 ;
        RECT 577.950 485.400 598.050 486.600 ;
        RECT 547.950 484.950 550.050 485.400 ;
        RECT 577.950 484.950 580.050 485.400 ;
        RECT 595.950 484.950 598.050 485.400 ;
        RECT 649.950 486.600 652.050 487.050 ;
        RECT 658.950 486.600 661.050 487.050 ;
        RECT 649.950 485.400 661.050 486.600 ;
        RECT 649.950 484.950 652.050 485.400 ;
        RECT 658.950 484.950 661.050 485.400 ;
        RECT 664.950 486.600 667.050 487.050 ;
        RECT 686.400 486.600 687.600 494.100 ;
        RECT 721.950 493.950 724.050 494.400 ;
        RECT 745.950 493.950 748.050 494.400 ;
        RECT 776.400 494.400 799.050 495.600 ;
        RECT 776.400 492.600 777.600 494.400 ;
        RECT 796.950 494.100 799.050 494.400 ;
        RECT 814.950 495.600 817.050 496.050 ;
        RECT 823.950 495.600 826.050 496.050 ;
        RECT 814.950 494.400 826.050 495.600 ;
        RECT 814.950 493.950 817.050 494.400 ;
        RECT 823.950 493.950 826.050 494.400 ;
        RECT 746.400 491.400 777.600 492.600 ;
        RECT 688.950 489.600 691.050 489.900 ;
        RECT 712.950 489.600 715.050 489.900 ;
        RECT 739.950 489.600 742.050 489.900 ;
        RECT 688.950 488.400 742.050 489.600 ;
        RECT 688.950 487.800 691.050 488.400 ;
        RECT 712.950 487.800 715.050 488.400 ;
        RECT 739.950 487.800 742.050 488.400 ;
        RECT 746.400 487.050 747.600 491.400 ;
        RECT 751.950 489.600 754.050 490.050 ;
        RECT 827.400 489.900 828.600 496.950 ;
        RECT 835.950 493.950 838.050 496.050 ;
        RECT 868.950 493.950 871.050 496.050 ;
        RECT 836.400 490.050 837.600 493.950 ;
        RECT 869.400 490.050 870.600 493.950 ;
        RECT 802.950 489.600 805.050 489.900 ;
        RECT 820.950 489.600 823.050 489.900 ;
        RECT 751.950 488.400 823.050 489.600 ;
        RECT 751.950 487.950 754.050 488.400 ;
        RECT 802.950 487.800 805.050 488.400 ;
        RECT 820.950 487.800 823.050 488.400 ;
        RECT 826.950 487.800 829.050 489.900 ;
        RECT 835.950 487.950 838.050 490.050 ;
        RECT 868.950 487.950 871.050 490.050 ;
        RECT 890.400 487.050 891.600 496.950 ;
        RECT 893.400 490.050 894.600 496.950 ;
        RECT 901.950 493.950 904.050 496.050 ;
        RECT 902.400 490.050 903.600 493.950 ;
        RECT 892.950 487.950 895.050 490.050 ;
        RECT 901.950 487.950 904.050 490.050 ;
        RECT 908.400 487.050 909.600 496.950 ;
        RECT 664.950 485.400 687.600 486.600 ;
        RECT 664.950 484.950 667.050 485.400 ;
        RECT 745.950 484.950 748.050 487.050 ;
        RECT 871.950 486.600 874.050 487.050 ;
        RECT 880.950 486.600 883.050 487.050 ;
        RECT 871.950 485.400 883.050 486.600 ;
        RECT 871.950 484.950 874.050 485.400 ;
        RECT 880.950 484.950 883.050 485.400 ;
        RECT 889.950 484.950 892.050 487.050 ;
        RECT 904.950 486.600 909.600 487.050 ;
        RECT 913.950 486.600 916.050 487.050 ;
        RECT 904.950 485.400 916.050 486.600 ;
        RECT 904.950 484.950 909.000 485.400 ;
        RECT 913.950 484.950 916.050 485.400 ;
        RECT 19.950 483.600 22.050 484.050 ;
        RECT 28.950 483.600 31.050 484.050 ;
        RECT 37.950 483.600 40.050 484.050 ;
        RECT 19.950 482.400 40.050 483.600 ;
        RECT 19.950 481.950 22.050 482.400 ;
        RECT 28.950 481.950 31.050 482.400 ;
        RECT 37.950 481.950 40.050 482.400 ;
        RECT 88.950 483.600 91.050 484.050 ;
        RECT 157.950 483.600 160.050 484.050 ;
        RECT 178.950 483.600 181.050 484.050 ;
        RECT 88.950 482.400 141.600 483.600 ;
        RECT 88.950 481.950 91.050 482.400 ;
        RECT 124.950 480.600 127.050 481.050 ;
        RECT 136.950 480.600 139.050 481.050 ;
        RECT 124.950 479.400 139.050 480.600 ;
        RECT 140.400 480.600 141.600 482.400 ;
        RECT 157.950 482.400 181.050 483.600 ;
        RECT 157.950 481.950 160.050 482.400 ;
        RECT 178.950 481.950 181.050 482.400 ;
        RECT 256.950 483.600 259.050 484.050 ;
        RECT 310.950 483.600 313.050 484.050 ;
        RECT 256.950 482.400 313.050 483.600 ;
        RECT 256.950 481.950 259.050 482.400 ;
        RECT 310.950 481.950 313.050 482.400 ;
        RECT 358.950 483.600 361.050 484.050 ;
        RECT 364.950 483.600 367.050 484.050 ;
        RECT 358.950 482.400 367.050 483.600 ;
        RECT 358.950 481.950 361.050 482.400 ;
        RECT 364.950 481.950 367.050 482.400 ;
        RECT 406.950 483.600 409.050 484.050 ;
        RECT 430.950 483.600 433.050 484.050 ;
        RECT 406.950 482.400 433.050 483.600 ;
        RECT 406.950 481.950 409.050 482.400 ;
        RECT 430.950 481.950 433.050 482.400 ;
        RECT 439.950 483.600 442.050 484.050 ;
        RECT 451.950 483.600 454.050 484.050 ;
        RECT 463.950 483.600 466.050 484.050 ;
        RECT 439.950 482.400 466.050 483.600 ;
        RECT 439.950 481.950 442.050 482.400 ;
        RECT 451.950 481.950 454.050 482.400 ;
        RECT 463.950 481.950 466.050 482.400 ;
        RECT 526.950 483.600 529.050 484.050 ;
        RECT 574.950 483.600 577.050 484.050 ;
        RECT 526.950 482.400 577.050 483.600 ;
        RECT 526.950 481.950 529.050 482.400 ;
        RECT 574.950 481.950 577.050 482.400 ;
        RECT 598.950 483.600 601.050 484.050 ;
        RECT 616.950 483.600 619.050 484.050 ;
        RECT 598.950 482.400 619.050 483.600 ;
        RECT 598.950 481.950 601.050 482.400 ;
        RECT 616.950 481.950 619.050 482.400 ;
        RECT 622.950 483.600 625.050 484.050 ;
        RECT 655.950 483.600 658.050 484.050 ;
        RECT 622.950 482.400 658.050 483.600 ;
        RECT 622.950 481.950 625.050 482.400 ;
        RECT 655.950 481.950 658.050 482.400 ;
        RECT 682.950 483.600 685.050 484.050 ;
        RECT 694.950 483.600 697.050 484.050 ;
        RECT 682.950 482.400 697.050 483.600 ;
        RECT 682.950 481.950 685.050 482.400 ;
        RECT 694.950 481.950 697.050 482.400 ;
        RECT 703.950 483.600 706.050 484.050 ;
        RECT 715.950 483.600 718.050 484.050 ;
        RECT 703.950 482.400 718.050 483.600 ;
        RECT 703.950 481.950 706.050 482.400 ;
        RECT 715.950 481.950 718.050 482.400 ;
        RECT 748.950 483.600 751.050 484.050 ;
        RECT 754.950 483.600 757.050 484.050 ;
        RECT 748.950 482.400 757.050 483.600 ;
        RECT 748.950 481.950 751.050 482.400 ;
        RECT 754.950 481.950 757.050 482.400 ;
        RECT 784.950 483.600 787.050 484.050 ;
        RECT 790.950 483.600 793.050 484.050 ;
        RECT 784.950 482.400 793.050 483.600 ;
        RECT 784.950 481.950 787.050 482.400 ;
        RECT 790.950 481.950 793.050 482.400 ;
        RECT 805.950 483.600 808.050 484.050 ;
        RECT 844.950 483.600 847.050 484.050 ;
        RECT 805.950 482.400 847.050 483.600 ;
        RECT 805.950 481.950 808.050 482.400 ;
        RECT 844.950 481.950 847.050 482.400 ;
        RECT 883.950 483.600 886.050 484.050 ;
        RECT 898.950 483.600 901.050 484.050 ;
        RECT 883.950 482.400 901.050 483.600 ;
        RECT 883.950 481.950 886.050 482.400 ;
        RECT 898.950 481.950 901.050 482.400 ;
        RECT 187.950 480.600 190.050 481.050 ;
        RECT 140.400 479.400 190.050 480.600 ;
        RECT 124.950 478.950 127.050 479.400 ;
        RECT 136.950 478.950 139.050 479.400 ;
        RECT 187.950 478.950 190.050 479.400 ;
        RECT 223.950 480.600 226.050 481.050 ;
        RECT 247.950 480.600 250.050 481.050 ;
        RECT 223.950 479.400 250.050 480.600 ;
        RECT 223.950 478.950 226.050 479.400 ;
        RECT 247.950 478.950 250.050 479.400 ;
        RECT 259.950 480.600 262.050 481.050 ;
        RECT 268.950 480.600 271.050 481.050 ;
        RECT 307.950 480.600 310.050 481.050 ;
        RECT 259.950 479.400 310.050 480.600 ;
        RECT 259.950 478.950 262.050 479.400 ;
        RECT 268.950 478.950 271.050 479.400 ;
        RECT 307.950 478.950 310.050 479.400 ;
        RECT 316.950 480.600 319.050 481.050 ;
        RECT 334.950 480.600 337.050 481.050 ;
        RECT 316.950 479.400 337.050 480.600 ;
        RECT 316.950 478.950 319.050 479.400 ;
        RECT 334.950 478.950 337.050 479.400 ;
        RECT 340.950 480.600 343.050 481.050 ;
        RECT 346.950 480.600 349.050 481.050 ;
        RECT 340.950 479.400 349.050 480.600 ;
        RECT 340.950 478.950 343.050 479.400 ;
        RECT 346.950 478.950 349.050 479.400 ;
        RECT 403.950 480.600 406.050 481.050 ;
        RECT 427.950 480.600 430.050 481.050 ;
        RECT 403.950 479.400 430.050 480.600 ;
        RECT 403.950 478.950 406.050 479.400 ;
        RECT 427.950 478.950 430.050 479.400 ;
        RECT 454.950 480.600 457.050 481.050 ;
        RECT 490.950 480.600 493.050 481.050 ;
        RECT 454.950 479.400 493.050 480.600 ;
        RECT 454.950 478.950 457.050 479.400 ;
        RECT 490.950 478.950 493.050 479.400 ;
        RECT 700.950 480.600 703.050 481.050 ;
        RECT 712.950 480.600 715.050 481.050 ;
        RECT 700.950 479.400 715.050 480.600 ;
        RECT 700.950 478.950 703.050 479.400 ;
        RECT 712.950 478.950 715.050 479.400 ;
        RECT 769.950 480.600 772.050 481.050 ;
        RECT 838.950 480.600 841.050 481.050 ;
        RECT 769.950 479.400 841.050 480.600 ;
        RECT 769.950 478.950 772.050 479.400 ;
        RECT 838.950 478.950 841.050 479.400 ;
        RECT 886.950 480.600 889.050 481.050 ;
        RECT 916.950 480.600 919.050 481.050 ;
        RECT 886.950 479.400 919.050 480.600 ;
        RECT 886.950 478.950 889.050 479.400 ;
        RECT 916.950 478.950 919.050 479.400 ;
        RECT 70.950 477.600 73.050 478.050 ;
        RECT 106.950 477.600 109.050 478.050 ;
        RECT 70.950 476.400 109.050 477.600 ;
        RECT 70.950 475.950 73.050 476.400 ;
        RECT 106.950 475.950 109.050 476.400 ;
        RECT 250.950 477.600 253.050 478.050 ;
        RECT 325.950 477.600 328.050 478.050 ;
        RECT 250.950 476.400 328.050 477.600 ;
        RECT 250.950 475.950 253.050 476.400 ;
        RECT 325.950 475.950 328.050 476.400 ;
        RECT 346.950 477.600 349.050 477.900 ;
        RECT 352.950 477.600 355.050 478.050 ;
        RECT 346.950 476.400 355.050 477.600 ;
        RECT 346.950 475.800 349.050 476.400 ;
        RECT 352.950 475.950 355.050 476.400 ;
        RECT 376.950 477.600 379.050 478.050 ;
        RECT 433.950 477.600 436.050 478.050 ;
        RECT 376.950 476.400 436.050 477.600 ;
        RECT 376.950 475.950 379.050 476.400 ;
        RECT 433.950 475.950 436.050 476.400 ;
        RECT 469.950 477.600 472.050 478.050 ;
        RECT 487.950 477.600 490.050 478.050 ;
        RECT 469.950 476.400 490.050 477.600 ;
        RECT 469.950 475.950 472.050 476.400 ;
        RECT 487.950 475.950 490.050 476.400 ;
        RECT 574.950 477.600 577.050 478.050 ;
        RECT 610.950 477.600 613.050 478.050 ;
        RECT 574.950 476.400 613.050 477.600 ;
        RECT 574.950 475.950 577.050 476.400 ;
        RECT 610.950 475.950 613.050 476.400 ;
        RECT 631.950 477.600 634.050 478.050 ;
        RECT 730.950 477.600 733.050 478.050 ;
        RECT 631.950 476.400 733.050 477.600 ;
        RECT 631.950 475.950 634.050 476.400 ;
        RECT 730.950 475.950 733.050 476.400 ;
        RECT 742.950 477.600 745.050 478.050 ;
        RECT 778.950 477.600 781.050 478.050 ;
        RECT 742.950 476.400 781.050 477.600 ;
        RECT 742.950 475.950 745.050 476.400 ;
        RECT 778.950 475.950 781.050 476.400 ;
        RECT 814.950 477.600 817.050 478.050 ;
        RECT 832.950 477.600 835.050 478.050 ;
        RECT 814.950 476.400 835.050 477.600 ;
        RECT 814.950 475.950 817.050 476.400 ;
        RECT 832.950 475.950 835.050 476.400 ;
        RECT 847.950 477.600 850.050 478.050 ;
        RECT 868.950 477.600 871.050 478.050 ;
        RECT 880.950 477.600 883.050 478.050 ;
        RECT 847.950 476.400 883.050 477.600 ;
        RECT 847.950 475.950 850.050 476.400 ;
        RECT 868.950 475.950 871.050 476.400 ;
        RECT 880.950 475.950 883.050 476.400 ;
        RECT 46.950 474.600 49.050 475.050 ;
        RECT 64.950 474.600 67.050 475.050 ;
        RECT 115.950 474.600 118.050 475.050 ;
        RECT 202.950 474.600 205.050 475.050 ;
        RECT 46.950 473.400 205.050 474.600 ;
        RECT 46.950 472.950 49.050 473.400 ;
        RECT 64.950 472.950 67.050 473.400 ;
        RECT 115.950 472.950 118.050 473.400 ;
        RECT 202.950 472.950 205.050 473.400 ;
        RECT 301.950 474.600 304.050 475.050 ;
        RECT 322.950 474.600 325.050 475.050 ;
        RECT 337.950 474.600 340.050 475.050 ;
        RECT 301.950 473.400 340.050 474.600 ;
        RECT 301.950 472.950 304.050 473.400 ;
        RECT 322.950 472.950 325.050 473.400 ;
        RECT 337.950 472.950 340.050 473.400 ;
        RECT 388.950 474.600 391.050 475.050 ;
        RECT 415.950 474.600 418.050 475.050 ;
        RECT 421.950 474.600 424.050 475.050 ;
        RECT 388.950 473.400 424.050 474.600 ;
        RECT 388.950 472.950 391.050 473.400 ;
        RECT 415.950 472.950 418.050 473.400 ;
        RECT 421.950 472.950 424.050 473.400 ;
        RECT 439.950 474.600 442.050 475.050 ;
        RECT 496.950 474.600 499.050 475.050 ;
        RECT 508.950 474.600 511.050 475.050 ;
        RECT 439.950 473.400 511.050 474.600 ;
        RECT 439.950 472.950 442.050 473.400 ;
        RECT 496.950 472.950 499.050 473.400 ;
        RECT 508.950 472.950 511.050 473.400 ;
        RECT 616.950 474.600 619.050 475.050 ;
        RECT 733.950 474.600 736.050 475.050 ;
        RECT 616.950 473.400 736.050 474.600 ;
        RECT 616.950 472.950 619.050 473.400 ;
        RECT 733.950 472.950 736.050 473.400 ;
        RECT 739.950 474.600 742.050 475.050 ;
        RECT 763.950 474.600 766.050 475.050 ;
        RECT 739.950 473.400 766.050 474.600 ;
        RECT 739.950 472.950 742.050 473.400 ;
        RECT 763.950 472.950 766.050 473.400 ;
        RECT 799.950 474.600 802.050 475.050 ;
        RECT 862.950 474.600 865.050 475.050 ;
        RECT 799.950 473.400 865.050 474.600 ;
        RECT 799.950 472.950 802.050 473.400 ;
        RECT 862.950 472.950 865.050 473.400 ;
        RECT 898.950 474.600 901.050 475.050 ;
        RECT 910.950 474.600 913.050 475.050 ;
        RECT 916.950 474.600 919.050 475.050 ;
        RECT 898.950 473.400 919.050 474.600 ;
        RECT 898.950 472.950 901.050 473.400 ;
        RECT 910.950 472.950 913.050 473.400 ;
        RECT 916.950 472.950 919.050 473.400 ;
        RECT 211.950 471.600 214.050 472.050 ;
        RECT 244.950 471.600 247.050 472.050 ;
        RECT 211.950 470.400 247.050 471.600 ;
        RECT 211.950 469.950 214.050 470.400 ;
        RECT 244.950 469.950 247.050 470.400 ;
        RECT 253.950 471.600 256.050 472.050 ;
        RECT 277.950 471.600 280.050 472.050 ;
        RECT 355.950 471.600 358.050 472.050 ;
        RECT 253.950 470.400 358.050 471.600 ;
        RECT 253.950 469.950 256.050 470.400 ;
        RECT 277.950 469.950 280.050 470.400 ;
        RECT 355.950 469.950 358.050 470.400 ;
        RECT 367.950 471.600 370.050 472.050 ;
        RECT 454.950 471.600 457.050 472.050 ;
        RECT 367.950 470.400 457.050 471.600 ;
        RECT 367.950 469.950 370.050 470.400 ;
        RECT 454.950 469.950 457.050 470.400 ;
        RECT 460.950 471.600 463.050 472.050 ;
        RECT 574.950 471.600 577.050 472.050 ;
        RECT 460.950 470.400 577.050 471.600 ;
        RECT 460.950 469.950 463.050 470.400 ;
        RECT 574.950 469.950 577.050 470.400 ;
        RECT 652.950 471.600 655.050 472.050 ;
        RECT 676.950 471.600 679.050 472.050 ;
        RECT 652.950 470.400 679.050 471.600 ;
        RECT 652.950 469.950 655.050 470.400 ;
        RECT 676.950 469.950 679.050 470.400 ;
        RECT 802.950 471.600 805.050 472.050 ;
        RECT 835.950 471.600 838.050 472.050 ;
        RECT 802.950 470.400 838.050 471.600 ;
        RECT 802.950 469.950 805.050 470.400 ;
        RECT 835.950 469.950 838.050 470.400 ;
        RECT 25.950 468.600 28.050 469.050 ;
        RECT 58.950 468.600 61.050 469.050 ;
        RECT 25.950 467.400 61.050 468.600 ;
        RECT 25.950 466.950 28.050 467.400 ;
        RECT 58.950 466.950 61.050 467.400 ;
        RECT 142.950 468.600 145.050 469.050 ;
        RECT 151.950 468.600 154.050 469.050 ;
        RECT 142.950 467.400 154.050 468.600 ;
        RECT 142.950 466.950 145.050 467.400 ;
        RECT 151.950 466.950 154.050 467.400 ;
        RECT 217.950 468.600 220.050 469.050 ;
        RECT 256.950 468.600 259.050 469.050 ;
        RECT 217.950 467.400 259.050 468.600 ;
        RECT 217.950 466.950 220.050 467.400 ;
        RECT 256.950 466.950 259.050 467.400 ;
        RECT 292.950 468.600 295.050 469.050 ;
        RECT 331.950 468.600 334.050 469.050 ;
        RECT 292.950 467.400 334.050 468.600 ;
        RECT 292.950 466.950 295.050 467.400 ;
        RECT 331.950 466.950 334.050 467.400 ;
        RECT 385.950 468.600 388.050 469.050 ;
        RECT 394.950 468.600 397.050 469.050 ;
        RECT 385.950 467.400 397.050 468.600 ;
        RECT 385.950 466.950 388.050 467.400 ;
        RECT 394.950 466.950 397.050 467.400 ;
        RECT 400.950 468.600 403.050 469.050 ;
        RECT 424.950 468.600 427.050 469.050 ;
        RECT 400.950 467.400 427.050 468.600 ;
        RECT 400.950 466.950 403.050 467.400 ;
        RECT 424.950 466.950 427.050 467.400 ;
        RECT 430.950 468.600 433.050 469.050 ;
        RECT 457.950 468.600 460.050 469.050 ;
        RECT 430.950 467.400 460.050 468.600 ;
        RECT 430.950 466.950 433.050 467.400 ;
        RECT 457.950 466.950 460.050 467.400 ;
        RECT 487.950 468.600 490.050 469.050 ;
        RECT 556.950 468.600 559.050 469.050 ;
        RECT 487.950 467.400 559.050 468.600 ;
        RECT 487.950 466.950 490.050 467.400 ;
        RECT 556.950 466.950 559.050 467.400 ;
        RECT 607.950 468.600 610.050 469.050 ;
        RECT 661.950 468.600 664.050 469.050 ;
        RECT 607.950 467.400 664.050 468.600 ;
        RECT 607.950 466.950 610.050 467.400 ;
        RECT 661.950 466.950 664.050 467.400 ;
        RECT 673.950 468.600 676.050 469.050 ;
        RECT 718.950 468.600 721.050 469.050 ;
        RECT 673.950 467.400 721.050 468.600 ;
        RECT 673.950 466.950 676.050 467.400 ;
        RECT 718.950 466.950 721.050 467.400 ;
        RECT 736.950 468.600 739.050 469.050 ;
        RECT 757.950 468.600 760.050 469.050 ;
        RECT 736.950 467.400 760.050 468.600 ;
        RECT 736.950 466.950 739.050 467.400 ;
        RECT 757.950 466.950 760.050 467.400 ;
        RECT 877.950 468.600 880.050 469.050 ;
        RECT 883.950 468.600 886.050 469.050 ;
        RECT 877.950 467.400 886.050 468.600 ;
        RECT 877.950 466.950 880.050 467.400 ;
        RECT 883.950 466.950 886.050 467.400 ;
        RECT 250.950 465.600 253.050 466.050 ;
        RECT 277.950 465.600 280.050 466.050 ;
        RECT 286.950 465.600 289.050 466.050 ;
        RECT 250.950 464.400 276.600 465.600 ;
        RECT 250.950 463.950 253.050 464.400 ;
        RECT 118.950 462.600 121.050 463.050 ;
        RECT 151.950 462.600 154.050 463.050 ;
        RECT 118.950 461.400 154.050 462.600 ;
        RECT 118.950 460.950 121.050 461.400 ;
        RECT 151.950 460.950 154.050 461.400 ;
        RECT 241.950 462.600 244.050 463.050 ;
        RECT 262.950 462.600 265.050 463.050 ;
        RECT 241.950 461.400 265.050 462.600 ;
        RECT 275.400 462.600 276.600 464.400 ;
        RECT 277.950 464.400 289.050 465.600 ;
        RECT 277.950 463.950 280.050 464.400 ;
        RECT 286.950 463.950 289.050 464.400 ;
        RECT 319.950 465.600 322.050 466.050 ;
        RECT 346.950 465.600 349.050 466.050 ;
        RECT 319.950 464.400 349.050 465.600 ;
        RECT 319.950 463.950 322.050 464.400 ;
        RECT 346.950 463.950 349.050 464.400 ;
        RECT 361.950 465.600 364.050 466.050 ;
        RECT 370.950 465.600 373.050 466.050 ;
        RECT 361.950 464.400 373.050 465.600 ;
        RECT 361.950 463.950 364.050 464.400 ;
        RECT 370.950 463.950 373.050 464.400 ;
        RECT 412.950 465.600 415.050 466.050 ;
        RECT 469.950 465.600 472.050 466.050 ;
        RECT 412.950 464.400 472.050 465.600 ;
        RECT 412.950 463.950 415.050 464.400 ;
        RECT 469.950 463.950 472.050 464.400 ;
        RECT 475.950 465.600 478.050 466.050 ;
        RECT 538.950 465.600 541.050 466.050 ;
        RECT 475.950 464.400 541.050 465.600 ;
        RECT 475.950 463.950 478.050 464.400 ;
        RECT 538.950 463.950 541.050 464.400 ;
        RECT 568.950 465.600 571.050 466.050 ;
        RECT 601.950 465.600 604.050 466.050 ;
        RECT 631.950 465.600 634.050 466.050 ;
        RECT 568.950 464.400 634.050 465.600 ;
        RECT 568.950 463.950 571.050 464.400 ;
        RECT 601.950 463.950 604.050 464.400 ;
        RECT 631.950 463.950 634.050 464.400 ;
        RECT 727.950 465.600 730.050 466.050 ;
        RECT 760.950 465.600 763.050 466.050 ;
        RECT 727.950 464.400 763.050 465.600 ;
        RECT 727.950 463.950 730.050 464.400 ;
        RECT 760.950 463.950 763.050 464.400 ;
        RECT 766.950 465.600 769.050 466.050 ;
        RECT 832.950 465.600 835.050 466.050 ;
        RECT 766.950 464.400 835.050 465.600 ;
        RECT 766.950 463.950 769.050 464.400 ;
        RECT 832.950 463.950 835.050 464.400 ;
        RECT 862.950 465.600 865.050 466.050 ;
        RECT 883.950 465.600 886.050 465.900 ;
        RECT 862.950 464.400 886.050 465.600 ;
        RECT 862.950 463.950 865.050 464.400 ;
        RECT 883.950 463.800 886.050 464.400 ;
        RECT 328.950 462.600 331.050 463.050 ;
        RECT 275.400 461.400 331.050 462.600 ;
        RECT 241.950 460.950 244.050 461.400 ;
        RECT 262.950 460.950 265.050 461.400 ;
        RECT 328.950 460.950 331.050 461.400 ;
        RECT 424.950 462.600 427.050 463.050 ;
        RECT 448.950 462.600 451.050 463.050 ;
        RECT 424.950 461.400 451.050 462.600 ;
        RECT 424.950 460.950 427.050 461.400 ;
        RECT 448.950 460.950 451.050 461.400 ;
        RECT 571.950 462.600 574.050 463.050 ;
        RECT 619.950 462.600 622.050 463.050 ;
        RECT 571.950 461.400 622.050 462.600 ;
        RECT 571.950 460.950 574.050 461.400 ;
        RECT 619.950 460.950 622.050 461.400 ;
        RECT 646.950 462.600 649.050 463.050 ;
        RECT 697.950 462.600 700.050 463.050 ;
        RECT 745.950 462.600 748.050 463.050 ;
        RECT 646.950 461.400 748.050 462.600 ;
        RECT 646.950 460.950 649.050 461.400 ;
        RECT 697.950 460.950 700.050 461.400 ;
        RECT 745.950 460.950 748.050 461.400 ;
        RECT 73.950 459.600 76.050 460.050 ;
        RECT 112.950 459.600 115.050 460.050 ;
        RECT 73.950 458.400 115.050 459.600 ;
        RECT 73.950 457.950 76.050 458.400 ;
        RECT 112.950 457.950 115.050 458.400 ;
        RECT 205.950 459.600 208.050 460.050 ;
        RECT 250.800 459.600 252.900 460.050 ;
        RECT 205.950 458.400 252.900 459.600 ;
        RECT 205.950 457.950 208.050 458.400 ;
        RECT 250.800 457.950 252.900 458.400 ;
        RECT 253.950 459.600 256.050 460.050 ;
        RECT 265.950 459.600 268.050 460.050 ;
        RECT 253.950 458.400 268.050 459.600 ;
        RECT 253.950 457.950 256.050 458.400 ;
        RECT 265.950 457.950 268.050 458.400 ;
        RECT 310.950 459.600 313.050 460.050 ;
        RECT 340.950 459.600 343.050 460.050 ;
        RECT 310.950 458.400 343.050 459.600 ;
        RECT 310.950 457.950 313.050 458.400 ;
        RECT 340.950 457.950 343.050 458.400 ;
        RECT 358.950 459.600 361.050 460.050 ;
        RECT 394.950 459.600 397.050 460.050 ;
        RECT 358.950 458.400 397.050 459.600 ;
        RECT 358.950 457.950 361.050 458.400 ;
        RECT 394.950 457.950 397.050 458.400 ;
        RECT 436.950 459.600 439.050 460.050 ;
        RECT 454.950 459.600 457.050 460.050 ;
        RECT 436.950 458.400 457.050 459.600 ;
        RECT 436.950 457.950 439.050 458.400 ;
        RECT 454.950 457.950 457.050 458.400 ;
        RECT 484.950 459.600 487.050 460.050 ;
        RECT 529.950 459.600 532.050 460.050 ;
        RECT 484.950 458.400 532.050 459.600 ;
        RECT 484.950 457.950 487.050 458.400 ;
        RECT 529.950 457.950 532.050 458.400 ;
        RECT 598.950 459.600 601.050 460.050 ;
        RECT 625.950 459.600 628.050 460.050 ;
        RECT 598.950 458.400 628.050 459.600 ;
        RECT 598.950 457.950 601.050 458.400 ;
        RECT 625.950 457.950 628.050 458.400 ;
        RECT 643.950 459.600 646.050 460.050 ;
        RECT 658.950 459.600 661.050 460.050 ;
        RECT 643.950 458.400 661.050 459.600 ;
        RECT 643.950 457.950 646.050 458.400 ;
        RECT 658.950 457.950 661.050 458.400 ;
        RECT 757.950 459.600 760.050 460.050 ;
        RECT 826.950 459.600 829.050 460.050 ;
        RECT 757.950 458.400 829.050 459.600 ;
        RECT 757.950 457.950 760.050 458.400 ;
        RECT 826.950 457.950 829.050 458.400 ;
        RECT 832.950 459.600 835.050 460.050 ;
        RECT 868.950 459.600 871.050 460.050 ;
        RECT 832.950 458.400 871.050 459.600 ;
        RECT 832.950 457.950 835.050 458.400 ;
        RECT 868.950 457.950 871.050 458.400 ;
        RECT 889.950 459.600 892.050 460.050 ;
        RECT 904.950 459.600 907.050 460.050 ;
        RECT 889.950 458.400 907.050 459.600 ;
        RECT 889.950 457.950 892.050 458.400 ;
        RECT 904.950 457.950 907.050 458.400 ;
        RECT 919.950 459.600 924.000 460.050 ;
        RECT 919.950 457.950 924.600 459.600 ;
        RECT 113.400 456.600 114.600 457.950 ;
        RECT 136.950 456.600 139.050 457.050 ;
        RECT 241.950 456.600 244.050 457.050 ;
        RECT 113.400 455.400 139.050 456.600 ;
        RECT 136.950 454.950 139.050 455.400 ;
        RECT 200.400 455.400 244.050 456.600 ;
        RECT 52.950 453.600 55.050 454.050 ;
        RECT 88.950 453.600 91.050 454.050 ;
        RECT 106.950 453.600 109.050 454.050 ;
        RECT 52.950 452.400 109.050 453.600 ;
        RECT 52.950 451.950 55.050 452.400 ;
        RECT 88.950 451.950 91.050 452.400 ;
        RECT 106.950 451.950 109.050 452.400 ;
        RECT 163.950 453.600 166.050 454.050 ;
        RECT 200.400 453.600 201.600 455.400 ;
        RECT 241.950 454.950 244.050 455.400 ;
        RECT 283.950 456.600 286.050 457.050 ;
        RECT 289.950 456.600 292.050 457.050 ;
        RECT 298.950 456.600 301.050 457.050 ;
        RECT 283.950 455.400 301.050 456.600 ;
        RECT 283.950 454.950 286.050 455.400 ;
        RECT 289.950 454.950 292.050 455.400 ;
        RECT 298.950 454.950 301.050 455.400 ;
        RECT 304.950 456.600 307.050 457.050 ;
        RECT 325.950 456.600 328.050 457.050 ;
        RECT 343.950 456.600 346.050 457.050 ;
        RECT 304.950 455.400 346.050 456.600 ;
        RECT 304.950 454.950 307.050 455.400 ;
        RECT 325.950 454.950 328.050 455.400 ;
        RECT 343.950 454.950 346.050 455.400 ;
        RECT 370.950 456.600 373.050 457.050 ;
        RECT 403.950 456.600 406.050 457.050 ;
        RECT 370.950 455.400 406.050 456.600 ;
        RECT 370.950 454.950 373.050 455.400 ;
        RECT 403.950 454.950 406.050 455.400 ;
        RECT 433.950 456.600 436.050 457.050 ;
        RECT 475.800 456.600 477.900 457.050 ;
        RECT 433.950 455.400 477.900 456.600 ;
        RECT 433.950 454.950 436.050 455.400 ;
        RECT 475.800 454.950 477.900 455.400 ;
        RECT 478.950 456.600 481.050 457.050 ;
        RECT 517.950 456.600 520.050 457.050 ;
        RECT 478.950 455.400 520.050 456.600 ;
        RECT 478.950 454.950 481.050 455.400 ;
        RECT 517.950 454.950 520.050 455.400 ;
        RECT 580.950 456.600 583.050 457.050 ;
        RECT 619.950 456.600 622.050 457.050 ;
        RECT 580.950 455.400 622.050 456.600 ;
        RECT 580.950 454.950 583.050 455.400 ;
        RECT 619.950 454.950 622.050 455.400 ;
        RECT 634.950 456.600 637.050 457.050 ;
        RECT 640.950 456.600 643.050 457.050 ;
        RECT 634.950 455.400 643.050 456.600 ;
        RECT 634.950 454.950 637.050 455.400 ;
        RECT 640.950 454.950 643.050 455.400 ;
        RECT 694.950 456.600 697.050 457.050 ;
        RECT 730.950 456.600 733.050 457.050 ;
        RECT 694.950 455.400 733.050 456.600 ;
        RECT 694.950 454.950 697.050 455.400 ;
        RECT 730.950 454.950 733.050 455.400 ;
        RECT 745.950 456.600 748.050 457.050 ;
        RECT 751.950 456.600 754.050 457.050 ;
        RECT 745.950 455.400 754.050 456.600 ;
        RECT 745.950 454.950 748.050 455.400 ;
        RECT 751.950 454.950 754.050 455.400 ;
        RECT 808.950 456.600 811.050 457.050 ;
        RECT 817.950 456.600 820.050 457.050 ;
        RECT 808.950 455.400 820.050 456.600 ;
        RECT 808.950 454.950 811.050 455.400 ;
        RECT 817.950 454.950 820.050 455.400 ;
        RECT 880.950 456.600 883.050 457.050 ;
        RECT 907.950 456.600 910.050 457.050 ;
        RECT 880.950 455.400 910.050 456.600 ;
        RECT 880.950 454.950 883.050 455.400 ;
        RECT 907.950 454.950 910.050 455.400 ;
        RECT 163.950 452.400 201.600 453.600 ;
        RECT 256.950 453.600 259.050 454.050 ;
        RECT 271.950 453.600 274.050 454.050 ;
        RECT 345.000 453.600 349.050 454.050 ;
        RECT 256.950 452.400 274.050 453.600 ;
        RECT 163.950 451.950 166.050 452.400 ;
        RECT 256.950 451.950 259.050 452.400 ;
        RECT 271.950 451.950 274.050 452.400 ;
        RECT 344.400 451.950 349.050 453.600 ;
        RECT 19.950 450.750 22.050 451.200 ;
        RECT 25.950 450.750 28.050 451.200 ;
        RECT 19.950 449.550 28.050 450.750 ;
        RECT 19.950 449.100 22.050 449.550 ;
        RECT 25.950 449.100 28.050 449.550 ;
        RECT 31.950 450.750 34.050 451.200 ;
        RECT 40.950 450.750 43.050 451.200 ;
        RECT 31.950 449.550 43.050 450.750 ;
        RECT 31.950 449.100 34.050 449.550 ;
        RECT 40.950 449.100 43.050 449.550 ;
        RECT 76.950 450.750 79.050 451.200 ;
        RECT 82.950 450.750 85.050 451.200 ;
        RECT 76.950 449.550 85.050 450.750 ;
        RECT 93.000 450.600 97.050 451.050 ;
        RECT 76.950 449.100 79.050 449.550 ;
        RECT 82.950 449.100 85.050 449.550 ;
        RECT 92.400 448.950 97.050 450.600 ;
        RECT 100.950 450.600 103.050 451.050 ;
        RECT 118.800 450.600 120.900 451.050 ;
        RECT 100.950 449.400 120.900 450.600 ;
        RECT 100.950 448.950 103.050 449.400 ;
        RECT 118.800 448.950 120.900 449.400 ;
        RECT 121.950 450.750 124.050 451.200 ;
        RECT 130.950 450.750 133.050 451.200 ;
        RECT 121.950 449.550 133.050 450.750 ;
        RECT 141.000 450.600 145.050 451.050 ;
        RECT 121.950 449.100 124.050 449.550 ;
        RECT 130.950 449.100 133.050 449.550 ;
        RECT 140.400 448.950 145.050 450.600 ;
        RECT 169.950 449.100 172.050 451.200 ;
        RECT 175.950 450.600 178.050 451.200 ;
        RECT 196.950 450.600 199.050 451.200 ;
        RECT 217.950 450.600 220.050 451.200 ;
        RECT 175.950 449.400 199.050 450.600 ;
        RECT 175.950 449.100 178.050 449.400 ;
        RECT 196.950 449.100 199.050 449.400 ;
        RECT 212.400 449.400 220.050 450.600 ;
        RECT 92.400 447.600 93.600 448.950 ;
        RECT 86.400 446.400 93.600 447.600 ;
        RECT 4.950 444.450 7.050 444.900 ;
        RECT 10.950 444.450 13.050 444.900 ;
        RECT 4.950 443.250 13.050 444.450 ;
        RECT 4.950 442.800 7.050 443.250 ;
        RECT 10.950 442.800 13.050 443.250 ;
        RECT 16.950 444.600 19.050 444.900 ;
        RECT 43.950 444.600 46.050 444.900 ;
        RECT 61.950 444.600 64.050 444.900 ;
        RECT 16.950 443.400 64.050 444.600 ;
        RECT 16.950 442.800 19.050 443.400 ;
        RECT 43.950 442.800 46.050 443.400 ;
        RECT 61.950 442.800 64.050 443.400 ;
        RECT 67.950 444.600 70.050 444.900 ;
        RECT 73.950 444.600 76.050 445.050 ;
        RECT 86.400 444.900 87.600 446.400 ;
        RECT 140.400 444.900 141.600 448.950 ;
        RECT 67.950 443.400 76.050 444.600 ;
        RECT 67.950 442.800 70.050 443.400 ;
        RECT 73.950 442.950 76.050 443.400 ;
        RECT 85.950 442.800 88.050 444.900 ;
        RECT 139.950 442.800 142.050 444.900 ;
        RECT 154.950 444.600 157.050 444.900 ;
        RECT 163.950 444.600 166.050 445.050 ;
        RECT 154.950 443.400 166.050 444.600 ;
        RECT 154.950 442.800 157.050 443.400 ;
        RECT 163.950 442.950 166.050 443.400 ;
        RECT 94.950 441.600 97.050 442.050 ;
        RECT 121.950 441.600 124.050 442.050 ;
        RECT 94.950 440.400 124.050 441.600 ;
        RECT 94.950 439.950 97.050 440.400 ;
        RECT 121.950 439.950 124.050 440.400 ;
        RECT 127.950 441.600 130.050 442.050 ;
        RECT 139.950 441.600 142.050 442.050 ;
        RECT 127.950 440.400 142.050 441.600 ;
        RECT 127.950 439.950 130.050 440.400 ;
        RECT 139.950 439.950 142.050 440.400 ;
        RECT 163.950 441.600 166.050 441.900 ;
        RECT 170.400 441.600 171.600 449.100 ;
        RECT 212.400 447.600 213.600 449.400 ;
        RECT 217.950 449.100 220.050 449.400 ;
        RECT 223.950 450.600 226.050 451.200 ;
        RECT 223.950 449.400 228.600 450.600 ;
        RECT 223.950 449.100 226.050 449.400 ;
        RECT 203.400 446.400 213.600 447.600 ;
        RECT 178.950 444.600 181.050 444.900 ;
        RECT 203.400 444.600 204.600 446.400 ;
        RECT 227.400 445.050 228.600 449.400 ;
        RECT 253.950 447.600 256.050 451.050 ;
        RECT 289.950 450.600 292.050 451.050 ;
        RECT 251.400 447.000 256.050 447.600 ;
        RECT 284.400 449.400 292.050 450.600 ;
        RECT 251.400 446.400 255.600 447.000 ;
        RECT 178.950 443.400 204.600 444.600 ;
        RECT 205.950 444.600 208.050 445.050 ;
        RECT 214.950 444.600 217.050 444.900 ;
        RECT 205.950 443.400 217.050 444.600 ;
        RECT 178.950 442.800 181.050 443.400 ;
        RECT 205.950 442.950 208.050 443.400 ;
        RECT 214.950 442.800 217.050 443.400 ;
        RECT 226.950 442.950 229.050 445.050 ;
        RECT 235.950 444.600 238.050 445.050 ;
        RECT 251.400 444.600 252.600 446.400 ;
        RECT 235.950 443.400 252.600 444.600 ;
        RECT 253.950 444.600 256.050 445.050 ;
        RECT 284.400 444.600 285.600 449.400 ;
        RECT 289.950 448.950 292.050 449.400 ;
        RECT 301.950 448.950 304.050 451.050 ;
        RECT 315.000 450.600 319.050 451.050 ;
        RECT 314.400 448.950 319.050 450.600 ;
        RECT 334.950 449.100 337.050 451.200 ;
        RECT 344.400 450.600 345.600 451.950 ;
        RECT 338.400 449.400 345.600 450.600 ;
        RECT 253.950 443.400 285.600 444.600 ;
        RECT 286.950 444.600 289.050 444.900 ;
        RECT 302.400 444.600 303.600 448.950 ;
        RECT 314.400 445.050 315.600 448.950 ;
        RECT 335.400 447.600 336.600 449.100 ;
        RECT 320.400 447.000 336.600 447.600 ;
        RECT 319.950 446.400 336.600 447.000 ;
        RECT 310.800 444.600 312.900 444.900 ;
        RECT 286.950 443.400 312.900 444.600 ;
        RECT 235.950 442.950 238.050 443.400 ;
        RECT 253.950 442.950 256.050 443.400 ;
        RECT 286.950 442.800 289.050 443.400 ;
        RECT 310.800 442.800 312.900 443.400 ;
        RECT 313.950 442.950 316.050 445.050 ;
        RECT 319.950 442.950 322.050 446.400 ;
        RECT 338.400 444.600 339.600 449.400 ;
        RECT 349.950 449.100 352.050 451.200 ;
        RECT 397.950 450.600 400.050 454.050 ;
        RECT 445.950 453.600 448.050 454.050 ;
        RECT 463.950 453.600 466.050 454.050 ;
        RECT 445.950 452.400 466.050 453.600 ;
        RECT 445.950 451.950 448.050 452.400 ;
        RECT 463.950 451.950 466.050 452.400 ;
        RECT 496.950 453.600 499.050 454.050 ;
        RECT 502.950 453.600 505.050 454.050 ;
        RECT 496.950 452.400 505.050 453.600 ;
        RECT 496.950 451.950 499.050 452.400 ;
        RECT 502.950 451.950 505.050 452.400 ;
        RECT 661.950 453.600 664.050 454.050 ;
        RECT 733.950 453.600 736.050 454.050 ;
        RECT 766.950 453.600 769.050 454.050 ;
        RECT 661.950 452.400 669.600 453.600 ;
        RECT 661.950 451.950 664.050 452.400 ;
        RECT 386.400 450.000 400.050 450.600 ;
        RECT 386.400 449.400 399.600 450.000 ;
        RECT 350.400 447.600 351.600 449.100 ;
        RECT 386.400 447.600 387.600 449.400 ;
        RECT 409.950 447.600 412.050 451.050 ;
        RECT 415.950 449.100 418.050 451.200 ;
        RECT 421.950 450.600 424.050 451.050 ;
        RECT 448.950 450.600 451.050 451.050 ;
        RECT 421.950 449.400 429.600 450.600 ;
        RECT 347.400 446.400 351.600 447.600 ;
        RECT 356.400 447.000 387.600 447.600 ;
        RECT 355.950 446.400 387.600 447.000 ;
        RECT 392.400 447.000 412.050 447.600 ;
        RECT 392.400 446.400 411.600 447.000 ;
        RECT 332.400 443.400 339.600 444.600 ;
        RECT 340.950 444.600 343.050 445.050 ;
        RECT 347.400 444.600 348.600 446.400 ;
        RECT 340.950 443.400 348.600 444.600 ;
        RECT 332.400 442.050 333.600 443.400 ;
        RECT 340.950 442.950 343.050 443.400 ;
        RECT 355.950 442.950 358.050 446.400 ;
        RECT 376.950 444.600 379.050 444.900 ;
        RECT 392.400 444.600 393.600 446.400 ;
        RECT 403.950 444.600 406.050 445.050 ;
        RECT 376.950 443.400 393.600 444.600 ;
        RECT 395.400 443.400 406.050 444.600 ;
        RECT 416.400 444.600 417.600 449.100 ;
        RECT 421.950 448.950 424.050 449.400 ;
        RECT 428.400 447.600 429.600 449.400 ;
        RECT 437.400 449.400 451.050 450.600 ;
        RECT 428.400 447.000 432.600 447.600 ;
        RECT 428.400 446.400 433.050 447.000 ;
        RECT 424.950 444.600 427.050 445.050 ;
        RECT 416.400 443.400 427.050 444.600 ;
        RECT 376.950 442.800 379.050 443.400 ;
        RECT 395.400 442.050 396.600 443.400 ;
        RECT 403.950 442.950 406.050 443.400 ;
        RECT 424.950 442.950 427.050 443.400 ;
        RECT 430.950 442.950 433.050 446.400 ;
        RECT 437.400 444.900 438.600 449.400 ;
        RECT 448.950 448.950 451.050 449.400 ;
        RECT 463.950 450.600 466.050 451.200 ;
        RECT 472.950 450.750 475.050 451.200 ;
        RECT 478.950 450.750 481.050 451.200 ;
        RECT 463.950 449.400 471.600 450.600 ;
        RECT 463.950 449.100 466.050 449.400 ;
        RECT 470.400 447.600 471.600 449.400 ;
        RECT 472.950 449.550 481.050 450.750 ;
        RECT 472.950 449.100 475.050 449.550 ;
        RECT 478.950 449.100 481.050 449.550 ;
        RECT 484.950 450.600 487.050 451.200 ;
        RECT 505.950 450.600 508.050 451.200 ;
        RECT 484.950 449.400 508.050 450.600 ;
        RECT 484.950 449.100 487.050 449.400 ;
        RECT 505.950 449.100 508.050 449.400 ;
        RECT 523.950 450.600 526.050 451.200 ;
        RECT 553.950 450.750 556.050 451.200 ;
        RECT 571.950 450.750 574.050 451.200 ;
        RECT 553.950 450.600 574.050 450.750 ;
        RECT 523.950 449.550 574.050 450.600 ;
        RECT 523.950 449.400 556.050 449.550 ;
        RECT 523.950 449.100 526.050 449.400 ;
        RECT 553.950 449.100 556.050 449.400 ;
        RECT 571.950 449.100 574.050 449.550 ;
        RECT 589.950 451.050 592.050 451.500 ;
        RECT 595.950 451.050 598.050 451.500 ;
        RECT 589.950 449.850 598.050 451.050 ;
        RECT 589.950 449.400 592.050 449.850 ;
        RECT 595.950 449.400 598.050 449.850 ;
        RECT 604.950 449.100 607.050 451.200 ;
        RECT 610.950 449.100 613.050 451.200 ;
        RECT 634.950 450.600 637.050 451.200 ;
        RECT 652.950 450.600 655.050 451.200 ;
        RECT 634.950 449.400 655.050 450.600 ;
        RECT 634.950 449.100 637.050 449.400 ;
        RECT 652.950 449.100 655.050 449.400 ;
        RECT 658.950 449.100 661.050 451.200 ;
        RECT 605.400 447.600 606.600 449.100 ;
        RECT 470.400 446.400 483.600 447.600 ;
        RECT 436.950 442.800 439.050 444.900 ;
        RECT 454.950 444.450 457.050 445.050 ;
        RECT 482.400 444.900 483.600 446.400 ;
        RECT 596.400 446.400 606.600 447.600 ;
        RECT 460.950 444.450 463.050 444.900 ;
        RECT 454.950 443.250 463.050 444.450 ;
        RECT 454.950 442.950 457.050 443.250 ;
        RECT 460.950 442.800 463.050 443.250 ;
        RECT 481.950 442.800 484.050 444.900 ;
        RECT 487.950 444.600 490.050 444.900 ;
        RECT 493.950 444.600 496.050 445.050 ;
        RECT 487.950 443.400 496.050 444.600 ;
        RECT 487.950 442.800 490.050 443.400 ;
        RECT 493.950 442.950 496.050 443.400 ;
        RECT 517.950 444.450 520.050 444.900 ;
        RECT 526.950 444.450 529.050 444.900 ;
        RECT 517.950 443.250 529.050 444.450 ;
        RECT 517.950 442.800 520.050 443.250 ;
        RECT 526.950 442.800 529.050 443.250 ;
        RECT 538.950 444.450 541.050 444.900 ;
        RECT 544.950 444.450 547.050 444.900 ;
        RECT 596.400 444.600 597.600 446.400 ;
        RECT 611.400 445.050 612.600 449.100 ;
        RECT 619.950 447.600 622.050 448.050 ;
        RECT 619.950 446.400 627.600 447.600 ;
        RECT 619.950 445.950 622.050 446.400 ;
        RECT 538.950 443.250 547.050 444.450 ;
        RECT 538.950 442.800 541.050 443.250 ;
        RECT 544.950 442.800 547.050 443.250 ;
        RECT 562.950 443.400 597.600 444.600 ;
        RECT 598.950 444.600 601.050 445.050 ;
        RECT 607.950 444.600 610.050 444.900 ;
        RECT 598.950 443.400 610.050 444.600 ;
        RECT 611.400 443.400 616.050 445.050 ;
        RECT 626.400 444.600 627.600 446.400 ;
        RECT 631.950 444.600 634.050 444.900 ;
        RECT 626.400 443.400 634.050 444.600 ;
        RECT 635.400 444.600 636.600 449.100 ;
        RECT 659.400 445.050 660.600 449.100 ;
        RECT 664.950 448.950 667.050 451.050 ;
        RECT 640.950 444.600 643.050 445.050 ;
        RECT 635.400 443.400 643.050 444.600 ;
        RECT 659.400 443.400 664.050 445.050 ;
        RECT 562.950 442.500 565.050 443.400 ;
        RECT 598.950 442.950 601.050 443.400 ;
        RECT 607.950 442.800 610.050 443.400 ;
        RECT 612.000 442.950 616.050 443.400 ;
        RECT 631.950 442.800 634.050 443.400 ;
        RECT 640.950 442.950 643.050 443.400 ;
        RECT 660.000 442.950 664.050 443.400 ;
        RECT 163.950 440.400 171.600 441.600 ;
        RECT 232.950 441.600 235.050 442.050 ;
        RECT 244.950 441.600 247.050 442.050 ;
        RECT 232.950 440.400 247.050 441.600 ;
        RECT 163.950 439.800 166.050 440.400 ;
        RECT 232.950 439.950 235.050 440.400 ;
        RECT 244.950 439.950 247.050 440.400 ;
        RECT 256.950 441.600 259.050 442.050 ;
        RECT 271.950 441.600 274.050 442.050 ;
        RECT 256.950 440.400 274.050 441.600 ;
        RECT 256.950 439.950 259.050 440.400 ;
        RECT 271.950 439.950 274.050 440.400 ;
        RECT 292.950 441.600 295.050 442.050 ;
        RECT 304.950 441.600 307.050 442.050 ;
        RECT 292.950 440.400 307.050 441.600 ;
        RECT 292.950 439.950 295.050 440.400 ;
        RECT 304.950 439.950 307.050 440.400 ;
        RECT 328.950 440.400 333.600 442.050 ;
        RECT 352.950 441.600 355.050 442.050 ;
        RECT 358.950 441.600 361.050 442.050 ;
        RECT 367.950 441.600 370.050 442.050 ;
        RECT 352.950 440.400 370.050 441.600 ;
        RECT 328.950 439.950 333.000 440.400 ;
        RECT 352.950 439.950 355.050 440.400 ;
        RECT 358.950 439.950 361.050 440.400 ;
        RECT 367.950 439.950 370.050 440.400 ;
        RECT 391.950 440.400 396.600 442.050 ;
        RECT 472.950 441.600 475.050 442.050 ;
        RECT 484.950 441.600 487.050 442.050 ;
        RECT 472.950 440.400 487.050 441.600 ;
        RECT 391.950 439.950 396.000 440.400 ;
        RECT 472.950 439.950 475.050 440.400 ;
        RECT 484.950 439.950 487.050 440.400 ;
        RECT 535.950 441.600 538.050 442.050 ;
        RECT 622.950 441.600 625.050 442.050 ;
        RECT 535.950 440.400 625.050 441.600 ;
        RECT 535.950 439.950 538.050 440.400 ;
        RECT 622.950 439.950 625.050 440.400 ;
        RECT 637.950 441.600 640.050 442.050 ;
        RECT 665.400 441.600 666.600 448.950 ;
        RECT 668.400 444.600 669.600 452.400 ;
        RECT 733.950 452.400 769.050 453.600 ;
        RECT 733.950 451.950 736.050 452.400 ;
        RECT 766.950 451.950 769.050 452.400 ;
        RECT 778.950 453.600 781.050 454.050 ;
        RECT 790.950 453.600 793.050 454.050 ;
        RECT 885.000 453.600 889.050 454.050 ;
        RECT 778.950 452.400 793.050 453.600 ;
        RECT 778.950 451.950 781.050 452.400 ;
        RECT 790.950 451.950 793.050 452.400 ;
        RECT 884.400 451.950 889.050 453.600 ;
        RECT 913.950 453.600 916.050 454.050 ;
        RECT 919.950 453.600 922.050 454.050 ;
        RECT 913.950 452.400 922.050 453.600 ;
        RECT 913.950 451.950 916.050 452.400 ;
        RECT 919.950 451.950 922.050 452.400 ;
        RECT 685.950 449.400 688.050 451.500 ;
        RECT 686.400 445.050 687.600 449.400 ;
        RECT 697.950 448.950 700.050 451.050 ;
        RECT 718.950 448.950 721.050 451.050 ;
        RECT 730.950 450.600 733.050 451.500 ;
        RECT 742.950 450.600 745.050 451.050 ;
        RECT 748.800 450.600 750.900 451.200 ;
        RECT 730.950 449.400 750.900 450.600 ;
        RECT 742.950 448.950 745.050 449.400 ;
        RECT 748.800 449.100 750.900 449.400 ;
        RECT 751.950 450.600 754.050 451.050 ;
        RECT 751.950 449.400 768.600 450.600 ;
        RECT 751.950 448.950 754.050 449.400 ;
        RECT 698.400 445.050 699.600 448.950 ;
        RECT 667.950 442.500 670.050 444.600 ;
        RECT 682.950 443.400 687.600 445.050 ;
        RECT 682.950 442.950 687.000 443.400 ;
        RECT 697.950 442.950 700.050 445.050 ;
        RECT 719.400 444.600 720.600 448.950 ;
        RECT 767.400 447.600 768.600 449.400 ;
        RECT 805.950 447.600 808.050 451.050 ;
        RECT 820.950 450.600 823.050 451.050 ;
        RECT 829.950 450.600 832.050 451.050 ;
        RECT 820.950 449.400 832.050 450.600 ;
        RECT 820.950 448.950 823.050 449.400 ;
        RECT 829.950 448.950 832.050 449.400 ;
        RECT 841.950 450.600 844.050 451.050 ;
        RECT 853.950 450.600 856.050 451.200 ;
        RECT 841.950 449.400 856.050 450.600 ;
        RECT 841.950 448.950 844.050 449.400 ;
        RECT 853.950 449.100 856.050 449.400 ;
        RECT 874.950 448.950 877.050 451.050 ;
        RECT 767.400 446.400 804.600 447.600 ;
        RECT 805.950 447.000 813.600 447.600 ;
        RECT 806.400 446.400 814.050 447.000 ;
        RECT 803.400 444.900 804.600 446.400 ;
        RECT 703.950 443.400 720.600 444.600 ;
        RECT 733.950 444.450 736.050 444.900 ;
        RECT 784.950 444.450 787.050 444.900 ;
        RECT 703.950 442.500 706.050 443.400 ;
        RECT 733.950 443.250 787.050 444.450 ;
        RECT 733.950 442.800 736.050 443.250 ;
        RECT 784.950 442.800 787.050 443.250 ;
        RECT 802.950 442.800 805.050 444.900 ;
        RECT 811.950 442.950 814.050 446.400 ;
        RECT 875.400 445.050 876.600 448.950 ;
        RECT 832.950 444.600 835.050 444.900 ;
        RECT 832.950 444.000 840.600 444.600 ;
        RECT 832.950 443.400 841.050 444.000 ;
        RECT 832.950 442.800 835.050 443.400 ;
        RECT 637.950 440.400 666.600 441.600 ;
        RECT 754.950 441.600 757.050 442.050 ;
        RECT 769.950 441.600 772.050 442.050 ;
        RECT 754.950 440.400 772.050 441.600 ;
        RECT 637.950 439.950 640.050 440.400 ;
        RECT 754.950 439.950 757.050 440.400 ;
        RECT 769.950 439.950 772.050 440.400 ;
        RECT 838.950 439.950 841.050 443.400 ;
        RECT 874.950 442.950 877.050 445.050 ;
        RECT 884.400 442.050 885.600 451.950 ;
        RECT 892.950 448.950 895.050 451.050 ;
        RECT 901.950 448.950 904.050 451.050 ;
        RECT 893.400 445.050 894.600 448.950 ;
        RECT 902.400 445.050 903.600 448.950 ;
        RECT 892.950 442.950 895.050 445.050 ;
        RECT 901.950 442.950 904.050 445.050 ;
        RECT 910.950 444.450 913.050 444.900 ;
        RECT 919.950 444.450 922.050 444.900 ;
        RECT 910.950 443.250 922.050 444.450 ;
        RECT 910.950 442.800 913.050 443.250 ;
        RECT 919.950 442.800 922.050 443.250 ;
        RECT 883.950 439.950 886.050 442.050 ;
        RECT 898.950 441.600 901.050 442.050 ;
        RECT 913.950 441.600 916.050 442.050 ;
        RECT 898.950 440.400 916.050 441.600 ;
        RECT 898.950 439.950 901.050 440.400 ;
        RECT 913.950 439.950 916.050 440.400 ;
        RECT 91.950 438.600 94.050 439.050 ;
        RECT 100.950 438.600 103.050 439.050 ;
        RECT 91.950 437.400 103.050 438.600 ;
        RECT 91.950 436.950 94.050 437.400 ;
        RECT 100.950 436.950 103.050 437.400 ;
        RECT 160.950 438.600 163.050 439.050 ;
        RECT 193.950 438.600 196.050 439.050 ;
        RECT 160.950 437.400 196.050 438.600 ;
        RECT 160.950 436.950 163.050 437.400 ;
        RECT 193.950 436.950 196.050 437.400 ;
        RECT 208.950 438.600 211.050 439.050 ;
        RECT 220.950 438.600 223.050 439.050 ;
        RECT 208.950 437.400 223.050 438.600 ;
        RECT 245.400 438.600 246.600 439.950 ;
        RECT 259.950 438.600 262.050 439.050 ;
        RECT 245.400 437.400 262.050 438.600 ;
        RECT 208.950 436.950 211.050 437.400 ;
        RECT 220.950 436.950 223.050 437.400 ;
        RECT 259.950 436.950 262.050 437.400 ;
        RECT 325.950 438.600 328.050 439.050 ;
        RECT 334.950 438.600 337.050 439.050 ;
        RECT 325.950 437.400 337.050 438.600 ;
        RECT 325.950 436.950 328.050 437.400 ;
        RECT 334.950 436.950 337.050 437.400 ;
        RECT 364.950 438.600 367.050 439.050 ;
        RECT 370.950 438.600 373.050 439.050 ;
        RECT 364.950 437.400 373.050 438.600 ;
        RECT 364.950 436.950 367.050 437.400 ;
        RECT 370.950 436.950 373.050 437.400 ;
        RECT 406.950 438.600 409.050 439.050 ;
        RECT 418.950 438.600 421.050 439.050 ;
        RECT 406.950 437.400 421.050 438.600 ;
        RECT 406.950 436.950 409.050 437.400 ;
        RECT 418.950 436.950 421.050 437.400 ;
        RECT 451.950 438.600 454.050 439.050 ;
        RECT 460.950 438.600 463.050 439.050 ;
        RECT 466.950 438.600 469.050 439.050 ;
        RECT 451.950 437.400 469.050 438.600 ;
        RECT 451.950 436.950 454.050 437.400 ;
        RECT 460.950 436.950 463.050 437.400 ;
        RECT 466.950 436.950 469.050 437.400 ;
        RECT 643.950 438.600 646.050 439.050 ;
        RECT 649.950 438.600 652.050 439.050 ;
        RECT 643.950 437.400 652.050 438.600 ;
        RECT 643.950 436.950 646.050 437.400 ;
        RECT 649.950 436.950 652.050 437.400 ;
        RECT 655.950 438.600 658.050 439.050 ;
        RECT 682.950 438.600 685.050 439.050 ;
        RECT 655.950 437.400 685.050 438.600 ;
        RECT 655.950 436.950 658.050 437.400 ;
        RECT 682.950 436.950 685.050 437.400 ;
        RECT 760.950 438.600 763.050 439.050 ;
        RECT 766.950 438.600 769.050 439.050 ;
        RECT 760.950 437.400 769.050 438.600 ;
        RECT 760.950 436.950 763.050 437.400 ;
        RECT 766.950 436.950 769.050 437.400 ;
        RECT 877.950 438.600 880.050 439.050 ;
        RECT 889.950 438.600 892.050 439.050 ;
        RECT 877.950 437.400 892.050 438.600 ;
        RECT 877.950 436.950 880.050 437.400 ;
        RECT 889.950 436.950 892.050 437.400 ;
        RECT 916.950 438.600 919.050 439.050 ;
        RECT 923.400 438.600 924.600 457.950 ;
        RECT 916.950 437.400 924.600 438.600 ;
        RECT 916.950 436.950 919.050 437.400 ;
        RECT 19.950 435.600 22.050 436.050 ;
        RECT 40.950 435.600 43.050 436.050 ;
        RECT 85.950 435.600 88.050 436.050 ;
        RECT 19.950 434.400 88.050 435.600 ;
        RECT 19.950 433.950 22.050 434.400 ;
        RECT 40.950 433.950 43.050 434.400 ;
        RECT 85.950 433.950 88.050 434.400 ;
        RECT 250.950 435.600 253.050 436.050 ;
        RECT 274.950 435.600 277.050 436.050 ;
        RECT 250.950 434.400 277.050 435.600 ;
        RECT 250.950 433.950 253.050 434.400 ;
        RECT 274.950 433.950 277.050 434.400 ;
        RECT 361.950 435.600 364.050 436.050 ;
        RECT 373.950 435.600 376.050 436.050 ;
        RECT 361.950 434.400 376.050 435.600 ;
        RECT 361.950 433.950 364.050 434.400 ;
        RECT 373.950 433.950 376.050 434.400 ;
        RECT 418.950 435.600 421.050 435.900 ;
        RECT 427.950 435.600 430.050 436.050 ;
        RECT 418.950 434.400 430.050 435.600 ;
        RECT 418.950 433.800 421.050 434.400 ;
        RECT 427.950 433.950 430.050 434.400 ;
        RECT 475.950 435.600 478.050 436.050 ;
        RECT 493.950 435.600 496.050 436.050 ;
        RECT 559.950 435.600 562.050 436.050 ;
        RECT 475.950 434.400 562.050 435.600 ;
        RECT 475.950 433.950 478.050 434.400 ;
        RECT 493.950 433.950 496.050 434.400 ;
        RECT 559.950 433.950 562.050 434.400 ;
        RECT 598.950 435.600 601.050 436.050 ;
        RECT 616.950 435.600 619.050 436.050 ;
        RECT 598.950 434.400 619.050 435.600 ;
        RECT 598.950 433.950 601.050 434.400 ;
        RECT 616.950 433.950 619.050 434.400 ;
        RECT 679.950 435.600 682.050 436.050 ;
        RECT 733.950 435.600 736.050 436.050 ;
        RECT 679.950 434.400 736.050 435.600 ;
        RECT 679.950 433.950 682.050 434.400 ;
        RECT 733.950 433.950 736.050 434.400 ;
        RECT 772.950 435.600 775.050 436.050 ;
        RECT 811.950 435.600 814.050 436.050 ;
        RECT 772.950 434.400 814.050 435.600 ;
        RECT 772.950 433.950 775.050 434.400 ;
        RECT 811.950 433.950 814.050 434.400 ;
        RECT 862.950 435.600 865.050 436.050 ;
        RECT 904.950 435.600 907.050 436.050 ;
        RECT 862.950 434.400 907.050 435.600 ;
        RECT 862.950 433.950 865.050 434.400 ;
        RECT 904.950 433.950 907.050 434.400 ;
        RECT 58.950 432.600 61.050 433.050 ;
        RECT 121.950 432.600 124.050 433.050 ;
        RECT 58.950 431.400 124.050 432.600 ;
        RECT 58.950 430.950 61.050 431.400 ;
        RECT 121.950 430.950 124.050 431.400 ;
        RECT 133.950 432.600 136.050 433.050 ;
        RECT 169.950 432.600 172.050 433.050 ;
        RECT 172.950 432.600 175.050 433.050 ;
        RECT 133.950 431.400 175.050 432.600 ;
        RECT 133.950 430.950 136.050 431.400 ;
        RECT 169.950 430.950 172.050 431.400 ;
        RECT 172.950 430.950 175.050 431.400 ;
        RECT 184.950 432.600 187.050 433.050 ;
        RECT 199.950 432.600 202.050 433.050 ;
        RECT 184.950 431.400 202.050 432.600 ;
        RECT 184.950 430.950 187.050 431.400 ;
        RECT 199.950 430.950 202.050 431.400 ;
        RECT 232.950 432.600 235.050 433.050 ;
        RECT 244.950 432.600 247.050 433.050 ;
        RECT 232.950 431.400 247.050 432.600 ;
        RECT 232.950 430.950 235.050 431.400 ;
        RECT 244.950 430.950 247.050 431.400 ;
        RECT 280.950 432.600 283.050 433.050 ;
        RECT 301.950 432.600 304.050 433.050 ;
        RECT 280.950 431.400 304.050 432.600 ;
        RECT 280.950 430.950 283.050 431.400 ;
        RECT 301.950 430.950 304.050 431.400 ;
        RECT 322.950 432.600 325.050 433.050 ;
        RECT 334.950 432.600 337.050 433.050 ;
        RECT 322.950 431.400 337.050 432.600 ;
        RECT 322.950 430.950 325.050 431.400 ;
        RECT 334.950 430.950 337.050 431.400 ;
        RECT 379.950 432.600 382.050 433.050 ;
        RECT 442.950 432.600 445.050 433.050 ;
        RECT 379.950 431.400 445.050 432.600 ;
        RECT 379.950 430.950 382.050 431.400 ;
        RECT 442.950 430.950 445.050 431.400 ;
        RECT 565.950 432.600 568.050 433.050 ;
        RECT 571.950 432.600 574.050 433.050 ;
        RECT 565.950 431.400 574.050 432.600 ;
        RECT 565.950 430.950 568.050 431.400 ;
        RECT 571.950 430.950 574.050 431.400 ;
        RECT 613.950 432.600 616.050 433.050 ;
        RECT 640.950 432.600 643.050 433.050 ;
        RECT 613.950 431.400 643.050 432.600 ;
        RECT 613.950 430.950 616.050 431.400 ;
        RECT 640.950 430.950 643.050 431.400 ;
        RECT 649.950 432.600 652.050 433.050 ;
        RECT 664.950 432.600 667.050 433.050 ;
        RECT 649.950 431.400 667.050 432.600 ;
        RECT 649.950 430.950 652.050 431.400 ;
        RECT 664.950 430.950 667.050 431.400 ;
        RECT 778.950 432.600 781.050 433.050 ;
        RECT 784.950 432.600 787.050 433.050 ;
        RECT 802.950 432.600 805.050 433.050 ;
        RECT 778.950 431.400 805.050 432.600 ;
        RECT 778.950 430.950 781.050 431.400 ;
        RECT 784.950 430.950 787.050 431.400 ;
        RECT 802.950 430.950 805.050 431.400 ;
        RECT 829.950 432.600 832.050 433.050 ;
        RECT 841.950 432.600 844.050 433.050 ;
        RECT 829.950 431.400 844.050 432.600 ;
        RECT 829.950 430.950 832.050 431.400 ;
        RECT 841.950 430.950 844.050 431.400 ;
        RECT 31.950 429.600 34.050 430.050 ;
        RECT 37.950 429.600 40.050 430.050 ;
        RECT 76.950 429.600 79.050 430.050 ;
        RECT 31.950 428.400 79.050 429.600 ;
        RECT 31.950 427.950 34.050 428.400 ;
        RECT 37.950 427.950 40.050 428.400 ;
        RECT 76.950 427.950 79.050 428.400 ;
        RECT 241.950 429.600 244.050 430.050 ;
        RECT 281.400 429.600 282.600 430.950 ;
        RECT 241.950 428.400 282.600 429.600 ;
        RECT 307.950 429.600 310.050 430.050 ;
        RECT 325.950 429.600 328.050 430.050 ;
        RECT 307.950 428.400 328.050 429.600 ;
        RECT 241.950 427.950 244.050 428.400 ;
        RECT 307.950 427.950 310.050 428.400 ;
        RECT 325.950 427.950 328.050 428.400 ;
        RECT 349.950 429.600 352.050 430.050 ;
        RECT 358.950 429.600 361.050 430.050 ;
        RECT 349.950 428.400 361.050 429.600 ;
        RECT 349.950 427.950 352.050 428.400 ;
        RECT 358.950 427.950 361.050 428.400 ;
        RECT 397.950 429.600 400.050 430.050 ;
        RECT 430.950 429.600 433.050 430.050 ;
        RECT 502.950 429.600 505.050 430.050 ;
        RECT 397.950 428.400 433.050 429.600 ;
        RECT 397.950 427.950 400.050 428.400 ;
        RECT 430.950 427.950 433.050 428.400 ;
        RECT 455.400 428.400 505.050 429.600 ;
        RECT 82.950 426.600 85.050 427.050 ;
        RECT 109.950 426.600 112.050 427.050 ;
        RECT 82.950 425.400 112.050 426.600 ;
        RECT 82.950 424.950 85.050 425.400 ;
        RECT 109.950 424.950 112.050 425.400 ;
        RECT 157.950 426.600 160.050 427.050 ;
        RECT 187.950 426.600 190.050 427.050 ;
        RECT 157.950 425.400 190.050 426.600 ;
        RECT 157.950 424.950 160.050 425.400 ;
        RECT 187.950 424.950 190.050 425.400 ;
        RECT 247.950 426.600 250.050 427.050 ;
        RECT 313.950 426.600 316.050 427.050 ;
        RECT 247.950 425.400 316.050 426.600 ;
        RECT 247.950 424.950 250.050 425.400 ;
        RECT 313.950 424.950 316.050 425.400 ;
        RECT 331.950 426.600 334.050 427.050 ;
        RECT 337.950 426.600 340.050 427.050 ;
        RECT 346.950 426.600 349.050 427.050 ;
        RECT 331.950 425.400 340.050 426.600 ;
        RECT 331.950 424.950 334.050 425.400 ;
        RECT 337.950 424.950 340.050 425.400 ;
        RECT 341.400 425.400 349.050 426.600 ;
        RECT 25.950 423.600 28.050 424.050 ;
        RECT 49.950 423.600 52.050 424.050 ;
        RECT 25.950 422.400 52.050 423.600 ;
        RECT 25.950 421.950 28.050 422.400 ;
        RECT 49.950 421.950 52.050 422.400 ;
        RECT 73.950 423.600 76.050 424.050 ;
        RECT 145.950 423.600 148.050 424.050 ;
        RECT 73.950 422.400 148.050 423.600 ;
        RECT 73.950 421.950 76.050 422.400 ;
        RECT 145.950 421.950 148.050 422.400 ;
        RECT 199.950 423.600 202.050 424.050 ;
        RECT 232.950 423.600 235.050 424.050 ;
        RECT 199.950 422.400 235.050 423.600 ;
        RECT 199.950 421.950 202.050 422.400 ;
        RECT 232.950 421.950 235.050 422.400 ;
        RECT 238.950 423.600 241.050 424.050 ;
        RECT 307.950 423.600 310.050 424.050 ;
        RECT 319.950 423.600 322.050 424.050 ;
        RECT 341.400 423.600 342.600 425.400 ;
        RECT 346.950 424.950 349.050 425.400 ;
        RECT 409.950 426.600 412.050 427.050 ;
        RECT 455.400 426.600 456.600 428.400 ;
        RECT 502.950 427.950 505.050 428.400 ;
        RECT 508.950 429.600 511.050 430.050 ;
        RECT 517.950 429.600 520.050 430.050 ;
        RECT 508.950 428.400 520.050 429.600 ;
        RECT 508.950 427.950 511.050 428.400 ;
        RECT 517.950 427.950 520.050 428.400 ;
        RECT 550.950 429.600 553.050 430.050 ;
        RECT 559.950 429.600 562.050 430.050 ;
        RECT 550.950 428.400 562.050 429.600 ;
        RECT 550.950 427.950 553.050 428.400 ;
        RECT 559.950 427.950 562.050 428.400 ;
        RECT 625.950 429.600 628.050 430.050 ;
        RECT 637.950 429.600 640.050 430.050 ;
        RECT 688.950 429.600 691.050 430.050 ;
        RECT 625.950 428.400 640.050 429.600 ;
        RECT 625.950 427.950 628.050 428.400 ;
        RECT 637.950 427.950 640.050 428.400 ;
        RECT 680.400 428.400 691.050 429.600 ;
        RECT 680.400 427.050 681.600 428.400 ;
        RECT 688.950 427.950 691.050 428.400 ;
        RECT 700.950 429.600 703.050 430.050 ;
        RECT 712.950 429.600 715.050 430.050 ;
        RECT 700.950 428.400 715.050 429.600 ;
        RECT 700.950 427.950 703.050 428.400 ;
        RECT 712.950 427.950 715.050 428.400 ;
        RECT 724.950 429.600 727.050 430.050 ;
        RECT 769.950 429.600 772.050 430.050 ;
        RECT 724.950 428.400 772.050 429.600 ;
        RECT 724.950 427.950 727.050 428.400 ;
        RECT 769.950 427.950 772.050 428.400 ;
        RECT 880.950 429.600 883.050 430.050 ;
        RECT 886.950 429.600 889.050 430.050 ;
        RECT 880.950 428.400 889.050 429.600 ;
        RECT 880.950 427.950 883.050 428.400 ;
        RECT 886.950 427.950 889.050 428.400 ;
        RECT 892.950 429.600 895.050 430.050 ;
        RECT 919.950 429.600 922.050 430.050 ;
        RECT 892.950 428.400 922.050 429.600 ;
        RECT 892.950 427.950 895.050 428.400 ;
        RECT 919.950 427.950 922.050 428.400 ;
        RECT 409.950 425.400 456.600 426.600 ;
        RECT 475.950 426.600 478.050 427.050 ;
        RECT 604.950 426.600 607.050 427.050 ;
        RECT 679.950 426.600 682.050 427.050 ;
        RECT 475.950 425.400 607.050 426.600 ;
        RECT 409.950 424.950 412.050 425.400 ;
        RECT 475.950 424.950 478.050 425.400 ;
        RECT 604.950 424.950 607.050 425.400 ;
        RECT 635.400 425.400 682.050 426.600 ;
        RECT 238.950 422.400 310.050 423.600 ;
        RECT 238.950 421.950 241.050 422.400 ;
        RECT 307.950 421.950 310.050 422.400 ;
        RECT 317.400 422.400 342.600 423.600 ;
        RECT 343.950 423.600 346.050 424.050 ;
        RECT 376.950 423.600 379.050 424.050 ;
        RECT 382.950 423.600 385.050 424.050 ;
        RECT 343.950 422.400 375.600 423.600 ;
        RECT 115.950 420.600 118.050 421.050 ;
        RECT 127.950 420.600 130.050 421.050 ;
        RECT 115.950 419.400 130.050 420.600 ;
        RECT 115.950 418.950 118.050 419.400 ;
        RECT 127.950 418.950 130.050 419.400 ;
        RECT 175.950 420.600 178.050 421.050 ;
        RECT 193.950 420.600 196.050 421.050 ;
        RECT 175.950 419.400 196.050 420.600 ;
        RECT 175.950 418.950 178.050 419.400 ;
        RECT 193.950 418.950 196.050 419.400 ;
        RECT 223.950 420.600 226.050 421.050 ;
        RECT 268.950 420.600 271.050 421.050 ;
        RECT 317.400 420.600 318.600 422.400 ;
        RECT 319.950 421.950 322.050 422.400 ;
        RECT 343.950 421.950 346.050 422.400 ;
        RECT 223.950 420.000 231.600 420.600 ;
        RECT 223.950 419.400 232.050 420.000 ;
        RECT 223.950 418.950 226.050 419.400 ;
        RECT 7.950 417.600 10.050 418.050 ;
        RECT 13.950 417.600 16.050 418.200 ;
        RECT 7.950 416.400 16.050 417.600 ;
        RECT 7.950 415.950 10.050 416.400 ;
        RECT 13.950 416.100 16.050 416.400 ;
        RECT 31.950 417.600 36.000 418.050 ;
        RECT 43.950 417.600 46.050 418.200 ;
        RECT 64.950 417.600 67.050 418.200 ;
        RECT 82.950 417.600 85.050 418.200 ;
        RECT 31.950 415.950 36.600 417.600 ;
        RECT 43.950 416.400 63.600 417.600 ;
        RECT 43.950 416.100 46.050 416.400 ;
        RECT 35.400 411.900 36.600 415.950 ;
        RECT 62.400 411.900 63.600 416.400 ;
        RECT 64.950 416.400 85.050 417.600 ;
        RECT 64.950 416.100 67.050 416.400 ;
        RECT 82.950 416.100 85.050 416.400 ;
        RECT 88.950 417.600 91.050 418.200 ;
        RECT 100.950 417.600 103.050 418.050 ;
        RECT 109.950 417.600 112.050 418.200 ;
        RECT 88.950 416.400 93.600 417.600 ;
        RECT 88.950 416.100 91.050 416.400 ;
        RECT 22.950 411.600 25.050 411.900 ;
        RECT 34.950 411.600 37.050 411.900 ;
        RECT 22.950 410.400 37.050 411.600 ;
        RECT 22.950 409.800 25.050 410.400 ;
        RECT 34.950 409.800 37.050 410.400 ;
        RECT 61.950 409.800 64.050 411.900 ;
        RECT 73.950 411.450 76.050 411.900 ;
        RECT 85.950 411.450 88.050 411.900 ;
        RECT 73.950 410.250 88.050 411.450 ;
        RECT 92.400 411.600 93.600 416.400 ;
        RECT 100.950 416.400 112.050 417.600 ;
        RECT 100.950 415.950 103.050 416.400 ;
        RECT 109.950 416.100 112.050 416.400 ;
        RECT 124.950 415.950 127.050 418.050 ;
        RECT 142.950 417.600 145.050 418.050 ;
        RECT 148.950 417.600 151.050 418.200 ;
        RECT 163.950 417.600 166.050 418.050 ;
        RECT 142.950 416.400 166.050 417.600 ;
        RECT 142.950 415.950 145.050 416.400 ;
        RECT 148.950 416.100 151.050 416.400 ;
        RECT 125.400 412.050 126.600 415.950 ;
        RECT 155.400 414.600 156.600 416.400 ;
        RECT 163.950 415.950 166.050 416.400 ;
        RECT 193.950 417.600 196.050 418.200 ;
        RECT 214.950 417.600 217.050 418.200 ;
        RECT 193.950 416.400 217.050 417.600 ;
        RECT 193.950 416.100 196.050 416.400 ;
        RECT 214.950 416.100 217.050 416.400 ;
        RECT 229.950 415.950 232.050 419.400 ;
        RECT 268.950 419.400 318.600 420.600 ;
        RECT 325.950 420.600 328.050 421.050 ;
        RECT 340.950 420.600 343.050 421.050 ;
        RECT 325.950 419.400 343.050 420.600 ;
        RECT 374.400 420.600 375.600 422.400 ;
        RECT 376.950 422.400 385.050 423.600 ;
        RECT 376.950 421.950 379.050 422.400 ;
        RECT 382.950 421.950 385.050 422.400 ;
        RECT 433.950 423.600 436.050 424.050 ;
        RECT 445.950 423.600 448.050 424.050 ;
        RECT 433.950 422.400 448.050 423.600 ;
        RECT 433.950 421.950 436.050 422.400 ;
        RECT 445.950 421.950 448.050 422.400 ;
        RECT 562.950 423.600 565.050 424.050 ;
        RECT 589.950 423.600 592.050 424.050 ;
        RECT 635.400 423.600 636.600 425.400 ;
        RECT 679.950 424.950 682.050 425.400 ;
        RECT 709.950 426.600 712.050 427.050 ;
        RECT 715.950 426.600 718.050 427.050 ;
        RECT 709.950 425.400 718.050 426.600 ;
        RECT 709.950 424.950 712.050 425.400 ;
        RECT 715.950 424.950 718.050 425.400 ;
        RECT 820.950 426.600 823.050 427.050 ;
        RECT 832.950 426.600 835.050 427.050 ;
        RECT 820.950 425.400 835.050 426.600 ;
        RECT 820.950 424.950 823.050 425.400 ;
        RECT 832.950 424.950 835.050 425.400 ;
        RECT 841.950 426.600 844.050 427.050 ;
        RECT 856.950 426.600 859.050 427.050 ;
        RECT 841.950 425.400 859.050 426.600 ;
        RECT 841.950 424.950 844.050 425.400 ;
        RECT 856.950 424.950 859.050 425.400 ;
        RECT 562.950 422.400 592.050 423.600 ;
        RECT 562.950 421.950 565.050 422.400 ;
        RECT 589.950 421.950 592.050 422.400 ;
        RECT 626.400 422.400 636.600 423.600 ;
        RECT 637.950 423.600 640.050 424.050 ;
        RECT 646.950 423.600 649.050 424.050 ;
        RECT 637.950 422.400 649.050 423.600 ;
        RECT 409.950 420.600 412.050 421.050 ;
        RECT 374.400 419.400 412.050 420.600 ;
        RECT 268.950 418.950 271.050 419.400 ;
        RECT 325.950 418.950 328.050 419.400 ;
        RECT 340.950 418.950 343.050 419.400 ;
        RECT 409.950 418.950 412.050 419.400 ;
        RECT 496.950 420.600 499.050 421.050 ;
        RECT 511.950 420.600 514.050 421.050 ;
        RECT 496.950 419.400 514.050 420.600 ;
        RECT 496.950 418.950 499.050 419.400 ;
        RECT 511.950 418.950 514.050 419.400 ;
        RECT 595.950 418.950 598.050 421.050 ;
        RECT 616.950 420.600 619.050 421.050 ;
        RECT 626.400 420.600 627.600 422.400 ;
        RECT 637.950 421.950 640.050 422.400 ;
        RECT 646.950 421.950 649.050 422.400 ;
        RECT 676.950 423.600 679.050 424.050 ;
        RECT 682.950 423.600 685.050 424.050 ;
        RECT 676.950 422.400 685.050 423.600 ;
        RECT 676.950 421.950 679.050 422.400 ;
        RECT 682.950 421.950 685.050 422.400 ;
        RECT 697.950 423.600 700.050 424.050 ;
        RECT 706.950 423.600 709.050 424.050 ;
        RECT 697.950 422.400 709.050 423.600 ;
        RECT 697.950 421.950 700.050 422.400 ;
        RECT 706.950 421.950 709.050 422.400 ;
        RECT 721.950 423.600 724.050 424.050 ;
        RECT 736.950 423.600 739.050 424.050 ;
        RECT 775.950 423.600 778.050 423.900 ;
        RECT 721.950 422.400 739.050 423.600 ;
        RECT 721.950 421.950 724.050 422.400 ;
        RECT 736.950 421.950 739.050 422.400 ;
        RECT 752.400 422.400 778.050 423.600 ;
        RECT 752.400 420.600 753.600 422.400 ;
        RECT 775.950 421.800 778.050 422.400 ;
        RECT 787.950 423.600 790.050 424.050 ;
        RECT 814.950 423.600 817.050 424.050 ;
        RECT 787.950 422.400 817.050 423.600 ;
        RECT 787.950 421.950 790.050 422.400 ;
        RECT 814.950 421.950 817.050 422.400 ;
        RECT 868.950 423.600 871.050 424.050 ;
        RECT 874.950 423.600 877.050 424.050 ;
        RECT 868.950 422.400 877.050 423.600 ;
        RECT 868.950 421.950 871.050 422.400 ;
        RECT 874.950 421.950 877.050 422.400 ;
        RECT 901.950 423.600 904.050 424.050 ;
        RECT 907.950 423.600 910.050 424.050 ;
        RECT 901.950 422.400 910.050 423.600 ;
        RECT 901.950 421.950 904.050 422.400 ;
        RECT 907.950 421.950 910.050 422.400 ;
        RECT 616.950 419.400 627.600 420.600 ;
        RECT 740.400 419.400 753.600 420.600 ;
        RECT 616.950 418.950 619.050 419.400 ;
        RECT 235.950 415.950 238.050 418.050 ;
        RECT 265.950 417.750 268.050 418.200 ;
        RECT 274.950 417.750 277.050 418.200 ;
        RECT 265.950 416.550 277.050 417.750 ;
        RECT 265.950 416.100 268.050 416.550 ;
        RECT 274.950 416.100 277.050 416.550 ;
        RECT 155.400 413.400 159.600 414.600 ;
        RECT 112.950 411.600 115.050 411.900 ;
        RECT 92.400 410.400 115.050 411.600 ;
        RECT 73.950 409.800 76.050 410.250 ;
        RECT 85.950 409.800 88.050 410.250 ;
        RECT 112.950 409.800 115.050 410.400 ;
        RECT 124.950 409.950 127.050 412.050 ;
        RECT 151.950 411.600 154.050 411.900 ;
        RECT 146.400 411.000 154.050 411.600 ;
        RECT 145.950 410.400 154.050 411.000 ;
        RECT 158.400 411.600 159.600 413.400 ;
        RECT 236.400 412.050 237.600 415.950 ;
        RECT 277.950 414.600 280.050 415.050 ;
        RECT 295.950 414.600 298.050 418.050 ;
        RECT 313.950 417.750 316.050 418.050 ;
        RECT 319.950 417.750 322.050 418.200 ;
        RECT 313.950 416.550 322.050 417.750 ;
        RECT 313.950 415.950 316.050 416.550 ;
        RECT 319.950 416.100 322.050 416.550 ;
        RECT 352.950 414.600 355.050 418.050 ;
        RECT 361.950 417.600 364.050 418.200 ;
        RECT 391.950 417.600 394.050 418.050 ;
        RECT 403.950 417.600 406.050 418.200 ;
        RECT 424.950 417.600 427.050 418.200 ;
        RECT 361.950 416.400 390.600 417.600 ;
        RECT 361.950 416.100 364.050 416.400 ;
        RECT 248.400 413.400 270.600 414.600 ;
        RECT 166.950 411.600 169.050 411.900 ;
        RECT 158.400 410.400 169.050 411.600 ;
        RECT 16.950 408.600 19.050 409.050 ;
        RECT 46.950 408.600 49.050 409.050 ;
        RECT 52.950 408.600 55.050 409.050 ;
        RECT 16.950 407.400 55.050 408.600 ;
        RECT 16.950 406.950 19.050 407.400 ;
        RECT 46.950 406.950 49.050 407.400 ;
        RECT 52.950 406.950 55.050 407.400 ;
        RECT 145.950 406.950 148.050 410.400 ;
        RECT 151.950 409.800 154.050 410.400 ;
        RECT 166.950 409.800 169.050 410.400 ;
        RECT 223.950 411.450 226.050 411.900 ;
        RECT 229.950 411.450 232.050 412.050 ;
        RECT 223.950 410.250 232.050 411.450 ;
        RECT 223.950 409.800 226.050 410.250 ;
        RECT 229.950 409.950 232.050 410.250 ;
        RECT 235.950 409.950 238.050 412.050 ;
        RECT 241.950 411.600 244.050 411.900 ;
        RECT 248.400 411.600 249.600 413.400 ;
        RECT 241.950 410.400 249.600 411.600 ;
        RECT 253.950 411.600 256.050 412.050 ;
        RECT 269.400 411.900 270.600 413.400 ;
        RECT 277.950 414.000 298.050 414.600 ;
        RECT 347.400 414.000 355.050 414.600 ;
        RECT 389.400 414.600 390.600 416.400 ;
        RECT 391.950 416.400 406.050 417.600 ;
        RECT 391.950 415.950 394.050 416.400 ;
        RECT 403.950 416.100 406.050 416.400 ;
        RECT 407.400 416.400 427.050 417.600 ;
        RECT 394.950 414.600 397.050 415.050 ;
        RECT 407.400 414.600 408.600 416.400 ;
        RECT 424.950 416.100 427.050 416.400 ;
        RECT 436.950 417.600 439.050 418.050 ;
        RECT 451.950 417.600 454.050 418.200 ;
        RECT 436.950 416.400 454.050 417.600 ;
        RECT 436.950 415.950 439.050 416.400 ;
        RECT 451.950 416.100 454.050 416.400 ;
        RECT 502.950 417.600 505.050 418.200 ;
        RECT 508.950 417.600 511.050 418.050 ;
        RECT 502.950 416.400 511.050 417.600 ;
        RECT 502.950 416.100 505.050 416.400 ;
        RECT 277.950 413.400 297.600 414.000 ;
        RECT 347.400 413.400 354.600 414.000 ;
        RECT 389.400 413.400 393.600 414.600 ;
        RECT 277.950 412.950 280.050 413.400 ;
        RECT 262.950 411.600 265.050 411.900 ;
        RECT 253.950 410.400 265.050 411.600 ;
        RECT 241.950 409.800 244.050 410.400 ;
        RECT 253.950 409.950 256.050 410.400 ;
        RECT 262.950 409.800 265.050 410.400 ;
        RECT 268.950 409.800 271.050 411.900 ;
        RECT 298.950 411.600 301.050 411.900 ;
        RECT 316.950 411.600 319.050 412.050 ;
        RECT 347.400 411.600 348.600 413.400 ;
        RECT 298.950 411.000 303.600 411.600 ;
        RECT 298.950 410.400 304.050 411.000 ;
        RECT 298.950 409.800 301.050 410.400 ;
        RECT 250.950 408.600 253.050 409.050 ;
        RECT 259.800 408.600 261.900 409.050 ;
        RECT 250.950 407.400 261.900 408.600 ;
        RECT 250.950 406.950 253.050 407.400 ;
        RECT 259.800 406.950 261.900 407.400 ;
        RECT 262.950 408.600 265.050 409.050 ;
        RECT 280.950 408.600 283.050 409.050 ;
        RECT 262.950 407.400 283.050 408.600 ;
        RECT 262.950 406.950 265.050 407.400 ;
        RECT 280.950 406.950 283.050 407.400 ;
        RECT 301.950 406.950 304.050 410.400 ;
        RECT 316.950 410.400 348.600 411.600 ;
        RECT 349.950 411.600 352.050 412.050 ;
        RECT 364.950 411.600 367.050 411.900 ;
        RECT 349.950 410.400 367.050 411.600 ;
        RECT 316.950 409.950 319.050 410.400 ;
        RECT 349.950 409.950 352.050 410.400 ;
        RECT 364.950 409.800 367.050 410.400 ;
        RECT 392.400 411.600 393.600 413.400 ;
        RECT 394.950 413.400 408.600 414.600 ;
        RECT 394.950 412.950 397.050 413.400 ;
        RECT 503.400 412.050 504.600 416.100 ;
        RECT 508.950 415.950 511.050 416.400 ;
        RECT 523.950 417.600 526.050 418.200 ;
        RECT 541.950 417.600 544.050 418.200 ;
        RECT 523.950 416.400 544.050 417.600 ;
        RECT 523.950 416.100 526.050 416.400 ;
        RECT 541.950 416.100 544.050 416.400 ;
        RECT 547.950 417.600 550.050 418.200 ;
        RECT 556.950 417.600 559.050 418.050 ;
        RECT 547.950 416.400 559.050 417.600 ;
        RECT 547.950 416.100 550.050 416.400 ;
        RECT 556.950 415.950 559.050 416.400 ;
        RECT 565.950 415.950 568.050 418.050 ;
        RECT 571.950 417.750 574.050 418.200 ;
        RECT 580.950 417.750 583.050 418.200 ;
        RECT 571.950 416.550 583.050 417.750 ;
        RECT 571.950 416.100 574.050 416.550 ;
        RECT 580.950 416.100 583.050 416.550 ;
        RECT 400.950 411.600 403.050 411.900 ;
        RECT 392.400 410.400 403.050 411.600 ;
        RECT 322.950 408.600 325.050 409.050 ;
        RECT 361.950 408.600 364.050 409.050 ;
        RECT 322.950 407.400 364.050 408.600 ;
        RECT 322.950 406.950 325.050 407.400 ;
        RECT 361.950 406.950 364.050 407.400 ;
        RECT 376.950 408.600 379.050 409.050 ;
        RECT 392.400 408.600 393.600 410.400 ;
        RECT 400.950 409.800 403.050 410.400 ;
        RECT 406.950 411.450 409.050 411.900 ;
        RECT 415.950 411.450 418.050 411.900 ;
        RECT 406.950 410.250 418.050 411.450 ;
        RECT 406.950 409.800 409.050 410.250 ;
        RECT 415.950 409.800 418.050 410.250 ;
        RECT 427.950 411.600 430.050 411.900 ;
        RECT 433.950 411.600 436.050 412.050 ;
        RECT 427.950 410.400 436.050 411.600 ;
        RECT 427.950 409.800 430.050 410.400 ;
        RECT 433.950 409.950 436.050 410.400 ;
        RECT 448.950 411.450 451.050 411.900 ;
        RECT 484.950 411.450 487.050 411.900 ;
        RECT 448.950 410.250 487.050 411.450 ;
        RECT 448.950 409.800 451.050 410.250 ;
        RECT 484.950 409.800 487.050 410.250 ;
        RECT 499.950 410.400 504.600 412.050 ;
        RECT 566.400 411.600 567.600 415.950 ;
        RECT 596.400 412.050 597.600 418.950 ;
        RECT 613.950 415.950 616.050 418.050 ;
        RECT 622.950 417.600 625.050 418.050 ;
        RECT 628.950 417.600 631.050 418.200 ;
        RECT 622.950 416.400 631.050 417.600 ;
        RECT 622.950 415.950 625.050 416.400 ;
        RECT 628.950 416.100 631.050 416.400 ;
        RECT 634.950 417.600 637.050 418.200 ;
        RECT 640.950 417.600 643.050 418.050 ;
        RECT 667.950 417.600 670.050 418.050 ;
        RECT 676.950 417.600 679.050 418.200 ;
        RECT 634.950 416.400 639.600 417.600 ;
        RECT 634.950 416.100 637.050 416.400 ;
        RECT 568.950 411.600 571.050 411.900 ;
        RECT 566.400 410.400 571.050 411.600 ;
        RECT 499.950 409.950 504.000 410.400 ;
        RECT 568.950 409.800 571.050 410.400 ;
        RECT 574.950 411.450 577.050 411.900 ;
        RECT 580.950 411.450 583.050 412.050 ;
        RECT 586.950 411.450 589.050 411.900 ;
        RECT 574.950 410.250 589.050 411.450 ;
        RECT 596.400 410.400 601.050 412.050 ;
        RECT 574.950 409.800 577.050 410.250 ;
        RECT 580.950 409.950 583.050 410.250 ;
        RECT 586.950 409.800 589.050 410.250 ;
        RECT 597.000 409.950 601.050 410.400 ;
        RECT 610.950 411.600 613.050 411.900 ;
        RECT 614.400 411.600 615.600 415.950 ;
        RECT 610.950 410.400 615.600 411.600 ;
        RECT 638.400 412.050 639.600 416.400 ;
        RECT 640.950 416.400 657.600 417.600 ;
        RECT 640.950 415.950 643.050 416.400 ;
        RECT 638.400 410.400 643.050 412.050 ;
        RECT 656.400 411.900 657.600 416.400 ;
        RECT 667.950 416.400 679.050 417.600 ;
        RECT 667.950 415.950 670.050 416.400 ;
        RECT 676.950 416.100 679.050 416.400 ;
        RECT 703.950 415.950 706.050 418.050 ;
        RECT 715.950 417.600 718.050 418.200 ;
        RECT 713.400 416.400 718.050 417.600 ;
        RECT 704.400 412.050 705.600 415.950 ;
        RECT 713.400 412.050 714.600 416.400 ;
        RECT 715.950 416.100 718.050 416.400 ;
        RECT 724.950 415.950 727.050 418.050 ;
        RECT 725.400 412.050 726.600 415.950 ;
        RECT 610.950 409.800 613.050 410.400 ;
        RECT 639.000 409.950 643.050 410.400 ;
        RECT 655.950 409.800 658.050 411.900 ;
        RECT 685.950 411.600 688.050 412.050 ;
        RECT 697.950 411.600 700.050 411.900 ;
        RECT 685.950 410.400 700.050 411.600 ;
        RECT 685.950 409.950 688.050 410.400 ;
        RECT 697.950 409.800 700.050 410.400 ;
        RECT 703.950 409.950 706.050 412.050 ;
        RECT 712.950 409.950 715.050 412.050 ;
        RECT 724.950 409.950 727.050 412.050 ;
        RECT 740.400 411.600 741.600 419.400 ;
        RECT 754.950 417.600 757.050 421.050 ;
        RECT 772.950 420.600 775.050 421.050 ;
        RECT 761.400 420.000 775.050 420.600 ;
        RECT 760.950 419.400 775.050 420.000 ;
        RECT 754.950 417.000 759.600 417.600 ;
        RECT 755.400 416.400 759.600 417.000 ;
        RECT 758.400 412.050 759.600 416.400 ;
        RECT 760.950 415.950 763.050 419.400 ;
        RECT 772.950 418.950 775.050 419.400 ;
        RECT 817.950 420.600 820.050 421.050 ;
        RECT 832.950 420.600 835.050 420.900 ;
        RECT 841.950 420.600 844.050 421.050 ;
        RECT 817.950 419.400 844.050 420.600 ;
        RECT 817.950 418.950 820.050 419.400 ;
        RECT 832.950 418.800 835.050 419.400 ;
        RECT 841.950 418.950 844.050 419.400 ;
        RECT 787.950 417.600 790.050 418.050 ;
        RECT 764.400 416.400 790.050 417.600 ;
        RECT 736.950 410.400 741.600 411.600 ;
        RECT 736.950 409.500 739.050 410.400 ;
        RECT 757.950 409.950 760.050 412.050 ;
        RECT 376.950 407.400 393.600 408.600 ;
        RECT 496.950 408.600 499.050 409.050 ;
        RECT 520.950 408.600 523.050 409.050 ;
        RECT 496.950 407.400 523.050 408.600 ;
        RECT 376.950 406.950 379.050 407.400 ;
        RECT 496.950 406.950 499.050 407.400 ;
        RECT 520.950 406.950 523.050 407.400 ;
        RECT 721.950 408.600 724.050 409.050 ;
        RECT 727.950 408.600 730.050 409.050 ;
        RECT 742.950 408.600 745.050 409.050 ;
        RECT 764.400 408.900 765.600 416.400 ;
        RECT 787.950 415.950 790.050 416.400 ;
        RECT 793.950 417.600 796.050 418.200 ;
        RECT 802.950 417.600 805.050 417.900 ;
        RECT 820.950 417.600 823.050 418.200 ;
        RECT 793.950 416.400 805.050 417.600 ;
        RECT 793.950 416.100 796.050 416.400 ;
        RECT 802.950 415.800 805.050 416.400 ;
        RECT 812.400 416.400 823.050 417.600 ;
        RECT 812.400 412.050 813.600 416.400 ;
        RECT 820.950 416.100 823.050 416.400 ;
        RECT 883.950 415.950 886.050 418.050 ;
        RECT 772.950 411.600 775.050 411.900 ;
        RECT 796.950 411.600 799.050 411.900 ;
        RECT 772.950 410.400 799.050 411.600 ;
        RECT 772.950 409.800 775.050 410.400 ;
        RECT 796.950 409.800 799.050 410.400 ;
        RECT 811.950 409.950 814.050 412.050 ;
        RECT 823.950 411.450 826.050 411.900 ;
        RECT 832.950 411.450 835.050 411.900 ;
        RECT 823.950 410.250 835.050 411.450 ;
        RECT 823.950 409.800 826.050 410.250 ;
        RECT 832.950 409.800 835.050 410.250 ;
        RECT 871.950 411.600 874.050 412.050 ;
        RECT 880.950 411.600 883.050 411.900 ;
        RECT 871.950 410.400 883.050 411.600 ;
        RECT 884.400 411.600 885.600 415.950 ;
        RECT 901.950 411.600 904.050 411.900 ;
        RECT 884.400 410.400 904.050 411.600 ;
        RECT 871.950 409.950 874.050 410.400 ;
        RECT 880.950 409.800 883.050 410.400 ;
        RECT 901.950 409.800 904.050 410.400 ;
        RECT 721.950 407.400 745.050 408.600 ;
        RECT 721.950 406.950 724.050 407.400 ;
        RECT 727.950 406.950 730.050 407.400 ;
        RECT 742.950 406.950 745.050 407.400 ;
        RECT 763.950 406.800 766.050 408.900 ;
        RECT 797.400 408.600 798.600 409.800 ;
        RECT 823.950 408.600 826.050 409.050 ;
        RECT 797.400 407.400 826.050 408.600 ;
        RECT 823.950 406.950 826.050 407.400 ;
        RECT 838.950 408.600 841.050 409.050 ;
        RECT 853.950 408.600 856.050 409.050 ;
        RECT 838.950 407.400 856.050 408.600 ;
        RECT 838.950 406.950 841.050 407.400 ;
        RECT 853.950 406.950 856.050 407.400 ;
        RECT 76.950 405.600 79.050 406.050 ;
        RECT 136.950 405.600 139.050 406.050 ;
        RECT 76.950 404.400 139.050 405.600 ;
        RECT 76.950 403.950 79.050 404.400 ;
        RECT 136.950 403.950 139.050 404.400 ;
        RECT 217.950 405.600 220.050 406.050 ;
        RECT 247.950 405.600 250.050 406.050 ;
        RECT 217.950 404.400 250.050 405.600 ;
        RECT 217.950 403.950 220.050 404.400 ;
        RECT 247.950 403.950 250.050 404.400 ;
        RECT 274.950 405.600 277.050 406.050 ;
        RECT 283.950 405.600 286.050 406.050 ;
        RECT 274.950 404.400 286.050 405.600 ;
        RECT 274.950 403.950 277.050 404.400 ;
        RECT 283.950 403.950 286.050 404.400 ;
        RECT 337.950 405.600 340.050 406.050 ;
        RECT 364.950 405.600 367.050 406.050 ;
        RECT 337.950 404.400 367.050 405.600 ;
        RECT 337.950 403.950 340.050 404.400 ;
        RECT 364.950 403.950 367.050 404.400 ;
        RECT 379.950 405.600 382.050 406.050 ;
        RECT 412.950 405.600 415.050 406.050 ;
        RECT 379.950 404.400 415.050 405.600 ;
        RECT 379.950 403.950 382.050 404.400 ;
        RECT 412.950 403.950 415.050 404.400 ;
        RECT 421.950 405.600 424.050 406.050 ;
        RECT 436.950 405.600 439.050 406.050 ;
        RECT 442.950 405.600 445.050 406.050 ;
        RECT 421.950 404.400 445.050 405.600 ;
        RECT 421.950 403.950 424.050 404.400 ;
        RECT 436.950 403.950 439.050 404.400 ;
        RECT 442.950 403.950 445.050 404.400 ;
        RECT 577.950 405.600 580.050 406.050 ;
        RECT 589.950 405.600 592.050 406.050 ;
        RECT 577.950 404.400 592.050 405.600 ;
        RECT 577.950 403.950 580.050 404.400 ;
        RECT 589.950 403.950 592.050 404.400 ;
        RECT 604.950 405.600 607.050 406.050 ;
        RECT 631.950 405.600 634.050 406.050 ;
        RECT 604.950 404.400 634.050 405.600 ;
        RECT 604.950 403.950 607.050 404.400 ;
        RECT 631.950 403.950 634.050 404.400 ;
        RECT 661.950 405.600 664.050 406.050 ;
        RECT 685.950 405.600 688.050 406.050 ;
        RECT 718.950 405.600 721.050 406.050 ;
        RECT 661.950 404.400 688.050 405.600 ;
        RECT 661.950 403.950 664.050 404.400 ;
        RECT 685.950 403.950 688.050 404.400 ;
        RECT 689.400 404.400 721.050 405.600 ;
        RECT 1.950 402.600 4.050 403.050 ;
        RECT 22.950 402.600 25.050 403.050 ;
        RECT 1.950 401.400 25.050 402.600 ;
        RECT 1.950 400.950 4.050 401.400 ;
        RECT 22.950 400.950 25.050 401.400 ;
        RECT 43.950 402.600 46.050 403.050 ;
        RECT 49.950 402.600 52.050 403.050 ;
        RECT 43.950 401.400 52.050 402.600 ;
        RECT 43.950 400.950 46.050 401.400 ;
        RECT 49.950 400.950 52.050 401.400 ;
        RECT 148.950 402.600 151.050 403.050 ;
        RECT 160.950 402.600 163.050 403.050 ;
        RECT 172.950 402.600 175.050 403.050 ;
        RECT 211.950 402.600 214.050 403.050 ;
        RECT 148.950 401.400 214.050 402.600 ;
        RECT 148.950 400.950 151.050 401.400 ;
        RECT 160.950 400.950 163.050 401.400 ;
        RECT 172.950 400.950 175.050 401.400 ;
        RECT 211.950 400.950 214.050 401.400 ;
        RECT 301.950 402.600 304.050 403.050 ;
        RECT 367.950 402.600 370.050 403.050 ;
        RECT 373.950 402.600 376.050 403.050 ;
        RECT 301.950 401.400 376.050 402.600 ;
        RECT 301.950 400.950 304.050 401.400 ;
        RECT 367.950 400.950 370.050 401.400 ;
        RECT 373.950 400.950 376.050 401.400 ;
        RECT 382.950 402.600 385.050 403.050 ;
        RECT 394.950 402.600 397.050 403.050 ;
        RECT 382.950 401.400 397.050 402.600 ;
        RECT 382.950 400.950 385.050 401.400 ;
        RECT 394.950 400.950 397.050 401.400 ;
        RECT 445.950 402.600 448.050 403.050 ;
        RECT 490.950 402.600 493.050 403.050 ;
        RECT 445.950 401.400 493.050 402.600 ;
        RECT 445.950 400.950 448.050 401.400 ;
        RECT 490.950 400.950 493.050 401.400 ;
        RECT 541.950 402.600 544.050 403.050 ;
        RECT 562.950 402.600 565.050 403.050 ;
        RECT 541.950 401.400 565.050 402.600 ;
        RECT 541.950 400.950 544.050 401.400 ;
        RECT 562.950 400.950 565.050 401.400 ;
        RECT 637.950 402.600 640.050 403.050 ;
        RECT 689.400 402.600 690.600 404.400 ;
        RECT 718.950 403.950 721.050 404.400 ;
        RECT 778.950 405.600 781.050 406.050 ;
        RECT 802.950 405.600 805.050 406.050 ;
        RECT 778.950 404.400 805.050 405.600 ;
        RECT 778.950 403.950 781.050 404.400 ;
        RECT 802.950 403.950 805.050 404.400 ;
        RECT 721.950 402.600 724.050 403.050 ;
        RECT 637.950 401.400 690.600 402.600 ;
        RECT 704.400 401.400 724.050 402.600 ;
        RECT 637.950 400.950 640.050 401.400 ;
        RECT 100.950 399.600 103.050 400.050 ;
        RECT 277.950 399.600 280.050 400.050 ;
        RECT 283.950 399.600 286.050 400.050 ;
        RECT 100.950 398.400 267.600 399.600 ;
        RECT 100.950 397.950 103.050 398.400 ;
        RECT 31.950 396.600 34.050 397.050 ;
        RECT 244.950 396.600 247.050 397.050 ;
        RECT 31.950 395.400 247.050 396.600 ;
        RECT 266.400 396.600 267.600 398.400 ;
        RECT 277.950 398.400 286.050 399.600 ;
        RECT 277.950 397.950 280.050 398.400 ;
        RECT 283.950 397.950 286.050 398.400 ;
        RECT 322.950 399.600 325.050 400.050 ;
        RECT 385.950 399.600 388.050 400.050 ;
        RECT 403.950 399.600 406.050 400.050 ;
        RECT 322.950 398.400 388.050 399.600 ;
        RECT 389.400 399.000 406.050 399.600 ;
        RECT 322.950 397.950 325.050 398.400 ;
        RECT 385.950 397.950 388.050 398.400 ;
        RECT 388.950 398.400 406.050 399.000 ;
        RECT 340.950 396.600 343.050 397.050 ;
        RECT 355.950 396.600 358.050 397.050 ;
        RECT 266.400 395.400 358.050 396.600 ;
        RECT 31.950 394.950 34.050 395.400 ;
        RECT 244.950 394.950 247.050 395.400 ;
        RECT 340.950 394.950 343.050 395.400 ;
        RECT 355.950 394.950 358.050 395.400 ;
        RECT 388.950 394.950 391.050 398.400 ;
        RECT 403.950 397.950 406.050 398.400 ;
        RECT 418.950 399.600 421.050 400.050 ;
        RECT 433.950 399.600 436.050 400.050 ;
        RECT 418.950 398.400 436.050 399.600 ;
        RECT 418.950 397.950 421.050 398.400 ;
        RECT 433.950 397.950 436.050 398.400 ;
        RECT 442.950 399.600 445.050 400.050 ;
        RECT 463.950 399.600 466.050 400.050 ;
        RECT 442.950 398.400 466.050 399.600 ;
        RECT 442.950 397.950 445.050 398.400 ;
        RECT 463.950 397.950 466.050 398.400 ;
        RECT 577.950 399.600 580.050 400.050 ;
        RECT 598.950 399.600 601.050 400.050 ;
        RECT 704.400 399.600 705.600 401.400 ;
        RECT 721.950 400.950 724.050 401.400 ;
        RECT 736.950 402.600 739.050 403.050 ;
        RECT 742.950 402.600 745.050 403.050 ;
        RECT 736.950 401.400 745.050 402.600 ;
        RECT 736.950 400.950 739.050 401.400 ;
        RECT 742.950 400.950 745.050 401.400 ;
        RECT 577.950 398.400 705.600 399.600 ;
        RECT 838.950 399.600 841.050 400.050 ;
        RECT 847.950 399.600 850.050 400.050 ;
        RECT 901.950 399.600 904.050 400.050 ;
        RECT 910.950 399.600 913.050 400.050 ;
        RECT 838.950 398.400 913.050 399.600 ;
        RECT 577.950 397.950 580.050 398.400 ;
        RECT 598.950 397.950 601.050 398.400 ;
        RECT 838.950 397.950 841.050 398.400 ;
        RECT 847.950 397.950 850.050 398.400 ;
        RECT 901.950 397.950 904.050 398.400 ;
        RECT 910.950 397.950 913.050 398.400 ;
        RECT 406.950 396.600 409.050 397.050 ;
        RECT 496.950 396.600 499.050 397.050 ;
        RECT 406.950 395.400 499.050 396.600 ;
        RECT 406.950 394.950 409.050 395.400 ;
        RECT 496.950 394.950 499.050 395.400 ;
        RECT 505.950 396.600 508.050 397.050 ;
        RECT 544.950 396.600 547.050 397.050 ;
        RECT 505.950 395.400 547.050 396.600 ;
        RECT 505.950 394.950 508.050 395.400 ;
        RECT 544.950 394.950 547.050 395.400 ;
        RECT 706.950 396.600 709.050 397.050 ;
        RECT 742.950 396.600 745.050 397.050 ;
        RECT 706.950 395.400 745.050 396.600 ;
        RECT 706.950 394.950 709.050 395.400 ;
        RECT 742.950 394.950 745.050 395.400 ;
        RECT 817.950 396.600 820.050 397.050 ;
        RECT 871.950 396.600 874.050 397.050 ;
        RECT 817.950 395.400 874.050 396.600 ;
        RECT 817.950 394.950 820.050 395.400 ;
        RECT 871.950 394.950 874.050 395.400 ;
        RECT 97.950 393.600 100.050 394.050 ;
        RECT 109.950 393.600 112.050 394.050 ;
        RECT 97.950 392.400 112.050 393.600 ;
        RECT 97.950 391.950 100.050 392.400 ;
        RECT 109.950 391.950 112.050 392.400 ;
        RECT 121.950 393.600 124.050 394.050 ;
        RECT 190.950 393.600 193.050 394.050 ;
        RECT 121.950 392.400 193.050 393.600 ;
        RECT 121.950 391.950 124.050 392.400 ;
        RECT 190.950 391.950 193.050 392.400 ;
        RECT 304.950 393.600 307.050 394.050 ;
        RECT 331.950 393.600 334.050 394.050 ;
        RECT 304.950 392.400 334.050 393.600 ;
        RECT 304.950 391.950 307.050 392.400 ;
        RECT 331.950 391.950 334.050 392.400 ;
        RECT 382.950 393.600 385.050 394.050 ;
        RECT 403.950 393.600 406.050 394.050 ;
        RECT 382.950 392.400 406.050 393.600 ;
        RECT 382.950 391.950 385.050 392.400 ;
        RECT 403.950 391.950 406.050 392.400 ;
        RECT 625.950 393.600 628.050 394.050 ;
        RECT 667.950 393.600 670.050 394.050 ;
        RECT 625.950 392.400 670.050 393.600 ;
        RECT 625.950 391.950 628.050 392.400 ;
        RECT 667.950 391.950 670.050 392.400 ;
        RECT 694.950 393.600 697.050 394.050 ;
        RECT 769.950 393.600 772.050 394.050 ;
        RECT 784.950 393.600 787.050 394.050 ;
        RECT 694.950 392.400 787.050 393.600 ;
        RECT 694.950 391.950 697.050 392.400 ;
        RECT 769.950 391.950 772.050 392.400 ;
        RECT 784.950 391.950 787.050 392.400 ;
        RECT 886.950 393.600 889.050 394.050 ;
        RECT 901.950 393.600 904.050 394.050 ;
        RECT 886.950 392.400 904.050 393.600 ;
        RECT 886.950 391.950 889.050 392.400 ;
        RECT 901.950 391.950 904.050 392.400 ;
        RECT 7.950 390.600 10.050 391.050 ;
        RECT 76.950 390.600 79.050 391.050 ;
        RECT 7.950 389.400 79.050 390.600 ;
        RECT 7.950 388.950 10.050 389.400 ;
        RECT 76.950 388.950 79.050 389.400 ;
        RECT 130.950 390.600 133.050 391.050 ;
        RECT 196.950 390.600 199.050 391.050 ;
        RECT 130.950 389.400 199.050 390.600 ;
        RECT 130.950 388.950 133.050 389.400 ;
        RECT 196.950 388.950 199.050 389.400 ;
        RECT 253.950 390.600 256.050 391.050 ;
        RECT 271.950 390.600 274.050 391.050 ;
        RECT 253.950 389.400 274.050 390.600 ;
        RECT 253.950 388.950 256.050 389.400 ;
        RECT 271.950 388.950 274.050 389.400 ;
        RECT 277.950 390.600 280.050 391.050 ;
        RECT 286.950 390.600 289.050 391.050 ;
        RECT 277.950 389.400 289.050 390.600 ;
        RECT 277.950 388.950 280.050 389.400 ;
        RECT 286.950 388.950 289.050 389.400 ;
        RECT 310.950 390.600 313.050 391.050 ;
        RECT 346.950 390.600 349.050 391.050 ;
        RECT 310.950 389.400 349.050 390.600 ;
        RECT 310.950 388.950 313.050 389.400 ;
        RECT 346.950 388.950 349.050 389.400 ;
        RECT 361.950 390.600 364.050 391.050 ;
        RECT 427.950 390.600 430.050 391.050 ;
        RECT 361.950 389.400 430.050 390.600 ;
        RECT 361.950 388.950 364.050 389.400 ;
        RECT 427.950 388.950 430.050 389.400 ;
        RECT 466.950 390.600 469.050 391.050 ;
        RECT 493.950 390.600 496.050 391.050 ;
        RECT 466.950 389.400 496.050 390.600 ;
        RECT 466.950 388.950 469.050 389.400 ;
        RECT 493.950 388.950 496.050 389.400 ;
        RECT 505.950 390.600 508.050 391.050 ;
        RECT 535.950 390.600 538.050 391.050 ;
        RECT 505.950 389.400 538.050 390.600 ;
        RECT 505.950 388.950 508.050 389.400 ;
        RECT 535.950 388.950 538.050 389.400 ;
        RECT 562.950 390.600 565.050 391.050 ;
        RECT 691.950 390.600 694.050 391.050 ;
        RECT 562.950 389.400 694.050 390.600 ;
        RECT 562.950 388.950 565.050 389.400 ;
        RECT 691.950 388.950 694.050 389.400 ;
        RECT 739.950 390.600 742.050 391.050 ;
        RECT 760.950 390.600 763.050 391.050 ;
        RECT 739.950 389.400 763.050 390.600 ;
        RECT 739.950 388.950 742.050 389.400 ;
        RECT 760.950 388.950 763.050 389.400 ;
        RECT 880.950 390.600 883.050 391.050 ;
        RECT 919.950 390.600 922.050 391.050 ;
        RECT 880.950 389.400 922.050 390.600 ;
        RECT 880.950 388.950 883.050 389.400 ;
        RECT 919.950 388.950 922.050 389.400 ;
        RECT 1.950 387.600 4.050 388.050 ;
        RECT 106.950 387.600 109.050 388.050 ;
        RECT 1.950 386.400 109.050 387.600 ;
        RECT 1.950 385.950 4.050 386.400 ;
        RECT 106.950 385.950 109.050 386.400 ;
        RECT 208.950 387.600 211.050 388.050 ;
        RECT 232.950 387.600 235.050 388.050 ;
        RECT 208.950 386.400 235.050 387.600 ;
        RECT 208.950 385.950 211.050 386.400 ;
        RECT 232.950 385.950 235.050 386.400 ;
        RECT 247.950 387.600 250.050 388.050 ;
        RECT 268.950 387.600 271.050 388.050 ;
        RECT 247.950 386.400 271.050 387.600 ;
        RECT 247.950 385.950 250.050 386.400 ;
        RECT 268.950 385.950 271.050 386.400 ;
        RECT 319.950 387.600 322.050 388.050 ;
        RECT 361.950 387.600 364.050 387.900 ;
        RECT 319.950 386.400 364.050 387.600 ;
        RECT 319.950 385.950 322.050 386.400 ;
        RECT 361.950 385.800 364.050 386.400 ;
        RECT 403.950 387.600 406.050 388.050 ;
        RECT 418.950 387.600 421.050 388.050 ;
        RECT 403.950 386.400 421.050 387.600 ;
        RECT 403.950 385.950 406.050 386.400 ;
        RECT 418.950 385.950 421.050 386.400 ;
        RECT 439.950 387.600 442.050 388.050 ;
        RECT 457.950 387.600 460.050 388.050 ;
        RECT 439.950 386.400 460.050 387.600 ;
        RECT 439.950 385.950 442.050 386.400 ;
        RECT 457.950 385.950 460.050 386.400 ;
        RECT 610.950 387.600 613.050 388.050 ;
        RECT 649.950 387.600 652.050 388.050 ;
        RECT 658.950 387.600 661.050 388.050 ;
        RECT 610.950 386.400 661.050 387.600 ;
        RECT 610.950 385.950 613.050 386.400 ;
        RECT 649.950 385.950 652.050 386.400 ;
        RECT 658.950 385.950 661.050 386.400 ;
        RECT 862.950 387.600 865.050 388.050 ;
        RECT 886.950 387.600 889.050 388.050 ;
        RECT 862.950 386.400 889.050 387.600 ;
        RECT 862.950 385.950 865.050 386.400 ;
        RECT 886.950 385.950 889.050 386.400 ;
        RECT 898.950 387.600 901.050 388.050 ;
        RECT 907.950 387.600 910.050 388.050 ;
        RECT 898.950 386.400 910.050 387.600 ;
        RECT 898.950 385.950 901.050 386.400 ;
        RECT 907.950 385.950 910.050 386.400 ;
        RECT 40.950 384.600 43.050 385.050 ;
        RECT 70.950 384.600 73.050 385.050 ;
        RECT 94.950 384.600 97.050 385.050 ;
        RECT 40.950 383.400 97.050 384.600 ;
        RECT 40.950 382.950 43.050 383.400 ;
        RECT 70.950 382.950 73.050 383.400 ;
        RECT 94.950 382.950 97.050 383.400 ;
        RECT 106.950 384.600 109.050 384.900 ;
        RECT 124.950 384.600 127.050 385.050 ;
        RECT 106.950 383.400 127.050 384.600 ;
        RECT 106.950 382.800 109.050 383.400 ;
        RECT 124.950 382.950 127.050 383.400 ;
        RECT 145.950 384.600 148.050 385.050 ;
        RECT 205.950 384.600 208.050 385.050 ;
        RECT 235.950 384.600 238.050 385.050 ;
        RECT 145.950 383.400 238.050 384.600 ;
        RECT 145.950 382.950 148.050 383.400 ;
        RECT 205.950 382.950 208.050 383.400 ;
        RECT 235.950 382.950 238.050 383.400 ;
        RECT 271.950 384.600 274.050 385.050 ;
        RECT 334.950 384.600 337.050 385.050 ;
        RECT 271.950 383.400 337.050 384.600 ;
        RECT 271.950 382.950 274.050 383.400 ;
        RECT 334.950 382.950 337.050 383.400 ;
        RECT 364.950 384.600 367.050 385.050 ;
        RECT 400.950 384.600 403.050 385.050 ;
        RECT 364.950 383.400 403.050 384.600 ;
        RECT 364.950 382.950 367.050 383.400 ;
        RECT 400.950 382.950 403.050 383.400 ;
        RECT 427.950 384.600 430.050 385.050 ;
        RECT 499.950 384.600 502.050 385.050 ;
        RECT 427.950 383.400 502.050 384.600 ;
        RECT 427.950 382.950 430.050 383.400 ;
        RECT 499.950 382.950 502.050 383.400 ;
        RECT 565.950 384.600 568.050 385.050 ;
        RECT 592.950 384.600 595.050 385.050 ;
        RECT 658.950 384.600 661.050 384.900 ;
        RECT 673.950 384.600 676.050 385.050 ;
        RECT 712.950 384.600 715.050 385.050 ;
        RECT 748.950 384.600 751.050 385.050 ;
        RECT 565.950 383.400 751.050 384.600 ;
        RECT 565.950 382.950 568.050 383.400 ;
        RECT 592.950 382.950 595.050 383.400 ;
        RECT 658.950 382.800 661.050 383.400 ;
        RECT 673.950 382.950 676.050 383.400 ;
        RECT 712.950 382.950 715.050 383.400 ;
        RECT 748.950 382.950 751.050 383.400 ;
        RECT 781.950 384.600 784.050 385.050 ;
        RECT 799.950 384.600 802.050 385.050 ;
        RECT 781.950 383.400 802.050 384.600 ;
        RECT 781.950 382.950 784.050 383.400 ;
        RECT 799.950 382.950 802.050 383.400 ;
        RECT 805.950 384.600 808.050 385.050 ;
        RECT 829.950 384.600 832.050 385.050 ;
        RECT 874.950 384.600 877.050 385.050 ;
        RECT 805.950 383.400 832.050 384.600 ;
        RECT 805.950 382.950 808.050 383.400 ;
        RECT 829.950 382.950 832.050 383.400 ;
        RECT 866.400 383.400 877.050 384.600 ;
        RECT 866.400 382.050 867.600 383.400 ;
        RECT 874.950 382.950 877.050 383.400 ;
        RECT 37.950 381.600 40.050 382.050 ;
        RECT 133.950 381.600 136.050 382.050 ;
        RECT 37.950 380.400 136.050 381.600 ;
        RECT 37.950 379.950 40.050 380.400 ;
        RECT 133.950 379.950 136.050 380.400 ;
        RECT 154.950 381.600 157.050 382.050 ;
        RECT 166.950 381.600 169.050 382.050 ;
        RECT 154.950 380.400 169.050 381.600 ;
        RECT 154.950 379.950 157.050 380.400 ;
        RECT 166.950 379.950 169.050 380.400 ;
        RECT 175.950 381.600 178.050 382.050 ;
        RECT 238.950 381.600 241.050 382.050 ;
        RECT 262.950 381.600 265.050 382.050 ;
        RECT 175.950 380.400 213.600 381.600 ;
        RECT 175.950 379.950 178.050 380.400 ;
        RECT 212.400 379.050 213.600 380.400 ;
        RECT 238.950 380.400 265.050 381.600 ;
        RECT 238.950 379.950 241.050 380.400 ;
        RECT 262.950 379.950 265.050 380.400 ;
        RECT 274.950 381.600 277.050 382.050 ;
        RECT 319.950 381.600 322.050 382.050 ;
        RECT 274.950 380.400 322.050 381.600 ;
        RECT 274.950 379.950 277.050 380.400 ;
        RECT 319.950 379.950 322.050 380.400 ;
        RECT 343.950 381.600 346.050 382.050 ;
        RECT 376.950 381.600 379.050 382.050 ;
        RECT 343.950 380.400 379.050 381.600 ;
        RECT 343.950 379.950 346.050 380.400 ;
        RECT 376.950 379.950 379.050 380.400 ;
        RECT 490.950 381.600 493.050 382.050 ;
        RECT 502.950 381.600 505.050 382.050 ;
        RECT 490.950 380.400 505.050 381.600 ;
        RECT 490.950 379.950 493.050 380.400 ;
        RECT 502.950 379.950 505.050 380.400 ;
        RECT 511.950 381.600 514.050 382.050 ;
        RECT 562.950 381.600 565.050 382.050 ;
        RECT 511.950 380.400 565.050 381.600 ;
        RECT 511.950 379.950 514.050 380.400 ;
        RECT 562.950 379.950 565.050 380.400 ;
        RECT 601.950 381.600 604.050 382.050 ;
        RECT 613.950 381.600 616.050 382.050 ;
        RECT 601.950 380.400 616.050 381.600 ;
        RECT 601.950 379.950 604.050 380.400 ;
        RECT 613.950 379.950 616.050 380.400 ;
        RECT 646.950 381.600 649.050 382.050 ;
        RECT 667.950 381.600 670.050 382.050 ;
        RECT 646.950 380.400 670.050 381.600 ;
        RECT 646.950 379.950 649.050 380.400 ;
        RECT 667.950 379.950 670.050 380.400 ;
        RECT 691.950 381.600 694.050 382.050 ;
        RECT 745.950 381.600 748.050 382.050 ;
        RECT 691.950 380.400 748.050 381.600 ;
        RECT 691.950 379.950 694.050 380.400 ;
        RECT 745.950 379.950 748.050 380.400 ;
        RECT 787.950 381.600 790.050 382.050 ;
        RECT 814.950 381.600 817.050 382.050 ;
        RECT 865.950 381.600 868.050 382.050 ;
        RECT 787.950 380.400 817.050 381.600 ;
        RECT 787.950 379.950 790.050 380.400 ;
        RECT 814.950 379.950 817.050 380.400 ;
        RECT 845.400 380.400 868.050 381.600 ;
        RECT 4.950 378.600 7.050 379.050 ;
        RECT 31.950 378.600 34.050 379.050 ;
        RECT 4.950 377.400 34.050 378.600 ;
        RECT 4.950 376.950 7.050 377.400 ;
        RECT 31.950 376.950 34.050 377.400 ;
        RECT 58.950 378.600 61.050 379.050 ;
        RECT 112.950 378.600 115.050 379.050 ;
        RECT 121.950 378.600 124.050 379.050 ;
        RECT 58.950 377.400 124.050 378.600 ;
        RECT 58.950 376.950 61.050 377.400 ;
        RECT 112.950 376.950 115.050 377.400 ;
        RECT 121.950 376.950 124.050 377.400 ;
        RECT 139.950 378.600 142.050 379.050 ;
        RECT 169.950 378.600 172.050 379.050 ;
        RECT 139.950 377.400 172.050 378.600 ;
        RECT 139.950 376.950 142.050 377.400 ;
        RECT 169.950 376.950 172.050 377.400 ;
        RECT 211.950 378.600 214.050 379.050 ;
        RECT 271.950 378.600 274.050 379.050 ;
        RECT 211.950 377.400 274.050 378.600 ;
        RECT 211.950 376.950 214.050 377.400 ;
        RECT 271.950 376.950 274.050 377.400 ;
        RECT 376.950 378.600 379.050 378.900 ;
        RECT 406.950 378.600 409.050 379.050 ;
        RECT 376.950 377.400 409.050 378.600 ;
        RECT 376.950 376.800 379.050 377.400 ;
        RECT 406.950 376.950 409.050 377.400 ;
        RECT 424.950 378.600 427.050 379.050 ;
        RECT 460.950 378.600 463.050 379.050 ;
        RECT 424.950 377.400 463.050 378.600 ;
        RECT 424.950 376.950 427.050 377.400 ;
        RECT 460.950 376.950 463.050 377.400 ;
        RECT 673.950 378.600 676.050 379.050 ;
        RECT 694.950 378.600 697.050 379.050 ;
        RECT 673.950 377.400 697.050 378.600 ;
        RECT 673.950 376.950 676.050 377.400 ;
        RECT 694.950 376.950 697.050 377.400 ;
        RECT 775.950 378.600 778.050 379.050 ;
        RECT 845.400 378.600 846.600 380.400 ;
        RECT 865.950 379.950 868.050 380.400 ;
        RECT 907.950 381.600 910.050 382.050 ;
        RECT 919.950 381.600 922.050 382.050 ;
        RECT 907.950 380.400 922.050 381.600 ;
        RECT 907.950 379.950 910.050 380.400 ;
        RECT 919.950 379.950 922.050 380.400 ;
        RECT 775.950 377.400 846.600 378.600 ;
        RECT 775.950 376.950 778.050 377.400 ;
        RECT 178.950 375.600 181.050 376.050 ;
        RECT 187.950 375.600 190.050 376.050 ;
        RECT 178.950 374.400 190.050 375.600 ;
        RECT 178.950 373.950 181.050 374.400 ;
        RECT 187.950 373.950 190.050 374.400 ;
        RECT 223.950 375.600 226.050 376.050 ;
        RECT 256.950 375.600 259.050 376.050 ;
        RECT 223.950 374.400 259.050 375.600 ;
        RECT 223.950 373.950 226.050 374.400 ;
        RECT 256.950 373.950 259.050 374.400 ;
        RECT 265.950 375.600 268.050 376.050 ;
        RECT 292.950 375.600 295.050 376.050 ;
        RECT 313.950 375.600 316.050 376.050 ;
        RECT 265.950 374.400 295.050 375.600 ;
        RECT 265.950 373.950 268.050 374.400 ;
        RECT 292.950 373.950 295.050 374.400 ;
        RECT 305.400 374.400 316.050 375.600 ;
        RECT 10.950 372.600 13.050 373.200 ;
        RECT 19.950 372.600 22.050 373.200 ;
        RECT 37.950 372.600 40.050 373.200 ;
        RECT 10.950 371.400 18.600 372.600 ;
        RECT 10.950 371.100 13.050 371.400 ;
        RECT 17.400 367.050 18.600 371.400 ;
        RECT 19.950 371.400 40.050 372.600 ;
        RECT 19.950 371.100 22.050 371.400 ;
        RECT 37.950 371.100 40.050 371.400 ;
        RECT 52.950 372.600 55.050 373.200 ;
        RECT 67.950 372.600 70.050 373.050 ;
        RECT 76.950 372.600 79.050 373.200 ;
        RECT 52.950 371.400 79.050 372.600 ;
        RECT 52.950 371.100 55.050 371.400 ;
        RECT 67.950 370.950 70.050 371.400 ;
        RECT 76.950 371.100 79.050 371.400 ;
        RECT 94.950 371.100 97.050 373.200 ;
        RECT 100.950 371.100 103.050 373.200 ;
        RECT 151.950 372.750 154.050 373.200 ;
        RECT 157.950 372.750 160.050 373.200 ;
        RECT 151.950 371.550 160.050 372.750 ;
        RECT 151.950 371.100 154.050 371.550 ;
        RECT 157.950 371.100 160.050 371.550 ;
        RECT 184.950 372.750 187.050 373.050 ;
        RECT 196.950 372.750 199.050 373.200 ;
        RECT 184.950 371.550 199.050 372.750 ;
        RECT 85.950 369.600 88.050 370.050 ;
        RECT 95.400 369.600 96.600 371.100 ;
        RECT 85.950 368.400 96.600 369.600 ;
        RECT 85.950 367.950 88.050 368.400 ;
        RECT 101.400 367.050 102.600 371.100 ;
        RECT 184.950 370.950 187.050 371.550 ;
        RECT 196.950 371.100 199.050 371.550 ;
        RECT 241.950 372.750 244.050 373.200 ;
        RECT 253.950 372.750 256.050 373.200 ;
        RECT 241.950 371.550 256.050 372.750 ;
        RECT 241.950 371.100 244.050 371.550 ;
        RECT 253.950 371.100 256.050 371.550 ;
        RECT 262.950 370.950 265.050 373.050 ;
        RECT 271.950 372.600 274.050 373.200 ;
        RECT 283.800 372.600 285.900 373.050 ;
        RECT 271.950 371.400 285.900 372.600 ;
        RECT 271.950 371.100 274.050 371.400 ;
        RECT 16.950 364.950 19.050 367.050 ;
        RECT 101.400 365.400 106.050 367.050 ;
        RECT 102.000 364.950 106.050 365.400 ;
        RECT 154.950 366.600 157.050 367.050 ;
        RECT 199.950 366.600 202.050 366.900 ;
        RECT 154.950 365.400 202.050 366.600 ;
        RECT 154.950 364.950 157.050 365.400 ;
        RECT 199.950 364.800 202.050 365.400 ;
        RECT 205.950 366.600 208.050 367.050 ;
        RECT 253.950 366.600 256.050 367.050 ;
        RECT 263.400 366.900 264.600 370.950 ;
        RECT 272.400 369.600 273.600 371.100 ;
        RECT 283.800 370.950 285.900 371.400 ;
        RECT 286.950 371.100 289.050 373.200 ;
        RECT 272.400 368.400 282.600 369.600 ;
        RECT 205.950 365.400 256.050 366.600 ;
        RECT 205.950 364.950 208.050 365.400 ;
        RECT 253.950 364.950 256.050 365.400 ;
        RECT 262.950 366.450 265.050 366.900 ;
        RECT 274.950 366.450 277.050 366.900 ;
        RECT 262.950 365.250 277.050 366.450 ;
        RECT 262.950 364.800 265.050 365.250 ;
        RECT 274.950 364.800 277.050 365.250 ;
        RECT 7.950 363.600 10.050 364.050 ;
        RECT 25.800 363.600 27.900 364.050 ;
        RECT 7.950 362.400 27.900 363.600 ;
        RECT 7.950 361.950 10.050 362.400 ;
        RECT 25.800 361.950 27.900 362.400 ;
        RECT 28.950 363.600 31.050 364.050 ;
        RECT 61.950 363.600 64.050 364.050 ;
        RECT 28.950 362.400 64.050 363.600 ;
        RECT 28.950 361.950 31.050 362.400 ;
        RECT 61.950 361.950 64.050 362.400 ;
        RECT 100.950 363.600 103.050 364.050 ;
        RECT 106.950 363.600 109.050 364.050 ;
        RECT 100.950 362.400 109.050 363.600 ;
        RECT 100.950 361.950 103.050 362.400 ;
        RECT 106.950 361.950 109.050 362.400 ;
        RECT 151.950 363.600 154.050 364.050 ;
        RECT 157.950 363.600 160.050 364.050 ;
        RECT 151.950 362.400 160.050 363.600 ;
        RECT 151.950 361.950 154.050 362.400 ;
        RECT 157.950 361.950 160.050 362.400 ;
        RECT 226.950 363.600 229.050 364.050 ;
        RECT 244.950 363.600 247.050 364.050 ;
        RECT 226.950 362.400 247.050 363.600 ;
        RECT 226.950 361.950 229.050 362.400 ;
        RECT 244.950 361.950 247.050 362.400 ;
        RECT 256.950 363.600 259.050 364.050 ;
        RECT 268.950 363.600 271.050 364.050 ;
        RECT 256.950 362.400 271.050 363.600 ;
        RECT 281.400 363.600 282.600 368.400 ;
        RECT 287.400 367.050 288.600 371.100 ;
        RECT 298.950 369.600 301.050 370.050 ;
        RECT 305.400 369.600 306.600 374.400 ;
        RECT 313.950 373.950 316.050 374.400 ;
        RECT 319.950 375.600 322.050 376.050 ;
        RECT 328.950 375.600 331.050 376.050 ;
        RECT 352.950 375.600 355.050 376.050 ;
        RECT 394.950 375.600 397.050 376.050 ;
        RECT 319.950 374.400 355.050 375.600 ;
        RECT 319.950 373.950 322.050 374.400 ;
        RECT 328.950 373.950 331.050 374.400 ;
        RECT 352.950 373.950 355.050 374.400 ;
        RECT 380.400 374.400 397.050 375.600 ;
        RECT 322.950 369.600 325.050 373.050 ;
        RECT 331.950 370.950 334.050 373.050 ;
        RECT 337.950 372.600 342.000 373.050 ;
        RECT 337.950 370.950 342.600 372.600 ;
        RECT 349.950 370.950 352.050 373.050 ;
        RECT 364.950 372.600 367.050 373.050 ;
        RECT 370.950 372.600 373.050 373.050 ;
        RECT 364.950 371.400 373.050 372.600 ;
        RECT 364.950 370.950 367.050 371.400 ;
        RECT 370.950 370.950 373.050 371.400 ;
        RECT 298.950 368.400 306.600 369.600 ;
        RECT 314.400 369.000 325.050 369.600 ;
        RECT 314.400 368.400 324.600 369.000 ;
        RECT 298.950 367.950 301.050 368.400 ;
        RECT 283.950 365.400 288.600 367.050 ;
        RECT 295.950 366.600 298.050 367.050 ;
        RECT 301.950 366.600 304.050 367.050 ;
        RECT 314.400 366.900 315.600 368.400 ;
        RECT 295.950 365.400 304.050 366.600 ;
        RECT 283.950 364.950 288.000 365.400 ;
        RECT 295.950 364.950 298.050 365.400 ;
        RECT 301.950 364.950 304.050 365.400 ;
        RECT 313.950 364.800 316.050 366.900 ;
        RECT 332.400 366.600 333.600 370.950 ;
        RECT 337.950 366.600 340.050 367.050 ;
        RECT 332.400 365.400 340.050 366.600 ;
        RECT 337.950 364.950 340.050 365.400 ;
        RECT 286.950 363.600 289.050 364.050 ;
        RECT 281.400 362.400 289.050 363.600 ;
        RECT 256.950 361.950 259.050 362.400 ;
        RECT 268.950 361.950 271.050 362.400 ;
        RECT 286.950 361.950 289.050 362.400 ;
        RECT 331.950 363.600 334.050 364.050 ;
        RECT 341.400 363.600 342.600 370.950 ;
        RECT 350.400 367.050 351.600 370.950 ;
        RECT 349.950 364.950 352.050 367.050 ;
        RECT 380.400 366.900 381.600 374.400 ;
        RECT 394.950 373.950 397.050 374.400 ;
        RECT 412.950 375.600 415.050 376.050 ;
        RECT 454.950 375.600 457.050 376.050 ;
        RECT 493.950 375.600 496.050 376.050 ;
        RECT 412.950 374.400 457.050 375.600 ;
        RECT 412.950 373.950 415.050 374.400 ;
        RECT 454.950 373.950 457.050 374.400 ;
        RECT 473.400 374.400 496.050 375.600 ;
        RECT 391.950 372.750 394.050 373.200 ;
        RECT 400.950 372.750 403.050 373.200 ;
        RECT 391.950 371.550 403.050 372.750 ;
        RECT 391.950 371.100 394.050 371.550 ;
        RECT 400.950 371.100 403.050 371.550 ;
        RECT 406.950 369.600 409.050 373.050 ;
        RECT 433.950 372.600 436.050 373.050 ;
        RECT 445.950 372.600 448.050 373.050 ;
        RECT 433.950 371.400 448.050 372.600 ;
        RECT 433.950 370.950 436.050 371.400 ;
        RECT 445.950 370.950 448.050 371.400 ;
        RECT 451.950 371.100 454.050 373.200 ;
        RECT 439.950 369.600 442.050 370.050 ;
        RECT 406.950 369.000 442.050 369.600 ;
        RECT 407.400 368.400 442.050 369.000 ;
        RECT 439.950 367.950 442.050 368.400 ;
        RECT 452.400 367.050 453.600 371.100 ;
        RECT 358.950 366.450 361.050 366.900 ;
        RECT 364.950 366.450 367.050 366.900 ;
        RECT 358.950 365.250 367.050 366.450 ;
        RECT 358.950 364.800 361.050 365.250 ;
        RECT 364.950 364.800 367.050 365.250 ;
        RECT 379.950 364.800 382.050 366.900 ;
        RECT 412.950 366.300 415.050 366.750 ;
        RECT 418.800 366.300 420.900 366.750 ;
        RECT 412.950 365.100 420.900 366.300 ;
        RECT 412.950 364.650 415.050 365.100 ;
        RECT 418.800 364.650 420.900 365.100 ;
        RECT 421.950 366.600 424.050 367.050 ;
        RECT 421.950 366.000 438.600 366.600 ;
        RECT 421.950 365.400 439.050 366.000 ;
        RECT 421.950 364.950 424.050 365.400 ;
        RECT 331.950 362.400 342.600 363.600 ;
        RECT 331.950 361.950 334.050 362.400 ;
        RECT 436.950 361.950 439.050 365.400 ;
        RECT 448.950 365.400 453.600 367.050 ;
        RECT 460.950 366.600 463.050 366.900 ;
        RECT 473.400 366.600 474.600 374.400 ;
        RECT 493.950 373.950 496.050 374.400 ;
        RECT 523.950 375.600 526.050 376.050 ;
        RECT 532.950 375.600 535.050 376.050 ;
        RECT 523.950 374.400 535.050 375.600 ;
        RECT 523.950 373.950 526.050 374.400 ;
        RECT 532.950 373.950 535.050 374.400 ;
        RECT 604.950 375.600 607.050 376.050 ;
        RECT 616.950 375.600 619.050 376.050 ;
        RECT 622.950 375.600 625.050 376.050 ;
        RECT 604.950 374.400 625.050 375.600 ;
        RECT 604.950 373.950 607.050 374.400 ;
        RECT 616.950 373.950 619.050 374.400 ;
        RECT 622.950 373.950 625.050 374.400 ;
        RECT 682.950 375.600 685.050 376.050 ;
        RECT 688.950 375.600 691.050 376.200 ;
        RECT 724.950 375.600 727.050 376.050 ;
        RECT 730.950 375.600 733.050 376.050 ;
        RECT 682.950 374.400 691.050 375.600 ;
        RECT 682.950 373.950 685.050 374.400 ;
        RECT 688.950 374.100 691.050 374.400 ;
        RECT 713.400 374.400 733.050 375.600 ;
        RECT 475.950 372.600 478.050 373.200 ;
        RECT 517.950 372.600 520.050 373.200 ;
        RECT 475.950 371.400 492.600 372.600 ;
        RECT 475.950 371.100 478.050 371.400 ;
        RECT 491.400 366.900 492.600 371.400 ;
        RECT 517.950 371.400 522.600 372.600 ;
        RECT 517.950 371.100 520.050 371.400 ;
        RECT 521.400 367.050 522.600 371.400 ;
        RECT 535.950 371.100 538.050 373.200 ;
        RECT 559.950 372.600 562.050 373.050 ;
        RECT 574.950 372.600 577.050 373.050 ;
        RECT 583.950 372.600 586.050 373.200 ;
        RECT 559.950 371.400 577.050 372.600 ;
        RECT 526.950 369.600 529.050 370.050 ;
        RECT 536.400 369.600 537.600 371.100 ;
        RECT 559.950 370.950 562.050 371.400 ;
        RECT 574.950 370.950 577.050 371.400 ;
        RECT 578.400 371.400 586.050 372.600 ;
        RECT 578.400 369.600 579.600 371.400 ;
        RECT 583.950 371.100 586.050 371.400 ;
        RECT 610.950 370.950 613.050 373.050 ;
        RECT 631.950 372.750 634.050 373.200 ;
        RECT 640.950 372.750 643.050 373.200 ;
        RECT 631.950 371.550 643.050 372.750 ;
        RECT 658.950 372.600 661.050 373.050 ;
        RECT 631.950 371.100 634.050 371.550 ;
        RECT 640.950 371.100 643.050 371.550 ;
        RECT 650.400 371.400 661.050 372.600 ;
        RECT 526.950 368.400 537.600 369.600 ;
        RECT 569.400 368.400 579.600 369.600 ;
        RECT 526.950 367.950 529.050 368.400 ;
        RECT 460.950 365.400 474.600 366.600 ;
        RECT 448.950 364.950 453.000 365.400 ;
        RECT 460.950 364.800 463.050 365.400 ;
        RECT 490.950 364.800 493.050 366.900 ;
        RECT 520.950 364.950 523.050 367.050 ;
        RECT 550.950 366.600 553.050 367.050 ;
        RECT 569.400 366.900 570.600 368.400 ;
        RECT 611.400 366.900 612.600 370.950 ;
        RECT 562.950 366.600 565.050 366.900 ;
        RECT 550.950 365.400 565.050 366.600 ;
        RECT 550.950 364.950 553.050 365.400 ;
        RECT 562.950 364.800 565.050 365.400 ;
        RECT 568.950 364.800 571.050 366.900 ;
        RECT 601.950 366.450 604.050 366.900 ;
        RECT 610.950 366.450 613.050 366.900 ;
        RECT 601.950 365.250 613.050 366.450 ;
        RECT 601.950 364.800 604.050 365.250 ;
        RECT 610.950 364.800 613.050 365.250 ;
        RECT 616.950 366.600 619.050 367.050 ;
        RECT 650.400 366.900 651.600 371.400 ;
        RECT 658.950 370.950 661.050 371.400 ;
        RECT 667.950 372.600 670.050 373.200 ;
        RECT 667.950 371.400 678.600 372.600 ;
        RECT 667.950 371.100 670.050 371.400 ;
        RECT 677.400 370.050 678.600 371.400 ;
        RECT 688.950 370.950 691.050 373.050 ;
        RECT 713.400 372.600 714.600 374.400 ;
        RECT 724.950 373.950 727.050 374.400 ;
        RECT 730.950 373.950 733.050 374.400 ;
        RECT 757.950 373.950 760.050 376.050 ;
        RECT 823.950 375.600 826.050 376.050 ;
        RECT 832.950 375.600 835.050 376.050 ;
        RECT 823.950 374.400 835.050 375.600 ;
        RECT 823.950 373.950 826.050 374.400 ;
        RECT 832.950 373.950 835.050 374.400 ;
        RECT 868.950 375.600 873.000 376.050 ;
        RECT 877.950 375.600 880.050 376.050 ;
        RECT 889.950 375.600 892.050 376.050 ;
        RECT 868.950 373.950 873.600 375.600 ;
        RECT 877.950 374.400 892.050 375.600 ;
        RECT 877.950 373.950 880.050 374.400 ;
        RECT 889.950 373.950 892.050 374.400 ;
        RECT 701.400 371.400 714.600 372.600 ;
        RECT 715.950 372.600 718.050 373.200 ;
        RECT 715.950 371.400 723.600 372.600 ;
        RECT 677.400 368.400 682.050 370.050 ;
        RECT 678.000 367.950 682.050 368.400 ;
        RECT 616.950 365.400 642.600 366.600 ;
        RECT 616.950 364.950 619.050 365.400 ;
        RECT 454.950 363.600 457.050 364.050 ;
        RECT 460.950 363.600 463.050 363.750 ;
        RECT 454.950 362.400 463.050 363.600 ;
        RECT 454.950 361.950 457.050 362.400 ;
        RECT 112.950 360.600 115.050 361.050 ;
        RECT 127.950 360.600 130.050 361.050 ;
        RECT 112.950 359.400 130.050 360.600 ;
        RECT 112.950 358.950 115.050 359.400 ;
        RECT 127.950 358.950 130.050 359.400 ;
        RECT 133.950 360.600 136.050 361.050 ;
        RECT 163.950 360.600 166.050 361.050 ;
        RECT 133.950 359.400 166.050 360.600 ;
        RECT 133.950 358.950 136.050 359.400 ;
        RECT 163.950 358.950 166.050 359.400 ;
        RECT 169.950 360.600 172.050 361.050 ;
        RECT 205.950 360.600 208.050 361.050 ;
        RECT 259.950 360.600 262.050 361.050 ;
        RECT 169.950 359.400 208.050 360.600 ;
        RECT 169.950 358.950 172.050 359.400 ;
        RECT 205.950 358.950 208.050 359.400 ;
        RECT 251.400 359.400 262.050 360.600 ;
        RECT 251.400 358.050 252.600 359.400 ;
        RECT 259.950 358.950 262.050 359.400 ;
        RECT 280.950 360.600 283.050 361.050 ;
        RECT 289.950 360.600 292.050 361.050 ;
        RECT 280.950 359.400 292.050 360.600 ;
        RECT 280.950 358.950 283.050 359.400 ;
        RECT 289.950 358.950 292.050 359.400 ;
        RECT 307.950 360.600 310.050 361.050 ;
        RECT 332.400 360.600 333.600 361.950 ;
        RECT 460.950 361.650 463.050 362.400 ;
        RECT 496.950 363.600 499.050 364.050 ;
        RECT 526.950 363.600 529.050 364.050 ;
        RECT 496.950 362.400 529.050 363.600 ;
        RECT 496.950 361.950 499.050 362.400 ;
        RECT 526.950 361.950 529.050 362.400 ;
        RECT 607.950 363.600 610.050 364.050 ;
        RECT 622.950 363.600 625.050 364.050 ;
        RECT 607.950 362.400 625.050 363.600 ;
        RECT 641.400 363.600 642.600 365.400 ;
        RECT 649.950 364.800 652.050 366.900 ;
        RECT 655.950 366.450 658.050 366.900 ;
        RECT 661.950 366.450 664.050 366.900 ;
        RECT 655.950 365.250 664.050 366.450 ;
        RECT 655.950 364.800 658.050 365.250 ;
        RECT 661.950 364.800 664.050 365.250 ;
        RECT 670.950 366.600 673.050 366.900 ;
        RECT 689.400 366.600 690.600 370.950 ;
        RECT 670.950 365.400 690.600 366.600 ;
        RECT 697.950 366.600 700.050 366.900 ;
        RECT 701.400 366.600 702.600 371.400 ;
        RECT 715.950 371.100 718.050 371.400 ;
        RECT 722.400 370.050 723.600 371.400 ;
        RECT 748.950 370.950 751.050 373.050 ;
        RECT 722.400 368.400 727.050 370.050 ;
        RECT 723.000 367.950 727.050 368.400 ;
        RECT 749.400 367.050 750.600 370.950 ;
        RECT 697.950 365.400 702.600 366.600 ;
        RECT 670.950 364.800 673.050 365.400 ;
        RECT 697.950 364.800 700.050 365.400 ;
        RECT 748.950 364.950 751.050 367.050 ;
        RECT 758.400 366.900 759.600 373.950 ;
        RECT 760.950 371.100 763.050 373.200 ;
        RECT 769.950 372.600 774.000 373.050 ;
        RECT 793.950 372.600 796.050 373.200 ;
        RECT 761.400 367.050 762.600 371.100 ;
        RECT 769.950 370.950 774.600 372.600 ;
        RECT 757.950 364.800 760.050 366.900 ;
        RECT 761.400 365.400 766.050 367.050 ;
        RECT 773.400 366.900 774.600 370.950 ;
        RECT 791.400 371.400 796.050 372.600 ;
        RECT 791.400 367.050 792.600 371.400 ;
        RECT 793.950 371.100 796.050 371.400 ;
        RECT 799.950 371.100 802.050 373.200 ;
        RECT 762.000 364.950 766.050 365.400 ;
        RECT 772.950 364.800 775.050 366.900 ;
        RECT 790.950 364.950 793.050 367.050 ;
        RECT 800.400 364.050 801.600 371.100 ;
        RECT 805.950 369.600 808.050 373.050 ;
        RECT 811.950 372.600 814.050 373.050 ;
        RECT 811.950 371.400 819.600 372.600 ;
        RECT 811.950 370.950 814.050 371.400 ;
        RECT 803.400 369.000 808.050 369.600 ;
        RECT 803.400 368.400 807.600 369.000 ;
        RECT 803.400 366.900 804.600 368.400 ;
        RECT 818.400 366.900 819.600 371.400 ;
        RECT 826.950 369.600 829.050 373.050 ;
        RECT 856.950 370.950 859.050 373.050 ;
        RECT 821.400 369.000 829.050 369.600 ;
        RECT 820.950 368.400 828.600 369.000 ;
        RECT 802.950 364.800 805.050 366.900 ;
        RECT 817.800 364.800 819.900 366.900 ;
        RECT 820.950 364.950 823.050 368.400 ;
        RECT 829.950 366.600 832.050 367.050 ;
        RECT 841.950 366.600 844.050 366.900 ;
        RECT 829.950 365.400 844.050 366.600 ;
        RECT 829.950 364.950 832.050 365.400 ;
        RECT 841.950 364.800 844.050 365.400 ;
        RECT 850.950 366.600 853.050 367.050 ;
        RECT 857.400 366.600 858.600 370.950 ;
        RECT 872.400 369.600 873.600 373.950 ;
        RECT 898.950 370.950 901.050 373.050 ;
        RECT 910.950 370.950 913.050 373.050 ;
        RECT 872.400 369.000 882.600 369.600 ;
        RECT 872.400 368.400 883.050 369.000 ;
        RECT 850.950 365.400 858.600 366.600 ;
        RECT 868.950 366.450 871.050 366.900 ;
        RECT 874.950 366.450 877.050 366.900 ;
        RECT 850.950 364.950 853.050 365.400 ;
        RECT 868.950 365.250 877.050 366.450 ;
        RECT 868.950 364.800 871.050 365.250 ;
        RECT 874.950 364.800 877.050 365.250 ;
        RECT 880.950 364.950 883.050 368.400 ;
        RECT 899.400 367.050 900.600 370.950 ;
        RECT 911.400 367.050 912.600 370.950 ;
        RECT 898.950 364.950 901.050 367.050 ;
        RECT 910.950 364.950 913.050 367.050 ;
        RECT 652.950 363.600 655.050 364.050 ;
        RECT 641.400 362.400 655.050 363.600 ;
        RECT 607.950 361.950 610.050 362.400 ;
        RECT 622.950 361.950 625.050 362.400 ;
        RECT 652.950 361.950 655.050 362.400 ;
        RECT 706.950 363.600 709.050 364.050 ;
        RECT 712.950 363.600 715.050 364.050 ;
        RECT 706.950 362.400 715.050 363.600 ;
        RECT 706.950 361.950 709.050 362.400 ;
        RECT 712.950 361.950 715.050 362.400 ;
        RECT 787.950 363.600 790.050 364.050 ;
        RECT 796.800 363.600 798.900 364.050 ;
        RECT 787.950 362.400 798.900 363.600 ;
        RECT 787.950 361.950 790.050 362.400 ;
        RECT 796.800 361.950 798.900 362.400 ;
        RECT 799.950 361.950 802.050 364.050 ;
        RECT 832.950 363.600 835.050 364.050 ;
        RECT 838.950 363.600 841.050 364.050 ;
        RECT 832.950 362.400 841.050 363.600 ;
        RECT 832.950 361.950 835.050 362.400 ;
        RECT 838.950 361.950 841.050 362.400 ;
        RECT 307.950 359.400 333.600 360.600 ;
        RECT 349.950 360.600 352.050 361.050 ;
        RECT 406.950 360.600 409.050 361.050 ;
        RECT 349.950 359.400 409.050 360.600 ;
        RECT 307.950 358.950 310.050 359.400 ;
        RECT 349.950 358.950 352.050 359.400 ;
        RECT 406.950 358.950 409.050 359.400 ;
        RECT 445.950 360.600 448.050 361.050 ;
        RECT 532.950 360.600 535.050 361.050 ;
        RECT 445.950 359.400 535.050 360.600 ;
        RECT 445.950 358.950 448.050 359.400 ;
        RECT 532.950 358.950 535.050 359.400 ;
        RECT 586.950 360.600 589.050 361.050 ;
        RECT 742.950 360.600 745.050 361.050 ;
        RECT 760.950 360.600 763.050 361.050 ;
        RECT 586.950 359.400 763.050 360.600 ;
        RECT 586.950 358.950 589.050 359.400 ;
        RECT 742.950 358.950 745.050 359.400 ;
        RECT 760.950 358.950 763.050 359.400 ;
        RECT 883.950 360.600 886.050 361.050 ;
        RECT 901.950 360.600 904.050 361.050 ;
        RECT 883.950 359.400 904.050 360.600 ;
        RECT 883.950 358.950 886.050 359.400 ;
        RECT 901.950 358.950 904.050 359.400 ;
        RECT 907.950 360.600 910.050 361.050 ;
        RECT 913.950 360.600 916.050 361.050 ;
        RECT 907.950 359.400 916.050 360.600 ;
        RECT 907.950 358.950 910.050 359.400 ;
        RECT 913.950 358.950 916.050 359.400 ;
        RECT 4.950 357.600 7.050 358.050 ;
        RECT 13.950 357.600 16.050 358.050 ;
        RECT 4.950 356.400 16.050 357.600 ;
        RECT 4.950 355.950 7.050 356.400 ;
        RECT 13.950 355.950 16.050 356.400 ;
        RECT 37.950 357.600 40.050 358.050 ;
        RECT 43.950 357.600 46.050 358.050 ;
        RECT 37.950 356.400 46.050 357.600 ;
        RECT 37.950 355.950 40.050 356.400 ;
        RECT 43.950 355.950 46.050 356.400 ;
        RECT 70.950 357.600 73.050 358.050 ;
        RECT 79.950 357.600 82.050 358.050 ;
        RECT 91.950 357.600 94.050 358.050 ;
        RECT 106.950 357.600 109.050 358.050 ;
        RECT 166.950 357.600 169.050 358.050 ;
        RECT 70.950 356.400 169.050 357.600 ;
        RECT 70.950 355.950 73.050 356.400 ;
        RECT 79.950 355.950 82.050 356.400 ;
        RECT 91.950 355.950 94.050 356.400 ;
        RECT 106.950 355.950 109.050 356.400 ;
        RECT 166.950 355.950 169.050 356.400 ;
        RECT 172.950 357.600 175.050 358.050 ;
        RECT 184.950 357.600 187.050 358.050 ;
        RECT 172.950 356.400 187.050 357.600 ;
        RECT 172.950 355.950 175.050 356.400 ;
        RECT 184.950 355.950 187.050 356.400 ;
        RECT 238.950 357.600 241.050 358.050 ;
        RECT 250.950 357.600 253.050 358.050 ;
        RECT 238.950 356.400 253.050 357.600 ;
        RECT 238.950 355.950 241.050 356.400 ;
        RECT 250.950 355.950 253.050 356.400 ;
        RECT 259.950 357.600 262.050 357.900 ;
        RECT 277.950 357.600 280.050 358.050 ;
        RECT 259.950 356.400 280.050 357.600 ;
        RECT 259.950 355.800 262.050 356.400 ;
        RECT 277.950 355.950 280.050 356.400 ;
        RECT 292.950 357.600 295.050 358.050 ;
        RECT 346.950 357.600 349.050 358.050 ;
        RECT 292.950 356.400 349.050 357.600 ;
        RECT 292.950 355.950 295.050 356.400 ;
        RECT 346.950 355.950 349.050 356.400 ;
        RECT 373.950 357.600 376.050 358.050 ;
        RECT 427.950 357.600 430.050 358.050 ;
        RECT 469.950 357.600 472.050 358.050 ;
        RECT 373.950 356.400 472.050 357.600 ;
        RECT 373.950 355.950 376.050 356.400 ;
        RECT 427.950 355.950 430.050 356.400 ;
        RECT 469.950 355.950 472.050 356.400 ;
        RECT 592.950 357.600 595.050 358.050 ;
        RECT 601.950 357.600 604.050 358.050 ;
        RECT 592.950 356.400 604.050 357.600 ;
        RECT 592.950 355.950 595.050 356.400 ;
        RECT 601.950 355.950 604.050 356.400 ;
        RECT 652.950 357.600 655.050 358.050 ;
        RECT 697.950 357.600 700.050 358.050 ;
        RECT 652.950 356.400 700.050 357.600 ;
        RECT 652.950 355.950 655.050 356.400 ;
        RECT 697.950 355.950 700.050 356.400 ;
        RECT 736.950 357.600 739.050 358.050 ;
        RECT 766.950 357.600 769.050 358.050 ;
        RECT 736.950 356.400 769.050 357.600 ;
        RECT 736.950 355.950 739.050 356.400 ;
        RECT 766.950 355.950 769.050 356.400 ;
        RECT 787.950 357.600 790.050 358.050 ;
        RECT 904.950 357.600 907.050 358.050 ;
        RECT 787.950 356.400 907.050 357.600 ;
        RECT 787.950 355.950 790.050 356.400 ;
        RECT 904.950 355.950 907.050 356.400 ;
        RECT 109.950 354.600 112.050 355.050 ;
        RECT 118.950 354.600 121.050 355.050 ;
        RECT 160.800 354.600 162.900 355.050 ;
        RECT 109.950 353.400 162.900 354.600 ;
        RECT 109.950 352.950 112.050 353.400 ;
        RECT 118.950 352.950 121.050 353.400 ;
        RECT 160.800 352.950 162.900 353.400 ;
        RECT 163.950 354.600 166.050 355.050 ;
        RECT 220.950 354.600 223.050 355.050 ;
        RECT 163.950 353.400 223.050 354.600 ;
        RECT 163.950 352.950 166.050 353.400 ;
        RECT 220.950 352.950 223.050 353.400 ;
        RECT 232.950 354.600 235.050 355.050 ;
        RECT 295.950 354.600 298.050 355.050 ;
        RECT 232.950 353.400 298.050 354.600 ;
        RECT 232.950 352.950 235.050 353.400 ;
        RECT 295.950 352.950 298.050 353.400 ;
        RECT 301.950 354.600 304.050 355.050 ;
        RECT 313.800 354.600 315.900 355.050 ;
        RECT 301.950 353.400 315.900 354.600 ;
        RECT 301.950 352.950 304.050 353.400 ;
        RECT 313.800 352.950 315.900 353.400 ;
        RECT 316.950 354.600 319.050 355.050 ;
        RECT 373.950 354.600 376.050 354.900 ;
        RECT 388.950 354.600 391.050 355.050 ;
        RECT 316.950 353.400 391.050 354.600 ;
        RECT 316.950 352.950 319.050 353.400 ;
        RECT 373.950 352.800 376.050 353.400 ;
        RECT 388.950 352.950 391.050 353.400 ;
        RECT 397.950 354.600 400.050 355.050 ;
        RECT 424.950 354.600 427.050 355.050 ;
        RECT 397.950 353.400 427.050 354.600 ;
        RECT 397.950 352.950 400.050 353.400 ;
        RECT 424.950 352.950 427.050 353.400 ;
        RECT 445.950 354.600 448.050 355.050 ;
        RECT 466.950 354.600 469.050 355.050 ;
        RECT 445.950 353.400 469.050 354.600 ;
        RECT 445.950 352.950 448.050 353.400 ;
        RECT 466.950 352.950 469.050 353.400 ;
        RECT 628.950 354.600 631.050 355.050 ;
        RECT 649.950 354.600 652.050 355.050 ;
        RECT 628.950 353.400 652.050 354.600 ;
        RECT 628.950 352.950 631.050 353.400 ;
        RECT 649.950 352.950 652.050 353.400 ;
        RECT 745.950 354.600 748.050 355.050 ;
        RECT 793.950 354.600 796.050 355.050 ;
        RECT 745.950 353.400 796.050 354.600 ;
        RECT 745.950 352.950 748.050 353.400 ;
        RECT 793.950 352.950 796.050 353.400 ;
        RECT 823.950 354.600 826.050 355.050 ;
        RECT 895.950 354.600 898.050 355.050 ;
        RECT 823.950 353.400 898.050 354.600 ;
        RECT 823.950 352.950 826.050 353.400 ;
        RECT 895.950 352.950 898.050 353.400 ;
        RECT 913.950 354.600 916.050 355.050 ;
        RECT 919.950 354.600 922.050 355.050 ;
        RECT 913.950 353.400 922.050 354.600 ;
        RECT 913.950 352.950 916.050 353.400 ;
        RECT 919.950 352.950 922.050 353.400 ;
        RECT 10.950 351.600 13.050 352.050 ;
        RECT 16.950 351.600 19.050 352.050 ;
        RECT 10.950 350.400 19.050 351.600 ;
        RECT 10.950 349.950 13.050 350.400 ;
        RECT 16.950 349.950 19.050 350.400 ;
        RECT 28.950 351.600 31.050 352.050 ;
        RECT 43.950 351.600 46.050 352.050 ;
        RECT 52.950 351.600 55.050 352.050 ;
        RECT 28.950 350.400 55.050 351.600 ;
        RECT 28.950 349.950 31.050 350.400 ;
        RECT 43.950 349.950 46.050 350.400 ;
        RECT 52.950 349.950 55.050 350.400 ;
        RECT 58.950 351.600 61.050 352.050 ;
        RECT 85.950 351.600 88.050 352.050 ;
        RECT 136.950 351.600 139.050 352.050 ;
        RECT 142.950 351.600 145.050 352.050 ;
        RECT 58.950 350.400 145.050 351.600 ;
        RECT 58.950 349.950 61.050 350.400 ;
        RECT 85.950 349.950 88.050 350.400 ;
        RECT 136.950 349.950 139.050 350.400 ;
        RECT 142.950 349.950 145.050 350.400 ;
        RECT 199.950 351.600 202.050 352.050 ;
        RECT 208.950 351.600 211.050 352.050 ;
        RECT 199.950 350.400 211.050 351.600 ;
        RECT 199.950 349.950 202.050 350.400 ;
        RECT 208.950 349.950 211.050 350.400 ;
        RECT 217.950 351.600 220.050 352.050 ;
        RECT 247.950 351.600 250.050 352.050 ;
        RECT 217.950 350.400 250.050 351.600 ;
        RECT 217.950 349.950 220.050 350.400 ;
        RECT 247.950 349.950 250.050 350.400 ;
        RECT 253.950 351.600 256.050 352.050 ;
        RECT 280.950 351.600 283.050 352.050 ;
        RECT 286.950 351.600 289.050 352.050 ;
        RECT 352.950 351.600 355.050 352.050 ;
        RECT 253.950 350.400 273.600 351.600 ;
        RECT 253.950 349.950 256.050 350.400 ;
        RECT 272.400 349.050 273.600 350.400 ;
        RECT 280.950 350.400 355.050 351.600 ;
        RECT 280.950 349.950 283.050 350.400 ;
        RECT 286.950 349.950 289.050 350.400 ;
        RECT 352.950 349.950 355.050 350.400 ;
        RECT 400.950 351.600 403.050 352.050 ;
        RECT 541.950 351.600 544.050 352.050 ;
        RECT 400.950 350.400 544.050 351.600 ;
        RECT 400.950 349.950 403.050 350.400 ;
        RECT 541.950 349.950 544.050 350.400 ;
        RECT 547.950 351.600 550.050 352.050 ;
        RECT 559.950 351.600 562.050 352.050 ;
        RECT 547.950 350.400 562.050 351.600 ;
        RECT 547.950 349.950 550.050 350.400 ;
        RECT 559.950 349.950 562.050 350.400 ;
        RECT 142.950 348.600 145.050 348.900 ;
        RECT 154.950 348.600 157.050 349.050 ;
        RECT 142.950 347.400 157.050 348.600 ;
        RECT 142.950 346.800 145.050 347.400 ;
        RECT 154.950 346.950 157.050 347.400 ;
        RECT 175.950 348.600 178.050 349.050 ;
        RECT 190.950 348.600 193.050 349.050 ;
        RECT 211.950 348.600 214.050 349.050 ;
        RECT 253.950 348.600 256.050 348.900 ;
        RECT 175.950 347.400 256.050 348.600 ;
        RECT 175.950 346.950 178.050 347.400 ;
        RECT 190.950 346.950 193.050 347.400 ;
        RECT 211.950 346.950 214.050 347.400 ;
        RECT 253.950 346.800 256.050 347.400 ;
        RECT 271.950 348.600 274.050 349.050 ;
        RECT 316.950 348.600 319.050 349.050 ;
        RECT 271.950 347.400 319.050 348.600 ;
        RECT 271.950 346.950 274.050 347.400 ;
        RECT 316.950 346.950 319.050 347.400 ;
        RECT 370.950 348.600 373.050 349.050 ;
        RECT 388.950 348.600 391.050 349.050 ;
        RECT 370.950 347.400 391.050 348.600 ;
        RECT 370.950 346.950 373.050 347.400 ;
        RECT 388.950 346.950 391.050 347.400 ;
        RECT 424.950 348.600 427.050 349.050 ;
        RECT 448.950 348.600 451.050 349.050 ;
        RECT 454.950 348.600 457.050 349.050 ;
        RECT 505.950 348.600 508.050 349.050 ;
        RECT 526.950 348.600 529.050 349.050 ;
        RECT 424.950 347.400 457.050 348.600 ;
        RECT 424.950 346.950 427.050 347.400 ;
        RECT 448.950 346.950 451.050 347.400 ;
        RECT 454.950 346.950 457.050 347.400 ;
        RECT 458.400 347.400 529.050 348.600 ;
        RECT 574.950 348.600 577.050 352.050 ;
        RECT 607.950 351.600 610.050 352.050 ;
        RECT 640.950 351.600 643.050 352.050 ;
        RECT 607.950 350.400 643.050 351.600 ;
        RECT 607.950 349.950 610.050 350.400 ;
        RECT 640.950 349.950 643.050 350.400 ;
        RECT 670.950 351.600 673.050 352.050 ;
        RECT 679.950 351.600 682.050 352.050 ;
        RECT 670.950 350.400 682.050 351.600 ;
        RECT 670.950 349.950 673.050 350.400 ;
        RECT 679.950 349.950 682.050 350.400 ;
        RECT 706.950 351.600 709.050 352.050 ;
        RECT 721.950 351.600 724.050 352.050 ;
        RECT 706.950 350.400 724.050 351.600 ;
        RECT 706.950 349.950 709.050 350.400 ;
        RECT 721.950 349.950 724.050 350.400 ;
        RECT 748.950 351.600 751.050 352.050 ;
        RECT 757.950 351.600 760.050 352.050 ;
        RECT 748.950 350.400 760.050 351.600 ;
        RECT 748.950 349.950 751.050 350.400 ;
        RECT 757.950 349.950 760.050 350.400 ;
        RECT 766.950 351.600 769.050 352.050 ;
        RECT 787.950 351.600 790.050 352.050 ;
        RECT 766.950 350.400 790.050 351.600 ;
        RECT 766.950 349.950 769.050 350.400 ;
        RECT 787.950 349.950 790.050 350.400 ;
        RECT 802.950 351.600 805.050 352.050 ;
        RECT 820.950 351.600 823.050 352.050 ;
        RECT 802.950 350.400 823.050 351.600 ;
        RECT 802.950 349.950 805.050 350.400 ;
        RECT 820.950 349.950 823.050 350.400 ;
        RECT 838.950 351.600 841.050 352.050 ;
        RECT 847.950 351.600 850.050 352.050 ;
        RECT 838.950 350.400 850.050 351.600 ;
        RECT 838.950 349.950 841.050 350.400 ;
        RECT 847.950 349.950 850.050 350.400 ;
        RECT 616.950 348.600 619.050 349.050 ;
        RECT 574.950 348.000 619.050 348.600 ;
        RECT 575.400 347.400 619.050 348.000 ;
        RECT 16.950 345.600 19.050 346.050 ;
        RECT 37.950 345.600 40.050 346.050 ;
        RECT 16.950 344.400 40.050 345.600 ;
        RECT 16.950 343.950 19.050 344.400 ;
        RECT 37.950 343.950 40.050 344.400 ;
        RECT 55.950 345.600 58.050 346.050 ;
        RECT 124.950 345.600 127.050 346.050 ;
        RECT 172.950 345.600 175.050 346.050 ;
        RECT 55.950 344.400 69.600 345.600 ;
        RECT 55.950 343.950 58.050 344.400 ;
        RECT 68.400 343.050 69.600 344.400 ;
        RECT 124.950 344.400 175.050 345.600 ;
        RECT 124.950 343.950 127.050 344.400 ;
        RECT 172.950 343.950 175.050 344.400 ;
        RECT 178.950 345.600 181.050 346.050 ;
        RECT 247.950 345.600 250.050 346.050 ;
        RECT 262.950 345.600 265.050 346.050 ;
        RECT 178.950 344.400 216.600 345.600 ;
        RECT 178.950 343.950 181.050 344.400 ;
        RECT 215.400 343.050 216.600 344.400 ;
        RECT 247.950 344.400 265.050 345.600 ;
        RECT 247.950 343.950 250.050 344.400 ;
        RECT 262.950 343.950 265.050 344.400 ;
        RECT 268.950 345.600 271.050 346.050 ;
        RECT 301.950 345.600 304.050 346.050 ;
        RECT 268.950 344.400 304.050 345.600 ;
        RECT 268.950 343.950 271.050 344.400 ;
        RECT 301.950 343.950 304.050 344.400 ;
        RECT 328.950 345.600 331.050 346.050 ;
        RECT 361.800 345.600 363.900 346.050 ;
        RECT 328.950 344.400 363.900 345.600 ;
        RECT 328.950 343.950 331.050 344.400 ;
        RECT 361.800 343.950 363.900 344.400 ;
        RECT 364.950 345.600 367.050 346.050 ;
        RECT 406.950 345.600 409.050 346.050 ;
        RECT 364.950 344.400 409.050 345.600 ;
        RECT 364.950 343.950 367.050 344.400 ;
        RECT 406.950 343.950 409.050 344.400 ;
        RECT 421.950 345.600 424.050 346.050 ;
        RECT 458.400 345.600 459.600 347.400 ;
        RECT 505.950 346.950 508.050 347.400 ;
        RECT 526.950 346.950 529.050 347.400 ;
        RECT 616.950 346.950 619.050 347.400 ;
        RECT 622.950 348.600 625.050 349.050 ;
        RECT 628.950 348.600 631.050 349.050 ;
        RECT 643.950 348.600 646.050 349.050 ;
        RECT 622.950 347.400 646.050 348.600 ;
        RECT 622.950 346.950 625.050 347.400 ;
        RECT 628.950 346.950 631.050 347.400 ;
        RECT 643.950 346.950 646.050 347.400 ;
        RECT 721.950 348.600 724.050 348.900 ;
        RECT 763.950 348.600 766.050 349.050 ;
        RECT 772.950 348.600 775.050 349.050 ;
        RECT 790.950 348.600 793.050 349.050 ;
        RECT 835.950 348.600 838.050 349.050 ;
        RECT 721.950 347.400 838.050 348.600 ;
        RECT 721.950 346.800 724.050 347.400 ;
        RECT 763.950 346.950 766.050 347.400 ;
        RECT 772.950 346.950 775.050 347.400 ;
        RECT 790.950 346.950 793.050 347.400 ;
        RECT 835.950 346.950 838.050 347.400 ;
        RECT 877.950 348.600 880.050 349.050 ;
        RECT 886.950 348.600 889.050 349.050 ;
        RECT 877.950 347.400 889.050 348.600 ;
        RECT 877.950 346.950 880.050 347.400 ;
        RECT 886.950 346.950 889.050 347.400 ;
        RECT 892.950 348.600 895.050 349.050 ;
        RECT 901.950 348.600 904.050 349.050 ;
        RECT 892.950 347.400 904.050 348.600 ;
        RECT 892.950 346.950 895.050 347.400 ;
        RECT 901.950 346.950 904.050 347.400 ;
        RECT 907.950 348.600 910.050 349.050 ;
        RECT 916.950 348.600 919.050 349.050 ;
        RECT 907.950 347.400 919.050 348.600 ;
        RECT 907.950 346.950 910.050 347.400 ;
        RECT 916.950 346.950 919.050 347.400 ;
        RECT 421.950 344.400 459.600 345.600 ;
        RECT 529.950 345.600 532.050 346.050 ;
        RECT 580.950 345.600 583.050 346.050 ;
        RECT 529.950 344.400 583.050 345.600 ;
        RECT 421.950 343.950 424.050 344.400 ;
        RECT 529.950 343.950 532.050 344.400 ;
        RECT 580.950 343.950 583.050 344.400 ;
        RECT 40.950 340.950 43.050 343.050 ;
        RECT 46.950 342.600 49.050 343.050 ;
        RECT 52.950 342.600 55.050 343.050 ;
        RECT 46.950 341.400 55.050 342.600 ;
        RECT 46.950 340.950 49.050 341.400 ;
        RECT 52.950 340.950 55.050 341.400 ;
        RECT 67.950 342.600 70.050 343.050 ;
        RECT 76.950 342.600 79.050 343.050 ;
        RECT 67.950 341.400 79.050 342.600 ;
        RECT 67.950 340.950 70.050 341.400 ;
        RECT 76.950 340.950 79.050 341.400 ;
        RECT 100.950 342.600 103.050 343.050 ;
        RECT 112.950 342.600 115.050 343.050 ;
        RECT 100.950 341.400 115.050 342.600 ;
        RECT 100.950 340.950 103.050 341.400 ;
        RECT 112.950 340.950 115.050 341.400 ;
        RECT 124.950 342.600 127.050 342.900 ;
        RECT 130.950 342.600 133.050 343.050 ;
        RECT 124.950 341.400 133.050 342.600 ;
        RECT 22.950 339.750 25.050 340.200 ;
        RECT 34.950 339.750 37.050 340.200 ;
        RECT 22.950 338.550 37.050 339.750 ;
        RECT 22.950 338.100 25.050 338.550 ;
        RECT 34.950 338.100 37.050 338.550 ;
        RECT 13.950 333.450 16.050 333.900 ;
        RECT 34.950 333.450 37.050 333.900 ;
        RECT 13.950 332.250 37.050 333.450 ;
        RECT 13.950 331.800 16.050 332.250 ;
        RECT 34.950 331.800 37.050 332.250 ;
        RECT 41.400 331.050 42.600 340.950 ;
        RECT 124.950 340.800 127.050 341.400 ;
        RECT 130.950 340.950 133.050 341.400 ;
        RECT 214.950 342.600 217.050 343.050 ;
        RECT 223.950 342.600 226.050 343.050 ;
        RECT 244.950 342.600 247.050 343.050 ;
        RECT 214.950 341.400 247.050 342.600 ;
        RECT 214.950 340.950 217.050 341.400 ;
        RECT 223.950 340.950 226.050 341.400 ;
        RECT 244.950 340.950 247.050 341.400 ;
        RECT 277.800 340.950 279.900 343.050 ;
        RECT 289.950 342.600 292.050 343.050 ;
        RECT 301.950 342.600 304.050 342.900 ;
        RECT 289.950 341.400 304.050 342.600 ;
        RECT 289.950 340.950 292.050 341.400 ;
        RECT 58.950 339.600 63.000 340.050 ;
        RECT 64.950 339.600 67.050 340.200 ;
        RECT 91.950 339.600 94.050 340.200 ;
        RECT 97.950 339.600 100.050 340.050 ;
        RECT 58.950 337.950 63.600 339.600 ;
        RECT 64.950 338.400 69.600 339.600 ;
        RECT 64.950 338.100 67.050 338.400 ;
        RECT 62.400 333.900 63.600 337.950 ;
        RECT 46.950 333.450 49.050 333.900 ;
        RECT 55.950 333.450 58.050 333.900 ;
        RECT 46.950 332.250 58.050 333.450 ;
        RECT 46.950 331.800 49.050 332.250 ;
        RECT 55.950 331.800 58.050 332.250 ;
        RECT 61.950 331.800 64.050 333.900 ;
        RECT 68.400 331.050 69.600 338.400 ;
        RECT 91.950 338.400 100.050 339.600 ;
        RECT 91.950 338.100 94.050 338.400 ;
        RECT 97.950 337.950 100.050 338.400 ;
        RECT 103.950 339.600 106.050 340.050 ;
        RECT 151.950 339.600 154.050 340.200 ;
        RECT 103.950 338.400 154.050 339.600 ;
        RECT 103.950 337.950 106.050 338.400 ;
        RECT 151.950 338.100 154.050 338.400 ;
        RECT 157.950 339.600 160.050 340.200 ;
        RECT 175.950 339.600 178.050 340.200 ;
        RECT 157.950 338.400 178.050 339.600 ;
        RECT 157.950 338.100 160.050 338.400 ;
        RECT 175.950 338.100 178.050 338.400 ;
        RECT 181.950 339.600 184.050 340.200 ;
        RECT 199.950 339.600 202.050 340.200 ;
        RECT 256.950 339.750 259.050 340.200 ;
        RECT 265.950 339.750 268.050 340.200 ;
        RECT 181.950 338.400 225.600 339.600 ;
        RECT 181.950 338.100 184.050 338.400 ;
        RECT 199.950 338.100 202.050 338.400 ;
        RECT 104.400 334.050 105.600 337.950 ;
        RECT 76.950 333.450 79.050 333.900 ;
        RECT 82.950 333.450 85.050 333.900 ;
        RECT 76.950 332.250 85.050 333.450 ;
        RECT 76.950 331.800 79.050 332.250 ;
        RECT 82.950 331.800 85.050 332.250 ;
        RECT 103.950 331.950 106.050 334.050 ;
        RECT 115.950 333.600 118.050 333.900 ;
        RECT 133.950 333.600 136.050 333.900 ;
        RECT 115.950 332.400 136.050 333.600 ;
        RECT 115.950 331.800 118.050 332.400 ;
        RECT 133.950 331.800 136.050 332.400 ;
        RECT 139.950 333.600 142.050 334.050 ;
        RECT 145.950 333.600 148.050 334.050 ;
        RECT 139.950 332.400 148.050 333.600 ;
        RECT 139.950 331.950 142.050 332.400 ;
        RECT 145.950 331.950 148.050 332.400 ;
        RECT 184.950 333.450 187.050 333.900 ;
        RECT 190.950 333.450 193.050 333.900 ;
        RECT 184.950 332.250 193.050 333.450 ;
        RECT 184.950 331.800 187.050 332.250 ;
        RECT 190.950 331.800 193.050 332.250 ;
        RECT 196.950 333.600 199.050 333.900 ;
        RECT 220.950 333.600 223.050 333.900 ;
        RECT 196.950 332.400 223.050 333.600 ;
        RECT 224.400 333.600 225.600 338.400 ;
        RECT 256.950 338.550 268.050 339.750 ;
        RECT 256.950 338.100 259.050 338.550 ;
        RECT 265.950 338.100 268.050 338.550 ;
        RECT 278.250 334.050 279.450 340.950 ;
        RECT 301.950 340.800 304.050 341.400 ;
        RECT 283.950 336.600 286.050 340.050 ;
        RECT 292.950 337.950 295.050 340.050 ;
        RECT 313.950 339.600 316.050 340.200 ;
        RECT 322.800 339.600 324.900 340.050 ;
        RECT 313.950 338.400 324.900 339.600 ;
        RECT 313.950 338.100 316.050 338.400 ;
        RECT 322.800 337.950 324.900 338.400 ;
        RECT 325.950 339.600 328.050 339.900 ;
        RECT 337.950 339.600 340.050 343.050 ;
        RECT 343.950 342.600 346.050 343.050 ;
        RECT 355.950 342.600 358.050 343.050 ;
        RECT 343.950 341.400 358.050 342.600 ;
        RECT 343.950 340.950 346.050 341.400 ;
        RECT 355.950 340.950 358.050 341.400 ;
        RECT 511.950 342.600 514.050 343.050 ;
        RECT 523.950 342.600 526.050 343.050 ;
        RECT 511.950 341.400 526.050 342.600 ;
        RECT 511.950 340.950 514.050 341.400 ;
        RECT 523.950 340.950 526.050 341.400 ;
        RECT 532.950 342.600 535.050 343.050 ;
        RECT 538.950 342.600 541.050 343.050 ;
        RECT 532.950 341.400 541.050 342.600 ;
        RECT 532.950 340.950 535.050 341.400 ;
        RECT 538.950 340.950 541.050 341.400 ;
        RECT 589.950 342.600 592.050 343.050 ;
        RECT 613.950 342.600 616.050 343.050 ;
        RECT 631.950 342.600 634.050 343.050 ;
        RECT 589.950 341.400 609.600 342.600 ;
        RECT 589.950 340.950 592.050 341.400 ;
        RECT 325.950 339.000 340.050 339.600 ;
        RECT 433.950 339.750 436.050 340.200 ;
        RECT 439.950 339.750 442.050 340.200 ;
        RECT 325.950 338.400 339.600 339.000 ;
        RECT 433.950 338.550 442.050 339.750 ;
        RECT 281.400 336.000 286.050 336.600 ;
        RECT 281.400 335.400 285.600 336.000 ;
        RECT 281.400 334.050 282.600 335.400 ;
        RECT 293.400 334.050 294.600 337.950 ;
        RECT 325.950 337.800 328.050 338.400 ;
        RECT 433.950 338.100 436.050 338.550 ;
        RECT 439.950 338.100 442.050 338.550 ;
        RECT 448.950 339.750 451.050 340.200 ;
        RECT 460.950 339.750 463.050 340.200 ;
        RECT 448.950 338.550 463.050 339.750 ;
        RECT 448.950 338.100 451.050 338.550 ;
        RECT 460.950 338.100 463.050 338.550 ;
        RECT 475.950 339.600 478.050 340.200 ;
        RECT 490.950 339.600 493.050 340.050 ;
        RECT 475.950 338.400 493.050 339.600 ;
        RECT 475.950 338.100 478.050 338.400 ;
        RECT 490.950 337.950 493.050 338.400 ;
        RECT 502.950 339.750 505.050 340.200 ;
        RECT 508.950 339.750 511.050 340.200 ;
        RECT 502.950 338.550 511.050 339.750 ;
        RECT 502.950 338.100 505.050 338.550 ;
        RECT 508.950 338.100 511.050 338.550 ;
        RECT 364.950 336.600 367.050 337.050 ;
        RECT 299.400 336.000 367.050 336.600 ;
        RECT 298.950 335.400 367.050 336.000 ;
        RECT 226.800 333.600 228.900 333.900 ;
        RECT 224.400 332.400 228.900 333.600 ;
        RECT 196.950 331.800 199.050 332.400 ;
        RECT 220.950 331.800 223.050 332.400 ;
        RECT 226.800 331.800 228.900 332.400 ;
        RECT 229.950 333.600 232.050 334.050 ;
        RECT 247.950 333.600 250.050 333.900 ;
        RECT 229.950 332.400 250.050 333.600 ;
        RECT 229.950 331.950 232.050 332.400 ;
        RECT 247.950 331.800 250.050 332.400 ;
        RECT 277.800 331.950 279.900 334.050 ;
        RECT 280.950 333.600 283.050 334.050 ;
        RECT 286.950 333.600 289.050 333.900 ;
        RECT 280.950 332.400 289.050 333.600 ;
        RECT 280.950 331.950 283.050 332.400 ;
        RECT 286.950 331.800 289.050 332.400 ;
        RECT 292.950 331.950 295.050 334.050 ;
        RECT 298.950 331.950 301.050 335.400 ;
        RECT 364.950 334.950 367.050 335.400 ;
        RECT 310.950 333.600 313.050 333.900 ;
        RECT 406.950 333.600 409.050 337.050 ;
        RECT 520.950 336.600 523.050 340.050 ;
        RECT 541.950 339.600 544.050 340.200 ;
        RECT 547.950 339.600 550.050 340.500 ;
        RECT 576.000 339.600 580.050 340.050 ;
        RECT 541.950 338.400 550.050 339.600 ;
        RECT 541.950 338.100 544.050 338.400 ;
        RECT 575.400 337.950 580.050 339.600 ;
        RECT 595.950 339.750 598.050 340.200 ;
        RECT 604.950 339.750 607.050 340.200 ;
        RECT 595.950 338.550 607.050 339.750 ;
        RECT 595.950 338.100 598.050 338.550 ;
        RECT 604.950 338.100 607.050 338.550 ;
        RECT 520.950 336.000 528.600 336.600 ;
        RECT 521.400 335.400 529.050 336.000 ;
        RECT 412.950 333.600 415.050 334.050 ;
        RECT 310.950 333.000 330.450 333.600 ;
        RECT 406.950 333.000 415.050 333.600 ;
        RECT 310.950 332.400 331.050 333.000 ;
        RECT 407.400 332.400 415.050 333.000 ;
        RECT 310.950 331.800 313.050 332.400 ;
        RECT 328.950 331.050 331.050 332.400 ;
        RECT 412.950 331.950 415.050 332.400 ;
        RECT 436.950 333.600 439.050 333.900 ;
        RECT 448.950 333.600 451.050 334.050 ;
        RECT 436.950 332.400 451.050 333.600 ;
        RECT 436.950 331.800 439.050 332.400 ;
        RECT 448.950 331.950 451.050 332.400 ;
        RECT 526.950 331.950 529.050 335.400 ;
        RECT 575.400 333.600 576.600 337.950 ;
        RECT 580.950 336.600 583.050 336.900 ;
        RECT 608.400 336.600 609.600 341.400 ;
        RECT 613.950 341.400 634.050 342.600 ;
        RECT 613.950 340.950 616.050 341.400 ;
        RECT 631.950 340.950 634.050 341.400 ;
        RECT 637.950 342.600 640.050 343.050 ;
        RECT 730.950 342.600 733.050 343.050 ;
        RECT 637.950 341.400 733.050 342.600 ;
        RECT 637.950 340.950 640.050 341.400 ;
        RECT 730.950 340.950 733.050 341.400 ;
        RECT 745.950 342.600 748.050 343.050 ;
        RECT 751.950 342.600 754.050 343.050 ;
        RECT 745.950 341.400 754.050 342.600 ;
        RECT 745.950 340.950 748.050 341.400 ;
        RECT 751.950 340.950 754.050 341.400 ;
        RECT 760.950 342.600 763.050 343.050 ;
        RECT 781.950 342.600 784.050 343.050 ;
        RECT 760.950 341.400 784.050 342.600 ;
        RECT 760.950 340.950 763.050 341.400 ;
        RECT 781.950 340.950 784.050 341.400 ;
        RECT 835.950 340.950 838.050 343.050 ;
        RECT 898.950 342.600 901.050 343.050 ;
        RECT 907.950 342.600 910.050 343.050 ;
        RECT 898.950 341.400 910.050 342.600 ;
        RECT 898.950 340.950 901.050 341.400 ;
        RECT 907.950 340.950 910.050 341.400 ;
        RECT 637.950 338.100 640.050 340.200 ;
        RECT 638.400 336.600 639.600 338.100 ;
        RECT 646.950 336.600 649.050 340.050 ;
        RECT 652.950 339.600 655.050 340.050 ;
        RECT 664.950 339.750 667.050 340.200 ;
        RECT 685.950 339.750 688.050 340.200 ;
        RECT 652.950 338.400 663.600 339.600 ;
        RECT 652.950 337.950 655.050 338.400 ;
        RECT 580.950 335.400 600.600 336.600 ;
        RECT 608.400 335.400 639.600 336.600 ;
        RECT 641.400 336.000 649.050 336.600 ;
        RECT 662.400 336.600 663.600 338.400 ;
        RECT 664.950 338.550 688.050 339.750 ;
        RECT 693.000 339.600 697.050 340.050 ;
        RECT 664.950 338.100 667.050 338.550 ;
        RECT 685.950 338.100 688.050 338.550 ;
        RECT 692.400 337.950 697.050 339.600 ;
        RECT 715.950 339.750 718.050 340.200 ;
        RECT 724.950 339.750 727.050 340.200 ;
        RECT 715.950 338.550 727.050 339.750 ;
        RECT 715.950 338.100 718.050 338.550 ;
        RECT 724.950 338.100 727.050 338.550 ;
        RECT 799.950 337.950 802.050 340.050 ;
        RECT 814.950 339.600 817.050 340.200 ;
        RECT 826.950 339.750 829.050 340.200 ;
        RECT 832.950 339.750 835.050 340.200 ;
        RECT 826.950 339.600 835.050 339.750 ;
        RECT 814.950 338.550 835.050 339.600 ;
        RECT 814.950 338.400 829.050 338.550 ;
        RECT 814.950 338.100 817.050 338.400 ;
        RECT 826.950 338.100 829.050 338.400 ;
        RECT 832.950 338.100 835.050 338.550 ;
        RECT 662.400 336.000 672.600 336.600 ;
        RECT 641.400 335.400 648.600 336.000 ;
        RECT 662.400 335.400 673.050 336.000 ;
        RECT 580.950 334.800 583.050 335.400 ;
        RECT 583.950 333.600 586.050 334.050 ;
        RECT 599.400 333.900 600.600 335.400 ;
        RECT 592.950 333.600 595.050 333.900 ;
        RECT 574.950 331.500 577.050 333.600 ;
        RECT 583.950 332.400 595.050 333.600 ;
        RECT 583.950 331.950 586.050 332.400 ;
        RECT 592.950 331.800 595.050 332.400 ;
        RECT 598.950 331.800 601.050 333.900 ;
        RECT 619.950 333.600 622.050 333.900 ;
        RECT 635.400 333.600 636.600 335.400 ;
        RECT 641.400 333.900 642.600 335.400 ;
        RECT 619.950 332.400 636.600 333.600 ;
        RECT 619.950 331.800 622.050 332.400 ;
        RECT 640.950 331.800 643.050 333.900 ;
        RECT 670.950 331.950 673.050 335.400 ;
        RECT 692.400 333.600 693.600 337.950 ;
        RECT 763.950 336.600 766.050 337.050 ;
        RECT 755.400 335.400 766.050 336.600 ;
        RECT 755.400 333.900 756.600 335.400 ;
        RECT 763.950 334.950 766.050 335.400 ;
        RECT 800.400 334.050 801.600 337.950 ;
        RECT 691.950 331.500 694.050 333.600 ;
        RECT 754.950 331.800 757.050 333.900 ;
        RECT 782.400 332.400 795.600 333.600 ;
        RECT 41.400 329.400 46.050 331.050 ;
        RECT 42.000 328.950 46.050 329.400 ;
        RECT 64.950 329.400 69.600 331.050 ;
        RECT 205.950 330.600 208.050 331.050 ;
        RECT 214.950 330.600 217.050 331.050 ;
        RECT 205.950 329.400 217.050 330.600 ;
        RECT 64.950 328.950 69.000 329.400 ;
        RECT 205.950 328.950 208.050 329.400 ;
        RECT 214.950 328.950 217.050 329.400 ;
        RECT 262.950 330.600 265.050 331.050 ;
        RECT 268.950 330.600 271.050 331.050 ;
        RECT 262.950 329.400 271.050 330.600 ;
        RECT 262.950 328.950 265.050 329.400 ;
        RECT 268.950 328.950 271.050 329.400 ;
        RECT 328.800 330.000 331.050 331.050 ;
        RECT 352.950 330.600 355.050 331.050 ;
        RECT 382.950 330.600 385.050 331.050 ;
        RECT 328.800 328.950 330.900 330.000 ;
        RECT 352.950 329.400 385.050 330.600 ;
        RECT 352.950 328.950 355.050 329.400 ;
        RECT 382.950 328.950 385.050 329.400 ;
        RECT 409.950 330.600 412.050 331.050 ;
        RECT 415.950 330.600 418.050 331.050 ;
        RECT 409.950 329.400 418.050 330.600 ;
        RECT 409.950 328.950 412.050 329.400 ;
        RECT 415.950 328.950 418.050 329.400 ;
        RECT 457.950 330.600 460.050 331.050 ;
        RECT 472.950 330.600 475.050 331.050 ;
        RECT 457.950 329.400 475.050 330.600 ;
        RECT 457.950 328.950 460.050 329.400 ;
        RECT 472.950 328.950 475.050 329.400 ;
        RECT 490.950 330.600 493.050 331.050 ;
        RECT 529.950 330.600 532.050 331.050 ;
        RECT 490.950 329.400 532.050 330.600 ;
        RECT 490.950 328.950 493.050 329.400 ;
        RECT 529.950 328.950 532.050 329.400 ;
        RECT 769.950 330.600 772.050 331.050 ;
        RECT 782.400 330.600 783.600 332.400 ;
        RECT 769.950 329.400 783.600 330.600 ;
        RECT 794.400 330.600 795.600 332.400 ;
        RECT 799.950 331.950 802.050 334.050 ;
        RECT 836.400 333.900 837.600 340.950 ;
        RECT 838.950 339.600 841.050 340.200 ;
        RECT 865.950 339.600 868.050 340.050 ;
        RECT 838.950 338.400 843.600 339.600 ;
        RECT 838.950 338.100 841.050 338.400 ;
        RECT 817.950 333.600 820.050 333.900 ;
        RECT 803.400 332.400 820.050 333.600 ;
        RECT 803.400 330.600 804.600 332.400 ;
        RECT 817.950 331.800 820.050 332.400 ;
        RECT 835.950 331.800 838.050 333.900 ;
        RECT 842.400 331.050 843.600 338.400 ;
        RECT 865.950 338.400 873.600 339.600 ;
        RECT 865.950 337.950 868.050 338.400 ;
        RECT 872.400 334.050 873.600 338.400 ;
        RECT 886.950 337.950 889.050 340.050 ;
        RECT 901.950 337.950 904.050 340.050 ;
        RECT 887.400 334.050 888.600 337.950 ;
        RECT 902.400 334.050 903.600 337.950 ;
        RECT 871.950 331.950 874.050 334.050 ;
        RECT 886.950 331.950 889.050 334.050 ;
        RECT 901.950 331.950 904.050 334.050 ;
        RECT 794.400 329.400 804.600 330.600 ;
        RECT 838.950 329.400 843.600 331.050 ;
        RECT 769.950 328.950 772.050 329.400 ;
        RECT 838.950 328.950 843.000 329.400 ;
        RECT 34.950 327.600 37.050 328.050 ;
        RECT 49.950 327.600 52.050 328.050 ;
        RECT 34.950 326.400 52.050 327.600 ;
        RECT 34.950 325.950 37.050 326.400 ;
        RECT 49.950 325.950 52.050 326.400 ;
        RECT 88.950 327.600 91.050 328.050 ;
        RECT 103.950 327.600 106.050 328.050 ;
        RECT 88.950 326.400 106.050 327.600 ;
        RECT 88.950 325.950 91.050 326.400 ;
        RECT 103.950 325.950 106.050 326.400 ;
        RECT 109.950 327.600 112.050 328.050 ;
        RECT 127.950 327.600 130.050 328.050 ;
        RECT 109.950 326.400 130.050 327.600 ;
        RECT 109.950 325.950 112.050 326.400 ;
        RECT 127.950 325.950 130.050 326.400 ;
        RECT 160.950 327.600 163.050 328.050 ;
        RECT 172.950 327.600 175.050 328.050 ;
        RECT 196.950 327.600 199.050 328.050 ;
        RECT 160.950 326.400 199.050 327.600 ;
        RECT 160.950 325.950 163.050 326.400 ;
        RECT 172.950 325.950 175.050 326.400 ;
        RECT 196.950 325.950 199.050 326.400 ;
        RECT 247.950 327.600 250.050 328.050 ;
        RECT 256.950 327.600 259.050 328.050 ;
        RECT 247.950 326.400 259.050 327.600 ;
        RECT 247.950 325.950 250.050 326.400 ;
        RECT 256.950 325.950 259.050 326.400 ;
        RECT 283.950 327.600 286.050 328.050 ;
        RECT 340.950 327.600 343.050 328.050 ;
        RECT 283.950 326.400 343.050 327.600 ;
        RECT 283.950 325.950 286.050 326.400 ;
        RECT 340.950 325.950 343.050 326.400 ;
        RECT 349.950 327.600 352.050 328.050 ;
        RECT 394.950 327.600 397.050 328.050 ;
        RECT 349.950 326.400 397.050 327.600 ;
        RECT 349.950 325.950 352.050 326.400 ;
        RECT 394.950 325.950 397.050 326.400 ;
        RECT 475.950 327.600 478.050 328.050 ;
        RECT 484.950 327.600 487.050 328.050 ;
        RECT 475.950 326.400 487.050 327.600 ;
        RECT 475.950 325.950 478.050 326.400 ;
        RECT 484.950 325.950 487.050 326.400 ;
        RECT 538.950 327.600 541.050 328.050 ;
        RECT 586.950 327.600 589.050 328.050 ;
        RECT 538.950 326.400 589.050 327.600 ;
        RECT 538.950 325.950 541.050 326.400 ;
        RECT 586.950 325.950 589.050 326.400 ;
        RECT 592.950 327.600 595.050 328.050 ;
        RECT 601.950 327.600 604.050 328.050 ;
        RECT 592.950 326.400 604.050 327.600 ;
        RECT 592.950 325.950 595.050 326.400 ;
        RECT 601.950 325.950 604.050 326.400 ;
        RECT 727.950 327.600 730.050 328.050 ;
        RECT 754.950 327.600 757.050 328.050 ;
        RECT 727.950 326.400 757.050 327.600 ;
        RECT 727.950 325.950 730.050 326.400 ;
        RECT 754.950 325.950 757.050 326.400 ;
        RECT 826.950 327.600 829.050 328.050 ;
        RECT 859.950 327.600 862.050 328.050 ;
        RECT 826.950 326.400 862.050 327.600 ;
        RECT 826.950 325.950 829.050 326.400 ;
        RECT 859.950 325.950 862.050 326.400 ;
        RECT 67.950 324.600 70.050 325.050 ;
        RECT 110.400 324.600 111.600 325.950 ;
        RECT 67.950 323.400 111.600 324.600 ;
        RECT 166.950 324.600 169.050 325.050 ;
        RECT 178.950 324.600 181.050 325.050 ;
        RECT 166.950 323.400 181.050 324.600 ;
        RECT 67.950 322.950 70.050 323.400 ;
        RECT 166.950 322.950 169.050 323.400 ;
        RECT 178.950 322.950 181.050 323.400 ;
        RECT 190.950 324.600 193.050 325.050 ;
        RECT 208.950 324.600 211.050 325.050 ;
        RECT 190.950 323.400 211.050 324.600 ;
        RECT 190.950 322.950 193.050 323.400 ;
        RECT 208.950 322.950 211.050 323.400 ;
        RECT 238.950 324.600 241.050 325.050 ;
        RECT 259.950 324.600 262.050 325.050 ;
        RECT 238.950 323.400 262.050 324.600 ;
        RECT 238.950 322.950 241.050 323.400 ;
        RECT 259.950 322.950 262.050 323.400 ;
        RECT 304.950 324.600 307.050 325.050 ;
        RECT 334.950 324.600 337.050 325.050 ;
        RECT 304.950 323.400 337.050 324.600 ;
        RECT 304.950 322.950 307.050 323.400 ;
        RECT 334.950 322.950 337.050 323.400 ;
        RECT 343.950 324.600 346.050 325.050 ;
        RECT 352.950 324.600 355.050 325.050 ;
        RECT 343.950 323.400 355.050 324.600 ;
        RECT 343.950 322.950 346.050 323.400 ;
        RECT 352.950 322.950 355.050 323.400 ;
        RECT 361.950 324.600 364.050 325.050 ;
        RECT 391.950 324.600 394.050 325.050 ;
        RECT 361.950 323.400 394.050 324.600 ;
        RECT 361.950 322.950 364.050 323.400 ;
        RECT 391.950 322.950 394.050 323.400 ;
        RECT 445.950 324.600 448.050 325.050 ;
        RECT 487.950 324.600 490.050 325.050 ;
        RECT 445.950 323.400 490.050 324.600 ;
        RECT 445.950 322.950 448.050 323.400 ;
        RECT 487.950 322.950 490.050 323.400 ;
        RECT 556.950 324.600 559.050 325.050 ;
        RECT 580.950 324.600 583.050 325.050 ;
        RECT 556.950 323.400 583.050 324.600 ;
        RECT 556.950 322.950 559.050 323.400 ;
        RECT 580.950 322.950 583.050 323.400 ;
        RECT 589.950 324.600 592.050 325.050 ;
        RECT 655.950 324.600 658.050 325.050 ;
        RECT 589.950 323.400 658.050 324.600 ;
        RECT 589.950 322.950 592.050 323.400 ;
        RECT 655.950 322.950 658.050 323.400 ;
        RECT 688.950 324.600 691.050 325.050 ;
        RECT 718.950 324.600 721.050 325.050 ;
        RECT 688.950 323.400 721.050 324.600 ;
        RECT 688.950 322.950 691.050 323.400 ;
        RECT 718.950 322.950 721.050 323.400 ;
        RECT 814.950 324.600 817.050 325.050 ;
        RECT 847.950 324.600 850.050 325.050 ;
        RECT 814.950 323.400 850.050 324.600 ;
        RECT 814.950 322.950 817.050 323.400 ;
        RECT 847.950 322.950 850.050 323.400 ;
        RECT 31.950 321.600 34.050 322.050 ;
        RECT 115.950 321.600 118.050 322.050 ;
        RECT 229.950 321.600 232.050 322.050 ;
        RECT 31.950 320.400 118.050 321.600 ;
        RECT 31.950 319.950 34.050 320.400 ;
        RECT 115.950 319.950 118.050 320.400 ;
        RECT 212.400 320.400 232.050 321.600 ;
        RECT 19.950 318.600 22.050 319.050 ;
        RECT 28.950 318.600 31.050 319.050 ;
        RECT 19.950 317.400 31.050 318.600 ;
        RECT 19.950 316.950 22.050 317.400 ;
        RECT 28.950 316.950 31.050 317.400 ;
        RECT 40.950 318.600 43.050 319.050 ;
        RECT 88.950 318.600 91.050 319.050 ;
        RECT 40.950 317.400 91.050 318.600 ;
        RECT 40.950 316.950 43.050 317.400 ;
        RECT 88.950 316.950 91.050 317.400 ;
        RECT 196.950 318.600 199.050 319.050 ;
        RECT 212.400 318.600 213.600 320.400 ;
        RECT 229.950 319.950 232.050 320.400 ;
        RECT 241.950 321.600 244.050 322.050 ;
        RECT 250.950 321.600 253.050 322.050 ;
        RECT 241.950 320.400 253.050 321.600 ;
        RECT 241.950 319.950 244.050 320.400 ;
        RECT 250.950 319.950 253.050 320.400 ;
        RECT 295.950 321.600 298.050 321.900 ;
        RECT 364.950 321.600 367.050 322.050 ;
        RECT 442.950 321.600 445.050 322.050 ;
        RECT 295.950 320.400 348.600 321.600 ;
        RECT 295.950 319.800 298.050 320.400 ;
        RECT 196.950 317.400 213.600 318.600 ;
        RECT 347.400 318.600 348.600 320.400 ;
        RECT 364.950 320.400 445.050 321.600 ;
        RECT 364.950 319.950 367.050 320.400 ;
        RECT 442.950 319.950 445.050 320.400 ;
        RECT 565.950 321.600 568.050 322.050 ;
        RECT 577.950 321.600 580.050 322.050 ;
        RECT 565.950 320.400 580.050 321.600 ;
        RECT 565.950 319.950 568.050 320.400 ;
        RECT 577.950 319.950 580.050 320.400 ;
        RECT 691.950 321.600 694.050 322.050 ;
        RECT 724.950 321.600 727.050 322.050 ;
        RECT 691.950 320.400 727.050 321.600 ;
        RECT 691.950 319.950 694.050 320.400 ;
        RECT 724.950 319.950 727.050 320.400 ;
        RECT 361.950 318.600 364.050 319.050 ;
        RECT 370.950 318.600 373.050 319.050 ;
        RECT 347.400 317.400 373.050 318.600 ;
        RECT 196.950 316.950 199.050 317.400 ;
        RECT 361.950 316.950 364.050 317.400 ;
        RECT 370.950 316.950 373.050 317.400 ;
        RECT 586.950 318.600 589.050 319.050 ;
        RECT 610.950 318.600 613.050 319.050 ;
        RECT 586.950 317.400 613.050 318.600 ;
        RECT 586.950 316.950 589.050 317.400 ;
        RECT 610.950 316.950 613.050 317.400 ;
        RECT 667.950 318.600 670.050 319.050 ;
        RECT 673.950 318.600 676.050 319.050 ;
        RECT 667.950 317.400 676.050 318.600 ;
        RECT 667.950 316.950 670.050 317.400 ;
        RECT 673.950 316.950 676.050 317.400 ;
        RECT 811.950 318.600 814.050 319.050 ;
        RECT 865.950 318.600 868.050 319.050 ;
        RECT 811.950 317.400 868.050 318.600 ;
        RECT 811.950 316.950 814.050 317.400 ;
        RECT 865.950 316.950 868.050 317.400 ;
        RECT 256.950 315.600 259.050 316.050 ;
        RECT 274.950 315.600 277.050 316.050 ;
        RECT 298.800 315.600 300.900 316.050 ;
        RECT 245.400 314.400 255.600 315.600 ;
        RECT 238.950 312.600 241.050 313.050 ;
        RECT 245.400 312.600 246.600 314.400 ;
        RECT 238.950 311.400 246.600 312.600 ;
        RECT 254.400 312.600 255.600 314.400 ;
        RECT 256.950 314.400 300.900 315.600 ;
        RECT 256.950 313.950 259.050 314.400 ;
        RECT 274.950 313.950 277.050 314.400 ;
        RECT 298.800 313.950 300.900 314.400 ;
        RECT 301.950 315.600 304.050 316.050 ;
        RECT 355.950 315.600 358.050 316.050 ;
        RECT 301.950 314.400 358.050 315.600 ;
        RECT 301.950 313.950 304.050 314.400 ;
        RECT 355.950 313.950 358.050 314.400 ;
        RECT 382.950 315.600 385.050 316.050 ;
        RECT 400.950 315.600 403.050 316.050 ;
        RECT 382.950 314.400 403.050 315.600 ;
        RECT 382.950 313.950 385.050 314.400 ;
        RECT 400.950 313.950 403.050 314.400 ;
        RECT 649.950 315.600 652.050 316.050 ;
        RECT 691.950 315.600 694.050 316.050 ;
        RECT 649.950 314.400 694.050 315.600 ;
        RECT 649.950 313.950 652.050 314.400 ;
        RECT 691.950 313.950 694.050 314.400 ;
        RECT 706.950 315.600 709.050 316.050 ;
        RECT 739.950 315.600 742.050 316.050 ;
        RECT 706.950 314.400 742.050 315.600 ;
        RECT 706.950 313.950 709.050 314.400 ;
        RECT 739.950 313.950 742.050 314.400 ;
        RECT 766.950 315.600 769.050 316.050 ;
        RECT 805.950 315.600 808.050 316.050 ;
        RECT 766.950 314.400 808.050 315.600 ;
        RECT 766.950 313.950 769.050 314.400 ;
        RECT 805.950 313.950 808.050 314.400 ;
        RECT 835.950 315.600 838.050 316.050 ;
        RECT 877.950 315.600 880.050 316.050 ;
        RECT 835.950 314.400 880.050 315.600 ;
        RECT 835.950 313.950 838.050 314.400 ;
        RECT 877.950 313.950 880.050 314.400 ;
        RECT 295.950 312.600 298.050 313.050 ;
        RECT 254.400 311.400 298.050 312.600 ;
        RECT 238.950 310.950 241.050 311.400 ;
        RECT 295.950 310.950 298.050 311.400 ;
        RECT 316.950 312.600 319.050 313.050 ;
        RECT 322.950 312.600 325.050 313.050 ;
        RECT 316.950 311.400 325.050 312.600 ;
        RECT 316.950 310.950 319.050 311.400 ;
        RECT 322.950 310.950 325.050 311.400 ;
        RECT 379.950 312.600 382.050 313.050 ;
        RECT 412.950 312.600 415.050 313.050 ;
        RECT 517.950 312.600 520.050 313.050 ;
        RECT 379.950 311.400 520.050 312.600 ;
        RECT 379.950 310.950 382.050 311.400 ;
        RECT 412.950 310.950 415.050 311.400 ;
        RECT 517.950 310.950 520.050 311.400 ;
        RECT 538.950 312.600 541.050 313.050 ;
        RECT 598.950 312.600 601.050 313.050 ;
        RECT 631.950 312.600 634.050 313.050 ;
        RECT 538.950 311.400 634.050 312.600 ;
        RECT 538.950 310.950 541.050 311.400 ;
        RECT 598.950 310.950 601.050 311.400 ;
        RECT 631.950 310.950 634.050 311.400 ;
        RECT 661.950 312.600 664.050 313.050 ;
        RECT 688.950 312.600 691.050 313.050 ;
        RECT 661.950 311.400 691.050 312.600 ;
        RECT 661.950 310.950 664.050 311.400 ;
        RECT 688.950 310.950 691.050 311.400 ;
        RECT 787.950 312.600 790.050 313.050 ;
        RECT 802.950 312.600 805.050 313.050 ;
        RECT 787.950 311.400 805.050 312.600 ;
        RECT 787.950 310.950 790.050 311.400 ;
        RECT 802.950 310.950 805.050 311.400 ;
        RECT 43.950 309.600 46.050 310.050 ;
        RECT 88.950 309.600 91.050 310.050 ;
        RECT 43.950 308.400 91.050 309.600 ;
        RECT 43.950 307.950 46.050 308.400 ;
        RECT 88.950 307.950 91.050 308.400 ;
        RECT 154.950 309.600 157.050 310.050 ;
        RECT 211.950 309.600 214.050 310.050 ;
        RECT 154.950 308.400 214.050 309.600 ;
        RECT 154.950 307.950 157.050 308.400 ;
        RECT 211.950 307.950 214.050 308.400 ;
        RECT 229.950 309.600 232.050 310.050 ;
        RECT 235.950 309.600 238.050 310.050 ;
        RECT 229.950 308.400 238.050 309.600 ;
        RECT 229.950 307.950 232.050 308.400 ;
        RECT 235.950 307.950 238.050 308.400 ;
        RECT 247.950 309.600 250.050 310.050 ;
        RECT 334.950 309.600 337.050 310.050 ;
        RECT 247.950 308.400 337.050 309.600 ;
        RECT 247.950 307.950 250.050 308.400 ;
        RECT 334.950 307.950 337.050 308.400 ;
        RECT 508.950 309.600 511.050 310.050 ;
        RECT 712.950 309.600 715.050 310.050 ;
        RECT 508.950 308.400 715.050 309.600 ;
        RECT 508.950 307.950 511.050 308.400 ;
        RECT 712.950 307.950 715.050 308.400 ;
        RECT 760.950 309.600 763.050 310.050 ;
        RECT 793.950 309.600 796.050 310.050 ;
        RECT 760.950 308.400 796.050 309.600 ;
        RECT 760.950 307.950 763.050 308.400 ;
        RECT 793.950 307.950 796.050 308.400 ;
        RECT 808.950 309.600 811.050 310.050 ;
        RECT 835.950 309.600 838.050 310.050 ;
        RECT 808.950 308.400 838.050 309.600 ;
        RECT 808.950 307.950 811.050 308.400 ;
        RECT 835.950 307.950 838.050 308.400 ;
        RECT 850.950 309.600 853.050 310.050 ;
        RECT 889.950 309.600 892.050 310.050 ;
        RECT 850.950 308.400 892.050 309.600 ;
        RECT 850.950 307.950 853.050 308.400 ;
        RECT 889.950 307.950 892.050 308.400 ;
        RECT 133.950 306.600 136.050 307.050 ;
        RECT 202.950 306.600 205.050 307.050 ;
        RECT 133.950 305.400 205.050 306.600 ;
        RECT 133.950 304.950 136.050 305.400 ;
        RECT 202.950 304.950 205.050 305.400 ;
        RECT 217.950 306.600 220.050 307.050 ;
        RECT 238.800 306.600 240.900 307.050 ;
        RECT 217.950 305.400 240.900 306.600 ;
        RECT 217.950 304.950 220.050 305.400 ;
        RECT 238.800 304.950 240.900 305.400 ;
        RECT 532.950 306.600 535.050 307.050 ;
        RECT 547.950 306.600 550.050 307.050 ;
        RECT 706.950 306.600 709.050 307.050 ;
        RECT 532.950 305.400 550.050 306.600 ;
        RECT 532.950 304.950 535.050 305.400 ;
        RECT 547.950 304.950 550.050 305.400 ;
        RECT 680.400 305.400 709.050 306.600 ;
        RECT 13.950 303.600 16.050 304.050 ;
        RECT 43.950 303.600 46.050 304.050 ;
        RECT 13.950 302.400 46.050 303.600 ;
        RECT 13.950 301.950 16.050 302.400 ;
        RECT 43.950 301.950 46.050 302.400 ;
        RECT 79.950 303.600 82.050 304.050 ;
        RECT 91.950 303.600 94.050 304.050 ;
        RECT 79.950 302.400 94.050 303.600 ;
        RECT 79.950 301.950 82.050 302.400 ;
        RECT 91.950 301.950 94.050 302.400 ;
        RECT 103.950 303.600 106.050 304.050 ;
        RECT 115.950 303.600 118.050 304.050 ;
        RECT 103.950 302.400 118.050 303.600 ;
        RECT 103.950 301.950 106.050 302.400 ;
        RECT 115.950 301.950 118.050 302.400 ;
        RECT 310.950 303.600 313.050 304.050 ;
        RECT 349.950 303.600 352.050 304.050 ;
        RECT 310.950 302.400 352.050 303.600 ;
        RECT 310.950 301.950 313.050 302.400 ;
        RECT 118.950 300.600 121.050 301.050 ;
        RECT 136.950 300.600 139.050 301.050 ;
        RECT 118.950 299.400 139.050 300.600 ;
        RECT 118.950 298.950 121.050 299.400 ;
        RECT 136.950 298.950 139.050 299.400 ;
        RECT 148.950 300.600 151.050 301.050 ;
        RECT 220.950 300.600 223.050 301.050 ;
        RECT 256.950 300.600 259.050 301.050 ;
        RECT 148.950 299.400 174.600 300.600 ;
        RECT 148.950 298.950 151.050 299.400 ;
        RECT 173.400 298.050 174.600 299.400 ;
        RECT 220.950 299.400 259.050 300.600 ;
        RECT 220.950 298.950 223.050 299.400 ;
        RECT 256.950 298.950 259.050 299.400 ;
        RECT 322.950 298.800 325.050 302.400 ;
        RECT 349.950 301.950 352.050 302.400 ;
        RECT 367.950 303.600 370.050 304.050 ;
        RECT 406.950 303.600 409.050 304.050 ;
        RECT 481.950 303.600 484.050 304.050 ;
        RECT 622.950 303.600 625.050 304.050 ;
        RECT 680.400 303.600 681.600 305.400 ;
        RECT 706.950 304.950 709.050 305.400 ;
        RECT 367.950 302.400 507.600 303.600 ;
        RECT 367.950 301.950 370.050 302.400 ;
        RECT 406.950 301.950 409.050 302.400 ;
        RECT 481.950 301.950 484.050 302.400 ;
        RECT 506.400 301.050 507.600 302.400 ;
        RECT 622.950 302.400 657.600 303.600 ;
        RECT 622.950 301.950 625.050 302.400 ;
        RECT 334.950 300.600 337.050 301.050 ;
        RECT 343.950 300.600 346.050 301.050 ;
        RECT 358.950 300.600 361.050 301.050 ;
        RECT 334.950 299.400 342.600 300.600 ;
        RECT 334.950 298.950 337.050 299.400 ;
        RECT 58.950 297.600 61.050 298.050 ;
        RECT 73.950 297.600 76.050 298.050 ;
        RECT 115.950 297.600 118.050 298.050 ;
        RECT 58.950 296.400 118.050 297.600 ;
        RECT 58.950 295.950 61.050 296.400 ;
        RECT 73.950 295.950 76.050 296.400 ;
        RECT 115.950 295.950 118.050 296.400 ;
        RECT 172.950 297.600 175.050 298.050 ;
        RECT 196.950 297.600 199.050 298.050 ;
        RECT 172.950 296.400 199.050 297.600 ;
        RECT 172.950 295.950 175.050 296.400 ;
        RECT 196.950 295.950 199.050 296.400 ;
        RECT 310.950 297.600 313.050 298.050 ;
        RECT 316.950 297.600 319.050 298.050 ;
        RECT 310.950 296.400 319.050 297.600 ;
        RECT 341.400 297.600 342.600 299.400 ;
        RECT 343.950 299.400 361.050 300.600 ;
        RECT 343.950 298.950 346.050 299.400 ;
        RECT 358.950 298.950 361.050 299.400 ;
        RECT 364.950 297.600 367.050 301.050 ;
        RECT 379.950 300.600 382.050 301.050 ;
        RECT 502.800 300.600 504.900 301.050 ;
        RECT 379.950 299.400 504.900 300.600 ;
        RECT 379.950 298.950 382.050 299.400 ;
        RECT 502.800 298.950 504.900 299.400 ;
        RECT 505.950 300.600 508.050 301.050 ;
        RECT 526.950 300.600 529.050 301.050 ;
        RECT 505.950 299.400 529.050 300.600 ;
        RECT 505.950 298.950 508.050 299.400 ;
        RECT 526.950 298.950 529.050 299.400 ;
        RECT 637.950 300.600 640.050 301.050 ;
        RECT 646.950 300.600 649.050 301.050 ;
        RECT 637.950 299.400 649.050 300.600 ;
        RECT 656.400 300.600 657.600 302.400 ;
        RECT 677.400 302.400 681.600 303.600 ;
        RECT 682.950 303.600 685.050 304.050 ;
        RECT 691.950 303.600 694.050 304.050 ;
        RECT 682.950 302.400 694.050 303.600 ;
        RECT 670.950 300.600 673.050 300.900 ;
        RECT 656.400 299.400 673.050 300.600 ;
        RECT 637.950 298.950 640.050 299.400 ;
        RECT 646.950 298.950 649.050 299.400 ;
        RECT 670.950 298.800 673.050 299.400 ;
        RECT 677.400 298.050 678.600 302.400 ;
        RECT 682.950 301.950 685.050 302.400 ;
        RECT 691.950 301.950 694.050 302.400 ;
        RECT 730.950 303.600 733.050 304.050 ;
        RECT 817.950 303.600 820.050 304.050 ;
        RECT 730.950 302.400 820.050 303.600 ;
        RECT 730.950 301.950 733.050 302.400 ;
        RECT 817.950 301.950 820.050 302.400 ;
        RECT 865.950 303.600 868.050 304.050 ;
        RECT 892.950 303.600 895.050 304.050 ;
        RECT 904.950 303.600 907.050 304.050 ;
        RECT 865.950 302.400 907.050 303.600 ;
        RECT 865.950 301.950 868.050 302.400 ;
        RECT 892.950 301.950 895.050 302.400 ;
        RECT 904.950 301.950 907.050 302.400 ;
        RECT 775.950 300.600 778.050 301.050 ;
        RECT 808.950 300.600 811.050 301.050 ;
        RECT 775.950 299.400 811.050 300.600 ;
        RECT 775.950 298.950 778.050 299.400 ;
        RECT 808.950 298.950 811.050 299.400 ;
        RECT 844.950 300.600 847.050 301.050 ;
        RECT 850.950 300.600 853.050 301.050 ;
        RECT 844.950 299.400 853.050 300.600 ;
        RECT 844.950 298.950 847.050 299.400 ;
        RECT 850.950 298.950 853.050 299.400 ;
        RECT 341.400 297.000 367.050 297.600 ;
        RECT 388.950 297.600 391.050 298.050 ;
        RECT 427.950 297.600 430.050 298.050 ;
        RECT 341.400 296.400 366.600 297.000 ;
        RECT 388.950 296.400 430.050 297.600 ;
        RECT 310.950 295.950 313.050 296.400 ;
        RECT 316.950 295.950 319.050 296.400 ;
        RECT 388.950 295.950 391.050 296.400 ;
        RECT 427.950 295.950 430.050 296.400 ;
        RECT 532.950 297.600 535.050 298.050 ;
        RECT 544.950 297.600 547.050 298.050 ;
        RECT 586.950 297.600 589.050 298.050 ;
        RECT 532.950 296.400 547.050 297.600 ;
        RECT 532.950 295.950 535.050 296.400 ;
        RECT 544.950 295.950 547.050 296.400 ;
        RECT 551.400 296.400 589.050 297.600 ;
        RECT 677.400 296.400 682.050 298.050 ;
        RECT 16.950 293.100 19.050 295.200 ;
        RECT 17.400 286.050 18.600 293.100 ;
        RECT 25.950 292.950 28.050 295.050 ;
        RECT 37.950 293.100 40.050 295.200 ;
        RECT 43.950 294.600 46.050 295.200 ;
        RECT 43.950 293.400 48.600 294.600 ;
        RECT 43.950 293.100 46.050 293.400 ;
        RECT 26.400 289.050 27.600 292.950 ;
        RECT 25.950 286.950 28.050 289.050 ;
        RECT 31.950 288.600 34.050 289.050 ;
        RECT 38.400 288.600 39.600 293.100 ;
        RECT 47.400 289.050 48.600 293.400 ;
        RECT 52.950 292.950 55.050 295.050 ;
        RECT 64.950 294.600 67.050 295.200 ;
        RECT 79.950 294.600 82.050 295.200 ;
        RECT 64.950 293.400 82.050 294.600 ;
        RECT 64.950 293.100 67.050 293.400 ;
        RECT 79.950 293.100 82.050 293.400 ;
        RECT 94.800 294.000 96.900 295.050 ;
        RECT 97.950 294.600 100.050 295.200 ;
        RECT 112.950 294.600 115.050 295.050 ;
        RECT 94.800 292.950 97.050 294.000 ;
        RECT 97.950 293.400 115.050 294.600 ;
        RECT 97.950 293.100 100.050 293.400 ;
        RECT 112.950 292.950 115.050 293.400 ;
        RECT 121.950 293.100 124.050 295.200 ;
        RECT 127.950 293.100 130.050 295.200 ;
        RECT 53.400 289.050 54.600 292.950 ;
        RECT 94.950 291.600 97.050 292.950 ;
        RECT 122.400 291.600 123.600 293.100 ;
        RECT 94.950 291.000 99.600 291.600 ;
        RECT 119.400 291.000 123.600 291.600 ;
        RECT 95.400 290.400 99.600 291.000 ;
        RECT 98.400 289.050 99.600 290.400 ;
        RECT 31.950 287.400 39.600 288.600 ;
        RECT 31.950 286.950 34.050 287.400 ;
        RECT 46.950 286.950 49.050 289.050 ;
        RECT 52.950 286.950 55.050 289.050 ;
        RECT 61.950 288.600 64.050 288.900 ;
        RECT 76.950 288.600 79.050 288.900 ;
        RECT 61.950 288.450 79.050 288.600 ;
        RECT 88.950 288.450 91.050 288.900 ;
        RECT 61.950 287.400 91.050 288.450 ;
        RECT 61.950 286.800 64.050 287.400 ;
        RECT 76.950 287.250 91.050 287.400 ;
        RECT 76.950 286.800 79.050 287.250 ;
        RECT 88.950 286.800 91.050 287.250 ;
        RECT 94.950 288.600 99.600 289.050 ;
        RECT 118.950 290.400 123.600 291.000 ;
        RECT 100.950 288.600 103.050 288.900 ;
        RECT 94.950 287.400 103.050 288.600 ;
        RECT 94.950 286.950 99.000 287.400 ;
        RECT 100.950 286.800 103.050 287.400 ;
        RECT 118.950 286.950 121.050 290.400 ;
        RECT 128.400 286.050 129.600 293.100 ;
        RECT 133.950 291.600 136.050 295.050 ;
        RECT 142.950 294.750 145.050 295.200 ;
        RECT 154.950 294.750 157.050 295.200 ;
        RECT 142.950 293.550 157.050 294.750 ;
        RECT 142.950 293.100 145.050 293.550 ;
        RECT 154.950 293.100 157.050 293.550 ;
        RECT 166.950 293.100 169.050 295.200 ;
        RECT 184.950 294.750 187.050 295.200 ;
        RECT 190.950 294.750 193.050 295.200 ;
        RECT 184.950 293.550 193.050 294.750 ;
        RECT 201.000 294.600 205.050 295.050 ;
        RECT 184.950 293.100 187.050 293.550 ;
        RECT 190.950 293.100 193.050 293.550 ;
        RECT 131.400 291.000 136.050 291.600 ;
        RECT 131.400 290.400 135.600 291.000 ;
        RECT 131.400 288.900 132.600 290.400 ;
        RECT 130.950 286.800 133.050 288.900 ;
        RECT 136.950 288.600 139.050 289.050 ;
        RECT 145.950 288.600 148.050 288.900 ;
        RECT 136.950 287.400 148.050 288.600 ;
        RECT 136.950 286.950 139.050 287.400 ;
        RECT 145.950 286.800 148.050 287.400 ;
        RECT 151.950 288.600 154.050 288.900 ;
        RECT 167.400 288.600 168.600 293.100 ;
        RECT 200.400 292.950 205.050 294.600 ;
        RECT 223.950 294.600 226.050 295.050 ;
        RECT 229.950 294.600 232.050 295.200 ;
        RECT 223.950 293.400 232.050 294.600 ;
        RECT 223.950 292.950 226.050 293.400 ;
        RECT 229.950 293.100 232.050 293.400 ;
        RECT 241.950 294.750 244.050 295.200 ;
        RECT 253.950 294.750 256.050 295.200 ;
        RECT 241.950 293.550 256.050 294.750 ;
        RECT 241.950 293.100 244.050 293.550 ;
        RECT 253.950 293.100 256.050 293.550 ;
        RECT 277.950 294.600 280.050 295.050 ;
        RECT 289.950 294.600 292.050 295.200 ;
        RECT 313.950 294.600 316.050 295.200 ;
        RECT 277.950 293.400 288.600 294.600 ;
        RECT 277.950 292.950 280.050 293.400 ;
        RECT 200.400 288.900 201.600 292.950 ;
        RECT 287.400 291.600 288.600 293.400 ;
        RECT 289.950 293.400 316.050 294.600 ;
        RECT 289.950 293.100 292.050 293.400 ;
        RECT 313.950 293.100 316.050 293.400 ;
        RECT 319.950 294.750 322.050 295.200 ;
        RECT 334.950 294.750 337.050 295.200 ;
        RECT 319.950 294.600 337.050 294.750 ;
        RECT 370.800 294.600 372.900 295.050 ;
        RECT 319.950 293.550 372.900 294.600 ;
        RECT 319.950 293.100 322.050 293.550 ;
        RECT 334.950 293.400 372.900 293.550 ;
        RECT 334.950 293.100 337.050 293.400 ;
        RECT 370.800 292.950 372.900 293.400 ;
        RECT 376.950 294.750 379.050 295.200 ;
        RECT 385.950 294.750 388.050 295.200 ;
        RECT 376.950 293.550 388.050 294.750 ;
        RECT 376.950 293.100 379.050 293.550 ;
        RECT 385.950 293.100 388.050 293.550 ;
        RECT 400.950 293.100 403.050 295.200 ;
        RECT 436.950 294.750 439.050 295.200 ;
        RECT 442.950 294.750 445.050 295.200 ;
        RECT 436.950 293.550 445.050 294.750 ;
        RECT 436.950 293.100 439.050 293.550 ;
        RECT 442.950 293.100 445.050 293.550 ;
        RECT 451.950 294.750 454.050 295.200 ;
        RECT 460.950 294.750 463.050 295.200 ;
        RECT 451.950 293.550 463.050 294.750 ;
        RECT 451.950 293.100 454.050 293.550 ;
        RECT 460.950 293.100 463.050 293.550 ;
        RECT 487.950 294.750 490.050 295.200 ;
        RECT 493.950 294.750 496.050 295.200 ;
        RECT 487.950 293.550 496.050 294.750 ;
        RECT 487.950 293.100 490.050 293.550 ;
        RECT 493.950 293.100 496.050 293.550 ;
        RECT 502.950 294.750 505.050 295.200 ;
        RECT 511.950 294.750 514.050 295.200 ;
        RECT 502.950 294.600 514.050 294.750 ;
        RECT 551.400 294.600 552.600 296.400 ;
        RECT 586.950 295.950 589.050 296.400 ;
        RECT 678.000 295.950 682.050 296.400 ;
        RECT 694.950 297.600 697.050 298.050 ;
        RECT 709.950 297.600 712.050 298.050 ;
        RECT 694.950 296.400 712.050 297.600 ;
        RECT 694.950 295.950 697.050 296.400 ;
        RECT 709.950 295.950 712.050 296.400 ;
        RECT 733.950 297.600 736.050 298.050 ;
        RECT 745.950 297.600 748.050 298.050 ;
        RECT 733.950 296.400 748.050 297.600 ;
        RECT 733.950 295.950 736.050 296.400 ;
        RECT 745.950 295.950 748.050 296.400 ;
        RECT 751.950 297.600 754.050 298.050 ;
        RECT 763.950 297.600 766.050 298.050 ;
        RECT 751.950 296.400 766.050 297.600 ;
        RECT 751.950 295.950 754.050 296.400 ;
        RECT 763.950 295.950 766.050 296.400 ;
        RECT 829.950 297.600 832.050 298.050 ;
        RECT 838.950 297.600 841.050 298.050 ;
        RECT 829.950 296.400 841.050 297.600 ;
        RECT 829.950 295.950 832.050 296.400 ;
        RECT 838.950 295.950 841.050 296.400 ;
        RECT 868.950 297.600 871.050 298.050 ;
        RECT 877.950 297.600 880.050 298.050 ;
        RECT 868.950 296.400 880.050 297.600 ;
        RECT 868.950 295.950 871.050 296.400 ;
        RECT 877.950 295.950 880.050 296.400 ;
        RECT 502.950 293.550 552.600 294.600 ;
        RECT 502.950 293.100 505.050 293.550 ;
        RECT 511.950 293.400 552.600 293.550 ;
        RECT 553.950 294.600 556.050 295.200 ;
        RECT 568.950 294.600 571.050 295.200 ;
        RECT 553.950 293.400 571.050 294.600 ;
        RECT 511.950 293.100 514.050 293.400 ;
        RECT 553.950 293.100 556.050 293.400 ;
        RECT 568.950 293.100 571.050 293.400 ;
        RECT 574.950 294.750 577.050 295.200 ;
        RECT 583.950 294.750 586.050 295.200 ;
        RECT 574.950 293.550 586.050 294.750 ;
        RECT 574.950 293.100 577.050 293.550 ;
        RECT 583.950 293.100 586.050 293.550 ;
        RECT 592.950 293.100 595.050 295.200 ;
        RECT 346.950 291.600 349.050 292.050 ;
        RECT 287.400 290.400 349.050 291.600 ;
        RECT 346.950 289.950 349.050 290.400 ;
        RECT 401.400 289.050 402.600 293.100 ;
        RECT 412.950 291.600 415.050 292.050 ;
        RECT 593.400 291.600 594.600 293.100 ;
        RECT 631.950 292.950 634.050 295.050 ;
        RECT 640.950 293.100 643.050 295.200 ;
        RECT 658.950 293.100 661.050 295.200 ;
        RECT 664.950 293.100 667.050 295.200 ;
        RECT 688.950 294.600 691.050 295.050 ;
        RECT 697.950 294.600 700.050 295.050 ;
        RECT 688.950 293.400 700.050 294.600 ;
        RECT 412.950 290.400 447.600 291.600 ;
        RECT 412.950 289.950 415.050 290.400 ;
        RECT 151.950 287.400 168.600 288.600 ;
        RECT 175.950 288.600 178.050 288.900 ;
        RECT 199.950 288.600 202.050 288.900 ;
        RECT 175.950 287.400 202.050 288.600 ;
        RECT 151.950 286.800 154.050 287.400 ;
        RECT 175.950 286.800 178.050 287.400 ;
        RECT 199.950 286.800 202.050 287.400 ;
        RECT 244.950 288.600 247.050 289.050 ;
        RECT 292.950 288.600 295.050 288.900 ;
        RECT 244.950 287.400 295.050 288.600 ;
        RECT 244.950 286.950 247.050 287.400 ;
        RECT 292.950 286.800 295.050 287.400 ;
        RECT 364.950 288.450 367.050 288.900 ;
        RECT 373.950 288.450 376.050 288.900 ;
        RECT 364.950 287.250 376.050 288.450 ;
        RECT 364.950 286.800 367.050 287.250 ;
        RECT 373.950 286.800 376.050 287.250 ;
        RECT 397.950 287.400 402.600 289.050 ;
        RECT 446.400 288.900 447.600 290.400 ;
        RECT 542.400 290.400 594.600 291.600 ;
        RECT 397.950 286.950 402.000 287.400 ;
        RECT 445.950 286.800 448.050 288.900 ;
        RECT 472.950 288.600 475.050 289.050 ;
        RECT 478.950 288.600 481.050 288.900 ;
        RECT 472.950 288.450 481.050 288.600 ;
        RECT 484.950 288.450 487.050 288.900 ;
        RECT 472.950 287.400 487.050 288.450 ;
        RECT 472.950 286.950 475.050 287.400 ;
        RECT 478.950 287.250 487.050 287.400 ;
        RECT 478.950 286.800 481.050 287.250 ;
        RECT 484.950 286.800 487.050 287.250 ;
        RECT 529.950 288.600 532.050 288.900 ;
        RECT 542.400 288.600 543.600 290.400 ;
        RECT 529.950 287.400 543.600 288.600 ;
        RECT 544.950 288.450 547.050 288.900 ;
        RECT 556.950 288.450 559.050 288.900 ;
        RECT 529.950 286.800 532.050 287.400 ;
        RECT 544.950 287.250 559.050 288.450 ;
        RECT 544.950 286.800 547.050 287.250 ;
        RECT 556.950 286.800 559.050 287.250 ;
        RECT 604.950 288.600 607.050 289.050 ;
        RECT 613.950 288.600 616.050 288.900 ;
        RECT 604.950 287.400 616.050 288.600 ;
        RECT 632.400 288.600 633.600 292.950 ;
        RECT 641.400 291.600 642.600 293.100 ;
        RECT 641.400 290.400 645.600 291.600 ;
        RECT 644.400 289.050 645.600 290.400 ;
        RECT 637.950 288.600 640.050 288.900 ;
        RECT 632.400 287.400 640.050 288.600 ;
        RECT 644.400 287.400 649.050 289.050 ;
        RECT 604.950 286.950 607.050 287.400 ;
        RECT 613.950 286.800 616.050 287.400 ;
        RECT 637.950 286.800 640.050 287.400 ;
        RECT 645.000 286.950 649.050 287.400 ;
        RECT 16.950 283.950 19.050 286.050 ;
        RECT 28.950 285.600 31.050 286.050 ;
        RECT 55.950 285.600 58.050 286.050 ;
        RECT 28.950 284.400 58.050 285.600 ;
        RECT 28.950 283.950 31.050 284.400 ;
        RECT 55.950 283.950 58.050 284.400 ;
        RECT 127.950 283.950 130.050 286.050 ;
        RECT 262.950 285.600 265.050 286.050 ;
        RECT 307.950 285.600 310.050 286.050 ;
        RECT 262.950 284.400 310.050 285.600 ;
        RECT 262.950 283.950 265.050 284.400 ;
        RECT 307.950 283.950 310.050 284.400 ;
        RECT 334.950 285.600 337.050 286.050 ;
        RECT 358.950 285.600 361.050 286.050 ;
        RECT 334.950 284.400 361.050 285.600 ;
        RECT 334.950 283.950 337.050 284.400 ;
        RECT 358.950 283.950 361.050 284.400 ;
        RECT 430.950 285.600 433.050 286.050 ;
        RECT 436.950 285.600 439.050 286.050 ;
        RECT 445.800 285.600 447.900 285.750 ;
        RECT 430.950 284.400 447.900 285.600 ;
        RECT 430.950 283.950 433.050 284.400 ;
        RECT 436.950 283.950 439.050 284.400 ;
        RECT 445.800 283.650 447.900 284.400 ;
        RECT 448.950 285.600 451.050 286.050 ;
        RECT 493.950 285.600 496.050 286.050 ;
        RECT 448.950 284.400 496.050 285.600 ;
        RECT 448.950 283.950 451.050 284.400 ;
        RECT 493.950 283.950 496.050 284.400 ;
        RECT 649.950 285.600 652.050 286.050 ;
        RECT 655.950 285.600 658.050 286.050 ;
        RECT 649.950 284.400 658.050 285.600 ;
        RECT 659.400 285.600 660.600 293.100 ;
        RECT 665.400 288.600 666.600 293.100 ;
        RECT 688.950 292.950 691.050 293.400 ;
        RECT 697.950 292.950 700.050 293.400 ;
        RECT 703.950 293.100 706.050 295.200 ;
        RECT 718.950 294.600 721.050 295.200 ;
        RECT 718.950 293.400 732.600 294.600 ;
        RECT 718.950 293.100 721.050 293.400 ;
        RECT 682.950 288.600 685.050 288.900 ;
        RECT 665.400 287.400 685.050 288.600 ;
        RECT 704.400 288.600 705.600 293.100 ;
        RECT 731.400 291.600 732.600 293.400 ;
        RECT 739.950 293.100 742.050 295.200 ;
        RECT 740.400 291.600 741.600 293.100 ;
        RECT 760.950 291.600 763.050 295.050 ;
        RECT 778.950 294.600 781.050 295.200 ;
        RECT 731.400 290.400 741.600 291.600 ;
        RECT 709.950 288.600 712.050 289.050 ;
        RECT 704.400 287.400 712.050 288.600 ;
        RECT 682.950 286.800 685.050 287.400 ;
        RECT 709.950 286.950 712.050 287.400 ;
        RECT 721.950 288.600 724.050 288.900 ;
        RECT 721.950 288.000 726.600 288.600 ;
        RECT 721.950 287.400 727.050 288.000 ;
        RECT 721.950 286.800 724.050 287.400 ;
        RECT 664.950 285.600 667.050 286.050 ;
        RECT 659.400 284.400 667.050 285.600 ;
        RECT 649.950 283.950 652.050 284.400 ;
        RECT 655.950 283.950 658.050 284.400 ;
        RECT 664.950 283.950 667.050 284.400 ;
        RECT 724.950 283.950 727.050 287.400 ;
        RECT 740.400 286.050 741.600 290.400 ;
        RECT 755.400 291.000 763.050 291.600 ;
        RECT 773.400 293.400 781.050 294.600 ;
        RECT 755.400 290.400 762.600 291.000 ;
        RECT 742.950 288.600 745.050 289.050 ;
        RECT 755.400 288.600 756.600 290.400 ;
        RECT 742.950 287.400 756.600 288.600 ;
        RECT 766.950 288.600 769.050 288.900 ;
        RECT 773.400 288.600 774.600 293.400 ;
        RECT 778.950 293.100 781.050 293.400 ;
        RECT 793.950 293.100 796.050 295.200 ;
        RECT 799.950 293.100 802.050 295.200 ;
        RECT 766.950 287.400 774.600 288.600 ;
        RECT 742.950 286.950 745.050 287.400 ;
        RECT 766.950 286.800 769.050 287.400 ;
        RECT 794.400 286.050 795.600 293.100 ;
        RECT 739.950 283.950 742.050 286.050 ;
        RECT 757.950 285.600 760.050 286.050 ;
        RECT 763.950 285.600 766.050 286.050 ;
        RECT 757.950 284.400 766.050 285.600 ;
        RECT 757.950 283.950 760.050 284.400 ;
        RECT 763.950 283.950 766.050 284.400 ;
        RECT 790.950 284.400 795.600 286.050 ;
        RECT 800.400 285.600 801.600 293.100 ;
        RECT 814.950 291.600 817.050 295.050 ;
        RECT 823.950 294.600 826.050 295.200 ;
        RECT 832.950 294.600 835.050 295.050 ;
        RECT 823.950 293.400 835.050 294.600 ;
        RECT 823.950 293.100 826.050 293.400 ;
        RECT 832.950 292.950 835.050 293.400 ;
        RECT 847.950 294.750 850.050 295.200 ;
        RECT 859.950 294.750 862.050 295.200 ;
        RECT 847.950 293.550 862.050 294.750 ;
        RECT 847.950 293.100 850.050 293.550 ;
        RECT 859.950 293.100 862.050 293.550 ;
        RECT 880.950 294.600 883.050 295.050 ;
        RECT 886.950 294.600 889.050 295.050 ;
        RECT 880.950 293.400 889.050 294.600 ;
        RECT 880.950 292.950 883.050 293.400 ;
        RECT 886.950 292.950 889.050 293.400 ;
        RECT 838.950 291.600 841.050 292.050 ;
        RECT 814.950 291.000 841.050 291.600 ;
        RECT 815.400 290.400 841.050 291.000 ;
        RECT 838.950 289.950 841.050 290.400 ;
        RECT 802.950 288.600 805.050 288.900 ;
        RECT 811.800 288.600 813.900 289.050 ;
        RECT 802.950 287.400 813.900 288.600 ;
        RECT 802.950 286.800 805.050 287.400 ;
        RECT 811.800 286.950 813.900 287.400 ;
        RECT 814.950 288.450 817.050 288.900 ;
        RECT 820.950 288.450 823.050 288.900 ;
        RECT 814.950 287.250 823.050 288.450 ;
        RECT 814.950 286.800 817.050 287.250 ;
        RECT 820.950 286.800 823.050 287.250 ;
        RECT 826.950 288.450 829.050 288.900 ;
        RECT 835.950 288.450 838.050 288.900 ;
        RECT 826.950 287.250 838.050 288.450 ;
        RECT 826.950 286.800 829.050 287.250 ;
        RECT 835.950 286.800 838.050 287.250 ;
        RECT 841.950 288.600 844.050 289.050 ;
        RECT 850.950 288.600 853.050 288.900 ;
        RECT 841.950 287.400 853.050 288.600 ;
        RECT 841.950 286.950 844.050 287.400 ;
        RECT 850.950 286.800 853.050 287.400 ;
        RECT 862.950 288.600 865.050 289.050 ;
        RECT 889.950 288.600 892.050 288.900 ;
        RECT 862.950 288.450 892.050 288.600 ;
        RECT 910.950 288.450 913.050 288.900 ;
        RECT 862.950 287.400 913.050 288.450 ;
        RECT 862.950 286.950 865.050 287.400 ;
        RECT 889.950 287.250 913.050 287.400 ;
        RECT 889.950 286.800 892.050 287.250 ;
        RECT 910.950 286.800 913.050 287.250 ;
        RECT 817.950 285.600 820.050 286.050 ;
        RECT 800.400 284.400 820.050 285.600 ;
        RECT 790.950 283.950 795.000 284.400 ;
        RECT 817.950 283.950 820.050 284.400 ;
        RECT 868.950 285.600 871.050 286.050 ;
        RECT 880.950 285.600 883.050 286.050 ;
        RECT 868.950 284.400 883.050 285.600 ;
        RECT 868.950 283.950 871.050 284.400 ;
        RECT 880.950 283.950 883.050 284.400 ;
        RECT 82.950 282.600 85.050 283.050 ;
        RECT 59.400 281.400 85.050 282.600 ;
        RECT 4.950 279.600 7.050 280.050 ;
        RECT 13.950 279.600 16.050 280.050 ;
        RECT 4.950 278.400 16.050 279.600 ;
        RECT 4.950 277.950 7.050 278.400 ;
        RECT 13.950 277.950 16.050 278.400 ;
        RECT 19.950 279.600 22.050 280.050 ;
        RECT 49.950 279.600 52.050 280.050 ;
        RECT 59.400 279.600 60.600 281.400 ;
        RECT 82.950 280.950 85.050 281.400 ;
        RECT 115.950 282.600 118.050 283.050 ;
        RECT 124.950 282.600 127.050 283.050 ;
        RECT 115.950 281.400 127.050 282.600 ;
        RECT 115.950 280.950 118.050 281.400 ;
        RECT 124.950 280.950 127.050 281.400 ;
        RECT 160.950 282.600 163.050 283.050 ;
        RECT 169.950 282.600 172.050 283.050 ;
        RECT 160.950 281.400 172.050 282.600 ;
        RECT 160.950 280.950 163.050 281.400 ;
        RECT 169.950 280.950 172.050 281.400 ;
        RECT 196.950 282.600 199.050 283.050 ;
        RECT 205.950 282.600 208.050 283.050 ;
        RECT 196.950 281.400 208.050 282.600 ;
        RECT 196.950 280.950 199.050 281.400 ;
        RECT 205.950 280.950 208.050 281.400 ;
        RECT 229.950 282.600 232.050 283.050 ;
        RECT 253.950 282.600 256.050 283.050 ;
        RECT 229.950 281.400 256.050 282.600 ;
        RECT 229.950 280.950 232.050 281.400 ;
        RECT 253.950 280.950 256.050 281.400 ;
        RECT 295.950 282.600 298.050 283.050 ;
        RECT 304.950 282.600 307.050 283.050 ;
        RECT 466.950 282.600 469.050 283.050 ;
        RECT 295.950 281.400 307.050 282.600 ;
        RECT 295.950 280.950 298.050 281.400 ;
        RECT 304.950 280.950 307.050 281.400 ;
        RECT 383.400 281.400 469.050 282.600 ;
        RECT 383.400 280.050 384.600 281.400 ;
        RECT 466.950 280.950 469.050 281.400 ;
        RECT 472.950 282.600 475.050 283.050 ;
        RECT 529.950 282.600 532.050 283.050 ;
        RECT 565.950 282.600 568.050 283.050 ;
        RECT 472.950 281.400 568.050 282.600 ;
        RECT 472.950 280.950 475.050 281.400 ;
        RECT 529.950 280.950 532.050 281.400 ;
        RECT 565.950 280.950 568.050 281.400 ;
        RECT 583.950 282.600 586.050 283.050 ;
        RECT 595.950 282.600 598.050 283.050 ;
        RECT 631.950 282.600 634.050 283.050 ;
        RECT 643.950 282.600 646.050 283.050 ;
        RECT 676.950 282.600 679.050 283.050 ;
        RECT 583.950 281.400 679.050 282.600 ;
        RECT 583.950 280.950 586.050 281.400 ;
        RECT 595.950 280.950 598.050 281.400 ;
        RECT 631.950 280.950 634.050 281.400 ;
        RECT 643.950 280.950 646.050 281.400 ;
        RECT 676.950 280.950 679.050 281.400 ;
        RECT 682.950 282.600 685.050 283.050 ;
        RECT 694.950 282.600 697.050 283.050 ;
        RECT 682.950 281.400 697.050 282.600 ;
        RECT 682.950 280.950 685.050 281.400 ;
        RECT 694.950 280.950 697.050 281.400 ;
        RECT 820.950 282.600 823.050 283.050 ;
        RECT 838.800 282.600 840.900 283.050 ;
        RECT 820.950 281.400 840.900 282.600 ;
        RECT 820.950 280.950 823.050 281.400 ;
        RECT 838.800 280.950 840.900 281.400 ;
        RECT 841.950 282.600 844.050 282.900 ;
        RECT 856.950 282.600 859.050 283.050 ;
        RECT 841.950 281.400 859.050 282.600 ;
        RECT 841.950 280.800 844.050 281.400 ;
        RECT 856.950 280.950 859.050 281.400 ;
        RECT 877.950 282.600 880.050 283.050 ;
        RECT 895.950 282.600 898.050 283.050 ;
        RECT 877.950 281.400 898.050 282.600 ;
        RECT 877.950 280.950 880.050 281.400 ;
        RECT 895.950 280.950 898.050 281.400 ;
        RECT 19.950 278.400 60.600 279.600 ;
        RECT 256.950 279.600 259.050 280.050 ;
        RECT 265.800 279.600 267.900 280.050 ;
        RECT 256.950 278.400 267.900 279.600 ;
        RECT 19.950 277.950 22.050 278.400 ;
        RECT 49.950 277.950 52.050 278.400 ;
        RECT 256.950 277.950 259.050 278.400 ;
        RECT 265.800 277.950 267.900 278.400 ;
        RECT 268.950 279.600 271.050 280.050 ;
        RECT 313.950 279.600 316.050 280.050 ;
        RECT 268.950 278.400 316.050 279.600 ;
        RECT 268.950 277.950 271.050 278.400 ;
        RECT 313.950 277.950 316.050 278.400 ;
        RECT 331.950 279.600 334.050 280.050 ;
        RECT 349.950 279.600 352.050 280.050 ;
        RECT 331.950 278.400 352.050 279.600 ;
        RECT 331.950 277.950 334.050 278.400 ;
        RECT 349.950 277.950 352.050 278.400 ;
        RECT 367.950 279.600 370.050 280.050 ;
        RECT 382.950 279.600 385.050 280.050 ;
        RECT 367.950 278.400 385.050 279.600 ;
        RECT 367.950 277.950 370.050 278.400 ;
        RECT 382.950 277.950 385.050 278.400 ;
        RECT 424.950 279.600 427.050 280.050 ;
        RECT 454.950 279.600 457.050 280.050 ;
        RECT 424.950 278.400 457.050 279.600 ;
        RECT 424.950 277.950 427.050 278.400 ;
        RECT 454.950 277.950 457.050 278.400 ;
        RECT 493.950 279.600 496.050 280.050 ;
        RECT 535.950 279.600 538.050 280.050 ;
        RECT 493.950 278.400 538.050 279.600 ;
        RECT 493.950 277.950 496.050 278.400 ;
        RECT 535.950 277.950 538.050 278.400 ;
        RECT 571.950 279.600 574.050 280.050 ;
        RECT 595.950 279.600 598.050 279.900 ;
        RECT 571.950 278.400 598.050 279.600 ;
        RECT 571.950 277.950 574.050 278.400 ;
        RECT 595.950 277.800 598.050 278.400 ;
        RECT 607.950 279.600 610.050 280.050 ;
        RECT 640.950 279.600 643.050 280.050 ;
        RECT 607.950 278.400 643.050 279.600 ;
        RECT 607.950 277.950 610.050 278.400 ;
        RECT 640.950 277.950 643.050 278.400 ;
        RECT 661.950 279.600 664.050 280.050 ;
        RECT 670.950 279.600 673.050 280.050 ;
        RECT 661.950 278.400 673.050 279.600 ;
        RECT 661.950 277.950 664.050 278.400 ;
        RECT 670.950 277.950 673.050 278.400 ;
        RECT 691.950 279.600 694.050 280.050 ;
        RECT 775.950 279.600 778.050 280.050 ;
        RECT 691.950 278.400 778.050 279.600 ;
        RECT 691.950 277.950 694.050 278.400 ;
        RECT 775.950 277.950 778.050 278.400 ;
        RECT 817.950 279.600 820.050 280.050 ;
        RECT 859.950 279.600 862.050 280.050 ;
        RECT 817.950 278.400 862.050 279.600 ;
        RECT 817.950 277.950 820.050 278.400 ;
        RECT 859.950 277.950 862.050 278.400 ;
        RECT 16.950 276.600 19.050 277.050 ;
        RECT 40.950 276.600 43.050 277.050 ;
        RECT 64.950 276.600 67.050 277.050 ;
        RECT 106.950 276.600 109.050 277.050 ;
        RECT 16.950 275.400 109.050 276.600 ;
        RECT 16.950 274.950 19.050 275.400 ;
        RECT 40.950 274.950 43.050 275.400 ;
        RECT 64.950 274.950 67.050 275.400 ;
        RECT 106.950 274.950 109.050 275.400 ;
        RECT 316.950 276.600 319.050 277.050 ;
        RECT 328.950 276.600 331.050 277.050 ;
        RECT 355.950 276.600 358.050 277.050 ;
        RECT 406.950 276.600 409.050 277.050 ;
        RECT 316.950 275.400 409.050 276.600 ;
        RECT 316.950 274.950 319.050 275.400 ;
        RECT 328.950 274.950 331.050 275.400 ;
        RECT 355.950 274.950 358.050 275.400 ;
        RECT 406.950 274.950 409.050 275.400 ;
        RECT 436.950 276.600 439.050 277.050 ;
        RECT 451.950 276.600 454.050 277.050 ;
        RECT 436.950 275.400 454.050 276.600 ;
        RECT 436.950 274.950 439.050 275.400 ;
        RECT 451.950 274.950 454.050 275.400 ;
        RECT 556.950 276.600 559.050 277.050 ;
        RECT 607.950 276.600 610.050 276.900 ;
        RECT 556.950 275.400 610.050 276.600 ;
        RECT 556.950 274.950 559.050 275.400 ;
        RECT 607.950 274.800 610.050 275.400 ;
        RECT 715.950 276.600 718.050 277.050 ;
        RECT 760.950 276.600 763.050 277.050 ;
        RECT 715.950 275.400 763.050 276.600 ;
        RECT 715.950 274.950 718.050 275.400 ;
        RECT 760.950 274.950 763.050 275.400 ;
        RECT 778.950 276.600 781.050 277.050 ;
        RECT 805.950 276.600 808.050 277.050 ;
        RECT 778.950 275.400 808.050 276.600 ;
        RECT 778.950 274.950 781.050 275.400 ;
        RECT 805.950 274.950 808.050 275.400 ;
        RECT 844.950 276.600 847.050 277.050 ;
        RECT 853.950 276.600 856.050 277.050 ;
        RECT 844.950 275.400 856.050 276.600 ;
        RECT 844.950 274.950 847.050 275.400 ;
        RECT 853.950 274.950 856.050 275.400 ;
        RECT 886.950 276.600 889.050 277.050 ;
        RECT 892.950 276.600 895.050 277.050 ;
        RECT 886.950 275.400 895.050 276.600 ;
        RECT 886.950 274.950 889.050 275.400 ;
        RECT 892.950 274.950 895.050 275.400 ;
        RECT 127.950 273.600 130.050 274.050 ;
        RECT 160.950 273.600 163.050 274.050 ;
        RECT 187.950 273.600 190.050 274.050 ;
        RECT 232.950 273.600 235.050 274.050 ;
        RECT 127.950 272.400 235.050 273.600 ;
        RECT 127.950 271.950 130.050 272.400 ;
        RECT 160.950 271.950 163.050 272.400 ;
        RECT 187.950 271.950 190.050 272.400 ;
        RECT 232.950 271.950 235.050 272.400 ;
        RECT 238.950 273.600 241.050 274.050 ;
        RECT 247.950 273.600 250.050 274.050 ;
        RECT 238.950 272.400 250.050 273.600 ;
        RECT 238.950 271.950 241.050 272.400 ;
        RECT 247.950 271.950 250.050 272.400 ;
        RECT 253.950 273.600 256.050 274.050 ;
        RECT 271.950 273.600 274.050 274.050 ;
        RECT 253.950 272.400 274.050 273.600 ;
        RECT 253.950 271.950 256.050 272.400 ;
        RECT 271.950 271.950 274.050 272.400 ;
        RECT 289.950 273.600 292.050 274.050 ;
        RECT 298.950 273.600 301.050 274.050 ;
        RECT 358.800 273.600 360.900 274.050 ;
        RECT 289.950 272.400 360.900 273.600 ;
        RECT 289.950 271.950 292.050 272.400 ;
        RECT 298.950 271.950 301.050 272.400 ;
        RECT 358.800 271.950 360.900 272.400 ;
        RECT 361.950 273.600 364.050 274.050 ;
        RECT 412.950 273.600 415.050 274.050 ;
        RECT 361.950 272.400 415.050 273.600 ;
        RECT 361.950 271.950 364.050 272.400 ;
        RECT 412.950 271.950 415.050 272.400 ;
        RECT 508.950 273.600 511.050 274.050 ;
        RECT 646.950 273.600 649.050 274.050 ;
        RECT 670.950 273.600 673.050 274.050 ;
        RECT 694.950 273.600 697.050 274.050 ;
        RECT 508.950 272.400 697.050 273.600 ;
        RECT 508.950 271.950 511.050 272.400 ;
        RECT 646.950 271.950 649.050 272.400 ;
        RECT 670.950 271.950 673.050 272.400 ;
        RECT 694.950 271.950 697.050 272.400 ;
        RECT 730.950 273.600 733.050 274.050 ;
        RECT 745.950 273.600 748.050 274.050 ;
        RECT 730.950 272.400 748.050 273.600 ;
        RECT 730.950 271.950 733.050 272.400 ;
        RECT 745.950 271.950 748.050 272.400 ;
        RECT 751.950 273.600 754.050 274.050 ;
        RECT 751.950 272.400 765.600 273.600 ;
        RECT 751.950 271.950 754.050 272.400 ;
        RECT 764.400 271.050 765.600 272.400 ;
        RECT 871.950 271.950 874.050 274.050 ;
        RECT 877.950 271.950 880.050 274.050 ;
        RECT 883.950 273.600 886.050 274.050 ;
        RECT 895.950 273.600 898.050 274.050 ;
        RECT 883.950 272.400 898.050 273.600 ;
        RECT 883.950 271.950 886.050 272.400 ;
        RECT 895.950 271.950 898.050 272.400 ;
        RECT 7.950 270.600 10.050 271.050 ;
        RECT 34.950 270.600 37.050 271.050 ;
        RECT 7.950 269.400 37.050 270.600 ;
        RECT 7.950 268.950 10.050 269.400 ;
        RECT 34.950 268.950 37.050 269.400 ;
        RECT 106.950 270.600 109.050 271.050 ;
        RECT 136.950 270.600 139.050 271.050 ;
        RECT 142.950 270.600 145.050 271.050 ;
        RECT 106.950 269.400 145.050 270.600 ;
        RECT 106.950 268.950 109.050 269.400 ;
        RECT 136.950 268.950 139.050 269.400 ;
        RECT 142.950 268.950 145.050 269.400 ;
        RECT 208.950 270.600 211.050 271.050 ;
        RECT 235.950 270.600 238.050 271.050 ;
        RECT 250.950 270.600 253.050 271.050 ;
        RECT 208.950 269.400 253.050 270.600 ;
        RECT 208.950 268.950 211.050 269.400 ;
        RECT 235.950 268.950 238.050 269.400 ;
        RECT 250.950 268.950 253.050 269.400 ;
        RECT 373.950 270.600 376.050 271.050 ;
        RECT 394.950 270.600 397.050 271.050 ;
        RECT 373.950 269.400 397.050 270.600 ;
        RECT 373.950 268.950 376.050 269.400 ;
        RECT 394.950 268.950 397.050 269.400 ;
        RECT 403.950 270.600 406.050 271.050 ;
        RECT 418.950 270.600 421.050 271.050 ;
        RECT 460.950 270.600 463.050 271.050 ;
        RECT 499.950 270.600 502.050 271.050 ;
        RECT 403.950 269.400 502.050 270.600 ;
        RECT 403.950 268.950 406.050 269.400 ;
        RECT 418.950 268.950 421.050 269.400 ;
        RECT 460.950 268.950 463.050 269.400 ;
        RECT 499.950 268.950 502.050 269.400 ;
        RECT 547.950 270.600 550.050 271.050 ;
        RECT 568.950 270.600 571.050 271.050 ;
        RECT 547.950 269.400 571.050 270.600 ;
        RECT 547.950 268.950 550.050 269.400 ;
        RECT 568.950 268.950 571.050 269.400 ;
        RECT 598.950 270.600 601.050 271.050 ;
        RECT 610.950 270.600 613.050 271.050 ;
        RECT 598.950 269.400 613.050 270.600 ;
        RECT 764.400 269.400 769.050 271.050 ;
        RECT 598.950 268.950 601.050 269.400 ;
        RECT 610.950 268.950 613.050 269.400 ;
        RECT 765.000 268.950 769.050 269.400 ;
        RECT 796.950 270.600 799.050 271.050 ;
        RECT 844.950 270.600 847.050 271.050 ;
        RECT 796.950 269.400 847.050 270.600 ;
        RECT 796.950 268.950 799.050 269.400 ;
        RECT 844.950 268.950 847.050 269.400 ;
        RECT 37.950 267.600 40.050 268.050 ;
        RECT 172.950 267.600 175.050 268.050 ;
        RECT 181.950 267.600 184.050 268.050 ;
        RECT 37.950 266.400 60.600 267.600 ;
        RECT 37.950 265.950 40.050 266.400 ;
        RECT 46.950 264.600 49.050 265.050 ;
        RECT 59.400 264.600 60.600 266.400 ;
        RECT 172.950 266.400 184.050 267.600 ;
        RECT 172.950 265.950 175.050 266.400 ;
        RECT 181.950 265.950 184.050 266.400 ;
        RECT 217.950 267.600 220.050 268.050 ;
        RECT 223.950 267.600 226.050 268.050 ;
        RECT 217.950 266.400 226.050 267.600 ;
        RECT 217.950 265.950 220.050 266.400 ;
        RECT 223.950 265.950 226.050 266.400 ;
        RECT 316.950 267.600 319.050 268.050 ;
        RECT 325.950 267.600 328.050 268.050 ;
        RECT 316.950 266.400 328.050 267.600 ;
        RECT 316.950 265.950 319.050 266.400 ;
        RECT 325.950 265.950 328.050 266.400 ;
        RECT 346.950 267.600 349.050 268.050 ;
        RECT 361.950 267.600 364.050 268.050 ;
        RECT 346.950 266.400 364.050 267.600 ;
        RECT 346.950 265.950 349.050 266.400 ;
        RECT 361.950 265.950 364.050 266.400 ;
        RECT 406.950 267.600 409.050 268.050 ;
        RECT 427.950 267.600 430.050 268.050 ;
        RECT 448.950 267.600 451.050 268.050 ;
        RECT 406.950 266.400 451.050 267.600 ;
        RECT 406.950 265.950 409.050 266.400 ;
        RECT 427.950 265.950 430.050 266.400 ;
        RECT 448.950 265.950 451.050 266.400 ;
        RECT 466.950 267.600 469.050 268.050 ;
        RECT 487.950 267.600 490.050 268.050 ;
        RECT 466.950 266.400 490.050 267.600 ;
        RECT 466.950 265.950 469.050 266.400 ;
        RECT 487.950 265.950 490.050 266.400 ;
        RECT 541.950 267.600 544.050 268.050 ;
        RECT 577.950 267.600 580.050 268.050 ;
        RECT 619.950 267.600 622.050 268.050 ;
        RECT 541.950 266.400 622.050 267.600 ;
        RECT 541.950 265.950 544.050 266.400 ;
        RECT 577.950 265.950 580.050 266.400 ;
        RECT 619.950 265.950 622.050 266.400 ;
        RECT 703.950 267.600 706.050 268.050 ;
        RECT 745.950 267.600 748.050 268.050 ;
        RECT 783.000 267.600 787.050 268.050 ;
        RECT 703.950 266.400 748.050 267.600 ;
        RECT 703.950 265.950 706.050 266.400 ;
        RECT 745.950 265.950 748.050 266.400 ;
        RECT 782.400 265.950 787.050 267.600 ;
        RECT 823.950 267.600 826.050 268.050 ;
        RECT 841.950 267.600 844.050 268.050 ;
        RECT 823.950 266.400 844.050 267.600 ;
        RECT 823.950 265.950 826.050 266.400 ;
        RECT 841.950 265.950 844.050 266.400 ;
        RECT 73.950 264.600 76.050 265.050 ;
        RECT 82.950 264.600 85.050 265.050 ;
        RECT 46.950 263.400 57.600 264.600 ;
        RECT 59.400 263.400 66.600 264.600 ;
        RECT 46.950 262.950 49.050 263.400 ;
        RECT 7.950 261.600 10.050 262.050 ;
        RECT 16.950 261.600 19.050 262.200 ;
        RECT 7.950 260.400 19.050 261.600 ;
        RECT 7.950 259.950 10.050 260.400 ;
        RECT 16.950 260.100 19.050 260.400 ;
        RECT 22.950 261.600 25.050 262.200 ;
        RECT 31.950 261.600 34.050 262.050 ;
        RECT 43.950 261.600 46.050 262.200 ;
        RECT 22.950 260.400 46.050 261.600 ;
        RECT 56.400 261.600 57.600 263.400 ;
        RECT 56.400 260.400 63.600 261.600 ;
        RECT 22.950 260.100 25.050 260.400 ;
        RECT 31.950 259.950 34.050 260.400 ;
        RECT 43.950 260.100 46.050 260.400 ;
        RECT 19.950 255.450 22.050 255.900 ;
        RECT 28.950 255.600 31.050 255.900 ;
        RECT 40.950 255.600 43.050 255.900 ;
        RECT 28.950 255.450 43.050 255.600 ;
        RECT 19.950 254.400 43.050 255.450 ;
        RECT 44.400 255.600 45.600 260.100 ;
        RECT 55.950 255.600 58.050 256.050 ;
        RECT 62.400 255.900 63.600 260.400 ;
        RECT 44.400 254.400 58.050 255.600 ;
        RECT 19.950 254.250 31.050 254.400 ;
        RECT 19.950 253.800 22.050 254.250 ;
        RECT 28.950 253.800 31.050 254.250 ;
        RECT 40.950 253.800 43.050 254.400 ;
        RECT 55.950 253.950 58.050 254.400 ;
        RECT 61.950 253.800 64.050 255.900 ;
        RECT 65.400 253.050 66.600 263.400 ;
        RECT 73.950 263.400 85.050 264.600 ;
        RECT 73.950 262.950 76.050 263.400 ;
        RECT 82.950 262.950 85.050 263.400 ;
        RECT 118.950 264.600 121.050 265.050 ;
        RECT 130.950 264.600 133.050 265.050 ;
        RECT 199.950 264.600 202.050 265.050 ;
        RECT 214.950 264.600 217.050 265.050 ;
        RECT 118.950 263.400 217.050 264.600 ;
        RECT 118.950 262.950 121.050 263.400 ;
        RECT 130.950 262.950 133.050 263.400 ;
        RECT 199.950 262.950 202.050 263.400 ;
        RECT 214.950 262.950 217.050 263.400 ;
        RECT 241.950 264.600 244.050 264.900 ;
        RECT 253.950 264.600 256.050 265.050 ;
        RECT 274.950 264.600 277.050 265.050 ;
        RECT 241.950 263.400 277.050 264.600 ;
        RECT 241.950 262.800 244.050 263.400 ;
        RECT 253.950 262.950 256.050 263.400 ;
        RECT 274.950 262.950 277.050 263.400 ;
        RECT 292.950 264.600 295.050 265.050 ;
        RECT 301.950 264.600 304.050 265.200 ;
        RECT 292.950 263.400 304.050 264.600 ;
        RECT 292.950 262.950 295.050 263.400 ;
        RECT 301.950 263.100 304.050 263.400 ;
        RECT 358.950 264.600 361.050 265.050 ;
        RECT 394.950 264.600 397.050 265.050 ;
        RECT 358.950 263.400 397.050 264.600 ;
        RECT 358.950 262.950 361.050 263.400 ;
        RECT 394.950 262.950 397.050 263.400 ;
        RECT 463.950 264.600 466.050 265.050 ;
        RECT 463.950 263.400 474.600 264.600 ;
        RECT 463.950 262.950 466.050 263.400 ;
        RECT 85.950 260.100 88.050 262.200 ;
        RECT 94.950 261.600 99.000 262.050 ;
        RECT 100.950 261.750 103.050 262.200 ;
        RECT 112.950 261.750 115.050 262.200 ;
        RECT 86.400 256.050 87.600 260.100 ;
        RECT 94.950 259.950 99.600 261.600 ;
        RECT 100.950 260.550 115.050 261.750 ;
        RECT 100.950 260.100 103.050 260.550 ;
        RECT 112.950 260.100 115.050 260.550 ;
        RECT 121.950 261.600 124.050 262.200 ;
        RECT 139.950 261.600 142.050 262.050 ;
        RECT 121.950 260.400 142.050 261.600 ;
        RECT 121.950 260.100 124.050 260.400 ;
        RECT 139.950 259.950 142.050 260.400 ;
        RECT 148.950 260.100 151.050 262.200 ;
        RECT 193.950 261.600 196.050 262.050 ;
        RECT 223.950 261.600 226.050 262.200 ;
        RECT 234.000 261.600 238.050 262.050 ;
        RECT 179.400 260.400 196.050 261.600 ;
        RECT 67.950 255.450 70.050 255.900 ;
        RECT 73.950 255.450 76.050 255.900 ;
        RECT 67.950 254.250 76.050 255.450 ;
        RECT 86.400 254.400 91.050 256.050 ;
        RECT 98.400 255.900 99.600 259.950 ;
        RECT 67.950 253.800 70.050 254.250 ;
        RECT 73.950 253.800 76.050 254.250 ;
        RECT 87.000 253.950 91.050 254.400 ;
        RECT 97.950 253.800 100.050 255.900 ;
        RECT 109.950 255.600 112.050 255.900 ;
        RECT 130.950 255.600 133.050 255.900 ;
        RECT 109.950 255.450 133.050 255.600 ;
        RECT 145.950 255.450 148.050 255.900 ;
        RECT 109.950 254.400 148.050 255.450 ;
        RECT 149.400 255.600 150.600 260.100 ;
        RECT 179.400 256.050 180.600 260.400 ;
        RECT 193.950 259.950 196.050 260.400 ;
        RECT 218.400 260.400 226.050 261.600 ;
        RECT 218.400 259.050 219.600 260.400 ;
        RECT 223.950 260.100 226.050 260.400 ;
        RECT 199.950 258.600 202.050 259.050 ;
        RECT 185.400 257.400 202.050 258.600 ;
        RECT 163.950 255.600 166.050 255.900 ;
        RECT 149.400 254.400 166.050 255.600 ;
        RECT 109.950 253.800 112.050 254.400 ;
        RECT 130.950 254.250 148.050 254.400 ;
        RECT 130.950 253.800 133.050 254.250 ;
        RECT 145.950 253.800 148.050 254.250 ;
        RECT 163.950 253.800 166.050 254.400 ;
        RECT 178.950 253.950 181.050 256.050 ;
        RECT 185.400 255.900 186.600 257.400 ;
        RECT 199.950 256.950 202.050 257.400 ;
        RECT 214.950 257.400 219.600 259.050 ;
        RECT 233.400 259.950 238.050 261.600 ;
        RECT 244.950 261.600 247.050 262.050 ;
        RECT 301.950 261.600 304.050 262.050 ;
        RECT 244.950 260.400 252.600 261.600 ;
        RECT 263.400 261.000 304.050 261.600 ;
        RECT 244.950 259.950 247.050 260.400 ;
        RECT 214.950 256.950 219.000 257.400 ;
        RECT 233.400 255.900 234.600 259.950 ;
        RECT 251.400 255.900 252.600 260.400 ;
        RECT 262.950 260.400 304.050 261.000 ;
        RECT 262.950 256.800 265.050 260.400 ;
        RECT 301.950 259.950 304.050 260.400 ;
        RECT 307.950 260.100 310.050 262.200 ;
        RECT 313.950 261.750 316.050 262.200 ;
        RECT 319.950 261.750 322.050 262.200 ;
        RECT 313.950 260.550 322.050 261.750 ;
        RECT 331.950 261.600 334.050 262.050 ;
        RECT 343.950 261.600 346.050 262.200 ;
        RECT 313.950 260.100 316.050 260.550 ;
        RECT 319.950 260.100 322.050 260.550 ;
        RECT 326.400 260.400 334.050 261.600 ;
        RECT 184.950 253.800 187.050 255.900 ;
        RECT 232.950 253.800 235.050 255.900 ;
        RECT 250.950 253.800 253.050 255.900 ;
        RECT 289.950 255.450 292.050 255.900 ;
        RECT 298.950 255.450 301.050 255.900 ;
        RECT 289.950 254.250 301.050 255.450 ;
        RECT 308.400 255.600 309.600 260.100 ;
        RECT 326.400 258.600 327.600 260.400 ;
        RECT 331.950 259.950 334.050 260.400 ;
        RECT 335.400 260.400 346.050 261.600 ;
        RECT 335.400 258.600 336.600 260.400 ;
        RECT 343.950 260.100 346.050 260.400 ;
        RECT 382.950 260.100 385.050 262.200 ;
        RECT 397.950 261.600 400.050 262.050 ;
        RECT 403.950 261.600 406.050 262.200 ;
        RECT 439.950 261.600 442.050 262.050 ;
        RECT 397.950 260.400 442.050 261.600 ;
        RECT 383.400 258.600 384.600 260.100 ;
        RECT 397.950 259.950 400.050 260.400 ;
        RECT 403.950 260.100 406.050 260.400 ;
        RECT 439.950 259.950 442.050 260.400 ;
        RECT 323.400 257.400 327.600 258.600 ;
        RECT 329.400 257.400 336.600 258.600 ;
        RECT 374.400 257.400 384.600 258.600 ;
        RECT 316.950 255.600 319.050 256.050 ;
        RECT 323.400 255.900 324.600 257.400 ;
        RECT 329.400 255.900 330.600 257.400 ;
        RECT 374.400 256.050 375.600 257.400 ;
        RECT 308.400 254.400 319.050 255.600 ;
        RECT 289.950 253.800 292.050 254.250 ;
        RECT 298.950 253.800 301.050 254.250 ;
        RECT 316.950 253.950 319.050 254.400 ;
        RECT 322.950 253.800 325.050 255.900 ;
        RECT 328.950 253.800 331.050 255.900 ;
        RECT 346.950 255.450 349.050 255.900 ;
        RECT 355.950 255.450 358.050 255.900 ;
        RECT 346.950 254.250 358.050 255.450 ;
        RECT 346.950 253.800 349.050 254.250 ;
        RECT 355.950 253.800 358.050 254.250 ;
        RECT 370.950 254.400 375.600 256.050 ;
        RECT 379.950 255.450 382.050 255.900 ;
        RECT 391.800 255.450 393.900 255.900 ;
        RECT 370.950 253.950 375.000 254.400 ;
        RECT 379.950 254.250 393.900 255.450 ;
        RECT 379.950 253.800 382.050 254.250 ;
        RECT 391.800 253.800 393.900 254.250 ;
        RECT 394.950 255.600 397.050 256.050 ;
        RECT 400.950 255.600 403.050 255.900 ;
        RECT 394.950 254.400 403.050 255.600 ;
        RECT 394.950 253.950 397.050 254.400 ;
        RECT 400.950 253.800 403.050 254.400 ;
        RECT 409.950 255.600 412.050 255.900 ;
        RECT 421.950 255.600 424.050 255.900 ;
        RECT 409.950 254.400 424.050 255.600 ;
        RECT 409.950 253.800 412.050 254.400 ;
        RECT 421.950 253.800 424.050 254.400 ;
        RECT 433.950 255.450 436.050 255.900 ;
        RECT 463.950 255.450 466.050 255.900 ;
        RECT 433.950 254.250 466.050 255.450 ;
        RECT 473.400 255.600 474.600 263.400 ;
        RECT 607.950 262.950 610.050 265.050 ;
        RECT 628.950 264.600 631.050 265.050 ;
        RECT 643.950 264.600 646.050 265.050 ;
        RECT 628.950 263.400 646.050 264.600 ;
        RECT 628.950 262.950 631.050 263.400 ;
        RECT 643.950 262.950 646.050 263.400 ;
        RECT 688.950 264.600 693.000 265.050 ;
        RECT 697.950 264.600 702.000 265.050 ;
        RECT 706.950 264.600 709.050 265.050 ;
        RECT 712.950 264.600 715.050 265.050 ;
        RECT 727.950 264.600 730.050 265.050 ;
        RECT 688.950 262.950 693.600 264.600 ;
        RECT 697.950 262.950 702.600 264.600 ;
        RECT 706.950 263.400 730.050 264.600 ;
        RECT 706.950 262.950 709.050 263.400 ;
        RECT 712.950 262.950 715.050 263.400 ;
        RECT 727.950 262.950 730.050 263.400 ;
        RECT 487.950 261.600 490.050 262.200 ;
        RECT 508.950 261.600 511.050 262.200 ;
        RECT 516.000 261.600 520.050 262.050 ;
        RECT 487.950 260.400 511.050 261.600 ;
        RECT 487.950 260.100 490.050 260.400 ;
        RECT 508.950 260.100 511.050 260.400 ;
        RECT 515.400 259.950 520.050 261.600 ;
        RECT 523.950 261.750 526.050 262.200 ;
        RECT 529.950 261.750 532.050 262.200 ;
        RECT 523.950 261.600 532.050 261.750 ;
        RECT 535.950 261.600 538.050 262.050 ;
        RECT 523.950 260.550 538.050 261.600 ;
        RECT 523.950 260.100 526.050 260.550 ;
        RECT 529.950 260.400 538.050 260.550 ;
        RECT 529.950 260.100 532.050 260.400 ;
        RECT 535.950 259.950 538.050 260.400 ;
        RECT 574.950 261.750 577.050 262.200 ;
        RECT 583.950 261.750 586.050 262.200 ;
        RECT 574.950 260.550 586.050 261.750 ;
        RECT 574.950 260.100 577.050 260.550 ;
        RECT 583.950 260.100 586.050 260.550 ;
        RECT 589.950 260.100 592.050 262.200 ;
        RECT 515.400 258.600 516.600 259.950 ;
        RECT 590.400 258.600 591.600 260.100 ;
        RECT 595.950 259.950 598.050 262.050 ;
        RECT 604.950 260.100 607.050 262.200 ;
        RECT 512.400 258.000 516.600 258.600 ;
        RECT 587.400 258.000 591.600 258.600 ;
        RECT 511.950 257.400 516.600 258.000 ;
        RECT 586.950 257.400 591.600 258.000 ;
        RECT 493.950 255.600 496.050 255.900 ;
        RECT 499.950 255.600 502.050 256.050 ;
        RECT 473.400 254.400 492.600 255.600 ;
        RECT 433.950 253.800 436.050 254.250 ;
        RECT 463.950 253.800 466.050 254.250 ;
        RECT 64.950 250.950 67.050 253.050 ;
        RECT 112.950 252.600 115.050 253.050 ;
        RECT 118.950 252.600 121.050 253.050 ;
        RECT 112.950 251.400 121.050 252.600 ;
        RECT 112.950 250.950 115.050 251.400 ;
        RECT 118.950 250.950 121.050 251.400 ;
        RECT 151.950 252.600 154.050 253.050 ;
        RECT 169.950 252.600 172.050 253.050 ;
        RECT 151.950 251.400 172.050 252.600 ;
        RECT 151.950 250.950 154.050 251.400 ;
        RECT 169.950 250.950 172.050 251.400 ;
        RECT 256.950 252.600 259.050 253.050 ;
        RECT 271.950 252.600 274.050 253.050 ;
        RECT 310.950 252.600 313.050 253.050 ;
        RECT 256.950 251.400 313.050 252.600 ;
        RECT 491.400 252.600 492.600 254.400 ;
        RECT 493.950 255.450 502.050 255.600 ;
        RECT 505.950 255.450 508.050 255.900 ;
        RECT 493.950 254.400 508.050 255.450 ;
        RECT 493.950 253.800 496.050 254.400 ;
        RECT 499.950 254.250 508.050 254.400 ;
        RECT 499.950 253.950 502.050 254.250 ;
        RECT 505.950 253.800 508.050 254.250 ;
        RECT 511.950 253.950 514.050 257.400 ;
        RECT 520.950 255.450 523.050 255.900 ;
        RECT 526.950 255.450 529.050 255.900 ;
        RECT 520.950 254.250 529.050 255.450 ;
        RECT 520.950 253.800 523.050 254.250 ;
        RECT 526.950 253.800 529.050 254.250 ;
        RECT 538.950 255.450 541.050 255.900 ;
        RECT 577.950 255.450 580.050 255.900 ;
        RECT 538.950 254.250 580.050 255.450 ;
        RECT 538.950 253.800 541.050 254.250 ;
        RECT 577.950 253.800 580.050 254.250 ;
        RECT 586.950 253.950 589.050 257.400 ;
        RECT 596.400 256.050 597.600 259.950 ;
        RECT 595.950 253.950 598.050 256.050 ;
        RECT 605.400 253.050 606.600 260.100 ;
        RECT 608.400 255.900 609.600 262.950 ;
        RECT 652.950 261.600 655.050 262.200 ;
        RECT 611.400 260.400 655.050 261.600 ;
        RECT 607.950 253.800 610.050 255.900 ;
        RECT 499.950 252.600 502.050 252.900 ;
        RECT 491.400 251.400 502.050 252.600 ;
        RECT 256.950 250.950 259.050 251.400 ;
        RECT 271.950 250.950 274.050 251.400 ;
        RECT 310.950 250.950 313.050 251.400 ;
        RECT 170.400 249.600 171.600 250.950 ;
        RECT 499.950 250.800 502.050 251.400 ;
        RECT 604.950 252.600 607.050 253.050 ;
        RECT 611.400 252.600 612.600 260.400 ;
        RECT 652.950 260.100 655.050 260.400 ;
        RECT 676.950 260.100 679.050 262.200 ;
        RECT 619.950 255.450 622.050 255.900 ;
        RECT 625.950 255.450 628.050 255.900 ;
        RECT 619.950 254.250 628.050 255.450 ;
        RECT 677.400 255.600 678.600 260.100 ;
        RECT 692.400 256.050 693.600 262.950 ;
        RECT 701.400 256.050 702.600 262.950 ;
        RECT 724.950 261.600 727.050 262.050 ;
        RECT 719.400 260.400 727.050 261.600 ;
        RECT 688.800 255.600 690.900 255.900 ;
        RECT 677.400 254.400 690.900 255.600 ;
        RECT 619.950 253.800 622.050 254.250 ;
        RECT 625.950 253.800 628.050 254.250 ;
        RECT 688.800 253.800 690.900 254.400 ;
        RECT 691.950 253.950 694.050 256.050 ;
        RECT 700.950 253.950 703.050 256.050 ;
        RECT 719.400 255.900 720.600 260.400 ;
        RECT 724.950 259.950 727.050 260.400 ;
        RECT 742.950 258.600 745.050 262.050 ;
        RECT 757.950 259.950 760.050 262.050 ;
        RECT 737.400 258.000 745.050 258.600 ;
        RECT 737.400 257.400 744.600 258.000 ;
        RECT 718.950 253.800 721.050 255.900 ;
        RECT 724.950 255.600 727.050 256.050 ;
        RECT 737.400 255.600 738.600 257.400 ;
        RECT 758.400 256.050 759.600 259.950 ;
        RECT 782.400 256.050 783.600 265.950 ;
        RECT 796.950 264.600 799.050 265.050 ;
        RECT 808.950 264.600 811.050 264.900 ;
        RECT 832.950 264.600 835.050 265.050 ;
        RECT 796.950 263.400 835.050 264.600 ;
        RECT 796.950 262.950 799.050 263.400 ;
        RECT 808.950 262.800 811.050 263.400 ;
        RECT 832.950 262.950 835.050 263.400 ;
        RECT 856.950 264.600 859.050 265.050 ;
        RECT 872.400 264.600 873.600 271.950 ;
        RECT 856.950 263.400 873.600 264.600 ;
        RECT 856.950 262.950 859.050 263.400 ;
        RECT 787.950 258.600 790.050 262.050 ;
        RECT 814.950 259.950 817.050 262.050 ;
        RECT 826.950 261.600 829.050 262.200 ;
        RECT 824.400 260.400 829.050 261.600 ;
        RECT 787.950 258.000 807.600 258.600 ;
        RECT 788.400 257.400 808.050 258.000 ;
        RECT 724.950 254.400 738.600 255.600 ;
        RECT 724.950 253.950 727.050 254.400 ;
        RECT 757.950 253.950 760.050 256.050 ;
        RECT 781.950 253.950 784.050 256.050 ;
        RECT 805.950 253.950 808.050 257.400 ;
        RECT 604.950 251.400 612.600 252.600 ;
        RECT 613.950 252.600 616.050 253.050 ;
        RECT 634.950 252.600 637.050 253.050 ;
        RECT 613.950 251.400 637.050 252.600 ;
        RECT 604.950 250.950 607.050 251.400 ;
        RECT 613.950 250.950 616.050 251.400 ;
        RECT 634.950 250.950 637.050 251.400 ;
        RECT 661.950 252.600 664.050 253.050 ;
        RECT 673.950 252.600 676.050 253.050 ;
        RECT 661.950 251.400 676.050 252.600 ;
        RECT 661.950 250.950 664.050 251.400 ;
        RECT 673.950 250.950 676.050 251.400 ;
        RECT 739.950 252.600 742.050 253.050 ;
        RECT 754.950 252.600 757.050 253.050 ;
        RECT 739.950 251.400 757.050 252.600 ;
        RECT 739.950 250.950 742.050 251.400 ;
        RECT 754.950 250.950 757.050 251.400 ;
        RECT 802.950 252.600 805.050 253.050 ;
        RECT 815.400 252.600 816.600 259.950 ;
        RECT 824.400 253.050 825.600 260.400 ;
        RECT 826.950 260.100 829.050 260.400 ;
        RECT 832.950 261.750 835.050 262.200 ;
        RECT 838.950 261.750 841.050 262.200 ;
        RECT 832.950 260.550 841.050 261.750 ;
        RECT 832.950 260.100 835.050 260.550 ;
        RECT 838.950 260.100 841.050 260.550 ;
        RECT 847.950 257.100 850.050 259.200 ;
        RECT 878.400 258.900 879.600 271.950 ;
        RECT 895.950 259.950 898.050 262.050 ;
        RECT 848.400 255.600 849.600 257.100 ;
        RECT 877.950 256.800 880.050 258.900 ;
        RECT 842.400 254.400 849.600 255.600 ;
        RECT 802.950 251.400 816.600 252.600 ;
        RECT 820.950 251.400 825.600 253.050 ;
        RECT 835.950 252.600 838.050 253.050 ;
        RECT 842.400 252.600 843.600 254.400 ;
        RECT 835.950 251.400 843.600 252.600 ;
        RECT 802.950 250.950 805.050 251.400 ;
        RECT 820.950 250.950 825.000 251.400 ;
        RECT 835.950 250.950 838.050 251.400 ;
        RECT 856.950 250.950 859.050 253.050 ;
        RECT 190.950 249.600 193.050 250.050 ;
        RECT 170.400 248.400 193.050 249.600 ;
        RECT 190.950 247.950 193.050 248.400 ;
        RECT 205.950 249.600 208.050 250.050 ;
        RECT 241.950 249.600 244.050 250.050 ;
        RECT 205.950 248.400 244.050 249.600 ;
        RECT 205.950 247.950 208.050 248.400 ;
        RECT 241.950 247.950 244.050 248.400 ;
        RECT 340.950 249.600 343.050 250.050 ;
        RECT 373.950 249.600 376.050 250.050 ;
        RECT 400.950 249.600 403.050 250.050 ;
        RECT 472.950 249.600 475.050 250.050 ;
        RECT 340.950 248.400 376.050 249.600 ;
        RECT 340.950 247.950 343.050 248.400 ;
        RECT 373.950 247.950 376.050 248.400 ;
        RECT 386.400 248.400 475.050 249.600 ;
        RECT 386.400 247.050 387.600 248.400 ;
        RECT 400.950 247.950 403.050 248.400 ;
        RECT 472.950 247.950 475.050 248.400 ;
        RECT 622.950 249.600 625.050 250.050 ;
        RECT 652.950 249.600 655.050 250.050 ;
        RECT 622.950 248.400 655.050 249.600 ;
        RECT 622.950 247.950 625.050 248.400 ;
        RECT 652.950 247.950 655.050 248.400 ;
        RECT 676.950 249.600 679.050 250.050 ;
        RECT 697.950 249.600 700.050 250.050 ;
        RECT 676.950 248.400 700.050 249.600 ;
        RECT 676.950 247.950 679.050 248.400 ;
        RECT 697.950 247.950 700.050 248.400 ;
        RECT 772.950 249.600 775.050 250.050 ;
        RECT 793.950 249.600 796.050 250.050 ;
        RECT 772.950 248.400 796.050 249.600 ;
        RECT 772.950 247.950 775.050 248.400 ;
        RECT 793.950 247.950 796.050 248.400 ;
        RECT 55.950 246.600 58.050 247.050 ;
        RECT 103.950 246.600 106.050 247.050 ;
        RECT 55.950 245.400 106.050 246.600 ;
        RECT 55.950 244.950 58.050 245.400 ;
        RECT 103.950 244.950 106.050 245.400 ;
        RECT 226.950 246.600 229.050 247.050 ;
        RECT 262.950 246.600 265.050 247.050 ;
        RECT 226.950 245.400 265.050 246.600 ;
        RECT 226.950 244.950 229.050 245.400 ;
        RECT 262.950 244.950 265.050 245.400 ;
        RECT 286.950 246.600 289.050 247.050 ;
        RECT 334.950 246.600 337.050 247.050 ;
        RECT 286.950 245.400 337.050 246.600 ;
        RECT 286.950 244.950 289.050 245.400 ;
        RECT 334.950 244.950 337.050 245.400 ;
        RECT 343.950 246.600 346.050 247.050 ;
        RECT 385.950 246.600 388.050 247.050 ;
        RECT 343.950 245.400 388.050 246.600 ;
        RECT 343.950 244.950 346.050 245.400 ;
        RECT 385.950 244.950 388.050 245.400 ;
        RECT 391.950 246.600 394.050 247.050 ;
        RECT 421.950 246.600 424.050 247.050 ;
        RECT 391.950 245.400 424.050 246.600 ;
        RECT 391.950 244.950 394.050 245.400 ;
        RECT 421.950 244.950 424.050 245.400 ;
        RECT 439.950 246.600 442.050 247.050 ;
        RECT 532.950 246.600 535.050 247.050 ;
        RECT 439.950 245.400 535.050 246.600 ;
        RECT 439.950 244.950 442.050 245.400 ;
        RECT 532.950 244.950 535.050 245.400 ;
        RECT 745.950 246.600 748.050 247.050 ;
        RECT 760.950 246.600 763.050 247.050 ;
        RECT 745.950 245.400 763.050 246.600 ;
        RECT 745.950 244.950 748.050 245.400 ;
        RECT 760.950 244.950 763.050 245.400 ;
        RECT 829.950 246.600 832.050 247.050 ;
        RECT 853.950 246.600 856.050 247.050 ;
        RECT 829.950 245.400 856.050 246.600 ;
        RECT 829.950 244.950 832.050 245.400 ;
        RECT 853.950 244.950 856.050 245.400 ;
        RECT 259.950 243.600 262.050 244.050 ;
        RECT 161.400 242.400 262.050 243.600 ;
        RECT 58.950 240.600 61.050 241.050 ;
        RECT 88.950 240.600 91.050 241.050 ;
        RECT 148.950 240.600 151.050 241.050 ;
        RECT 58.950 239.400 151.050 240.600 ;
        RECT 58.950 238.950 61.050 239.400 ;
        RECT 88.950 238.950 91.050 239.400 ;
        RECT 148.950 238.950 151.050 239.400 ;
        RECT 154.950 240.600 157.050 241.050 ;
        RECT 161.400 240.600 162.600 242.400 ;
        RECT 259.950 241.950 262.050 242.400 ;
        RECT 322.950 243.600 325.050 244.050 ;
        RECT 460.950 243.600 463.050 244.050 ;
        RECT 484.950 243.600 487.050 244.050 ;
        RECT 322.950 242.400 378.600 243.600 ;
        RECT 322.950 241.950 325.050 242.400 ;
        RECT 154.950 239.400 162.600 240.600 ;
        RECT 211.950 240.600 214.050 241.050 ;
        RECT 292.950 240.600 295.050 241.050 ;
        RECT 211.950 239.400 295.050 240.600 ;
        RECT 154.950 238.950 157.050 239.400 ;
        RECT 211.950 238.950 214.050 239.400 ;
        RECT 292.950 238.950 295.050 239.400 ;
        RECT 313.950 240.600 316.050 241.050 ;
        RECT 346.950 240.600 349.050 241.050 ;
        RECT 313.950 239.400 349.050 240.600 ;
        RECT 377.400 240.600 378.600 242.400 ;
        RECT 460.950 242.400 487.050 243.600 ;
        RECT 460.950 241.950 463.050 242.400 ;
        RECT 484.950 241.950 487.050 242.400 ;
        RECT 586.950 243.600 589.050 244.050 ;
        RECT 649.950 243.600 652.050 244.050 ;
        RECT 586.950 242.400 652.050 243.600 ;
        RECT 586.950 241.950 589.050 242.400 ;
        RECT 649.950 241.950 652.050 242.400 ;
        RECT 790.950 243.600 793.050 244.050 ;
        RECT 820.950 243.600 823.050 244.050 ;
        RECT 790.950 242.400 823.050 243.600 ;
        RECT 790.950 241.950 793.050 242.400 ;
        RECT 820.950 241.950 823.050 242.400 ;
        RECT 436.950 240.600 439.050 241.050 ;
        RECT 377.400 239.400 439.050 240.600 ;
        RECT 313.950 238.950 316.050 239.400 ;
        RECT 346.950 238.950 349.050 239.400 ;
        RECT 436.950 238.950 439.050 239.400 ;
        RECT 487.950 240.600 490.050 241.050 ;
        RECT 547.950 240.600 550.050 241.050 ;
        RECT 571.950 240.600 574.050 241.050 ;
        RECT 577.950 240.600 580.050 241.050 ;
        RECT 655.950 240.600 658.050 241.050 ;
        RECT 682.950 240.600 685.050 241.050 ;
        RECT 784.950 240.600 787.050 241.050 ;
        RECT 487.950 239.400 685.050 240.600 ;
        RECT 487.950 238.950 490.050 239.400 ;
        RECT 547.950 238.950 550.050 239.400 ;
        RECT 571.950 238.950 574.050 239.400 ;
        RECT 577.950 238.950 580.050 239.400 ;
        RECT 655.950 238.950 658.050 239.400 ;
        RECT 682.950 238.950 685.050 239.400 ;
        RECT 773.400 239.400 787.050 240.600 ;
        RECT 13.950 237.600 16.050 238.050 ;
        RECT 61.950 237.600 64.050 238.050 ;
        RECT 13.950 236.400 64.050 237.600 ;
        RECT 13.950 235.950 16.050 236.400 ;
        RECT 61.950 235.950 64.050 236.400 ;
        RECT 238.950 237.600 241.050 238.050 ;
        RECT 265.800 237.600 267.900 238.050 ;
        RECT 238.950 236.400 267.900 237.600 ;
        RECT 238.950 235.950 241.050 236.400 ;
        RECT 265.800 235.950 267.900 236.400 ;
        RECT 268.950 237.600 271.050 238.050 ;
        RECT 652.950 237.600 655.050 238.050 ;
        RECT 697.950 237.600 700.050 238.050 ;
        RECT 773.400 237.600 774.600 239.400 ;
        RECT 784.950 238.950 787.050 239.400 ;
        RECT 857.400 238.050 858.600 250.950 ;
        RECT 896.400 250.050 897.600 259.950 ;
        RECT 898.950 258.600 901.050 259.050 ;
        RECT 898.950 257.400 906.600 258.600 ;
        RECT 898.950 256.950 901.050 257.400 ;
        RECT 905.400 253.050 906.600 257.400 ;
        RECT 904.950 250.950 907.050 253.050 ;
        RECT 895.950 247.950 898.050 250.050 ;
        RECT 268.950 236.400 312.600 237.600 ;
        RECT 268.950 235.950 271.050 236.400 ;
        RECT 22.950 234.600 25.050 235.050 ;
        RECT 49.950 234.600 52.050 235.050 ;
        RECT 22.950 233.400 52.050 234.600 ;
        RECT 22.950 232.950 25.050 233.400 ;
        RECT 49.950 232.950 52.050 233.400 ;
        RECT 70.950 234.600 73.050 235.050 ;
        RECT 124.950 234.600 127.050 235.050 ;
        RECT 70.950 233.400 127.050 234.600 ;
        RECT 70.950 232.950 73.050 233.400 ;
        RECT 124.950 232.950 127.050 233.400 ;
        RECT 148.950 234.600 151.050 235.050 ;
        RECT 277.950 234.600 280.050 235.050 ;
        RECT 148.950 233.400 280.050 234.600 ;
        RECT 311.400 234.600 312.600 236.400 ;
        RECT 652.950 236.400 774.600 237.600 ;
        RECT 652.950 235.950 655.050 236.400 ;
        RECT 697.950 235.950 700.050 236.400 ;
        RECT 856.950 235.950 859.050 238.050 ;
        RECT 343.950 234.600 346.050 235.050 ;
        RECT 311.400 233.400 346.050 234.600 ;
        RECT 148.950 232.950 151.050 233.400 ;
        RECT 277.950 232.950 280.050 233.400 ;
        RECT 343.950 232.950 346.050 233.400 ;
        RECT 349.950 234.600 352.050 235.050 ;
        RECT 445.950 234.600 448.050 235.050 ;
        RECT 349.950 233.400 448.050 234.600 ;
        RECT 349.950 232.950 352.050 233.400 ;
        RECT 445.950 232.950 448.050 233.400 ;
        RECT 511.950 234.600 514.050 235.050 ;
        RECT 541.950 234.600 544.050 235.050 ;
        RECT 511.950 233.400 544.050 234.600 ;
        RECT 511.950 232.950 514.050 233.400 ;
        RECT 541.950 232.950 544.050 233.400 ;
        RECT 643.950 234.600 646.050 235.050 ;
        RECT 724.950 234.600 727.050 235.050 ;
        RECT 775.950 234.600 778.050 235.050 ;
        RECT 643.950 233.400 778.050 234.600 ;
        RECT 643.950 232.950 646.050 233.400 ;
        RECT 724.950 232.950 727.050 233.400 ;
        RECT 775.950 232.950 778.050 233.400 ;
        RECT 196.950 231.600 199.050 232.050 ;
        RECT 223.950 231.600 226.050 232.050 ;
        RECT 286.950 231.600 289.050 232.050 ;
        RECT 196.950 230.400 226.050 231.600 ;
        RECT 196.950 229.950 199.050 230.400 ;
        RECT 223.950 229.950 226.050 230.400 ;
        RECT 242.400 230.400 289.050 231.600 ;
        RECT 242.400 229.050 243.600 230.400 ;
        RECT 286.950 229.950 289.050 230.400 ;
        RECT 322.950 231.600 325.050 232.050 ;
        RECT 350.400 231.600 351.600 232.950 ;
        RECT 322.950 230.400 351.600 231.600 ;
        RECT 361.950 231.600 364.050 232.050 ;
        RECT 430.950 231.600 433.050 232.050 ;
        RECT 361.950 230.400 433.050 231.600 ;
        RECT 322.950 229.950 325.050 230.400 ;
        RECT 361.950 229.950 364.050 230.400 ;
        RECT 430.950 229.950 433.050 230.400 ;
        RECT 778.950 231.600 781.050 232.050 ;
        RECT 790.950 231.600 793.050 232.050 ;
        RECT 778.950 230.400 793.050 231.600 ;
        RECT 778.950 229.950 781.050 230.400 ;
        RECT 790.950 229.950 793.050 230.400 ;
        RECT 796.950 231.600 799.050 232.050 ;
        RECT 814.950 231.600 817.050 232.050 ;
        RECT 796.950 230.400 817.050 231.600 ;
        RECT 796.950 229.950 799.050 230.400 ;
        RECT 814.950 229.950 817.050 230.400 ;
        RECT 16.950 228.600 19.050 229.050 ;
        RECT 31.950 228.600 34.050 229.050 ;
        RECT 64.950 228.600 67.050 229.050 ;
        RECT 16.950 227.400 67.050 228.600 ;
        RECT 16.950 226.950 19.050 227.400 ;
        RECT 31.950 226.950 34.050 227.400 ;
        RECT 64.950 226.950 67.050 227.400 ;
        RECT 160.950 228.600 163.050 229.050 ;
        RECT 175.950 228.600 178.050 229.050 ;
        RECT 160.950 227.400 178.050 228.600 ;
        RECT 160.950 226.950 163.050 227.400 ;
        RECT 175.950 226.950 178.050 227.400 ;
        RECT 232.950 228.600 235.050 229.050 ;
        RECT 241.800 228.600 243.900 229.050 ;
        RECT 232.950 227.400 243.900 228.600 ;
        RECT 232.950 226.950 235.050 227.400 ;
        RECT 241.800 226.950 243.900 227.400 ;
        RECT 244.950 228.600 247.050 229.050 ;
        RECT 268.950 228.600 271.050 229.050 ;
        RECT 244.950 227.400 271.050 228.600 ;
        RECT 244.950 226.950 247.050 227.400 ;
        RECT 268.950 226.950 271.050 227.400 ;
        RECT 277.950 228.600 280.050 229.050 ;
        RECT 289.950 228.600 292.050 229.050 ;
        RECT 319.800 228.600 321.900 229.050 ;
        RECT 277.950 227.400 321.900 228.600 ;
        RECT 277.950 226.950 280.050 227.400 ;
        RECT 289.950 226.950 292.050 227.400 ;
        RECT 319.800 226.950 321.900 227.400 ;
        RECT 322.950 228.600 325.050 228.900 ;
        RECT 362.400 228.600 363.600 229.950 ;
        RECT 322.950 227.400 363.600 228.600 ;
        RECT 364.950 228.600 367.050 229.050 ;
        RECT 490.950 228.600 493.050 229.050 ;
        RECT 514.950 228.600 517.050 229.050 ;
        RECT 364.950 227.400 429.600 228.600 ;
        RECT 322.950 226.800 325.050 227.400 ;
        RECT 364.950 226.950 367.050 227.400 ;
        RECT 37.950 225.600 40.050 226.050 ;
        RECT 46.950 225.600 49.050 226.050 ;
        RECT 37.950 224.400 49.050 225.600 ;
        RECT 37.950 223.950 40.050 224.400 ;
        RECT 46.950 223.950 49.050 224.400 ;
        RECT 226.950 225.600 229.050 226.050 ;
        RECT 238.950 225.600 241.050 226.050 ;
        RECT 226.950 224.400 241.050 225.600 ;
        RECT 226.950 223.950 229.050 224.400 ;
        RECT 238.950 223.950 241.050 224.400 ;
        RECT 307.950 225.600 310.050 226.050 ;
        RECT 331.950 225.600 334.050 226.050 ;
        RECT 337.950 225.600 340.050 226.050 ;
        RECT 307.950 224.400 340.050 225.600 ;
        RECT 428.400 225.600 429.600 227.400 ;
        RECT 490.950 227.400 517.050 228.600 ;
        RECT 490.950 226.950 493.050 227.400 ;
        RECT 514.950 226.950 517.050 227.400 ;
        RECT 568.950 228.600 571.050 229.050 ;
        RECT 625.950 228.600 628.050 229.050 ;
        RECT 568.950 227.400 628.050 228.600 ;
        RECT 568.950 226.950 571.050 227.400 ;
        RECT 625.950 226.950 628.050 227.400 ;
        RECT 712.950 228.600 715.050 229.050 ;
        RECT 742.950 228.600 745.050 229.050 ;
        RECT 754.950 228.600 757.050 229.050 ;
        RECT 769.950 228.600 772.050 229.050 ;
        RECT 712.950 227.400 772.050 228.600 ;
        RECT 712.950 226.950 715.050 227.400 ;
        RECT 742.950 226.950 745.050 227.400 ;
        RECT 754.950 226.950 757.050 227.400 ;
        RECT 769.950 226.950 772.050 227.400 ;
        RECT 856.950 226.950 859.050 229.050 ;
        RECT 892.950 228.600 895.050 229.050 ;
        RECT 910.950 228.600 913.050 229.050 ;
        RECT 892.950 227.400 913.050 228.600 ;
        RECT 892.950 226.950 895.050 227.400 ;
        RECT 910.950 226.950 913.050 227.400 ;
        RECT 487.950 225.600 490.050 226.050 ;
        RECT 428.400 224.400 490.050 225.600 ;
        RECT 307.950 223.950 310.050 224.400 ;
        RECT 331.950 223.950 334.050 224.400 ;
        RECT 337.950 223.950 340.050 224.400 ;
        RECT 487.950 223.950 490.050 224.400 ;
        RECT 526.950 225.600 529.050 226.050 ;
        RECT 559.950 225.600 562.050 226.050 ;
        RECT 526.950 224.400 562.050 225.600 ;
        RECT 526.950 223.950 529.050 224.400 ;
        RECT 559.950 223.950 562.050 224.400 ;
        RECT 646.950 225.600 649.050 226.050 ;
        RECT 661.950 225.600 664.050 226.050 ;
        RECT 646.950 224.400 664.050 225.600 ;
        RECT 646.950 223.950 649.050 224.400 ;
        RECT 661.950 223.950 664.050 224.400 ;
        RECT 733.950 225.600 736.050 226.050 ;
        RECT 742.950 225.600 745.050 225.900 ;
        RECT 805.950 225.600 808.050 226.050 ;
        RECT 811.950 225.600 814.050 226.050 ;
        RECT 733.950 224.400 814.050 225.600 ;
        RECT 733.950 223.950 736.050 224.400 ;
        RECT 742.950 223.800 745.050 224.400 ;
        RECT 805.950 223.950 808.050 224.400 ;
        RECT 811.950 223.950 814.050 224.400 ;
        RECT 106.950 222.600 109.050 223.050 ;
        RECT 121.950 222.600 124.050 223.050 ;
        RECT 106.950 221.400 124.050 222.600 ;
        RECT 106.950 220.950 109.050 221.400 ;
        RECT 121.950 220.950 124.050 221.400 ;
        RECT 136.950 222.600 139.050 223.050 ;
        RECT 157.950 222.600 160.050 223.050 ;
        RECT 136.950 221.400 160.050 222.600 ;
        RECT 136.950 220.950 139.050 221.400 ;
        RECT 157.950 220.950 160.050 221.400 ;
        RECT 163.950 222.600 166.050 223.050 ;
        RECT 172.950 222.600 175.050 223.050 ;
        RECT 163.950 221.400 175.050 222.600 ;
        RECT 163.950 220.950 166.050 221.400 ;
        RECT 172.950 220.950 175.050 221.400 ;
        RECT 184.950 222.600 187.050 223.050 ;
        RECT 199.950 222.600 202.050 223.050 ;
        RECT 184.950 221.400 202.050 222.600 ;
        RECT 184.950 220.950 187.050 221.400 ;
        RECT 199.950 220.950 202.050 221.400 ;
        RECT 205.950 222.600 208.050 223.050 ;
        RECT 214.950 222.600 217.050 223.050 ;
        RECT 205.950 221.400 217.050 222.600 ;
        RECT 205.950 220.950 208.050 221.400 ;
        RECT 214.950 220.950 217.050 221.400 ;
        RECT 220.950 222.600 223.050 223.050 ;
        RECT 364.950 222.600 367.050 223.050 ;
        RECT 544.950 222.600 547.050 223.050 ;
        RECT 220.950 221.400 367.050 222.600 ;
        RECT 220.950 220.950 223.050 221.400 ;
        RECT 364.950 220.950 367.050 221.400 ;
        RECT 494.400 221.400 547.050 222.600 ;
        RECT 494.400 220.050 495.600 221.400 ;
        RECT 544.950 220.950 547.050 221.400 ;
        RECT 628.950 222.600 631.050 223.050 ;
        RECT 640.950 222.600 643.050 223.050 ;
        RECT 628.950 221.400 643.050 222.600 ;
        RECT 628.950 220.950 631.050 221.400 ;
        RECT 640.950 220.950 643.050 221.400 ;
        RECT 694.950 222.600 697.050 223.050 ;
        RECT 703.950 222.600 706.050 223.050 ;
        RECT 694.950 221.400 706.050 222.600 ;
        RECT 694.950 220.950 697.050 221.400 ;
        RECT 703.950 220.950 706.050 221.400 ;
        RECT 766.950 222.600 769.050 223.050 ;
        RECT 778.950 222.600 781.050 223.050 ;
        RECT 766.950 221.400 781.050 222.600 ;
        RECT 766.950 220.950 769.050 221.400 ;
        RECT 778.950 220.950 781.050 221.400 ;
        RECT 817.950 222.600 820.050 223.050 ;
        RECT 817.950 221.400 843.600 222.600 ;
        RECT 817.950 220.950 820.050 221.400 ;
        RECT 82.950 219.600 85.050 220.050 ;
        RECT 97.950 219.600 100.050 220.050 ;
        RECT 82.950 218.400 100.050 219.600 ;
        RECT 82.950 217.950 85.050 218.400 ;
        RECT 97.950 217.950 100.050 218.400 ;
        RECT 103.950 219.600 106.050 220.050 ;
        RECT 130.950 219.600 133.050 220.050 ;
        RECT 142.950 219.600 145.050 220.050 ;
        RECT 223.950 219.600 226.050 220.050 ;
        RECT 277.800 219.600 279.900 220.050 ;
        RECT 103.950 218.400 204.600 219.600 ;
        RECT 103.950 217.950 106.050 218.400 ;
        RECT 130.950 217.950 133.050 218.400 ;
        RECT 142.950 217.950 145.050 218.400 ;
        RECT 64.950 216.600 67.050 217.200 ;
        RECT 76.950 216.750 79.050 217.200 ;
        RECT 94.950 216.750 97.050 217.200 ;
        RECT 76.950 216.600 97.050 216.750 ;
        RECT 64.950 215.550 97.050 216.600 ;
        RECT 64.950 215.400 79.050 215.550 ;
        RECT 64.950 215.100 67.050 215.400 ;
        RECT 76.950 215.100 79.050 215.400 ;
        RECT 94.950 215.100 97.050 215.550 ;
        RECT 163.950 214.950 166.050 217.050 ;
        RECT 178.950 216.750 181.050 217.200 ;
        RECT 190.950 216.750 193.050 217.200 ;
        RECT 178.950 215.550 193.050 216.750 ;
        RECT 178.950 215.100 181.050 215.550 ;
        RECT 190.950 215.100 193.050 215.550 ;
        RECT 203.400 216.600 204.600 218.400 ;
        RECT 223.950 218.400 279.900 219.600 ;
        RECT 223.950 217.950 226.050 218.400 ;
        RECT 277.800 217.950 279.900 218.400 ;
        RECT 280.950 219.600 283.050 219.900 ;
        RECT 283.950 219.600 286.050 220.050 ;
        RECT 322.950 219.600 325.050 220.050 ;
        RECT 370.800 219.600 372.900 220.050 ;
        RECT 280.950 218.400 325.050 219.600 ;
        RECT 280.950 217.800 283.050 218.400 ;
        RECT 283.950 217.950 286.050 218.400 ;
        RECT 322.950 217.950 325.050 218.400 ;
        RECT 338.400 218.400 372.900 219.600 ;
        RECT 256.950 216.600 259.050 217.200 ;
        RECT 203.400 215.400 259.050 216.600 ;
        RECT 256.950 215.100 259.050 215.400 ;
        RECT 164.400 211.050 165.600 214.950 ;
        RECT 268.950 213.600 271.050 217.050 ;
        RECT 286.950 216.750 289.050 217.200 ;
        RECT 301.950 216.750 304.050 217.200 ;
        RECT 286.950 215.550 304.050 216.750 ;
        RECT 286.950 215.100 289.050 215.550 ;
        RECT 301.950 215.100 304.050 215.550 ;
        RECT 325.950 216.600 328.050 217.200 ;
        RECT 338.400 216.600 339.600 218.400 ;
        RECT 370.800 217.950 372.900 218.400 ;
        RECT 373.950 219.600 376.050 220.050 ;
        RECT 385.950 219.600 388.050 220.050 ;
        RECT 394.950 219.600 397.050 220.050 ;
        RECT 373.950 218.400 397.050 219.600 ;
        RECT 373.950 217.950 376.050 218.400 ;
        RECT 385.950 217.950 388.050 218.400 ;
        RECT 394.950 217.950 397.050 218.400 ;
        RECT 424.950 219.600 427.050 220.050 ;
        RECT 445.950 219.600 448.050 220.050 ;
        RECT 460.950 219.600 463.050 220.050 ;
        RECT 424.950 218.400 463.050 219.600 ;
        RECT 424.950 217.950 427.050 218.400 ;
        RECT 445.950 217.950 448.050 218.400 ;
        RECT 460.950 217.950 463.050 218.400 ;
        RECT 478.950 219.600 481.050 220.050 ;
        RECT 493.950 219.600 496.050 220.050 ;
        RECT 478.950 218.400 496.050 219.600 ;
        RECT 478.950 217.950 481.050 218.400 ;
        RECT 493.950 217.950 496.050 218.400 ;
        RECT 325.950 215.400 339.600 216.600 ;
        RECT 340.950 216.600 343.050 217.200 ;
        RECT 355.950 216.600 358.050 217.200 ;
        RECT 370.950 216.600 373.050 216.900 ;
        RECT 376.950 216.600 379.050 217.200 ;
        RECT 400.950 216.600 403.050 217.200 ;
        RECT 340.950 215.400 354.600 216.600 ;
        RECT 325.950 215.100 328.050 215.400 ;
        RECT 340.950 215.100 343.050 215.400 ;
        RECT 266.400 213.000 271.050 213.600 ;
        RECT 266.400 212.400 270.600 213.000 ;
        RECT 34.950 210.450 37.050 210.900 ;
        RECT 49.950 210.450 52.050 210.900 ;
        RECT 34.950 209.250 52.050 210.450 ;
        RECT 34.950 208.800 37.050 209.250 ;
        RECT 49.950 208.800 52.050 209.250 ;
        RECT 124.950 210.450 127.050 210.900 ;
        RECT 130.950 210.450 133.050 210.900 ;
        RECT 124.950 209.250 133.050 210.450 ;
        RECT 124.950 208.800 127.050 209.250 ;
        RECT 130.950 208.800 133.050 209.250 ;
        RECT 163.950 208.950 166.050 211.050 ;
        RECT 214.950 210.450 217.050 210.900 ;
        RECT 226.950 210.450 229.050 210.900 ;
        RECT 214.950 209.250 229.050 210.450 ;
        RECT 214.950 208.800 217.050 209.250 ;
        RECT 226.950 208.800 229.050 209.250 ;
        RECT 241.950 210.600 244.050 210.900 ;
        RECT 250.950 210.600 253.050 211.050 ;
        RECT 241.950 209.400 253.050 210.600 ;
        RECT 241.950 208.800 244.050 209.400 ;
        RECT 250.950 208.950 253.050 209.400 ;
        RECT 259.950 210.600 262.050 210.900 ;
        RECT 266.400 210.600 267.600 212.400 ;
        RECT 259.950 209.400 267.600 210.600 ;
        RECT 271.950 210.600 274.050 210.900 ;
        RECT 289.950 210.600 292.050 211.050 ;
        RECT 271.950 209.400 292.050 210.600 ;
        RECT 259.950 208.800 262.050 209.400 ;
        RECT 271.950 208.800 274.050 209.400 ;
        RECT 289.950 208.950 292.050 209.400 ;
        RECT 304.950 210.450 307.050 210.900 ;
        RECT 313.950 210.450 316.050 210.900 ;
        RECT 304.950 209.250 316.050 210.450 ;
        RECT 304.950 208.800 307.050 209.250 ;
        RECT 313.950 208.800 316.050 209.250 ;
        RECT 103.950 207.600 106.050 208.050 ;
        RECT 142.950 207.600 145.050 208.050 ;
        RECT 103.950 206.400 145.050 207.600 ;
        RECT 103.950 205.950 106.050 206.400 ;
        RECT 142.950 205.950 145.050 206.400 ;
        RECT 157.950 207.600 160.050 208.050 ;
        RECT 172.950 207.600 175.050 208.050 ;
        RECT 187.950 207.600 190.050 208.050 ;
        RECT 157.950 206.400 190.050 207.600 ;
        RECT 157.950 205.950 160.050 206.400 ;
        RECT 172.950 205.950 175.050 206.400 ;
        RECT 187.950 205.950 190.050 206.400 ;
        RECT 199.950 207.600 202.050 208.050 ;
        RECT 217.950 207.600 220.050 208.050 ;
        RECT 199.950 206.400 220.050 207.600 ;
        RECT 199.950 205.950 202.050 206.400 ;
        RECT 217.950 205.950 220.050 206.400 ;
        RECT 232.950 205.950 238.050 208.050 ;
        RECT 277.950 207.600 280.050 208.050 ;
        RECT 286.950 207.600 289.050 208.050 ;
        RECT 277.950 206.400 289.050 207.600 ;
        RECT 326.400 207.600 327.600 215.100 ;
        RECT 353.400 213.600 354.600 215.400 ;
        RECT 355.950 215.400 379.050 216.600 ;
        RECT 355.950 215.100 358.050 215.400 ;
        RECT 370.950 214.800 373.050 215.400 ;
        RECT 376.950 215.100 379.050 215.400 ;
        RECT 383.400 215.400 403.050 216.600 ;
        RECT 353.400 212.400 363.600 213.600 ;
        RECT 331.950 210.600 334.050 211.050 ;
        RECT 337.950 210.600 340.050 210.900 ;
        RECT 331.950 209.400 340.050 210.600 ;
        RECT 331.950 208.950 334.050 209.400 ;
        RECT 337.950 208.800 340.050 209.400 ;
        RECT 362.400 208.050 363.600 212.400 ;
        RECT 379.950 210.600 382.050 210.900 ;
        RECT 383.400 210.600 384.600 215.400 ;
        RECT 400.950 215.100 403.050 215.400 ;
        RECT 412.950 216.750 415.050 217.200 ;
        RECT 418.950 216.750 421.050 217.200 ;
        RECT 412.950 215.550 421.050 216.750 ;
        RECT 454.950 216.600 457.050 217.050 ;
        RECT 412.950 215.100 415.050 215.550 ;
        RECT 418.950 215.100 421.050 215.550 ;
        RECT 443.400 215.400 457.050 216.600 ;
        RECT 443.400 213.600 444.600 215.400 ;
        RECT 454.950 214.950 457.050 215.400 ;
        RECT 466.950 216.750 469.050 217.200 ;
        RECT 472.800 216.750 474.900 217.200 ;
        RECT 466.950 215.550 474.900 216.750 ;
        RECT 466.950 215.100 469.050 215.550 ;
        RECT 472.800 215.100 474.900 215.550 ;
        RECT 475.950 213.600 478.050 217.050 ;
        RECT 487.950 216.750 490.050 217.200 ;
        RECT 496.800 216.750 498.900 217.200 ;
        RECT 487.950 215.550 498.900 216.750 ;
        RECT 487.950 215.100 490.050 215.550 ;
        RECT 496.800 215.100 498.900 215.550 ;
        RECT 499.950 216.600 504.000 217.050 ;
        RECT 505.950 216.600 508.050 217.200 ;
        RECT 511.950 216.600 514.050 220.050 ;
        RECT 592.950 217.950 595.050 220.050 ;
        RECT 736.950 219.600 739.050 220.050 ;
        RECT 745.950 219.600 748.050 220.050 ;
        RECT 736.950 218.400 748.050 219.600 ;
        RECT 736.950 217.950 739.050 218.400 ;
        RECT 745.950 217.950 748.050 218.400 ;
        RECT 757.950 219.600 762.000 220.050 ;
        RECT 757.950 217.950 762.600 219.600 ;
        RECT 808.950 217.950 811.050 220.050 ;
        RECT 823.950 219.600 826.050 220.050 ;
        RECT 838.950 219.600 841.050 220.050 ;
        RECT 823.950 218.400 841.050 219.600 ;
        RECT 823.950 217.950 826.050 218.400 ;
        RECT 838.950 217.950 841.050 218.400 ;
        RECT 499.950 214.950 504.600 216.600 ;
        RECT 505.950 216.000 514.050 216.600 ;
        RECT 520.950 216.750 523.050 217.200 ;
        RECT 532.950 216.750 535.050 217.200 ;
        RECT 505.950 215.400 513.600 216.000 ;
        RECT 520.950 215.550 535.050 216.750 ;
        RECT 505.950 215.100 508.050 215.400 ;
        RECT 520.950 215.100 523.050 215.550 ;
        RECT 532.950 215.100 535.050 215.550 ;
        RECT 553.950 216.750 556.050 217.200 ;
        RECT 565.950 216.750 568.050 217.200 ;
        RECT 553.950 215.550 568.050 216.750 ;
        RECT 553.950 215.100 556.050 215.550 ;
        RECT 565.950 215.100 568.050 215.550 ;
        RECT 571.950 216.600 574.050 217.200 ;
        RECT 589.950 216.600 592.050 217.200 ;
        RECT 571.950 215.400 592.050 216.600 ;
        RECT 571.950 215.100 574.050 215.400 ;
        RECT 589.950 215.100 592.050 215.400 ;
        RECT 503.400 213.600 504.600 214.950 ;
        RECT 440.400 212.400 444.600 213.600 ;
        RECT 446.400 212.400 474.600 213.600 ;
        RECT 475.950 213.000 480.600 213.600 ;
        RECT 476.400 212.400 480.600 213.000 ;
        RECT 503.400 213.000 525.600 213.600 ;
        RECT 503.400 212.400 526.050 213.000 ;
        RECT 379.950 209.400 384.600 210.600 ;
        RECT 430.950 210.600 433.050 211.050 ;
        RECT 440.400 210.600 441.600 212.400 ;
        RECT 430.950 209.400 441.600 210.600 ;
        RECT 442.950 210.600 445.050 210.900 ;
        RECT 446.400 210.600 447.600 212.400 ;
        RECT 473.400 211.050 474.600 212.400 ;
        RECT 479.400 211.050 480.600 212.400 ;
        RECT 442.950 209.400 447.600 210.600 ;
        RECT 448.950 210.600 451.050 210.900 ;
        RECT 457.950 210.600 460.050 210.900 ;
        RECT 448.950 209.400 460.050 210.600 ;
        RECT 473.400 209.400 478.050 211.050 ;
        RECT 479.400 209.400 483.900 211.050 ;
        RECT 379.950 208.800 382.050 209.400 ;
        RECT 430.950 208.950 433.050 209.400 ;
        RECT 442.950 208.800 445.050 209.400 ;
        RECT 448.950 208.800 451.050 209.400 ;
        RECT 457.950 208.800 460.050 209.400 ;
        RECT 474.000 208.950 478.050 209.400 ;
        RECT 480.000 208.950 483.900 209.400 ;
        RECT 484.950 210.450 487.050 210.900 ;
        RECT 490.800 210.450 492.900 210.900 ;
        RECT 484.950 209.250 492.900 210.450 ;
        RECT 484.950 208.800 487.050 209.250 ;
        RECT 490.800 208.800 492.900 209.250 ;
        RECT 493.950 210.600 496.050 211.050 ;
        RECT 502.950 210.600 505.050 210.900 ;
        RECT 493.950 209.400 505.050 210.600 ;
        RECT 493.950 208.950 496.050 209.400 ;
        RECT 502.950 208.800 505.050 209.400 ;
        RECT 508.950 210.600 511.050 210.900 ;
        RECT 514.950 210.600 517.050 211.050 ;
        RECT 508.950 209.400 517.050 210.600 ;
        RECT 508.950 208.800 511.050 209.400 ;
        RECT 514.950 208.950 517.050 209.400 ;
        RECT 523.950 208.950 526.050 212.400 ;
        RECT 541.950 210.600 544.050 211.050 ;
        RECT 556.950 210.600 559.050 211.050 ;
        RECT 541.950 209.400 559.050 210.600 ;
        RECT 541.950 208.950 544.050 209.400 ;
        RECT 556.950 208.950 559.050 209.400 ;
        RECT 586.950 210.600 589.050 210.900 ;
        RECT 593.400 210.600 594.600 217.950 ;
        RECT 595.950 216.600 598.050 217.200 ;
        RECT 610.950 216.600 613.050 217.200 ;
        RECT 595.950 215.400 613.050 216.600 ;
        RECT 595.950 215.100 598.050 215.400 ;
        RECT 610.950 215.100 613.050 215.400 ;
        RECT 619.950 216.600 622.050 217.200 ;
        RECT 637.950 216.600 640.050 217.200 ;
        RECT 619.950 215.400 640.050 216.600 ;
        RECT 619.950 215.100 622.050 215.400 ;
        RECT 637.950 215.100 640.050 215.400 ;
        RECT 679.950 215.100 682.050 217.200 ;
        RECT 586.950 209.400 594.600 210.600 ;
        RECT 604.950 210.450 607.050 210.900 ;
        RECT 613.950 210.450 616.050 210.900 ;
        RECT 331.950 207.600 334.050 207.900 ;
        RECT 326.400 206.400 334.050 207.600 ;
        RECT 277.950 205.950 280.050 206.400 ;
        RECT 286.950 205.950 289.050 206.400 ;
        RECT 331.950 205.800 334.050 206.400 ;
        RECT 361.950 205.950 364.050 208.050 ;
        RECT 412.950 207.600 415.050 208.050 ;
        RECT 418.950 207.600 421.050 208.050 ;
        RECT 412.950 206.400 421.050 207.600 ;
        RECT 412.950 205.950 415.050 206.400 ;
        RECT 418.950 205.950 421.050 206.400 ;
        RECT 433.950 207.600 436.050 208.050 ;
        RECT 448.950 207.600 451.050 208.050 ;
        RECT 433.950 206.400 451.050 207.600 ;
        RECT 524.400 207.600 525.600 208.950 ;
        RECT 586.950 208.800 589.050 209.400 ;
        RECT 604.950 209.250 616.050 210.450 ;
        RECT 604.950 208.800 607.050 209.250 ;
        RECT 613.950 208.800 616.050 209.250 ;
        RECT 664.950 210.600 667.050 210.900 ;
        RECT 670.950 210.600 673.050 211.050 ;
        RECT 664.950 209.400 673.050 210.600 ;
        RECT 664.950 208.800 667.050 209.400 ;
        RECT 670.950 208.950 673.050 209.400 ;
        RECT 565.950 207.600 568.050 208.050 ;
        RECT 524.400 206.400 568.050 207.600 ;
        RECT 433.950 205.950 436.050 206.400 ;
        RECT 448.950 205.950 451.050 206.400 ;
        RECT 565.950 205.950 568.050 206.400 ;
        RECT 673.950 207.600 676.050 208.050 ;
        RECT 680.400 207.600 681.600 215.100 ;
        RECT 688.950 214.950 691.050 217.050 ;
        RECT 715.950 216.600 718.050 217.050 ;
        RECT 727.950 216.600 730.050 217.200 ;
        RECT 715.950 215.400 730.050 216.600 ;
        RECT 715.950 214.950 718.050 215.400 ;
        RECT 727.950 215.100 730.050 215.400 ;
        RECT 739.950 214.950 742.050 217.050 ;
        RECT 682.950 210.600 685.050 210.900 ;
        RECT 689.400 210.600 690.600 214.950 ;
        RECT 740.400 211.050 741.600 214.950 ;
        RECT 761.400 211.050 762.600 217.950 ;
        RECT 775.950 216.600 778.050 217.200 ;
        RECT 784.800 216.600 786.900 217.050 ;
        RECT 775.950 215.400 786.900 216.600 ;
        RECT 775.950 215.100 778.050 215.400 ;
        RECT 784.800 214.950 786.900 215.400 ;
        RECT 802.950 214.950 805.050 217.050 ;
        RECT 682.950 209.400 690.600 210.600 ;
        RECT 694.950 210.450 697.050 210.900 ;
        RECT 700.950 210.450 703.050 210.900 ;
        RECT 682.950 208.800 685.050 209.400 ;
        RECT 694.950 209.250 703.050 210.450 ;
        RECT 694.950 208.800 697.050 209.250 ;
        RECT 700.950 208.800 703.050 209.250 ;
        RECT 718.950 210.600 721.050 211.050 ;
        RECT 730.950 210.600 733.050 210.900 ;
        RECT 718.950 209.400 733.050 210.600 ;
        RECT 718.950 208.950 721.050 209.400 ;
        RECT 730.950 208.800 733.050 209.400 ;
        RECT 739.950 208.950 742.050 211.050 ;
        RECT 760.950 208.950 763.050 211.050 ;
        RECT 803.400 210.600 804.600 214.950 ;
        RECT 809.400 213.600 810.600 217.950 ;
        RECT 811.950 216.600 814.050 217.200 ;
        RECT 811.950 215.400 819.600 216.600 ;
        RECT 811.950 215.100 814.050 215.400 ;
        RECT 818.400 213.600 819.600 215.400 ;
        RECT 820.950 213.600 823.050 213.900 ;
        RECT 809.400 212.400 816.600 213.600 ;
        RECT 818.400 212.400 823.050 213.600 ;
        RECT 808.950 210.600 811.050 210.900 ;
        RECT 803.400 209.400 811.050 210.600 ;
        RECT 815.400 210.600 816.600 212.400 ;
        RECT 820.950 211.800 823.050 212.400 ;
        RECT 829.950 213.450 832.050 213.900 ;
        RECT 835.950 213.450 838.050 213.900 ;
        RECT 829.950 212.250 838.050 213.450 ;
        RECT 829.950 211.800 832.050 212.250 ;
        RECT 835.950 211.800 838.050 212.250 ;
        RECT 823.950 210.600 826.050 211.050 ;
        RECT 815.400 209.400 826.050 210.600 ;
        RECT 808.950 208.800 811.050 209.400 ;
        RECT 823.950 208.950 826.050 209.400 ;
        RECT 673.950 206.400 681.600 207.600 ;
        RECT 742.950 207.600 745.050 208.050 ;
        RECT 751.950 207.600 754.050 208.050 ;
        RECT 742.950 206.400 754.050 207.600 ;
        RECT 673.950 205.950 676.050 206.400 ;
        RECT 742.950 205.950 745.050 206.400 ;
        RECT 751.950 205.950 754.050 206.400 ;
        RECT 829.950 207.600 832.050 208.050 ;
        RECT 838.950 207.600 841.050 208.050 ;
        RECT 829.950 206.400 841.050 207.600 ;
        RECT 829.950 205.950 832.050 206.400 ;
        RECT 838.950 205.950 841.050 206.400 ;
        RECT 19.950 204.600 22.050 205.050 ;
        RECT 46.950 204.600 49.050 205.050 ;
        RECT 100.950 204.600 103.050 205.050 ;
        RECT 19.950 203.400 103.050 204.600 ;
        RECT 19.950 202.950 22.050 203.400 ;
        RECT 46.950 202.950 49.050 203.400 ;
        RECT 100.950 202.950 103.050 203.400 ;
        RECT 106.950 204.600 109.050 205.050 ;
        RECT 118.950 204.600 121.050 205.050 ;
        RECT 139.950 204.600 142.050 205.050 ;
        RECT 271.950 204.600 274.050 205.050 ;
        RECT 106.950 203.400 274.050 204.600 ;
        RECT 106.950 202.950 109.050 203.400 ;
        RECT 118.950 202.950 121.050 203.400 ;
        RECT 139.950 202.950 142.050 203.400 ;
        RECT 271.950 202.950 274.050 203.400 ;
        RECT 298.950 204.600 301.050 205.050 ;
        RECT 316.950 204.600 319.050 205.050 ;
        RECT 298.950 203.400 319.050 204.600 ;
        RECT 298.950 202.950 301.050 203.400 ;
        RECT 316.950 202.950 319.050 203.400 ;
        RECT 322.950 204.600 325.050 205.050 ;
        RECT 340.950 204.600 343.050 205.050 ;
        RECT 322.950 203.400 343.050 204.600 ;
        RECT 322.950 202.950 325.050 203.400 ;
        RECT 340.950 202.950 343.050 203.400 ;
        RECT 346.950 204.600 349.050 205.050 ;
        RECT 376.950 204.600 379.050 205.050 ;
        RECT 346.950 203.400 379.050 204.600 ;
        RECT 346.950 202.950 349.050 203.400 ;
        RECT 376.950 202.950 379.050 203.400 ;
        RECT 391.950 204.600 394.050 205.050 ;
        RECT 409.950 204.600 412.050 205.050 ;
        RECT 391.950 203.400 412.050 204.600 ;
        RECT 391.950 202.950 394.050 203.400 ;
        RECT 409.950 202.950 412.050 203.400 ;
        RECT 463.950 204.600 466.050 205.050 ;
        RECT 469.950 204.600 472.050 205.050 ;
        RECT 463.950 203.400 472.050 204.600 ;
        RECT 463.950 202.950 466.050 203.400 ;
        RECT 469.950 202.950 472.050 203.400 ;
        RECT 496.950 204.600 499.050 205.050 ;
        RECT 520.950 204.600 523.050 205.050 ;
        RECT 496.950 203.400 523.050 204.600 ;
        RECT 496.950 202.950 499.050 203.400 ;
        RECT 520.950 202.950 523.050 203.400 ;
        RECT 535.950 204.600 538.050 205.050 ;
        RECT 544.950 204.600 547.050 205.050 ;
        RECT 550.950 204.600 553.050 205.050 ;
        RECT 535.950 203.400 553.050 204.600 ;
        RECT 535.950 202.950 538.050 203.400 ;
        RECT 544.950 202.950 547.050 203.400 ;
        RECT 550.950 202.950 553.050 203.400 ;
        RECT 568.950 204.600 571.050 205.050 ;
        RECT 577.950 204.600 580.050 205.050 ;
        RECT 568.950 203.400 580.050 204.600 ;
        RECT 568.950 202.950 571.050 203.400 ;
        RECT 577.950 202.950 580.050 203.400 ;
        RECT 592.950 204.600 595.050 205.050 ;
        RECT 640.950 204.600 643.050 205.050 ;
        RECT 658.950 204.600 661.050 205.050 ;
        RECT 592.950 203.400 661.050 204.600 ;
        RECT 592.950 202.950 595.050 203.400 ;
        RECT 640.950 202.950 643.050 203.400 ;
        RECT 658.950 202.950 661.050 203.400 ;
        RECT 691.950 204.600 694.050 205.050 ;
        RECT 736.950 204.600 739.050 205.050 ;
        RECT 757.950 204.600 760.050 205.050 ;
        RECT 793.950 204.600 796.050 205.050 ;
        RECT 820.950 204.600 823.050 205.050 ;
        RECT 691.950 203.400 735.600 204.600 ;
        RECT 691.950 202.950 694.050 203.400 ;
        RECT 46.950 201.600 49.050 201.900 ;
        RECT 70.950 201.600 73.050 202.050 ;
        RECT 100.950 201.600 103.050 201.900 ;
        RECT 46.950 200.400 103.050 201.600 ;
        RECT 46.950 199.800 49.050 200.400 ;
        RECT 70.950 199.950 73.050 200.400 ;
        RECT 100.950 199.800 103.050 200.400 ;
        RECT 151.950 201.600 154.050 202.050 ;
        RECT 166.950 201.600 169.050 202.050 ;
        RECT 151.950 200.400 169.050 201.600 ;
        RECT 151.950 199.950 154.050 200.400 ;
        RECT 166.950 199.950 169.050 200.400 ;
        RECT 412.950 201.600 415.050 202.050 ;
        RECT 421.950 201.600 424.050 202.050 ;
        RECT 412.950 200.400 424.050 201.600 ;
        RECT 412.950 199.950 415.050 200.400 ;
        RECT 421.950 199.950 424.050 200.400 ;
        RECT 427.950 201.600 430.050 202.050 ;
        RECT 442.950 201.600 445.050 202.050 ;
        RECT 472.950 201.600 475.050 202.050 ;
        RECT 478.950 201.600 481.050 202.050 ;
        RECT 580.950 201.600 583.050 202.050 ;
        RECT 427.950 200.400 583.050 201.600 ;
        RECT 427.950 199.950 430.050 200.400 ;
        RECT 442.950 199.950 445.050 200.400 ;
        RECT 472.950 199.950 475.050 200.400 ;
        RECT 478.950 199.950 481.050 200.400 ;
        RECT 580.950 199.950 583.050 200.400 ;
        RECT 700.950 201.600 703.050 202.050 ;
        RECT 718.950 201.600 721.050 202.050 ;
        RECT 700.950 200.400 721.050 201.600 ;
        RECT 734.400 201.600 735.600 203.400 ;
        RECT 736.950 203.400 823.050 204.600 ;
        RECT 736.950 202.950 739.050 203.400 ;
        RECT 757.950 202.950 760.050 203.400 ;
        RECT 793.950 202.950 796.050 203.400 ;
        RECT 820.950 202.950 823.050 203.400 ;
        RECT 832.950 204.600 835.050 205.050 ;
        RECT 842.400 204.600 843.600 221.400 ;
        RECT 857.400 213.600 858.600 226.950 ;
        RECT 889.950 222.600 892.050 223.050 ;
        RECT 907.950 222.600 910.050 223.050 ;
        RECT 889.950 221.400 910.050 222.600 ;
        RECT 889.950 220.950 892.050 221.400 ;
        RECT 907.950 220.950 910.050 221.400 ;
        RECT 901.950 216.600 904.050 217.200 ;
        RECT 887.400 215.400 904.050 216.600 ;
        RECT 859.950 213.600 862.050 214.200 ;
        RECT 857.400 212.400 862.050 213.600 ;
        RECT 859.950 212.100 862.050 212.400 ;
        RECT 877.950 213.600 880.050 213.900 ;
        RECT 887.400 213.600 888.600 215.400 ;
        RECT 901.950 215.100 904.050 215.400 ;
        RECT 877.950 212.400 888.600 213.600 ;
        RECT 877.950 211.800 880.050 212.400 ;
        RECT 832.950 203.400 843.600 204.600 ;
        RECT 832.950 202.950 835.050 203.400 ;
        RECT 742.950 201.600 745.050 202.050 ;
        RECT 734.400 200.400 745.050 201.600 ;
        RECT 700.950 199.950 703.050 200.400 ;
        RECT 718.950 199.950 721.050 200.400 ;
        RECT 742.950 199.950 745.050 200.400 ;
        RECT 892.950 201.600 895.050 202.050 ;
        RECT 901.950 201.600 904.050 202.050 ;
        RECT 892.950 200.400 904.050 201.600 ;
        RECT 892.950 199.950 895.050 200.400 ;
        RECT 901.950 199.950 904.050 200.400 ;
        RECT 16.950 198.600 19.050 199.050 ;
        RECT 52.950 198.600 55.050 199.050 ;
        RECT 16.950 197.400 55.050 198.600 ;
        RECT 16.950 196.950 19.050 197.400 ;
        RECT 52.950 196.950 55.050 197.400 ;
        RECT 160.950 198.600 163.050 199.050 ;
        RECT 187.950 198.600 190.050 199.050 ;
        RECT 160.950 197.400 190.050 198.600 ;
        RECT 160.950 196.950 163.050 197.400 ;
        RECT 187.950 196.950 190.050 197.400 ;
        RECT 271.950 198.600 274.050 199.050 ;
        RECT 295.950 198.600 298.050 199.050 ;
        RECT 271.950 197.400 298.050 198.600 ;
        RECT 271.950 196.950 274.050 197.400 ;
        RECT 295.950 196.950 298.050 197.400 ;
        RECT 316.950 198.600 319.050 199.050 ;
        RECT 400.950 198.600 403.050 199.050 ;
        RECT 586.950 198.600 589.050 199.050 ;
        RECT 316.950 197.400 589.050 198.600 ;
        RECT 316.950 196.950 319.050 197.400 ;
        RECT 400.950 196.950 403.050 197.400 ;
        RECT 586.950 196.950 589.050 197.400 ;
        RECT 835.950 198.600 838.050 199.050 ;
        RECT 850.950 198.600 853.050 199.050 ;
        RECT 835.950 197.400 853.050 198.600 ;
        RECT 835.950 196.950 838.050 197.400 ;
        RECT 850.950 196.950 853.050 197.400 ;
        RECT 856.950 198.600 859.050 199.050 ;
        RECT 895.950 198.600 898.050 199.050 ;
        RECT 856.950 197.400 898.050 198.600 ;
        RECT 856.950 196.950 859.050 197.400 ;
        RECT 895.950 196.950 898.050 197.400 ;
        RECT 73.950 195.600 76.050 196.050 ;
        RECT 127.950 195.600 130.050 196.050 ;
        RECT 154.950 195.600 157.050 196.050 ;
        RECT 73.950 194.400 157.050 195.600 ;
        RECT 73.950 193.950 76.050 194.400 ;
        RECT 127.950 193.950 130.050 194.400 ;
        RECT 154.950 193.950 157.050 194.400 ;
        RECT 202.950 195.600 205.050 196.050 ;
        RECT 232.950 195.600 235.050 196.050 ;
        RECT 265.950 195.600 268.050 196.050 ;
        RECT 202.950 194.400 268.050 195.600 ;
        RECT 202.950 193.950 205.050 194.400 ;
        RECT 232.950 193.950 235.050 194.400 ;
        RECT 265.950 193.950 268.050 194.400 ;
        RECT 322.950 195.600 325.050 196.050 ;
        RECT 346.950 195.600 349.050 196.050 ;
        RECT 322.950 194.400 349.050 195.600 ;
        RECT 322.950 193.950 325.050 194.400 ;
        RECT 346.950 193.950 349.050 194.400 ;
        RECT 397.950 195.600 400.050 196.050 ;
        RECT 412.950 195.600 415.050 196.050 ;
        RECT 397.950 194.400 415.050 195.600 ;
        RECT 397.950 193.950 400.050 194.400 ;
        RECT 412.950 193.950 415.050 194.400 ;
        RECT 418.950 195.600 421.050 196.050 ;
        RECT 463.950 195.600 466.050 196.050 ;
        RECT 529.950 195.600 532.050 196.050 ;
        RECT 541.950 195.600 544.050 196.050 ;
        RECT 418.950 194.400 501.600 195.600 ;
        RECT 418.950 193.950 421.050 194.400 ;
        RECT 463.950 193.950 466.050 194.400 ;
        RECT 500.400 193.050 501.600 194.400 ;
        RECT 529.950 194.400 544.050 195.600 ;
        RECT 529.950 193.950 532.050 194.400 ;
        RECT 541.950 193.950 544.050 194.400 ;
        RECT 706.950 195.600 709.050 196.050 ;
        RECT 721.950 195.600 724.050 196.050 ;
        RECT 706.950 194.400 724.050 195.600 ;
        RECT 706.950 193.950 709.050 194.400 ;
        RECT 721.950 193.950 724.050 194.400 ;
        RECT 829.950 195.600 832.050 196.050 ;
        RECT 853.950 195.600 856.050 196.050 ;
        RECT 829.950 194.400 856.050 195.600 ;
        RECT 829.950 193.950 832.050 194.400 ;
        RECT 853.950 193.950 856.050 194.400 ;
        RECT 877.950 195.600 880.050 196.050 ;
        RECT 877.950 194.400 894.600 195.600 ;
        RECT 877.950 193.950 880.050 194.400 ;
        RECT 79.950 192.600 82.050 193.050 ;
        RECT 106.950 192.600 109.050 193.050 ;
        RECT 112.950 192.600 115.050 193.050 ;
        RECT 79.950 191.400 115.050 192.600 ;
        RECT 79.950 190.950 82.050 191.400 ;
        RECT 106.950 190.950 109.050 191.400 ;
        RECT 112.950 190.950 115.050 191.400 ;
        RECT 163.950 192.600 166.050 193.050 ;
        RECT 169.950 192.600 172.050 193.050 ;
        RECT 178.950 192.600 181.050 193.050 ;
        RECT 415.950 192.600 418.050 193.050 ;
        RECT 163.950 191.400 181.050 192.600 ;
        RECT 163.950 190.950 166.050 191.400 ;
        RECT 169.950 190.950 172.050 191.400 ;
        RECT 178.950 190.950 181.050 191.400 ;
        RECT 371.400 191.400 418.050 192.600 ;
        RECT 371.400 190.050 372.600 191.400 ;
        RECT 415.950 190.950 418.050 191.400 ;
        RECT 499.950 192.600 502.050 193.050 ;
        RECT 517.950 192.600 520.050 193.050 ;
        RECT 499.950 191.400 520.050 192.600 ;
        RECT 499.950 190.950 502.050 191.400 ;
        RECT 517.950 190.950 520.050 191.400 ;
        RECT 625.950 192.600 628.050 193.050 ;
        RECT 649.950 192.600 652.050 193.050 ;
        RECT 625.950 191.400 652.050 192.600 ;
        RECT 625.950 190.950 628.050 191.400 ;
        RECT 649.950 190.950 652.050 191.400 ;
        RECT 820.950 192.600 823.050 193.050 ;
        RECT 832.950 192.600 835.050 193.050 ;
        RECT 820.950 191.400 835.050 192.600 ;
        RECT 893.400 192.600 894.600 194.400 ;
        RECT 913.950 192.600 916.050 193.050 ;
        RECT 893.400 191.400 916.050 192.600 ;
        RECT 820.950 190.950 823.050 191.400 ;
        RECT 832.950 190.950 835.050 191.400 ;
        RECT 913.950 190.950 916.050 191.400 ;
        RECT 28.950 189.600 31.050 190.050 ;
        RECT 40.950 189.600 43.050 190.050 ;
        RECT 28.950 188.400 43.050 189.600 ;
        RECT 28.950 187.950 31.050 188.400 ;
        RECT 40.950 187.950 43.050 188.400 ;
        RECT 94.950 189.600 97.050 190.050 ;
        RECT 121.950 189.600 124.050 190.050 ;
        RECT 145.950 189.600 148.050 190.050 ;
        RECT 94.950 188.400 148.050 189.600 ;
        RECT 94.950 187.950 97.050 188.400 ;
        RECT 121.950 187.950 124.050 188.400 ;
        RECT 145.950 187.950 148.050 188.400 ;
        RECT 193.950 189.600 196.050 190.050 ;
        RECT 199.950 189.600 202.050 190.050 ;
        RECT 193.950 188.400 202.050 189.600 ;
        RECT 193.950 187.950 196.050 188.400 ;
        RECT 199.950 187.950 202.050 188.400 ;
        RECT 226.950 189.600 229.050 190.050 ;
        RECT 277.950 189.600 280.050 190.050 ;
        RECT 226.950 188.400 280.050 189.600 ;
        RECT 226.950 187.950 229.050 188.400 ;
        RECT 277.950 187.950 280.050 188.400 ;
        RECT 322.950 189.600 325.050 190.050 ;
        RECT 370.950 189.600 373.050 190.050 ;
        RECT 322.950 188.400 373.050 189.600 ;
        RECT 322.950 187.950 325.050 188.400 ;
        RECT 370.950 187.950 373.050 188.400 ;
        RECT 427.950 189.600 430.050 190.050 ;
        RECT 454.950 189.600 457.050 190.050 ;
        RECT 484.950 189.600 487.050 190.050 ;
        RECT 427.950 188.400 487.050 189.600 ;
        RECT 427.950 187.950 430.050 188.400 ;
        RECT 454.950 187.950 457.050 188.400 ;
        RECT 484.950 187.950 487.050 188.400 ;
        RECT 535.950 189.600 538.050 190.050 ;
        RECT 583.950 189.600 586.050 190.050 ;
        RECT 592.950 189.600 595.050 190.050 ;
        RECT 535.950 188.400 595.050 189.600 ;
        RECT 535.950 187.950 538.050 188.400 ;
        RECT 583.950 187.950 586.050 188.400 ;
        RECT 592.950 187.950 595.050 188.400 ;
        RECT 601.950 189.600 604.050 190.050 ;
        RECT 616.950 189.600 619.050 190.050 ;
        RECT 601.950 188.400 619.050 189.600 ;
        RECT 601.950 187.950 604.050 188.400 ;
        RECT 616.950 187.950 619.050 188.400 ;
        RECT 772.950 189.600 775.050 190.050 ;
        RECT 811.950 189.600 814.050 190.050 ;
        RECT 772.950 188.400 814.050 189.600 ;
        RECT 772.950 187.950 775.050 188.400 ;
        RECT 811.950 187.950 814.050 188.400 ;
        RECT 13.950 184.950 16.050 187.050 ;
        RECT 82.950 186.600 85.050 187.050 ;
        RECT 97.950 186.600 100.050 187.050 ;
        RECT 82.950 185.400 100.050 186.600 ;
        RECT 82.950 184.950 85.050 185.400 ;
        RECT 97.950 184.950 100.050 185.400 ;
        RECT 241.950 186.600 244.050 187.050 ;
        RECT 253.950 186.600 256.050 187.050 ;
        RECT 241.950 185.400 256.050 186.600 ;
        RECT 241.950 184.950 244.050 185.400 ;
        RECT 253.950 184.950 256.050 185.400 ;
        RECT 307.950 186.600 310.050 187.050 ;
        RECT 316.950 186.600 319.050 187.050 ;
        RECT 307.950 185.400 319.050 186.600 ;
        RECT 307.950 184.950 310.050 185.400 ;
        RECT 316.950 184.950 319.050 185.400 ;
        RECT 331.800 186.000 333.900 187.050 ;
        RECT 334.950 186.600 337.050 187.050 ;
        RECT 349.950 186.600 352.050 187.050 ;
        RECT 331.800 184.950 334.050 186.000 ;
        RECT 334.950 185.400 352.050 186.600 ;
        RECT 334.950 184.950 337.050 185.400 ;
        RECT 349.950 184.950 352.050 185.400 ;
        RECT 358.950 184.950 361.050 187.050 ;
        RECT 376.950 186.600 379.050 187.050 ;
        RECT 406.950 186.600 409.050 187.050 ;
        RECT 376.950 185.400 409.050 186.600 ;
        RECT 376.950 184.950 379.050 185.400 ;
        RECT 406.950 184.950 409.050 185.400 ;
        RECT 463.950 184.950 466.050 187.050 ;
        RECT 481.950 186.600 484.050 187.050 ;
        RECT 473.400 185.400 484.050 186.600 ;
        RECT 14.400 177.900 15.600 184.950 ;
        RECT 22.950 183.600 25.050 184.200 ;
        RECT 37.950 183.600 40.050 184.200 ;
        RECT 49.950 183.600 52.050 184.050 ;
        RECT 55.950 183.600 58.050 184.200 ;
        RECT 22.950 182.400 52.050 183.600 ;
        RECT 22.950 182.100 25.050 182.400 ;
        RECT 37.950 182.100 40.050 182.400 ;
        RECT 49.950 181.950 52.050 182.400 ;
        RECT 53.400 182.400 58.050 183.600 ;
        RECT 53.400 180.600 54.600 182.400 ;
        RECT 55.950 182.100 58.050 182.400 ;
        RECT 61.950 182.100 64.050 184.200 ;
        RECT 109.950 183.600 112.050 184.050 ;
        RECT 115.950 183.600 118.050 184.200 ;
        RECT 126.000 183.600 130.050 184.050 ;
        RECT 109.950 182.400 118.050 183.600 ;
        RECT 35.400 179.400 54.600 180.600 ;
        RECT 35.400 177.900 36.600 179.400 ;
        RECT 13.950 175.800 16.050 177.900 ;
        RECT 19.950 177.450 22.050 177.900 ;
        RECT 28.950 177.450 31.050 177.900 ;
        RECT 19.950 176.250 31.050 177.450 ;
        RECT 19.950 175.800 22.050 176.250 ;
        RECT 28.950 175.800 31.050 176.250 ;
        RECT 34.950 175.800 37.050 177.900 ;
        RECT 62.400 177.600 63.600 182.100 ;
        RECT 109.950 181.950 112.050 182.400 ;
        RECT 115.950 182.100 118.050 182.400 ;
        RECT 125.400 181.950 130.050 183.600 ;
        RECT 136.950 182.100 139.050 184.200 ;
        RECT 154.950 183.600 157.050 184.050 ;
        RECT 163.950 183.600 166.050 184.200 ;
        RECT 193.950 183.600 196.050 184.200 ;
        RECT 214.950 183.600 217.050 184.200 ;
        RECT 154.950 182.400 166.050 183.600 ;
        RECT 70.950 177.600 73.050 178.050 ;
        RECT 125.400 177.900 126.600 181.950 ;
        RECT 137.400 180.600 138.600 182.100 ;
        RECT 154.950 181.950 157.050 182.400 ;
        RECT 163.950 182.100 166.050 182.400 ;
        RECT 170.400 182.400 196.050 183.600 ;
        RECT 170.400 180.600 171.600 182.400 ;
        RECT 193.950 182.100 196.050 182.400 ;
        RECT 197.400 182.400 217.050 183.600 ;
        RECT 137.400 179.400 144.600 180.600 ;
        RECT 161.400 180.000 171.600 180.600 ;
        RECT 62.400 176.400 73.050 177.600 ;
        RECT 70.950 175.950 73.050 176.400 ;
        RECT 76.950 177.600 79.050 177.900 ;
        RECT 91.950 177.600 94.050 177.900 ;
        RECT 76.950 176.400 94.050 177.600 ;
        RECT 76.950 175.800 79.050 176.400 ;
        RECT 91.950 175.800 94.050 176.400 ;
        RECT 97.950 177.450 100.050 177.900 ;
        RECT 106.950 177.600 109.050 177.900 ;
        RECT 118.950 177.600 121.050 177.900 ;
        RECT 106.950 177.450 121.050 177.600 ;
        RECT 97.950 176.400 121.050 177.450 ;
        RECT 97.950 176.250 109.050 176.400 ;
        RECT 97.950 175.800 100.050 176.250 ;
        RECT 106.950 175.800 109.050 176.250 ;
        RECT 118.950 175.800 121.050 176.400 ;
        RECT 124.950 175.800 127.050 177.900 ;
        RECT 143.400 177.600 144.600 179.400 ;
        RECT 160.950 179.400 171.600 180.000 ;
        RECT 148.950 177.600 151.050 178.050 ;
        RECT 143.400 176.400 151.050 177.600 ;
        RECT 148.950 175.950 151.050 176.400 ;
        RECT 160.950 175.950 163.050 179.400 ;
        RECT 197.400 178.050 198.600 182.400 ;
        RECT 214.950 182.100 217.050 182.400 ;
        RECT 259.950 183.600 262.050 184.200 ;
        RECT 268.950 183.600 271.050 184.050 ;
        RECT 259.950 182.400 271.050 183.600 ;
        RECT 259.950 182.100 262.050 182.400 ;
        RECT 268.950 181.950 271.050 182.400 ;
        RECT 277.950 183.600 280.050 184.200 ;
        RECT 286.950 183.600 289.050 184.050 ;
        RECT 277.950 182.400 289.050 183.600 ;
        RECT 277.950 182.100 280.050 182.400 ;
        RECT 286.950 181.950 289.050 182.400 ;
        RECT 301.950 183.600 306.000 184.050 ;
        RECT 301.950 181.950 306.600 183.600 ;
        RECT 325.800 183.000 327.900 184.050 ;
        RECT 328.950 183.600 331.050 184.200 ;
        RECT 331.950 183.600 334.050 184.950 ;
        RECT 328.950 183.000 334.050 183.600 ;
        RECT 343.950 183.600 346.050 184.050 ;
        RECT 355.950 183.600 358.050 184.200 ;
        RECT 325.800 181.950 328.050 183.000 ;
        RECT 328.950 182.400 333.450 183.000 ;
        RECT 343.950 182.400 358.050 183.600 ;
        RECT 328.950 182.100 331.050 182.400 ;
        RECT 343.950 181.950 346.050 182.400 ;
        RECT 355.950 182.100 358.050 182.400 ;
        RECT 241.950 180.600 244.050 181.050 ;
        RECT 221.400 180.000 244.050 180.600 ;
        RECT 220.950 179.400 244.050 180.000 ;
        RECT 196.950 175.950 199.050 178.050 ;
        RECT 205.950 177.450 208.050 177.900 ;
        RECT 211.950 177.450 214.050 177.900 ;
        RECT 205.950 176.250 214.050 177.450 ;
        RECT 205.950 175.800 208.050 176.250 ;
        RECT 211.950 175.800 214.050 176.250 ;
        RECT 220.950 175.950 223.050 179.400 ;
        RECT 241.950 178.950 244.050 179.400 ;
        RECT 305.400 178.050 306.600 181.950 ;
        RECT 325.950 180.600 328.050 181.950 ;
        RECT 325.950 180.000 333.600 180.600 ;
        RECT 326.400 179.400 333.600 180.000 ;
        RECT 268.950 177.450 271.050 177.900 ;
        RECT 274.950 177.450 277.050 177.900 ;
        RECT 268.950 176.250 277.050 177.450 ;
        RECT 268.950 175.800 271.050 176.250 ;
        RECT 274.950 175.800 277.050 176.250 ;
        RECT 304.950 175.950 307.050 178.050 ;
        RECT 332.400 177.900 333.600 179.400 ;
        RECT 359.400 177.900 360.600 184.950 ;
        RECT 382.950 183.600 385.050 184.200 ;
        RECT 365.400 182.400 385.050 183.600 ;
        RECT 365.400 177.900 366.600 182.400 ;
        RECT 382.950 182.100 385.050 182.400 ;
        RECT 394.950 183.600 397.050 184.050 ;
        RECT 409.950 183.600 412.050 184.050 ;
        RECT 394.950 182.400 412.050 183.600 ;
        RECT 394.950 181.950 397.050 182.400 ;
        RECT 409.950 181.950 412.050 182.400 ;
        RECT 421.950 182.100 424.050 184.200 ;
        RECT 436.950 183.750 439.050 184.200 ;
        RECT 460.950 183.750 463.050 184.200 ;
        RECT 436.950 182.550 463.050 183.750 ;
        RECT 436.950 182.100 439.050 182.550 ;
        RECT 460.950 182.100 463.050 182.550 ;
        RECT 422.400 178.050 423.600 182.100 ;
        RECT 316.950 177.450 319.050 177.900 ;
        RECT 322.950 177.450 325.050 177.900 ;
        RECT 316.950 176.250 325.050 177.450 ;
        RECT 316.950 175.800 319.050 176.250 ;
        RECT 322.950 175.800 325.050 176.250 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 337.950 177.450 340.050 177.900 ;
        RECT 343.950 177.450 346.050 177.900 ;
        RECT 337.950 176.250 346.050 177.450 ;
        RECT 337.950 175.800 340.050 176.250 ;
        RECT 343.950 175.800 346.050 176.250 ;
        RECT 358.950 175.800 361.050 177.900 ;
        RECT 364.950 175.800 367.050 177.900 ;
        RECT 418.950 176.400 423.600 178.050 ;
        RECT 464.400 177.900 465.600 184.950 ;
        RECT 466.950 183.600 469.050 184.200 ;
        RECT 466.950 182.400 471.600 183.600 ;
        RECT 466.950 182.100 469.050 182.400 ;
        RECT 470.400 178.050 471.600 182.400 ;
        RECT 473.400 180.600 474.600 185.400 ;
        RECT 481.950 184.950 484.050 185.400 ;
        RECT 511.950 186.600 514.050 187.050 ;
        RECT 523.950 186.600 526.050 187.050 ;
        RECT 529.950 186.600 532.050 187.050 ;
        RECT 511.950 185.400 532.050 186.600 ;
        RECT 511.950 184.950 514.050 185.400 ;
        RECT 523.950 184.950 526.050 185.400 ;
        RECT 529.950 184.950 532.050 185.400 ;
        RECT 634.950 186.600 637.050 187.050 ;
        RECT 676.950 186.600 679.050 187.050 ;
        RECT 634.950 185.400 679.050 186.600 ;
        RECT 634.950 184.950 637.050 185.400 ;
        RECT 478.950 181.950 481.050 184.050 ;
        RECT 502.950 183.600 505.050 184.050 ;
        RECT 508.950 183.600 511.050 184.200 ;
        RECT 502.950 182.400 511.050 183.600 ;
        RECT 502.950 181.950 505.050 182.400 ;
        RECT 508.950 182.100 511.050 182.400 ;
        RECT 473.400 179.400 477.600 180.600 ;
        RECT 430.950 177.450 433.050 177.900 ;
        RECT 436.950 177.600 439.050 177.900 ;
        RECT 445.950 177.600 448.050 177.900 ;
        RECT 436.950 177.450 448.050 177.600 ;
        RECT 430.950 176.400 448.050 177.450 ;
        RECT 418.950 175.950 423.000 176.400 ;
        RECT 430.950 176.250 439.050 176.400 ;
        RECT 430.950 175.800 433.050 176.250 ;
        RECT 436.950 175.800 439.050 176.250 ;
        RECT 445.950 175.800 448.050 176.400 ;
        RECT 463.950 175.800 466.050 177.900 ;
        RECT 469.950 175.950 472.050 178.050 ;
        RECT 476.400 175.050 477.600 179.400 ;
        RECT 479.400 177.600 480.600 181.950 ;
        RECT 499.950 180.600 502.050 181.050 ;
        RECT 488.400 179.400 502.050 180.600 ;
        RECT 520.950 180.600 523.050 184.050 ;
        RECT 571.950 183.600 574.050 184.200 ;
        RECT 560.400 182.400 574.050 183.600 ;
        RECT 520.950 180.000 528.600 180.600 ;
        RECT 521.400 179.400 528.600 180.000 ;
        RECT 488.400 177.900 489.600 179.400 ;
        RECT 499.950 178.950 502.050 179.400 ;
        RECT 481.950 177.600 484.050 177.900 ;
        RECT 479.400 176.400 484.050 177.600 ;
        RECT 481.950 175.800 484.050 176.400 ;
        RECT 487.950 175.800 490.050 177.900 ;
        RECT 511.950 177.450 514.050 177.900 ;
        RECT 523.950 177.450 526.050 177.900 ;
        RECT 511.950 176.250 526.050 177.450 ;
        RECT 527.400 177.600 528.600 179.400 ;
        RECT 532.950 177.600 535.050 177.900 ;
        RECT 527.400 176.400 535.050 177.600 ;
        RECT 511.950 175.800 514.050 176.250 ;
        RECT 523.950 175.800 526.050 176.250 ;
        RECT 532.950 175.800 535.050 176.400 ;
        RECT 538.950 177.450 541.050 177.900 ;
        RECT 544.950 177.450 547.050 177.900 ;
        RECT 538.950 176.250 547.050 177.450 ;
        RECT 538.950 175.800 541.050 176.250 ;
        RECT 544.950 175.800 547.050 176.250 ;
        RECT 553.950 177.600 556.050 177.900 ;
        RECT 560.400 177.600 561.600 182.400 ;
        RECT 571.950 182.100 574.050 182.400 ;
        RECT 577.950 183.600 580.050 184.200 ;
        RECT 598.950 183.600 601.050 184.200 ;
        RECT 607.950 183.600 610.050 184.050 ;
        RECT 577.950 182.400 591.600 183.600 ;
        RECT 577.950 182.100 580.050 182.400 ;
        RECT 590.400 177.900 591.600 182.400 ;
        RECT 598.950 182.400 610.050 183.600 ;
        RECT 598.950 182.100 601.050 182.400 ;
        RECT 607.950 181.950 610.050 182.400 ;
        RECT 622.950 183.600 625.050 184.200 ;
        RECT 631.950 183.600 634.050 184.050 ;
        RECT 622.950 182.400 634.050 183.600 ;
        RECT 622.950 182.100 625.050 182.400 ;
        RECT 631.950 181.950 634.050 182.400 ;
        RECT 640.950 183.600 643.050 184.200 ;
        RECT 640.950 182.400 660.600 183.600 ;
        RECT 640.950 182.100 643.050 182.400 ;
        RECT 659.400 177.900 660.600 182.400 ;
        RECT 665.400 177.900 666.600 185.400 ;
        RECT 676.950 184.950 679.050 185.400 ;
        RECT 673.950 181.950 676.050 184.050 ;
        RECT 700.950 183.600 703.050 184.200 ;
        RECT 706.950 184.050 709.050 184.500 ;
        RECT 715.950 184.050 718.050 184.500 ;
        RECT 706.950 183.600 718.050 184.050 ;
        RECT 700.950 182.850 718.050 183.600 ;
        RECT 700.950 182.400 709.050 182.850 ;
        RECT 715.950 182.400 718.050 182.850 ;
        RECT 700.950 182.100 703.050 182.400 ;
        RECT 721.950 181.950 724.050 184.050 ;
        RECT 757.950 183.600 760.050 184.050 ;
        RECT 796.800 183.600 798.900 184.200 ;
        RECT 757.950 182.400 798.900 183.600 ;
        RECT 757.950 181.950 760.050 182.400 ;
        RECT 796.800 182.100 798.900 182.400 ;
        RECT 799.950 183.600 802.050 184.050 ;
        RECT 805.950 183.600 808.050 184.050 ;
        RECT 799.950 182.400 808.050 183.600 ;
        RECT 799.950 181.950 802.050 182.400 ;
        RECT 805.950 181.950 808.050 182.400 ;
        RECT 553.950 176.400 561.600 177.600 ;
        RECT 553.950 175.800 556.050 176.400 ;
        RECT 589.950 175.800 592.050 177.900 ;
        RECT 595.950 177.450 598.050 177.900 ;
        RECT 604.950 177.450 607.050 177.900 ;
        RECT 595.950 176.250 607.050 177.450 ;
        RECT 595.950 175.800 598.050 176.250 ;
        RECT 604.950 175.800 607.050 176.250 ;
        RECT 658.950 175.800 661.050 177.900 ;
        RECT 664.950 175.800 667.050 177.900 ;
        RECT 674.400 177.600 675.600 181.950 ;
        RECT 722.400 178.050 723.600 181.950 ;
        RECT 817.950 180.600 820.050 184.050 ;
        RECT 826.950 183.750 829.050 184.200 ;
        RECT 832.950 183.750 835.050 184.200 ;
        RECT 826.950 182.550 835.050 183.750 ;
        RECT 826.950 182.100 829.050 182.550 ;
        RECT 832.950 182.100 835.050 182.550 ;
        RECT 853.950 183.600 856.050 184.050 ;
        RECT 898.950 183.600 901.050 184.050 ;
        RECT 853.950 182.400 861.600 183.600 ;
        RECT 853.950 181.950 856.050 182.400 ;
        RECT 841.950 180.600 844.050 181.200 ;
        RECT 817.950 180.000 844.050 180.600 ;
        RECT 818.400 179.400 844.050 180.000 ;
        RECT 841.950 179.100 844.050 179.400 ;
        RECT 850.950 180.750 853.050 181.200 ;
        RECT 856.950 180.750 859.050 181.200 ;
        RECT 850.950 179.550 859.050 180.750 ;
        RECT 850.950 179.100 853.050 179.550 ;
        RECT 856.950 179.100 859.050 179.550 ;
        RECT 860.400 180.600 861.600 182.400 ;
        RECT 890.400 182.400 901.050 183.600 ;
        RECT 880.950 180.600 883.050 180.900 ;
        RECT 860.400 179.400 883.050 180.600 ;
        RECT 679.950 177.600 682.050 177.900 ;
        RECT 674.400 176.400 682.050 177.600 ;
        RECT 679.950 175.800 682.050 176.400 ;
        RECT 721.950 175.950 724.050 178.050 ;
        RECT 751.950 177.600 754.050 177.900 ;
        RECT 733.950 176.400 754.050 177.600 ;
        RECT 733.950 175.500 736.050 176.400 ;
        RECT 751.950 175.800 754.050 176.400 ;
        RECT 769.950 177.600 772.050 178.050 ;
        RECT 805.950 177.600 808.050 178.050 ;
        RECT 769.950 176.400 808.050 177.600 ;
        RECT 769.950 175.950 772.050 176.400 ;
        RECT 805.950 175.950 808.050 176.400 ;
        RECT 814.950 177.600 817.050 177.900 ;
        RECT 820.950 177.600 823.050 178.050 ;
        RECT 814.950 176.400 823.050 177.600 ;
        RECT 814.950 175.800 817.050 176.400 ;
        RECT 820.950 175.950 823.050 176.400 ;
        RECT 829.950 177.600 832.050 177.900 ;
        RECT 842.400 177.600 843.600 179.100 ;
        RECT 880.950 178.800 883.050 179.400 ;
        RECT 829.950 176.400 843.600 177.600 ;
        RECT 829.950 175.800 832.050 176.400 ;
        RECT 139.950 174.600 142.050 175.050 ;
        RECT 151.950 174.600 154.050 175.050 ;
        RECT 139.950 173.400 154.050 174.600 ;
        RECT 139.950 172.950 142.050 173.400 ;
        RECT 151.950 172.950 154.050 173.400 ;
        RECT 157.950 174.600 160.050 175.050 ;
        RECT 172.950 174.600 175.050 175.050 ;
        RECT 157.950 173.400 175.050 174.600 ;
        RECT 157.950 172.950 160.050 173.400 ;
        RECT 172.950 172.950 175.050 173.400 ;
        RECT 202.950 174.600 205.050 175.050 ;
        RECT 217.950 174.600 220.050 175.050 ;
        RECT 202.950 173.400 220.050 174.600 ;
        RECT 202.950 172.950 205.050 173.400 ;
        RECT 217.950 172.950 220.050 173.400 ;
        RECT 310.950 174.600 313.050 175.050 ;
        RECT 346.950 174.600 349.050 175.050 ;
        RECT 379.950 174.600 382.050 175.050 ;
        RECT 310.950 173.400 382.050 174.600 ;
        RECT 310.950 172.950 313.050 173.400 ;
        RECT 346.950 172.950 349.050 173.400 ;
        RECT 379.950 172.950 382.050 173.400 ;
        RECT 385.950 174.600 388.050 175.050 ;
        RECT 412.950 174.600 415.050 175.050 ;
        RECT 385.950 173.400 415.050 174.600 ;
        RECT 385.950 172.950 388.050 173.400 ;
        RECT 412.950 172.950 415.050 173.400 ;
        RECT 424.950 174.600 427.050 175.050 ;
        RECT 451.950 174.600 454.050 175.050 ;
        RECT 424.950 173.400 454.050 174.600 ;
        RECT 476.400 173.400 481.050 175.050 ;
        RECT 424.950 172.950 427.050 173.400 ;
        RECT 451.950 172.950 454.050 173.400 ;
        RECT 477.000 172.950 481.050 173.400 ;
        RECT 559.950 174.600 562.050 175.050 ;
        RECT 574.950 174.600 577.050 175.050 ;
        RECT 559.950 173.400 577.050 174.600 ;
        RECT 559.950 172.950 562.050 173.400 ;
        RECT 574.950 172.950 577.050 173.400 ;
        RECT 589.950 174.600 592.050 175.050 ;
        RECT 619.950 174.600 622.050 175.050 ;
        RECT 589.950 173.400 622.050 174.600 ;
        RECT 589.950 172.950 592.050 173.400 ;
        RECT 619.950 172.950 622.050 173.400 ;
        RECT 742.950 174.600 745.050 175.050 ;
        RECT 787.950 174.600 790.050 175.050 ;
        RECT 742.950 173.400 790.050 174.600 ;
        RECT 742.950 172.950 745.050 173.400 ;
        RECT 787.950 172.950 790.050 173.400 ;
        RECT 793.950 174.600 796.050 175.050 ;
        RECT 826.950 174.600 829.050 175.050 ;
        RECT 858.000 174.600 862.050 175.050 ;
        RECT 793.950 173.400 829.050 174.600 ;
        RECT 857.400 174.000 862.050 174.600 ;
        RECT 793.950 172.950 796.050 173.400 ;
        RECT 826.950 172.950 829.050 173.400 ;
        RECT 856.950 172.950 862.050 174.000 ;
        RECT 58.950 171.600 61.050 172.050 ;
        RECT 82.950 171.600 85.050 172.050 ;
        RECT 58.950 170.400 85.050 171.600 ;
        RECT 58.950 169.950 61.050 170.400 ;
        RECT 82.950 169.950 85.050 170.400 ;
        RECT 97.950 171.600 100.050 172.050 ;
        RECT 130.950 171.600 133.050 172.050 ;
        RECT 97.950 170.400 133.050 171.600 ;
        RECT 97.950 169.950 100.050 170.400 ;
        RECT 130.950 169.950 133.050 170.400 ;
        RECT 517.950 171.600 520.050 172.050 ;
        RECT 553.950 171.600 556.050 172.050 ;
        RECT 517.950 170.400 556.050 171.600 ;
        RECT 517.950 169.950 520.050 170.400 ;
        RECT 553.950 169.950 556.050 170.400 ;
        RECT 592.950 171.600 595.050 172.050 ;
        RECT 613.950 171.600 616.050 172.050 ;
        RECT 592.950 170.400 616.050 171.600 ;
        RECT 592.950 169.950 595.050 170.400 ;
        RECT 613.950 169.950 616.050 170.400 ;
        RECT 628.950 171.600 631.050 172.050 ;
        RECT 664.950 171.600 667.050 172.050 ;
        RECT 628.950 170.400 667.050 171.600 ;
        RECT 628.950 169.950 631.050 170.400 ;
        RECT 664.950 169.950 667.050 170.400 ;
        RECT 718.950 171.600 721.050 172.050 ;
        RECT 790.950 171.600 793.050 172.050 ;
        RECT 718.950 170.400 793.050 171.600 ;
        RECT 718.950 169.950 721.050 170.400 ;
        RECT 790.950 169.950 793.050 170.400 ;
        RECT 856.950 169.950 859.050 172.950 ;
        RECT 190.950 168.600 193.050 169.050 ;
        RECT 220.950 168.600 223.050 169.050 ;
        RECT 190.950 167.400 223.050 168.600 ;
        RECT 190.950 166.950 193.050 167.400 ;
        RECT 220.950 166.950 223.050 167.400 ;
        RECT 649.950 168.600 652.050 169.050 ;
        RECT 667.800 168.600 669.900 169.050 ;
        RECT 649.950 167.400 669.900 168.600 ;
        RECT 649.950 166.950 652.050 167.400 ;
        RECT 667.800 166.950 669.900 167.400 ;
        RECT 670.950 168.600 673.050 169.050 ;
        RECT 700.800 168.600 702.900 169.050 ;
        RECT 670.950 167.400 702.900 168.600 ;
        RECT 670.950 166.950 673.050 167.400 ;
        RECT 700.800 166.950 702.900 167.400 ;
        RECT 802.950 168.600 805.050 169.050 ;
        RECT 826.950 168.600 829.050 169.050 ;
        RECT 802.950 167.400 829.050 168.600 ;
        RECT 802.950 166.950 805.050 167.400 ;
        RECT 826.950 166.950 829.050 167.400 ;
        RECT 211.950 165.600 214.050 166.050 ;
        RECT 226.950 165.600 229.050 166.050 ;
        RECT 211.950 164.400 229.050 165.600 ;
        RECT 211.950 163.950 214.050 164.400 ;
        RECT 226.950 163.950 229.050 164.400 ;
        RECT 277.950 165.600 280.050 166.050 ;
        RECT 349.950 165.600 352.050 166.050 ;
        RECT 838.950 165.600 841.050 166.050 ;
        RECT 277.950 164.400 352.050 165.600 ;
        RECT 277.950 163.950 280.050 164.400 ;
        RECT 349.950 163.950 352.050 164.400 ;
        RECT 764.400 164.400 841.050 165.600 ;
        RECT 64.950 162.600 67.050 163.050 ;
        RECT 124.950 162.600 127.050 163.050 ;
        RECT 64.950 161.400 127.050 162.600 ;
        RECT 64.950 160.950 67.050 161.400 ;
        RECT 124.950 160.950 127.050 161.400 ;
        RECT 166.950 162.600 169.050 163.050 ;
        RECT 190.950 162.600 193.050 163.050 ;
        RECT 166.950 161.400 193.050 162.600 ;
        RECT 166.950 160.950 169.050 161.400 ;
        RECT 190.950 160.950 193.050 161.400 ;
        RECT 241.950 162.600 244.050 163.050 ;
        RECT 286.950 162.600 289.050 163.050 ;
        RECT 241.950 161.400 289.050 162.600 ;
        RECT 241.950 160.950 244.050 161.400 ;
        RECT 286.950 160.950 289.050 161.400 ;
        RECT 304.950 162.600 307.050 163.050 ;
        RECT 349.950 162.600 352.050 162.900 ;
        RECT 304.950 161.400 352.050 162.600 ;
        RECT 304.950 160.950 307.050 161.400 ;
        RECT 349.950 160.800 352.050 161.400 ;
        RECT 592.950 162.600 595.050 163.050 ;
        RECT 643.950 162.600 646.050 163.050 ;
        RECT 592.950 161.400 646.050 162.600 ;
        RECT 592.950 160.950 595.050 161.400 ;
        RECT 643.950 160.950 646.050 161.400 ;
        RECT 712.950 162.600 715.050 163.050 ;
        RECT 764.400 162.600 765.600 164.400 ;
        RECT 838.950 163.950 841.050 164.400 ;
        RECT 890.400 163.050 891.600 182.400 ;
        RECT 898.950 181.950 901.050 182.400 ;
        RECT 907.950 183.600 910.050 184.050 ;
        RECT 907.950 182.400 918.600 183.600 ;
        RECT 907.950 181.950 910.050 182.400 ;
        RECT 901.950 180.600 904.050 181.050 ;
        RECT 901.950 179.400 915.600 180.600 ;
        RECT 901.950 178.950 904.050 179.400 ;
        RECT 914.400 175.050 915.600 179.400 ;
        RECT 913.950 172.950 916.050 175.050 ;
        RECT 917.400 171.600 918.600 182.400 ;
        RECT 917.400 170.400 924.600 171.600 ;
        RECT 907.950 168.600 910.050 169.050 ;
        RECT 919.950 168.600 922.050 169.050 ;
        RECT 907.950 167.400 922.050 168.600 ;
        RECT 907.950 166.950 910.050 167.400 ;
        RECT 919.950 166.950 922.050 167.400 ;
        RECT 923.400 163.050 924.600 170.400 ;
        RECT 712.950 161.400 765.600 162.600 ;
        RECT 712.950 160.950 715.050 161.400 ;
        RECT 889.950 160.950 892.050 163.050 ;
        RECT 919.950 161.400 924.600 163.050 ;
        RECT 919.950 160.950 924.000 161.400 ;
        RECT 13.950 159.600 16.050 160.050 ;
        RECT 58.950 159.600 61.050 160.050 ;
        RECT 13.950 158.400 61.050 159.600 ;
        RECT 13.950 157.950 16.050 158.400 ;
        RECT 58.950 157.950 61.050 158.400 ;
        RECT 376.950 159.600 379.050 160.050 ;
        RECT 394.950 159.600 397.050 160.050 ;
        RECT 400.950 159.600 403.050 160.050 ;
        RECT 376.950 158.400 403.050 159.600 ;
        RECT 376.950 157.950 379.050 158.400 ;
        RECT 394.950 157.950 397.050 158.400 ;
        RECT 400.950 157.950 403.050 158.400 ;
        RECT 649.950 159.600 652.050 160.050 ;
        RECT 682.950 159.600 685.050 160.050 ;
        RECT 649.950 158.400 685.050 159.600 ;
        RECT 649.950 157.950 652.050 158.400 ;
        RECT 682.950 157.950 685.050 158.400 ;
        RECT 742.950 159.600 745.050 160.050 ;
        RECT 748.950 159.600 751.050 160.050 ;
        RECT 742.950 158.400 751.050 159.600 ;
        RECT 742.950 157.950 745.050 158.400 ;
        RECT 748.950 157.950 751.050 158.400 ;
        RECT 145.950 156.600 148.050 157.050 ;
        RECT 199.950 156.600 202.050 157.050 ;
        RECT 145.950 155.400 202.050 156.600 ;
        RECT 145.950 154.950 148.050 155.400 ;
        RECT 199.950 154.950 202.050 155.400 ;
        RECT 286.950 156.600 289.050 157.050 ;
        RECT 313.950 156.600 316.050 157.050 ;
        RECT 286.950 155.400 316.050 156.600 ;
        RECT 286.950 154.950 289.050 155.400 ;
        RECT 313.950 154.950 316.050 155.400 ;
        RECT 352.950 156.600 355.050 157.050 ;
        RECT 433.950 156.600 436.050 157.050 ;
        RECT 352.950 155.400 436.050 156.600 ;
        RECT 352.950 154.950 355.050 155.400 ;
        RECT 433.950 154.950 436.050 155.400 ;
        RECT 472.950 156.600 475.050 157.050 ;
        RECT 538.950 156.600 541.050 157.050 ;
        RECT 562.950 156.600 565.050 157.050 ;
        RECT 472.950 155.400 565.050 156.600 ;
        RECT 472.950 154.950 475.050 155.400 ;
        RECT 538.950 154.950 541.050 155.400 ;
        RECT 562.950 154.950 565.050 155.400 ;
        RECT 688.950 156.600 691.050 157.050 ;
        RECT 781.950 156.600 784.050 157.050 ;
        RECT 817.950 156.600 820.050 157.050 ;
        RECT 688.950 155.400 820.050 156.600 ;
        RECT 688.950 154.950 691.050 155.400 ;
        RECT 781.950 154.950 784.050 155.400 ;
        RECT 817.950 154.950 820.050 155.400 ;
        RECT 823.950 156.600 826.050 157.050 ;
        RECT 904.950 156.600 907.050 157.050 ;
        RECT 823.950 155.400 907.050 156.600 ;
        RECT 823.950 154.950 826.050 155.400 ;
        RECT 904.950 154.950 907.050 155.400 ;
        RECT 4.950 153.600 7.050 154.050 ;
        RECT 61.950 153.600 64.050 154.050 ;
        RECT 4.950 152.400 64.050 153.600 ;
        RECT 4.950 151.950 7.050 152.400 ;
        RECT 61.950 151.950 64.050 152.400 ;
        RECT 244.950 153.600 247.050 154.050 ;
        RECT 253.950 153.600 256.050 154.050 ;
        RECT 367.950 153.600 370.050 154.050 ;
        RECT 418.950 153.600 421.050 154.050 ;
        RECT 244.950 152.400 256.050 153.600 ;
        RECT 244.950 151.950 247.050 152.400 ;
        RECT 253.950 151.950 256.050 152.400 ;
        RECT 326.400 152.400 370.050 153.600 ;
        RECT 7.950 150.600 10.050 151.050 ;
        RECT 22.950 150.600 25.050 151.050 ;
        RECT 46.950 150.600 49.050 151.050 ;
        RECT 7.950 149.400 49.050 150.600 ;
        RECT 7.950 148.950 10.050 149.400 ;
        RECT 22.950 148.950 25.050 149.400 ;
        RECT 46.950 148.950 49.050 149.400 ;
        RECT 148.950 150.600 151.050 151.050 ;
        RECT 157.950 150.600 160.050 151.050 ;
        RECT 178.950 150.600 181.050 151.050 ;
        RECT 148.950 149.400 181.050 150.600 ;
        RECT 148.950 148.950 151.050 149.400 ;
        RECT 157.950 148.950 160.050 149.400 ;
        RECT 178.950 148.950 181.050 149.400 ;
        RECT 256.950 150.600 259.050 151.050 ;
        RECT 310.950 150.600 313.050 151.050 ;
        RECT 326.400 150.600 327.600 152.400 ;
        RECT 367.950 151.950 370.050 152.400 ;
        RECT 380.400 152.400 421.050 153.600 ;
        RECT 256.950 149.400 327.600 150.600 ;
        RECT 328.950 150.600 331.050 151.050 ;
        RECT 380.400 150.600 381.600 152.400 ;
        RECT 418.950 151.950 421.050 152.400 ;
        RECT 643.950 153.600 646.050 154.050 ;
        RECT 673.950 153.600 676.050 154.050 ;
        RECT 643.950 152.400 676.050 153.600 ;
        RECT 643.950 151.950 646.050 152.400 ;
        RECT 673.950 151.950 676.050 152.400 ;
        RECT 328.950 149.400 381.600 150.600 ;
        RECT 469.950 150.600 472.050 151.050 ;
        RECT 532.950 150.600 535.050 151.050 ;
        RECT 550.950 150.600 553.050 151.050 ;
        RECT 469.950 149.400 553.050 150.600 ;
        RECT 256.950 148.950 259.050 149.400 ;
        RECT 310.950 148.950 313.050 149.400 ;
        RECT 328.950 148.950 331.050 149.400 ;
        RECT 469.950 148.950 472.050 149.400 ;
        RECT 532.950 148.950 535.050 149.400 ;
        RECT 550.950 148.950 553.050 149.400 ;
        RECT 691.950 150.600 694.050 151.050 ;
        RECT 724.950 150.600 727.050 151.050 ;
        RECT 691.950 149.400 727.050 150.600 ;
        RECT 691.950 148.950 694.050 149.400 ;
        RECT 724.950 148.950 727.050 149.400 ;
        RECT 742.950 150.600 745.050 151.050 ;
        RECT 763.950 150.600 766.050 151.050 ;
        RECT 808.950 150.600 811.050 151.050 ;
        RECT 742.950 149.400 762.600 150.600 ;
        RECT 742.950 148.950 745.050 149.400 ;
        RECT 160.950 147.600 163.050 148.050 ;
        RECT 184.950 147.600 187.050 148.050 ;
        RECT 160.950 146.400 187.050 147.600 ;
        RECT 160.950 145.950 163.050 146.400 ;
        RECT 184.950 145.950 187.050 146.400 ;
        RECT 205.950 147.600 208.050 148.050 ;
        RECT 235.950 147.600 238.050 148.050 ;
        RECT 283.950 147.600 286.050 148.050 ;
        RECT 205.950 146.400 238.050 147.600 ;
        RECT 205.950 145.950 208.050 146.400 ;
        RECT 235.950 145.950 238.050 146.400 ;
        RECT 263.400 146.400 286.050 147.600 ;
        RECT 263.400 145.050 264.600 146.400 ;
        RECT 283.950 145.950 286.050 146.400 ;
        RECT 322.950 147.600 325.050 148.050 ;
        RECT 382.950 147.600 385.050 148.050 ;
        RECT 322.950 146.400 385.050 147.600 ;
        RECT 322.950 145.950 325.050 146.400 ;
        RECT 382.950 145.950 385.050 146.400 ;
        RECT 403.950 147.600 406.050 148.050 ;
        RECT 424.950 147.600 427.050 148.050 ;
        RECT 457.950 147.600 460.050 148.050 ;
        RECT 574.950 147.600 577.050 148.050 ;
        RECT 403.950 146.400 577.050 147.600 ;
        RECT 403.950 145.950 406.050 146.400 ;
        RECT 424.950 145.950 427.050 146.400 ;
        RECT 457.950 145.950 460.050 146.400 ;
        RECT 574.950 145.950 577.050 146.400 ;
        RECT 631.950 147.600 634.050 148.050 ;
        RECT 655.950 147.600 658.050 148.050 ;
        RECT 631.950 146.400 658.050 147.600 ;
        RECT 631.950 145.950 634.050 146.400 ;
        RECT 655.950 145.950 658.050 146.400 ;
        RECT 715.950 147.600 718.050 148.050 ;
        RECT 739.950 147.600 742.050 148.050 ;
        RECT 715.950 146.400 742.050 147.600 ;
        RECT 761.400 147.600 762.600 149.400 ;
        RECT 763.950 149.400 811.050 150.600 ;
        RECT 763.950 148.950 766.050 149.400 ;
        RECT 808.950 148.950 811.050 149.400 ;
        RECT 814.950 150.600 817.050 151.050 ;
        RECT 823.950 150.600 826.050 151.050 ;
        RECT 814.950 149.400 826.050 150.600 ;
        RECT 814.950 148.950 817.050 149.400 ;
        RECT 823.950 148.950 826.050 149.400 ;
        RECT 856.950 150.600 859.050 151.050 ;
        RECT 871.950 150.600 874.050 151.050 ;
        RECT 856.950 149.400 874.050 150.600 ;
        RECT 856.950 148.950 859.050 149.400 ;
        RECT 871.950 148.950 874.050 149.400 ;
        RECT 772.950 147.600 775.050 148.050 ;
        RECT 761.400 146.400 775.050 147.600 ;
        RECT 715.950 145.950 718.050 146.400 ;
        RECT 739.950 145.950 742.050 146.400 ;
        RECT 772.950 145.950 775.050 146.400 ;
        RECT 37.950 144.600 40.050 145.050 ;
        RECT 115.950 144.600 118.050 145.050 ;
        RECT 37.950 143.400 118.050 144.600 ;
        RECT 37.950 142.950 40.050 143.400 ;
        RECT 115.950 142.950 118.050 143.400 ;
        RECT 193.950 144.600 196.050 145.050 ;
        RECT 199.950 144.600 202.050 145.050 ;
        RECT 193.950 143.400 202.050 144.600 ;
        RECT 193.950 142.950 196.050 143.400 ;
        RECT 199.950 142.950 202.050 143.400 ;
        RECT 244.950 144.600 247.050 145.050 ;
        RECT 262.950 144.600 265.050 145.050 ;
        RECT 244.950 143.400 265.050 144.600 ;
        RECT 244.950 142.950 247.050 143.400 ;
        RECT 262.950 142.950 265.050 143.400 ;
        RECT 298.950 144.600 301.050 145.050 ;
        RECT 319.950 144.600 322.050 145.050 ;
        RECT 298.950 143.400 322.050 144.600 ;
        RECT 298.950 142.950 301.050 143.400 ;
        RECT 319.950 142.950 322.050 143.400 ;
        RECT 325.950 144.600 328.050 145.050 ;
        RECT 367.950 144.600 370.050 145.050 ;
        RECT 379.950 144.600 382.050 145.050 ;
        RECT 325.950 143.400 382.050 144.600 ;
        RECT 325.950 142.950 328.050 143.400 ;
        RECT 367.950 142.950 370.050 143.400 ;
        RECT 379.950 142.950 382.050 143.400 ;
        RECT 433.950 144.600 436.050 145.050 ;
        RECT 448.950 144.600 451.050 145.050 ;
        RECT 433.950 143.400 451.050 144.600 ;
        RECT 433.950 142.950 436.050 143.400 ;
        RECT 448.950 142.950 451.050 143.400 ;
        RECT 466.950 144.600 469.050 145.050 ;
        RECT 604.950 144.600 607.050 145.050 ;
        RECT 466.950 143.400 607.050 144.600 ;
        RECT 466.950 142.950 469.050 143.400 ;
        RECT 604.950 142.950 607.050 143.400 ;
        RECT 637.950 144.600 640.050 145.050 ;
        RECT 649.950 144.600 652.050 145.050 ;
        RECT 637.950 143.400 652.050 144.600 ;
        RECT 637.950 142.950 640.050 143.400 ;
        RECT 649.950 142.950 652.050 143.400 ;
        RECT 700.950 144.600 703.050 145.050 ;
        RECT 706.950 144.600 709.050 145.050 ;
        RECT 700.950 143.400 709.050 144.600 ;
        RECT 700.950 142.950 703.050 143.400 ;
        RECT 706.950 142.950 709.050 143.400 ;
        RECT 742.950 144.600 745.050 145.050 ;
        RECT 778.950 144.600 781.050 145.050 ;
        RECT 742.950 143.400 781.050 144.600 ;
        RECT 742.950 142.950 745.050 143.400 ;
        RECT 778.950 142.950 781.050 143.400 ;
        RECT 856.950 144.600 859.050 145.050 ;
        RECT 877.950 144.600 880.050 145.050 ;
        RECT 856.950 143.400 880.050 144.600 ;
        RECT 856.950 142.950 859.050 143.400 ;
        RECT 877.950 142.950 880.050 143.400 ;
        RECT 10.950 141.600 13.050 142.050 ;
        RECT 31.950 141.600 34.050 142.050 ;
        RECT 10.950 140.400 34.050 141.600 ;
        RECT 10.950 139.950 13.050 140.400 ;
        RECT 31.950 139.950 34.050 140.400 ;
        RECT 58.950 141.600 61.050 142.050 ;
        RECT 94.950 141.600 97.050 142.050 ;
        RECT 58.950 140.400 97.050 141.600 ;
        RECT 58.950 139.950 61.050 140.400 ;
        RECT 94.950 139.950 97.050 140.400 ;
        RECT 127.950 141.600 130.050 142.050 ;
        RECT 154.950 141.600 157.050 142.050 ;
        RECT 163.950 141.600 166.050 142.050 ;
        RECT 172.950 141.600 175.050 142.050 ;
        RECT 127.950 140.400 175.050 141.600 ;
        RECT 127.950 139.950 130.050 140.400 ;
        RECT 154.950 139.950 157.050 140.400 ;
        RECT 163.950 139.950 166.050 140.400 ;
        RECT 172.950 139.950 175.050 140.400 ;
        RECT 235.950 141.600 238.050 142.050 ;
        RECT 247.950 141.600 250.050 142.050 ;
        RECT 289.950 141.600 292.050 142.050 ;
        RECT 235.950 140.400 292.050 141.600 ;
        RECT 235.950 139.950 238.050 140.400 ;
        RECT 247.950 139.950 250.050 140.400 ;
        RECT 289.950 139.950 292.050 140.400 ;
        RECT 487.950 141.600 490.050 142.050 ;
        RECT 502.950 141.600 505.050 142.050 ;
        RECT 487.950 140.400 505.050 141.600 ;
        RECT 487.950 139.950 490.050 140.400 ;
        RECT 502.950 139.950 505.050 140.400 ;
        RECT 547.950 141.600 550.050 142.050 ;
        RECT 556.950 141.600 559.050 142.050 ;
        RECT 622.950 141.600 625.050 142.050 ;
        RECT 547.950 140.400 559.050 141.600 ;
        RECT 547.950 139.950 550.050 140.400 ;
        RECT 556.950 139.950 559.050 140.400 ;
        RECT 578.400 140.400 625.050 141.600 ;
        RECT 27.000 138.600 31.050 139.050 ;
        RECT 26.400 136.950 31.050 138.600 ;
        RECT 55.950 137.100 58.050 139.200 ;
        RECT 103.950 137.100 106.050 139.200 ;
        RECT 133.950 138.600 136.050 139.200 ;
        RECT 151.950 138.600 154.050 139.200 ;
        RECT 133.950 137.400 154.050 138.600 ;
        RECT 133.950 137.100 136.050 137.400 ;
        RECT 151.950 137.100 154.050 137.400 ;
        RECT 199.950 138.750 202.050 139.200 ;
        RECT 205.950 138.750 208.050 139.200 ;
        RECT 199.950 137.550 208.050 138.750 ;
        RECT 199.950 137.100 202.050 137.550 ;
        RECT 205.950 137.100 208.050 137.550 ;
        RECT 229.950 138.600 232.050 139.200 ;
        RECT 244.950 138.600 247.050 139.200 ;
        RECT 229.950 137.400 247.050 138.600 ;
        RECT 229.950 137.100 232.050 137.400 ;
        RECT 244.950 137.100 247.050 137.400 ;
        RECT 256.950 138.750 259.050 139.200 ;
        RECT 262.950 138.750 265.050 139.200 ;
        RECT 256.950 137.550 265.050 138.750 ;
        RECT 256.950 137.100 259.050 137.550 ;
        RECT 262.950 137.100 265.050 137.550 ;
        RECT 304.950 138.750 307.050 139.200 ;
        RECT 334.950 138.750 337.050 139.200 ;
        RECT 304.950 137.550 337.050 138.750 ;
        RECT 304.950 137.100 307.050 137.550 ;
        RECT 334.950 137.100 337.050 137.550 ;
        RECT 26.400 133.050 27.600 136.950 ;
        RECT 56.400 133.050 57.600 137.100 ;
        RECT 25.950 130.950 28.050 133.050 ;
        RECT 34.950 132.450 37.050 132.900 ;
        RECT 46.950 132.450 49.050 132.900 ;
        RECT 34.950 131.250 49.050 132.450 ;
        RECT 34.950 130.800 37.050 131.250 ;
        RECT 46.950 130.800 49.050 131.250 ;
        RECT 52.950 131.400 57.600 133.050 ;
        RECT 70.950 132.450 73.050 132.900 ;
        RECT 79.950 132.450 82.050 132.900 ;
        RECT 52.950 130.950 57.000 131.400 ;
        RECT 70.950 131.250 82.050 132.450 ;
        RECT 70.950 130.800 73.050 131.250 ;
        RECT 79.950 130.800 82.050 131.250 ;
        RECT 85.950 132.600 88.050 132.900 ;
        RECT 104.400 132.600 105.600 137.100 ;
        RECT 343.950 136.950 346.050 139.050 ;
        RECT 358.950 138.600 361.050 139.200 ;
        RECT 364.950 138.600 367.050 139.050 ;
        RECT 358.950 137.400 367.050 138.600 ;
        RECT 358.950 137.100 361.050 137.400 ;
        RECT 364.950 136.950 367.050 137.400 ;
        RECT 382.950 138.600 385.050 139.200 ;
        RECT 442.950 138.600 445.050 139.200 ;
        RECT 466.950 138.600 469.050 139.200 ;
        RECT 382.950 137.400 399.600 138.600 ;
        RECT 382.950 137.100 385.050 137.400 ;
        RECT 85.950 131.400 105.600 132.600 ;
        RECT 115.950 132.600 118.050 133.050 ;
        RECT 124.950 132.600 127.050 132.900 ;
        RECT 115.950 131.400 127.050 132.600 ;
        RECT 85.950 130.800 88.050 131.400 ;
        RECT 115.950 130.950 118.050 131.400 ;
        RECT 124.950 130.800 127.050 131.400 ;
        RECT 139.950 132.450 142.050 132.900 ;
        RECT 169.950 132.450 172.050 132.900 ;
        RECT 139.950 131.250 172.050 132.450 ;
        RECT 139.950 130.800 142.050 131.250 ;
        RECT 169.950 130.800 172.050 131.250 ;
        RECT 184.950 132.450 187.050 132.900 ;
        RECT 196.950 132.450 199.050 132.900 ;
        RECT 184.950 131.250 199.050 132.450 ;
        RECT 184.950 130.800 187.050 131.250 ;
        RECT 196.950 130.800 199.050 131.250 ;
        RECT 226.950 132.450 229.050 132.900 ;
        RECT 235.950 132.450 238.050 132.900 ;
        RECT 226.950 131.250 238.050 132.450 ;
        RECT 226.950 130.800 229.050 131.250 ;
        RECT 235.950 130.800 238.050 131.250 ;
        RECT 247.950 132.600 250.050 132.900 ;
        RECT 253.950 132.600 256.050 132.900 ;
        RECT 247.950 132.450 256.050 132.600 ;
        RECT 259.950 132.450 262.050 132.900 ;
        RECT 247.950 131.400 262.050 132.450 ;
        RECT 247.950 130.800 250.050 131.400 ;
        RECT 253.950 131.250 262.050 131.400 ;
        RECT 253.950 130.800 256.050 131.250 ;
        RECT 259.950 130.800 262.050 131.250 ;
        RECT 274.950 132.450 277.050 132.900 ;
        RECT 286.950 132.450 289.050 132.900 ;
        RECT 274.950 131.250 289.050 132.450 ;
        RECT 274.950 130.800 277.050 131.250 ;
        RECT 286.950 130.800 289.050 131.250 ;
        RECT 292.950 132.450 295.050 132.900 ;
        RECT 298.950 132.450 301.050 132.900 ;
        RECT 292.950 131.250 301.050 132.450 ;
        RECT 292.950 130.800 295.050 131.250 ;
        RECT 298.950 130.800 301.050 131.250 ;
        RECT 313.950 132.450 316.050 132.900 ;
        RECT 322.950 132.450 325.050 132.900 ;
        RECT 313.950 131.250 325.050 132.450 ;
        RECT 344.400 132.600 345.600 136.950 ;
        RECT 355.950 132.600 358.050 132.900 ;
        RECT 344.400 131.400 358.050 132.600 ;
        RECT 313.950 130.800 316.050 131.250 ;
        RECT 322.950 130.800 325.050 131.250 ;
        RECT 355.950 130.800 358.050 131.400 ;
        RECT 367.950 132.600 370.050 133.050 ;
        RECT 398.400 132.900 399.600 137.400 ;
        RECT 442.950 137.400 469.050 138.600 ;
        RECT 442.950 137.100 445.050 137.400 ;
        RECT 466.950 137.100 469.050 137.400 ;
        RECT 496.950 138.750 499.050 139.200 ;
        RECT 508.950 138.750 511.050 139.200 ;
        RECT 496.950 137.550 511.050 138.750 ;
        RECT 562.950 138.600 565.050 139.050 ;
        RECT 496.950 137.100 499.050 137.550 ;
        RECT 508.950 137.100 511.050 137.550 ;
        RECT 554.400 137.400 565.050 138.600 ;
        RECT 544.950 135.600 547.050 136.050 ;
        RECT 536.400 134.400 547.050 135.600 ;
        RECT 536.400 132.900 537.600 134.400 ;
        RECT 544.950 133.950 547.050 134.400 ;
        RECT 554.400 132.900 555.600 137.400 ;
        RECT 562.950 136.950 565.050 137.400 ;
        RECT 578.400 132.900 579.600 140.400 ;
        RECT 622.950 139.950 625.050 140.400 ;
        RECT 745.950 141.600 748.050 142.050 ;
        RECT 757.800 141.600 759.900 141.900 ;
        RECT 745.950 140.400 759.900 141.600 ;
        RECT 745.950 139.950 748.050 140.400 ;
        RECT 757.800 139.800 759.900 140.400 ;
        RECT 760.950 141.600 763.050 142.050 ;
        RECT 766.800 141.600 768.900 142.050 ;
        RECT 760.950 140.400 768.900 141.600 ;
        RECT 760.950 139.950 763.050 140.400 ;
        RECT 766.800 139.950 768.900 140.400 ;
        RECT 580.950 138.600 583.050 139.200 ;
        RECT 598.950 138.600 601.050 139.200 ;
        RECT 580.950 137.400 601.050 138.600 ;
        RECT 580.950 137.100 583.050 137.400 ;
        RECT 598.950 137.100 601.050 137.400 ;
        RECT 607.950 138.750 610.050 139.200 ;
        RECT 616.950 138.750 619.050 139.200 ;
        RECT 607.950 137.550 619.050 138.750 ;
        RECT 607.950 137.100 610.050 137.550 ;
        RECT 616.950 137.100 619.050 137.550 ;
        RECT 628.950 138.600 631.050 139.050 ;
        RECT 643.950 138.600 646.050 139.050 ;
        RECT 628.950 137.400 646.050 138.600 ;
        RECT 628.950 136.950 631.050 137.400 ;
        RECT 643.950 136.950 646.050 137.400 ;
        RECT 655.950 138.600 660.000 139.050 ;
        RECT 673.950 138.600 676.050 139.050 ;
        RECT 694.950 138.750 697.050 139.200 ;
        RECT 700.950 138.750 703.050 139.200 ;
        RECT 655.950 136.950 660.600 138.600 ;
        RECT 673.950 137.400 681.600 138.600 ;
        RECT 673.950 136.950 676.050 137.400 ;
        RECT 379.950 132.600 382.050 132.900 ;
        RECT 367.950 131.400 382.050 132.600 ;
        RECT 367.950 130.950 370.050 131.400 ;
        RECT 379.950 130.800 382.050 131.400 ;
        RECT 397.950 130.800 400.050 132.900 ;
        RECT 412.950 132.450 415.050 132.900 ;
        RECT 439.950 132.450 442.050 132.900 ;
        RECT 412.950 131.250 442.050 132.450 ;
        RECT 412.950 130.800 415.050 131.250 ;
        RECT 439.950 130.800 442.050 131.250 ;
        RECT 457.950 132.450 460.050 132.900 ;
        RECT 463.950 132.450 466.050 132.900 ;
        RECT 457.950 131.250 466.050 132.450 ;
        RECT 457.950 130.800 460.050 131.250 ;
        RECT 463.950 130.800 466.050 131.250 ;
        RECT 475.950 132.450 478.050 132.900 ;
        RECT 490.950 132.450 493.050 132.900 ;
        RECT 475.950 131.250 493.050 132.450 ;
        RECT 475.950 130.800 478.050 131.250 ;
        RECT 490.950 130.800 493.050 131.250 ;
        RECT 499.950 132.450 502.050 132.900 ;
        RECT 505.950 132.450 508.050 132.900 ;
        RECT 499.950 131.250 508.050 132.450 ;
        RECT 499.950 130.800 502.050 131.250 ;
        RECT 505.950 130.800 508.050 131.250 ;
        RECT 517.950 132.450 520.050 132.900 ;
        RECT 529.950 132.450 532.050 132.900 ;
        RECT 517.950 131.250 532.050 132.450 ;
        RECT 517.950 130.800 520.050 131.250 ;
        RECT 529.950 130.800 532.050 131.250 ;
        RECT 535.950 130.800 538.050 132.900 ;
        RECT 553.950 130.800 556.050 132.900 ;
        RECT 577.950 130.800 580.050 132.900 ;
        RECT 583.950 132.600 586.050 132.900 ;
        RECT 592.950 132.600 595.050 133.050 ;
        RECT 583.950 131.400 595.050 132.600 ;
        RECT 583.950 130.800 586.050 131.400 ;
        RECT 592.950 130.950 595.050 131.400 ;
        RECT 601.950 132.450 604.050 132.900 ;
        RECT 607.800 132.450 609.900 132.900 ;
        RECT 601.950 131.250 609.900 132.450 ;
        RECT 601.950 130.800 604.050 131.250 ;
        RECT 607.800 130.800 609.900 131.250 ;
        RECT 613.950 132.600 616.050 132.900 ;
        RECT 628.950 132.600 631.050 133.050 ;
        RECT 613.950 131.400 631.050 132.600 ;
        RECT 613.950 130.800 616.050 131.400 ;
        RECT 628.950 130.950 631.050 131.400 ;
        RECT 640.950 132.600 643.050 132.900 ;
        RECT 649.950 132.600 652.050 133.050 ;
        RECT 659.400 132.900 660.600 136.950 ;
        RECT 680.400 132.900 681.600 137.400 ;
        RECT 694.950 137.550 703.050 138.750 ;
        RECT 694.950 137.100 697.050 137.550 ;
        RECT 700.950 137.100 703.050 137.550 ;
        RECT 730.950 137.100 733.050 139.200 ;
        RECT 748.950 138.600 751.050 139.200 ;
        RECT 754.950 138.600 757.050 139.050 ;
        RECT 748.950 137.400 757.050 138.600 ;
        RECT 748.950 137.100 751.050 137.400 ;
        RECT 640.950 131.400 652.050 132.600 ;
        RECT 640.950 130.800 643.050 131.400 ;
        RECT 649.950 130.950 652.050 131.400 ;
        RECT 658.950 130.800 661.050 132.900 ;
        RECT 679.950 130.800 682.050 132.900 ;
        RECT 685.950 132.600 688.050 132.900 ;
        RECT 694.950 132.600 697.050 133.050 ;
        RECT 685.950 131.400 697.050 132.600 ;
        RECT 685.950 130.800 688.050 131.400 ;
        RECT 694.950 130.950 697.050 131.400 ;
        RECT 703.950 132.600 706.050 132.900 ;
        RECT 712.950 132.600 715.050 133.050 ;
        RECT 703.950 131.400 715.050 132.600 ;
        RECT 731.400 132.600 732.600 137.100 ;
        RECT 754.950 136.950 757.050 137.400 ;
        RECT 760.950 138.600 763.050 138.900 ;
        RECT 769.950 138.600 772.050 142.050 ;
        RECT 802.950 141.600 805.050 142.050 ;
        RECT 832.950 141.600 835.050 142.050 ;
        RECT 802.950 140.400 835.050 141.600 ;
        RECT 802.950 139.950 805.050 140.400 ;
        RECT 832.950 139.950 835.050 140.400 ;
        RECT 760.950 138.000 772.050 138.600 ;
        RECT 760.950 137.400 771.600 138.000 ;
        RECT 760.950 136.800 763.050 137.400 ;
        RECT 793.950 137.100 796.050 139.200 ;
        RECT 794.400 135.600 795.600 137.100 ;
        RECT 820.950 135.600 823.050 136.050 ;
        RECT 794.400 134.400 823.050 135.600 ;
        RECT 820.950 133.950 823.050 134.400 ;
        RECT 745.950 132.600 748.050 132.900 ;
        RECT 731.400 131.400 748.050 132.600 ;
        RECT 703.950 130.800 706.050 131.400 ;
        RECT 712.950 130.950 715.050 131.400 ;
        RECT 745.950 130.800 748.050 131.400 ;
        RECT 754.950 132.450 757.050 132.900 ;
        RECT 775.950 132.450 778.050 132.900 ;
        RECT 754.950 131.250 778.050 132.450 ;
        RECT 754.950 130.800 757.050 131.250 ;
        RECT 775.950 130.800 778.050 131.250 ;
        RECT 781.950 132.450 784.050 132.900 ;
        RECT 790.950 132.450 793.050 132.900 ;
        RECT 781.950 131.250 793.050 132.450 ;
        RECT 781.950 130.800 784.050 131.250 ;
        RECT 790.950 130.800 793.050 131.250 ;
        RECT 802.950 132.600 805.050 133.050 ;
        RECT 811.950 132.600 814.050 132.900 ;
        RECT 802.950 131.400 814.050 132.600 ;
        RECT 802.950 130.950 805.050 131.400 ;
        RECT 811.950 130.800 814.050 131.400 ;
        RECT 7.950 129.600 10.050 130.050 ;
        RECT 19.950 129.600 22.050 130.050 ;
        RECT 7.950 128.400 22.050 129.600 ;
        RECT 7.950 127.950 10.050 128.400 ;
        RECT 19.950 127.950 22.050 128.400 ;
        RECT 142.950 129.600 145.050 130.050 ;
        RECT 154.950 129.600 157.050 130.050 ;
        RECT 142.950 128.400 157.050 129.600 ;
        RECT 142.950 127.950 145.050 128.400 ;
        RECT 154.950 127.950 157.050 128.400 ;
        RECT 259.950 129.600 262.050 130.050 ;
        RECT 307.950 129.600 310.050 130.050 ;
        RECT 259.950 128.400 310.050 129.600 ;
        RECT 259.950 127.950 262.050 128.400 ;
        RECT 307.950 127.950 310.050 128.400 ;
        RECT 388.950 129.600 391.050 130.050 ;
        RECT 394.950 129.600 397.050 130.050 ;
        RECT 388.950 128.400 397.050 129.600 ;
        RECT 608.400 129.600 609.600 130.800 ;
        RECT 634.950 129.600 637.050 130.050 ;
        RECT 608.400 128.400 637.050 129.600 ;
        RECT 388.950 127.950 391.050 128.400 ;
        RECT 394.950 127.950 397.050 128.400 ;
        RECT 634.950 127.950 637.050 128.400 ;
        RECT 775.950 129.600 778.050 130.050 ;
        RECT 817.950 129.600 820.050 130.050 ;
        RECT 841.950 129.600 844.050 130.050 ;
        RECT 859.950 129.600 862.050 130.050 ;
        RECT 775.950 128.400 862.050 129.600 ;
        RECT 775.950 127.950 778.050 128.400 ;
        RECT 817.950 127.950 820.050 128.400 ;
        RECT 841.950 127.950 844.050 128.400 ;
        RECT 859.950 127.950 862.050 128.400 ;
        RECT 64.950 126.600 67.050 127.050 ;
        RECT 91.950 126.600 94.050 127.050 ;
        RECT 64.950 125.400 94.050 126.600 ;
        RECT 64.950 124.950 67.050 125.400 ;
        RECT 91.950 124.950 94.050 125.400 ;
        RECT 121.950 126.600 124.050 127.050 ;
        RECT 130.950 126.600 133.050 127.050 ;
        RECT 208.950 126.600 211.050 127.050 ;
        RECT 121.950 125.400 211.050 126.600 ;
        RECT 121.950 124.950 124.050 125.400 ;
        RECT 130.950 124.950 133.050 125.400 ;
        RECT 208.950 124.950 211.050 125.400 ;
        RECT 469.950 126.600 472.050 127.050 ;
        RECT 526.950 126.600 529.050 127.050 ;
        RECT 469.950 125.400 529.050 126.600 ;
        RECT 469.950 124.950 472.050 125.400 ;
        RECT 526.950 124.950 529.050 125.400 ;
        RECT 694.950 126.600 697.050 127.050 ;
        RECT 715.950 126.600 718.050 127.050 ;
        RECT 694.950 125.400 718.050 126.600 ;
        RECT 694.950 124.950 697.050 125.400 ;
        RECT 715.950 124.950 718.050 125.400 ;
        RECT 721.950 126.600 724.050 127.050 ;
        RECT 754.950 126.600 757.050 127.050 ;
        RECT 721.950 125.400 757.050 126.600 ;
        RECT 721.950 124.950 724.050 125.400 ;
        RECT 754.950 124.950 757.050 125.400 ;
        RECT 259.950 123.600 262.050 124.050 ;
        RECT 292.950 123.600 295.050 124.050 ;
        RECT 259.950 122.400 295.050 123.600 ;
        RECT 259.950 121.950 262.050 122.400 ;
        RECT 292.950 121.950 295.050 122.400 ;
        RECT 337.950 123.600 340.050 124.050 ;
        RECT 370.950 123.600 373.050 124.050 ;
        RECT 337.950 122.400 373.050 123.600 ;
        RECT 337.950 121.950 340.050 122.400 ;
        RECT 370.950 121.950 373.050 122.400 ;
        RECT 445.950 123.600 448.050 124.050 ;
        RECT 532.950 123.600 535.050 124.050 ;
        RECT 445.950 122.400 535.050 123.600 ;
        RECT 445.950 121.950 448.050 122.400 ;
        RECT 532.950 121.950 535.050 122.400 ;
        RECT 538.950 123.600 541.050 124.050 ;
        RECT 559.950 123.600 562.050 124.050 ;
        RECT 538.950 122.400 562.050 123.600 ;
        RECT 538.950 121.950 541.050 122.400 ;
        RECT 559.950 121.950 562.050 122.400 ;
        RECT 607.950 123.600 610.050 124.050 ;
        RECT 691.950 123.600 694.050 124.050 ;
        RECT 607.950 122.400 694.050 123.600 ;
        RECT 607.950 121.950 610.050 122.400 ;
        RECT 691.950 121.950 694.050 122.400 ;
        RECT 163.950 120.600 166.050 121.050 ;
        RECT 172.950 120.600 175.050 121.050 ;
        RECT 163.950 119.400 175.050 120.600 ;
        RECT 163.950 118.950 166.050 119.400 ;
        RECT 172.950 118.950 175.050 119.400 ;
        RECT 226.950 120.600 229.050 121.050 ;
        RECT 310.950 120.600 313.050 121.050 ;
        RECT 322.950 120.600 325.050 121.050 ;
        RECT 358.950 120.600 361.050 121.050 ;
        RECT 226.950 119.400 361.050 120.600 ;
        RECT 226.950 118.950 229.050 119.400 ;
        RECT 310.950 118.950 313.050 119.400 ;
        RECT 322.950 118.950 325.050 119.400 ;
        RECT 358.950 118.950 361.050 119.400 ;
        RECT 397.950 120.600 400.050 121.050 ;
        RECT 469.950 120.600 472.050 121.050 ;
        RECT 397.950 119.400 472.050 120.600 ;
        RECT 397.950 118.950 400.050 119.400 ;
        RECT 469.950 118.950 472.050 119.400 ;
        RECT 667.950 120.600 670.050 121.050 ;
        RECT 709.950 120.600 712.050 121.050 ;
        RECT 667.950 119.400 712.050 120.600 ;
        RECT 667.950 118.950 670.050 119.400 ;
        RECT 709.950 118.950 712.050 119.400 ;
        RECT 763.950 120.600 766.050 121.050 ;
        RECT 784.950 120.600 787.050 121.050 ;
        RECT 763.950 119.400 787.050 120.600 ;
        RECT 763.950 118.950 766.050 119.400 ;
        RECT 784.950 118.950 787.050 119.400 ;
        RECT 826.950 120.600 829.050 121.050 ;
        RECT 886.950 120.600 889.050 121.050 ;
        RECT 826.950 119.400 889.050 120.600 ;
        RECT 826.950 118.950 829.050 119.400 ;
        RECT 886.950 118.950 889.050 119.400 ;
        RECT 40.950 117.600 43.050 118.050 ;
        RECT 52.950 117.600 55.050 118.050 ;
        RECT 85.950 117.600 88.050 118.050 ;
        RECT 40.950 116.400 88.050 117.600 ;
        RECT 40.950 115.950 43.050 116.400 ;
        RECT 52.950 115.950 55.050 116.400 ;
        RECT 85.950 115.950 88.050 116.400 ;
        RECT 118.950 117.600 121.050 118.050 ;
        RECT 139.950 117.600 142.050 118.050 ;
        RECT 118.950 116.400 142.050 117.600 ;
        RECT 118.950 115.950 121.050 116.400 ;
        RECT 139.950 115.950 142.050 116.400 ;
        RECT 247.950 117.600 250.050 118.050 ;
        RECT 265.950 117.600 268.050 118.050 ;
        RECT 247.950 116.400 268.050 117.600 ;
        RECT 247.950 115.950 250.050 116.400 ;
        RECT 265.950 115.950 268.050 116.400 ;
        RECT 271.950 117.600 274.050 118.050 ;
        RECT 289.800 117.600 291.900 118.050 ;
        RECT 271.950 116.400 291.900 117.600 ;
        RECT 271.950 115.950 274.050 116.400 ;
        RECT 289.800 115.950 291.900 116.400 ;
        RECT 292.950 117.600 295.050 118.050 ;
        RECT 328.950 117.600 331.050 118.050 ;
        RECT 292.950 116.400 331.050 117.600 ;
        RECT 292.950 115.950 295.050 116.400 ;
        RECT 328.950 115.950 331.050 116.400 ;
        RECT 475.950 117.600 478.050 118.050 ;
        RECT 484.950 117.600 487.050 118.050 ;
        RECT 544.950 117.600 547.050 118.050 ;
        RECT 475.950 116.400 547.050 117.600 ;
        RECT 475.950 115.950 478.050 116.400 ;
        RECT 484.950 115.950 487.050 116.400 ;
        RECT 544.950 115.950 547.050 116.400 ;
        RECT 568.950 117.600 571.050 118.050 ;
        RECT 613.950 117.600 616.050 118.050 ;
        RECT 568.950 116.400 616.050 117.600 ;
        RECT 568.950 115.950 571.050 116.400 ;
        RECT 613.950 115.950 616.050 116.400 ;
        RECT 646.950 117.600 649.050 118.050 ;
        RECT 685.950 117.600 688.050 118.050 ;
        RECT 646.950 116.400 688.050 117.600 ;
        RECT 646.950 115.950 649.050 116.400 ;
        RECT 685.950 115.950 688.050 116.400 ;
        RECT 721.950 117.600 724.050 118.050 ;
        RECT 790.950 117.600 793.050 118.050 ;
        RECT 721.950 116.400 793.050 117.600 ;
        RECT 721.950 115.950 724.050 116.400 ;
        RECT 790.950 115.950 793.050 116.400 ;
        RECT 7.950 114.600 10.050 115.050 ;
        RECT 58.950 114.600 61.050 115.050 ;
        RECT 79.950 114.600 82.050 115.050 ;
        RECT 106.950 114.600 109.050 115.050 ;
        RECT 7.950 113.400 109.050 114.600 ;
        RECT 7.950 112.950 10.050 113.400 ;
        RECT 58.950 112.950 61.050 113.400 ;
        RECT 79.950 112.950 82.050 113.400 ;
        RECT 106.950 112.950 109.050 113.400 ;
        RECT 286.950 114.600 289.050 115.050 ;
        RECT 355.950 114.600 358.050 115.050 ;
        RECT 382.950 114.600 385.050 115.050 ;
        RECT 403.950 114.600 406.050 115.050 ;
        RECT 286.950 113.400 406.050 114.600 ;
        RECT 286.950 112.950 289.050 113.400 ;
        RECT 355.950 112.950 358.050 113.400 ;
        RECT 382.950 112.950 385.050 113.400 ;
        RECT 403.950 112.950 406.050 113.400 ;
        RECT 601.950 114.600 604.050 115.050 ;
        RECT 637.950 114.600 640.050 115.050 ;
        RECT 601.950 113.400 640.050 114.600 ;
        RECT 601.950 112.950 604.050 113.400 ;
        RECT 637.950 112.950 640.050 113.400 ;
        RECT 844.950 114.600 847.050 115.050 ;
        RECT 856.950 114.600 859.050 115.050 ;
        RECT 844.950 113.400 859.050 114.600 ;
        RECT 844.950 112.950 847.050 113.400 ;
        RECT 856.950 112.950 859.050 113.400 ;
        RECT 16.950 111.600 19.050 112.050 ;
        RECT 28.950 111.600 31.050 112.050 ;
        RECT 16.950 110.400 31.050 111.600 ;
        RECT 16.950 109.950 19.050 110.400 ;
        RECT 28.950 109.950 31.050 110.400 ;
        RECT 82.950 111.600 85.050 112.050 ;
        RECT 91.950 111.600 94.050 112.050 ;
        RECT 82.950 110.400 94.050 111.600 ;
        RECT 82.950 109.950 85.050 110.400 ;
        RECT 91.950 109.950 94.050 110.400 ;
        RECT 112.950 111.600 115.050 112.050 ;
        RECT 124.800 111.600 126.900 112.050 ;
        RECT 112.950 110.400 126.900 111.600 ;
        RECT 112.950 109.950 115.050 110.400 ;
        RECT 124.800 109.950 126.900 110.400 ;
        RECT 127.950 111.600 130.050 112.050 ;
        RECT 163.950 111.600 166.050 112.050 ;
        RECT 127.950 110.400 166.050 111.600 ;
        RECT 127.950 109.950 130.050 110.400 ;
        RECT 163.950 109.950 166.050 110.400 ;
        RECT 175.950 111.600 178.050 112.050 ;
        RECT 184.950 111.600 187.050 112.050 ;
        RECT 175.950 110.400 187.050 111.600 ;
        RECT 175.950 109.950 178.050 110.400 ;
        RECT 184.950 109.950 187.050 110.400 ;
        RECT 193.950 111.600 196.050 112.050 ;
        RECT 271.950 111.600 274.050 112.050 ;
        RECT 193.950 110.400 274.050 111.600 ;
        RECT 193.950 109.950 196.050 110.400 ;
        RECT 271.950 109.950 274.050 110.400 ;
        RECT 298.950 111.600 301.050 112.050 ;
        RECT 328.950 111.600 331.050 112.050 ;
        RECT 337.950 111.600 340.050 112.050 ;
        RECT 298.950 110.400 340.050 111.600 ;
        RECT 298.950 109.950 301.050 110.400 ;
        RECT 328.950 109.950 331.050 110.400 ;
        RECT 337.950 109.950 340.050 110.400 ;
        RECT 343.950 111.600 346.050 112.050 ;
        RECT 352.950 111.600 355.050 112.050 ;
        RECT 343.950 110.400 355.050 111.600 ;
        RECT 343.950 109.950 346.050 110.400 ;
        RECT 352.950 109.950 355.050 110.400 ;
        RECT 364.950 111.600 367.050 112.050 ;
        RECT 403.950 111.600 406.050 111.900 ;
        RECT 364.950 110.400 406.050 111.600 ;
        RECT 364.950 109.950 367.050 110.400 ;
        RECT 403.950 109.800 406.050 110.400 ;
        RECT 451.950 111.600 454.050 112.050 ;
        RECT 481.950 111.600 484.050 112.050 ;
        RECT 451.950 110.400 484.050 111.600 ;
        RECT 451.950 109.950 454.050 110.400 ;
        RECT 481.950 109.950 484.050 110.400 ;
        RECT 487.950 111.600 490.050 112.050 ;
        RECT 502.950 111.600 505.050 112.050 ;
        RECT 511.950 111.600 514.050 112.050 ;
        RECT 487.950 110.400 514.050 111.600 ;
        RECT 487.950 109.950 490.050 110.400 ;
        RECT 502.950 109.950 505.050 110.400 ;
        RECT 511.950 109.950 514.050 110.400 ;
        RECT 532.950 111.600 535.050 112.050 ;
        RECT 541.950 111.600 544.050 112.050 ;
        RECT 532.950 110.400 544.050 111.600 ;
        RECT 532.950 109.950 535.050 110.400 ;
        RECT 541.950 109.950 544.050 110.400 ;
        RECT 577.950 111.600 580.050 112.050 ;
        RECT 610.950 111.600 613.050 112.050 ;
        RECT 619.950 111.600 622.050 112.050 ;
        RECT 577.950 110.400 622.050 111.600 ;
        RECT 577.950 109.950 580.050 110.400 ;
        RECT 610.950 109.950 613.050 110.400 ;
        RECT 619.950 109.950 622.050 110.400 ;
        RECT 670.950 111.600 673.050 112.050 ;
        RECT 685.950 111.600 688.050 112.050 ;
        RECT 670.950 110.400 688.050 111.600 ;
        RECT 670.950 109.950 673.050 110.400 ;
        RECT 685.950 109.950 688.050 110.400 ;
        RECT 760.950 111.600 763.050 112.050 ;
        RECT 769.950 111.600 772.050 112.050 ;
        RECT 760.950 110.400 772.050 111.600 ;
        RECT 760.950 109.950 763.050 110.400 ;
        RECT 769.950 109.950 772.050 110.400 ;
        RECT 790.950 111.600 793.050 112.050 ;
        RECT 832.800 111.600 834.900 112.050 ;
        RECT 790.950 110.400 834.900 111.600 ;
        RECT 790.950 109.950 793.050 110.400 ;
        RECT 832.800 109.950 834.900 110.400 ;
        RECT 835.950 111.600 838.050 112.050 ;
        RECT 841.950 111.600 844.050 112.050 ;
        RECT 835.950 110.400 844.050 111.600 ;
        RECT 835.950 109.950 838.050 110.400 ;
        RECT 841.950 109.950 844.050 110.400 ;
        RECT 4.950 108.600 7.050 109.050 ;
        RECT 13.950 108.600 16.050 109.050 ;
        RECT 4.950 107.400 16.050 108.600 ;
        RECT 4.950 106.950 7.050 107.400 ;
        RECT 13.950 106.950 16.050 107.400 ;
        RECT 25.950 105.750 28.050 106.200 ;
        RECT 58.950 105.750 61.050 106.200 ;
        RECT 25.950 104.550 61.050 105.750 ;
        RECT 25.950 104.100 28.050 104.550 ;
        RECT 58.950 104.100 61.050 104.550 ;
        RECT 64.950 105.600 67.050 106.200 ;
        RECT 73.950 105.600 76.050 106.050 ;
        RECT 64.950 104.400 76.050 105.600 ;
        RECT 64.950 104.100 67.050 104.400 ;
        RECT 73.950 103.950 76.050 104.400 ;
        RECT 79.950 105.600 84.000 106.050 ;
        RECT 94.950 105.600 97.050 106.050 ;
        RECT 100.950 105.600 103.050 106.050 ;
        RECT 121.950 105.600 124.050 106.050 ;
        RECT 133.950 105.600 136.050 106.200 ;
        RECT 79.950 103.950 84.600 105.600 ;
        RECT 94.950 104.400 103.050 105.600 ;
        RECT 94.950 103.950 97.050 104.400 ;
        RECT 100.950 103.950 103.050 104.400 ;
        RECT 110.400 104.400 124.050 105.600 ;
        RECT 83.400 99.900 84.600 103.950 ;
        RECT 110.400 99.900 111.600 104.400 ;
        RECT 121.950 103.950 124.050 104.400 ;
        RECT 131.400 104.400 136.050 105.600 ;
        RECT 131.400 100.050 132.600 104.400 ;
        RECT 133.950 104.100 136.050 104.400 ;
        RECT 139.950 105.750 142.050 106.200 ;
        RECT 148.950 105.750 151.050 106.200 ;
        RECT 139.950 104.550 151.050 105.750 ;
        RECT 139.950 104.100 142.050 104.550 ;
        RECT 148.950 104.100 151.050 104.550 ;
        RECT 157.950 104.100 160.050 106.200 ;
        RECT 169.950 105.600 172.050 106.050 ;
        RECT 178.950 105.600 181.050 106.200 ;
        RECT 169.950 104.400 181.050 105.600 ;
        RECT 7.950 99.450 10.050 99.900 ;
        RECT 13.950 99.450 16.050 99.900 ;
        RECT 7.950 98.250 16.050 99.450 ;
        RECT 7.950 97.800 10.050 98.250 ;
        RECT 13.950 97.800 16.050 98.250 ;
        RECT 46.950 99.450 49.050 99.900 ;
        RECT 52.950 99.450 55.050 99.900 ;
        RECT 46.950 98.250 55.050 99.450 ;
        RECT 46.950 97.800 49.050 98.250 ;
        RECT 52.950 97.800 55.050 98.250 ;
        RECT 82.950 97.800 85.050 99.900 ;
        RECT 109.950 97.800 112.050 99.900 ;
        RECT 130.950 97.950 133.050 100.050 ;
        RECT 136.950 99.600 139.050 99.900 ;
        RECT 158.400 99.600 159.600 104.100 ;
        RECT 169.950 103.950 172.050 104.400 ;
        RECT 178.950 104.100 181.050 104.400 ;
        RECT 184.950 105.600 187.050 106.200 ;
        RECT 190.950 105.600 193.050 109.050 ;
        RECT 274.950 108.600 277.050 109.050 ;
        RECT 331.950 108.600 334.050 109.050 ;
        RECT 361.950 108.600 364.050 109.050 ;
        RECT 406.950 108.600 409.050 109.050 ;
        RECT 448.950 108.600 451.050 109.050 ;
        RECT 274.950 107.400 369.600 108.600 ;
        RECT 274.950 106.950 277.050 107.400 ;
        RECT 331.950 106.950 334.050 107.400 ;
        RECT 361.950 106.950 364.050 107.400 ;
        RECT 202.950 105.600 205.050 106.200 ;
        RECT 184.950 105.000 193.050 105.600 ;
        RECT 184.950 104.400 192.600 105.000 ;
        RECT 194.400 104.400 205.050 105.600 ;
        RECT 184.950 104.100 187.050 104.400 ;
        RECT 194.400 102.600 195.600 104.400 ;
        RECT 202.950 104.100 205.050 104.400 ;
        RECT 208.950 105.600 211.050 106.200 ;
        RECT 220.950 105.600 223.050 106.050 ;
        RECT 232.950 105.600 235.050 106.200 ;
        RECT 208.950 104.400 213.600 105.600 ;
        RECT 208.950 104.100 211.050 104.400 ;
        RECT 188.400 101.400 195.600 102.600 ;
        RECT 188.400 99.900 189.600 101.400 ;
        RECT 212.400 100.050 213.600 104.400 ;
        RECT 220.950 104.400 235.050 105.600 ;
        RECT 220.950 103.950 223.050 104.400 ;
        RECT 232.950 104.100 235.050 104.400 ;
        RECT 247.950 104.100 250.050 106.200 ;
        RECT 262.950 105.600 265.050 106.050 ;
        RECT 268.950 105.600 271.050 106.200 ;
        RECT 262.950 104.400 271.050 105.600 ;
        RECT 136.950 98.400 159.600 99.600 ;
        RECT 136.950 97.800 139.050 98.400 ;
        RECT 187.950 97.800 190.050 99.900 ;
        RECT 193.950 99.450 196.050 99.900 ;
        RECT 205.950 99.450 208.050 99.900 ;
        RECT 193.950 98.250 208.050 99.450 ;
        RECT 193.950 97.800 196.050 98.250 ;
        RECT 205.950 97.800 208.050 98.250 ;
        RECT 211.950 97.950 214.050 100.050 ;
        RECT 235.950 99.600 238.050 99.900 ;
        RECT 248.400 99.600 249.600 104.100 ;
        RECT 262.950 103.950 265.050 104.400 ;
        RECT 268.950 104.100 271.050 104.400 ;
        RECT 286.950 105.600 291.000 106.050 ;
        RECT 307.950 105.600 310.050 106.050 ;
        RECT 316.950 105.600 319.050 106.200 ;
        RECT 286.950 103.950 291.600 105.600 ;
        RECT 307.950 104.400 319.050 105.600 ;
        RECT 307.950 103.950 310.050 104.400 ;
        RECT 316.950 104.100 319.050 104.400 ;
        RECT 355.950 103.950 358.050 106.050 ;
        RECT 235.950 98.400 249.600 99.600 ;
        RECT 250.950 99.600 253.050 99.900 ;
        RECT 259.950 99.600 262.050 100.050 ;
        RECT 250.950 98.400 262.050 99.600 ;
        RECT 235.950 97.800 238.050 98.400 ;
        RECT 250.950 97.800 253.050 98.400 ;
        RECT 259.950 97.950 262.050 98.400 ;
        RECT 265.950 99.600 268.050 100.050 ;
        RECT 290.400 99.900 291.600 103.950 ;
        RECT 277.950 99.600 280.050 99.900 ;
        RECT 265.950 98.400 280.050 99.600 ;
        RECT 265.950 97.950 268.050 98.400 ;
        RECT 277.950 97.800 280.050 98.400 ;
        RECT 289.950 97.800 292.050 99.900 ;
        RECT 331.950 99.450 334.050 99.900 ;
        RECT 340.950 99.450 343.050 99.900 ;
        RECT 331.950 98.250 343.050 99.450 ;
        RECT 331.950 97.800 334.050 98.250 ;
        RECT 340.950 97.800 343.050 98.250 ;
        RECT 346.950 99.600 349.050 99.900 ;
        RECT 356.400 99.600 357.600 103.950 ;
        RECT 368.400 99.900 369.600 107.400 ;
        RECT 406.950 107.400 451.050 108.600 ;
        RECT 406.950 106.950 409.050 107.400 ;
        RECT 448.950 106.950 451.050 107.400 ;
        RECT 550.950 108.600 553.050 109.050 ;
        RECT 559.950 108.600 562.050 109.050 ;
        RECT 550.950 107.400 562.050 108.600 ;
        RECT 550.950 106.950 553.050 107.400 ;
        RECT 559.950 106.950 562.050 107.400 ;
        RECT 703.950 108.600 706.050 109.050 ;
        RECT 715.950 108.600 718.050 109.050 ;
        RECT 703.950 107.400 718.050 108.600 ;
        RECT 703.950 106.950 706.050 107.400 ;
        RECT 715.950 106.950 718.050 107.400 ;
        RECT 745.950 108.600 748.050 109.050 ;
        RECT 763.950 108.600 766.050 109.050 ;
        RECT 847.950 108.600 850.050 109.050 ;
        RECT 862.950 108.600 865.050 109.050 ;
        RECT 745.950 107.400 766.050 108.600 ;
        RECT 745.950 106.950 748.050 107.400 ;
        RECT 763.950 106.950 766.050 107.400 ;
        RECT 821.400 107.400 865.050 108.600 ;
        RECT 370.950 102.600 373.050 106.050 ;
        RECT 388.950 105.600 391.050 106.200 ;
        RECT 445.950 105.600 448.050 106.050 ;
        RECT 388.950 104.400 448.050 105.600 ;
        RECT 388.950 104.100 391.050 104.400 ;
        RECT 370.950 102.000 381.600 102.600 ;
        RECT 371.400 101.400 381.600 102.000 ;
        RECT 380.400 99.900 381.600 101.400 ;
        RECT 404.400 99.900 405.600 104.400 ;
        RECT 445.950 103.950 448.050 104.400 ;
        RECT 463.950 104.100 466.050 106.200 ;
        RECT 508.950 105.600 511.050 106.200 ;
        RECT 514.950 105.600 517.050 106.050 ;
        RECT 508.950 104.400 517.050 105.600 ;
        RECT 508.950 104.100 511.050 104.400 ;
        RECT 464.400 102.600 465.600 104.100 ;
        RECT 509.400 102.600 510.600 104.100 ;
        RECT 514.950 103.950 517.050 104.400 ;
        RECT 541.950 105.600 544.050 106.050 ;
        RECT 562.950 105.600 565.050 106.050 ;
        RECT 571.950 105.600 574.050 106.200 ;
        RECT 541.950 104.400 552.600 105.600 ;
        RECT 541.950 103.950 544.050 104.400 ;
        RECT 464.400 101.400 489.600 102.600 ;
        RECT 346.950 98.400 357.600 99.600 ;
        RECT 346.950 97.800 349.050 98.400 ;
        RECT 367.950 97.800 370.050 99.900 ;
        RECT 379.950 97.800 382.050 99.900 ;
        RECT 403.950 97.800 406.050 99.900 ;
        RECT 421.950 99.600 424.050 100.050 ;
        RECT 427.950 99.600 430.050 99.900 ;
        RECT 421.950 98.400 430.050 99.600 ;
        RECT 421.950 97.950 424.050 98.400 ;
        RECT 427.950 97.800 430.050 98.400 ;
        RECT 448.950 99.450 451.050 99.900 ;
        RECT 454.950 99.450 457.050 99.900 ;
        RECT 448.950 98.250 457.050 99.450 ;
        RECT 448.950 97.800 451.050 98.250 ;
        RECT 454.950 97.800 457.050 98.250 ;
        RECT 478.950 99.450 481.050 99.900 ;
        RECT 484.950 99.450 487.050 99.900 ;
        RECT 478.950 98.250 487.050 99.450 ;
        RECT 488.400 99.600 489.600 101.400 ;
        RECT 506.400 101.400 510.600 102.600 ;
        RECT 551.400 102.600 552.600 104.400 ;
        RECT 562.950 104.400 574.050 105.600 ;
        RECT 562.950 103.950 565.050 104.400 ;
        RECT 571.950 104.100 574.050 104.400 ;
        RECT 628.950 104.250 631.050 106.350 ;
        RECT 821.400 106.200 822.600 107.400 ;
        RECT 847.950 106.950 850.050 107.400 ;
        RECT 862.950 106.950 865.050 107.400 ;
        RECT 658.950 105.600 661.050 106.200 ;
        RECT 667.950 105.600 670.050 106.050 ;
        RECT 658.950 104.400 670.050 105.600 ;
        RECT 616.950 102.600 619.050 103.050 ;
        RECT 629.400 102.600 630.600 104.250 ;
        RECT 658.950 104.100 661.050 104.400 ;
        RECT 667.950 103.950 670.050 104.400 ;
        RECT 673.950 104.100 676.050 106.200 ;
        RECT 726.000 105.600 729.900 106.050 ;
        RECT 551.400 101.400 555.600 102.600 ;
        RECT 506.400 99.600 507.600 101.400 ;
        RECT 488.400 98.400 507.600 99.600 ;
        RECT 529.950 99.600 532.050 99.900 ;
        RECT 538.950 99.600 541.050 100.050 ;
        RECT 554.400 99.900 555.600 101.400 ;
        RECT 616.950 101.400 630.600 102.600 ;
        RECT 635.400 102.000 648.600 102.600 ;
        RECT 634.950 101.400 648.600 102.000 ;
        RECT 616.950 100.950 619.050 101.400 ;
        RECT 547.950 99.600 550.050 99.900 ;
        RECT 529.950 98.400 550.050 99.600 ;
        RECT 478.950 97.800 481.050 98.250 ;
        RECT 484.950 97.800 487.050 98.250 ;
        RECT 529.950 97.800 532.050 98.400 ;
        RECT 538.950 97.950 541.050 98.400 ;
        RECT 547.950 97.800 550.050 98.400 ;
        RECT 553.950 97.800 556.050 99.900 ;
        RECT 559.950 99.450 562.050 99.900 ;
        RECT 574.950 99.450 577.050 99.900 ;
        RECT 559.950 98.250 577.050 99.450 ;
        RECT 559.950 97.800 562.050 98.250 ;
        RECT 574.950 97.800 577.050 98.250 ;
        RECT 598.950 99.450 601.050 99.900 ;
        RECT 610.950 99.450 613.050 99.900 ;
        RECT 598.950 98.250 613.050 99.450 ;
        RECT 598.950 97.800 601.050 98.250 ;
        RECT 610.950 97.800 613.050 98.250 ;
        RECT 634.950 97.950 637.050 101.400 ;
        RECT 647.400 99.900 648.600 101.400 ;
        RECT 674.400 100.050 675.600 104.100 ;
        RECT 646.950 99.450 649.050 99.900 ;
        RECT 661.950 99.450 664.050 99.900 ;
        RECT 646.950 98.250 664.050 99.450 ;
        RECT 646.950 97.800 649.050 98.250 ;
        RECT 661.950 97.800 664.050 98.250 ;
        RECT 670.950 98.400 675.600 100.050 ;
        RECT 725.400 103.950 729.900 105.600 ;
        RECT 730.950 105.750 733.050 106.200 ;
        RECT 739.950 105.750 742.050 106.200 ;
        RECT 730.950 104.550 742.050 105.750 ;
        RECT 730.950 104.100 733.050 104.550 ;
        RECT 739.950 104.100 742.050 104.550 ;
        RECT 754.950 105.600 757.050 106.050 ;
        RECT 790.950 105.600 793.050 106.200 ;
        RECT 754.950 104.400 793.050 105.600 ;
        RECT 754.950 103.950 757.050 104.400 ;
        RECT 790.950 104.100 793.050 104.400 ;
        RECT 796.950 105.750 799.050 106.200 ;
        RECT 808.950 105.750 811.050 106.200 ;
        RECT 796.950 104.550 811.050 105.750 ;
        RECT 796.950 104.100 799.050 104.550 ;
        RECT 808.950 104.100 811.050 104.550 ;
        RECT 814.950 105.750 817.050 106.200 ;
        RECT 820.950 105.750 823.050 106.200 ;
        RECT 814.950 104.550 823.050 105.750 ;
        RECT 841.950 105.600 844.050 106.050 ;
        RECT 895.950 105.600 898.050 106.200 ;
        RECT 814.950 104.100 817.050 104.550 ;
        RECT 820.950 104.100 823.050 104.550 ;
        RECT 830.400 104.400 844.050 105.600 ;
        RECT 725.400 99.900 726.600 103.950 ;
        RECT 830.400 99.900 831.600 104.400 ;
        RECT 841.950 103.950 844.050 104.400 ;
        RECT 851.400 104.400 898.050 105.600 ;
        RECT 851.400 100.050 852.600 104.400 ;
        RECT 895.950 104.100 898.050 104.400 ;
        RECT 670.950 97.950 675.000 98.400 ;
        RECT 724.950 97.800 727.050 99.900 ;
        RECT 766.950 99.600 769.050 99.900 ;
        RECT 787.950 99.600 790.050 99.900 ;
        RECT 766.950 98.400 790.050 99.600 ;
        RECT 766.950 97.800 769.050 98.400 ;
        RECT 787.950 97.800 790.050 98.400 ;
        RECT 829.950 97.800 832.050 99.900 ;
        RECT 850.950 97.950 853.050 100.050 ;
        RECT 61.950 96.600 64.050 97.050 ;
        RECT 50.400 95.400 64.050 96.600 ;
        RECT 4.950 93.600 7.050 94.050 ;
        RECT 19.950 93.600 22.050 94.050 ;
        RECT 50.400 93.600 51.600 95.400 ;
        RECT 61.950 94.950 64.050 95.400 ;
        RECT 88.950 96.600 91.050 97.050 ;
        RECT 100.950 96.600 103.050 97.050 ;
        RECT 88.950 95.400 103.050 96.600 ;
        RECT 88.950 94.950 91.050 95.400 ;
        RECT 100.950 94.950 103.050 95.400 ;
        RECT 181.950 96.600 184.050 97.050 ;
        RECT 194.400 96.600 195.600 97.800 ;
        RECT 181.950 95.400 195.600 96.600 ;
        RECT 223.950 96.600 226.050 97.050 ;
        RECT 262.950 96.600 265.050 97.050 ;
        RECT 223.950 95.400 265.050 96.600 ;
        RECT 181.950 94.950 184.050 95.400 ;
        RECT 223.950 94.950 226.050 95.400 ;
        RECT 262.950 94.950 265.050 95.400 ;
        RECT 313.950 96.600 316.050 97.050 ;
        RECT 328.950 96.600 331.050 97.050 ;
        RECT 313.950 95.400 331.050 96.600 ;
        RECT 313.950 94.950 316.050 95.400 ;
        RECT 328.950 94.950 331.050 95.400 ;
        RECT 514.950 96.600 517.050 97.050 ;
        RECT 676.950 96.600 679.050 97.050 ;
        RECT 697.950 96.600 700.050 97.050 ;
        RECT 514.950 95.400 522.600 96.600 ;
        RECT 514.950 94.950 517.050 95.400 ;
        RECT 4.950 92.400 51.600 93.600 ;
        RECT 52.950 93.600 55.050 94.050 ;
        RECT 67.950 93.600 70.050 94.050 ;
        RECT 52.950 92.400 70.050 93.600 ;
        RECT 4.950 91.950 7.050 92.400 ;
        RECT 19.950 91.950 22.050 92.400 ;
        RECT 52.950 91.950 55.050 92.400 ;
        RECT 67.950 91.950 70.050 92.400 ;
        RECT 115.950 93.600 118.050 94.050 ;
        RECT 172.950 93.600 175.050 94.050 ;
        RECT 115.950 92.400 175.050 93.600 ;
        RECT 115.950 91.950 118.050 92.400 ;
        RECT 172.950 91.950 175.050 92.400 ;
        RECT 220.950 93.600 223.050 94.050 ;
        RECT 244.950 93.600 247.050 94.050 ;
        RECT 220.950 92.400 247.050 93.600 ;
        RECT 220.950 91.950 223.050 92.400 ;
        RECT 244.950 91.950 247.050 92.400 ;
        RECT 361.950 93.600 364.050 94.050 ;
        RECT 373.950 93.600 376.050 94.050 ;
        RECT 361.950 92.400 376.050 93.600 ;
        RECT 361.950 91.950 364.050 92.400 ;
        RECT 373.950 91.950 376.050 92.400 ;
        RECT 436.950 93.600 439.050 94.050 ;
        RECT 490.950 93.600 493.050 94.050 ;
        RECT 499.950 93.600 502.050 94.050 ;
        RECT 436.950 92.400 502.050 93.600 ;
        RECT 521.400 93.600 522.600 95.400 ;
        RECT 676.950 95.400 700.050 96.600 ;
        RECT 676.950 94.950 679.050 95.400 ;
        RECT 697.950 94.950 700.050 95.400 ;
        RECT 721.950 96.600 724.050 97.050 ;
        RECT 730.950 96.600 733.050 97.050 ;
        RECT 721.950 95.400 733.050 96.600 ;
        RECT 721.950 94.950 724.050 95.400 ;
        RECT 730.950 94.950 733.050 95.400 ;
        RECT 757.950 96.600 760.050 97.050 ;
        RECT 805.950 96.600 808.050 97.050 ;
        RECT 757.950 95.400 808.050 96.600 ;
        RECT 757.950 94.950 760.050 95.400 ;
        RECT 805.950 94.950 808.050 95.400 ;
        RECT 865.950 96.600 868.050 97.050 ;
        RECT 898.950 96.600 901.050 97.050 ;
        RECT 865.950 95.400 901.050 96.600 ;
        RECT 865.950 94.950 868.050 95.400 ;
        RECT 898.950 94.950 901.050 95.400 ;
        RECT 580.950 93.600 583.050 94.050 ;
        RECT 586.950 93.600 589.050 94.050 ;
        RECT 521.400 92.400 589.050 93.600 ;
        RECT 436.950 91.950 439.050 92.400 ;
        RECT 490.950 91.950 493.050 92.400 ;
        RECT 499.950 91.950 502.050 92.400 ;
        RECT 580.950 91.950 583.050 92.400 ;
        RECT 586.950 91.950 589.050 92.400 ;
        RECT 667.950 93.600 670.050 94.050 ;
        RECT 691.950 93.600 694.050 94.050 ;
        RECT 667.950 92.400 694.050 93.600 ;
        RECT 667.950 91.950 670.050 92.400 ;
        RECT 691.950 91.950 694.050 92.400 ;
        RECT 745.950 93.600 748.050 94.050 ;
        RECT 781.950 93.600 784.050 94.050 ;
        RECT 745.950 92.400 784.050 93.600 ;
        RECT 745.950 91.950 748.050 92.400 ;
        RECT 781.950 91.950 784.050 92.400 ;
        RECT 136.950 90.600 139.050 91.050 ;
        RECT 223.950 90.600 226.050 91.050 ;
        RECT 136.950 89.400 226.050 90.600 ;
        RECT 136.950 88.950 139.050 89.400 ;
        RECT 223.950 88.950 226.050 89.400 ;
        RECT 295.950 90.600 298.050 91.050 ;
        RECT 319.950 90.600 322.050 91.050 ;
        RECT 362.400 90.600 363.600 91.950 ;
        RECT 295.950 89.400 363.600 90.600 ;
        RECT 445.950 90.600 448.050 91.050 ;
        RECT 469.950 90.600 472.050 91.050 ;
        RECT 445.950 89.400 472.050 90.600 ;
        RECT 295.950 88.950 298.050 89.400 ;
        RECT 319.950 88.950 322.050 89.400 ;
        RECT 445.950 88.950 448.050 89.400 ;
        RECT 469.950 88.950 472.050 89.400 ;
        RECT 505.950 90.600 508.050 91.050 ;
        RECT 517.950 90.600 520.050 91.050 ;
        RECT 523.950 90.600 526.050 91.050 ;
        RECT 505.950 89.400 526.050 90.600 ;
        RECT 505.950 88.950 508.050 89.400 ;
        RECT 517.950 88.950 520.050 89.400 ;
        RECT 523.950 88.950 526.050 89.400 ;
        RECT 613.950 90.600 616.050 91.050 ;
        RECT 688.950 90.600 691.050 91.050 ;
        RECT 613.950 89.400 691.050 90.600 ;
        RECT 613.950 88.950 616.050 89.400 ;
        RECT 688.950 88.950 691.050 89.400 ;
        RECT 787.950 90.600 790.050 91.050 ;
        RECT 835.950 90.600 838.050 91.050 ;
        RECT 847.950 90.600 850.050 91.050 ;
        RECT 787.950 89.400 850.050 90.600 ;
        RECT 787.950 88.950 790.050 89.400 ;
        RECT 835.950 88.950 838.050 89.400 ;
        RECT 847.950 88.950 850.050 89.400 ;
        RECT 40.950 87.600 43.050 88.050 ;
        RECT 88.950 87.600 91.050 88.050 ;
        RECT 40.950 86.400 91.050 87.600 ;
        RECT 40.950 85.950 43.050 86.400 ;
        RECT 88.950 85.950 91.050 86.400 ;
        RECT 124.950 87.600 127.050 88.050 ;
        RECT 142.950 87.600 145.050 88.050 ;
        RECT 160.950 87.600 163.050 88.050 ;
        RECT 124.950 86.400 163.050 87.600 ;
        RECT 124.950 85.950 127.050 86.400 ;
        RECT 142.950 85.950 145.050 86.400 ;
        RECT 160.950 85.950 163.050 86.400 ;
        RECT 247.950 87.600 250.050 88.050 ;
        RECT 283.950 87.600 286.050 88.050 ;
        RECT 247.950 86.400 286.050 87.600 ;
        RECT 247.950 85.950 250.050 86.400 ;
        RECT 283.950 85.950 286.050 86.400 ;
        RECT 409.950 87.600 412.050 88.050 ;
        RECT 442.950 87.600 445.050 88.050 ;
        RECT 409.950 86.400 445.050 87.600 ;
        RECT 409.950 85.950 412.050 86.400 ;
        RECT 442.950 85.950 445.050 86.400 ;
        RECT 622.950 87.600 625.050 88.050 ;
        RECT 670.950 87.600 673.050 88.050 ;
        RECT 622.950 86.400 673.050 87.600 ;
        RECT 622.950 85.950 625.050 86.400 ;
        RECT 670.950 85.950 673.050 86.400 ;
        RECT 709.950 87.600 712.050 88.050 ;
        RECT 748.950 87.600 751.050 88.050 ;
        RECT 709.950 86.400 751.050 87.600 ;
        RECT 709.950 85.950 712.050 86.400 ;
        RECT 748.950 85.950 751.050 86.400 ;
        RECT 817.950 87.600 820.050 88.050 ;
        RECT 880.950 87.600 883.050 88.050 ;
        RECT 817.950 86.400 883.050 87.600 ;
        RECT 817.950 85.950 820.050 86.400 ;
        RECT 880.950 85.950 883.050 86.400 ;
        RECT 241.950 84.600 244.050 85.050 ;
        RECT 304.950 84.600 307.050 85.050 ;
        RECT 241.950 83.400 307.050 84.600 ;
        RECT 241.950 82.950 244.050 83.400 ;
        RECT 304.950 82.950 307.050 83.400 ;
        RECT 340.950 84.600 343.050 85.050 ;
        RECT 397.950 84.600 400.050 85.050 ;
        RECT 340.950 83.400 400.050 84.600 ;
        RECT 340.950 82.950 343.050 83.400 ;
        RECT 397.950 82.950 400.050 83.400 ;
        RECT 466.950 84.600 469.050 85.050 ;
        RECT 505.950 84.600 508.050 85.050 ;
        RECT 466.950 83.400 508.050 84.600 ;
        RECT 466.950 82.950 469.050 83.400 ;
        RECT 505.950 82.950 508.050 83.400 ;
        RECT 688.950 84.600 691.050 85.050 ;
        RECT 751.950 84.600 754.050 85.050 ;
        RECT 688.950 83.400 754.050 84.600 ;
        RECT 688.950 82.950 691.050 83.400 ;
        RECT 751.950 82.950 754.050 83.400 ;
        RECT 823.950 84.600 826.050 85.050 ;
        RECT 856.950 84.600 859.050 85.050 ;
        RECT 823.950 83.400 859.050 84.600 ;
        RECT 823.950 82.950 826.050 83.400 ;
        RECT 856.950 82.950 859.050 83.400 ;
        RECT 130.950 81.600 133.050 82.050 ;
        RECT 181.950 81.600 184.050 82.050 ;
        RECT 130.950 80.400 184.050 81.600 ;
        RECT 130.950 79.950 133.050 80.400 ;
        RECT 181.950 79.950 184.050 80.400 ;
        RECT 271.950 81.600 274.050 82.050 ;
        RECT 301.950 81.600 304.050 82.050 ;
        RECT 271.950 80.400 304.050 81.600 ;
        RECT 271.950 79.950 274.050 80.400 ;
        RECT 301.950 79.950 304.050 80.400 ;
        RECT 352.950 81.600 355.050 82.050 ;
        RECT 385.950 81.600 388.050 82.050 ;
        RECT 352.950 80.400 388.050 81.600 ;
        RECT 352.950 79.950 355.050 80.400 ;
        RECT 385.950 79.950 388.050 80.400 ;
        RECT 685.950 81.600 688.050 82.050 ;
        RECT 853.950 81.600 856.050 82.050 ;
        RECT 685.950 80.400 856.050 81.600 ;
        RECT 685.950 79.950 688.050 80.400 ;
        RECT 853.950 79.950 856.050 80.400 ;
        RECT 865.950 81.600 868.050 82.050 ;
        RECT 889.950 81.600 892.050 82.050 ;
        RECT 865.950 80.400 892.050 81.600 ;
        RECT 865.950 79.950 868.050 80.400 ;
        RECT 889.950 79.950 892.050 80.400 ;
        RECT 148.950 78.600 151.050 79.050 ;
        RECT 163.950 78.600 166.050 79.050 ;
        RECT 169.950 78.600 172.050 79.050 ;
        RECT 148.950 77.400 172.050 78.600 ;
        RECT 148.950 76.950 151.050 77.400 ;
        RECT 163.950 76.950 166.050 77.400 ;
        RECT 169.950 76.950 172.050 77.400 ;
        RECT 304.950 78.600 307.050 79.050 ;
        RECT 397.950 78.600 400.050 79.050 ;
        RECT 505.950 78.600 508.050 79.050 ;
        RECT 304.950 77.400 508.050 78.600 ;
        RECT 304.950 76.950 307.050 77.400 ;
        RECT 397.950 76.950 400.050 77.400 ;
        RECT 505.950 76.950 508.050 77.400 ;
        RECT 553.950 78.600 556.050 79.050 ;
        RECT 616.950 78.600 619.050 79.050 ;
        RECT 655.950 78.600 658.050 79.050 ;
        RECT 553.950 77.400 658.050 78.600 ;
        RECT 553.950 76.950 556.050 77.400 ;
        RECT 616.950 76.950 619.050 77.400 ;
        RECT 655.950 76.950 658.050 77.400 ;
        RECT 61.950 75.600 64.050 76.050 ;
        RECT 82.950 75.600 85.050 76.050 ;
        RECT 142.950 75.600 145.050 76.050 ;
        RECT 61.950 74.400 145.050 75.600 ;
        RECT 61.950 73.950 64.050 74.400 ;
        RECT 82.950 73.950 85.050 74.400 ;
        RECT 142.950 73.950 145.050 74.400 ;
        RECT 154.950 75.600 157.050 76.050 ;
        RECT 175.950 75.600 178.050 76.050 ;
        RECT 154.950 74.400 178.050 75.600 ;
        RECT 154.950 73.950 157.050 74.400 ;
        RECT 175.950 73.950 178.050 74.400 ;
        RECT 205.950 75.600 208.050 76.050 ;
        RECT 253.950 75.600 256.050 76.050 ;
        RECT 205.950 74.400 256.050 75.600 ;
        RECT 205.950 73.950 208.050 74.400 ;
        RECT 253.950 73.950 256.050 74.400 ;
        RECT 673.950 75.600 676.050 76.050 ;
        RECT 772.950 75.600 775.050 76.050 ;
        RECT 673.950 74.400 775.050 75.600 ;
        RECT 673.950 73.950 676.050 74.400 ;
        RECT 772.950 73.950 775.050 74.400 ;
        RECT 805.950 75.600 808.050 76.050 ;
        RECT 811.950 75.600 814.050 76.050 ;
        RECT 805.950 74.400 814.050 75.600 ;
        RECT 805.950 73.950 808.050 74.400 ;
        RECT 811.950 73.950 814.050 74.400 ;
        RECT 865.950 75.600 868.050 76.050 ;
        RECT 901.950 75.600 904.050 76.050 ;
        RECT 916.950 75.600 919.050 76.050 ;
        RECT 865.950 74.400 919.050 75.600 ;
        RECT 865.950 73.950 868.050 74.400 ;
        RECT 901.950 73.950 904.050 74.400 ;
        RECT 916.950 73.950 919.050 74.400 ;
        RECT 16.950 72.600 19.050 73.050 ;
        RECT 37.950 72.600 40.050 73.050 ;
        RECT 118.950 72.600 121.050 73.050 ;
        RECT 16.950 71.400 121.050 72.600 ;
        RECT 16.950 70.950 19.050 71.400 ;
        RECT 37.950 70.950 40.050 71.400 ;
        RECT 118.950 70.950 121.050 71.400 ;
        RECT 277.950 72.600 280.050 73.050 ;
        RECT 352.950 72.600 355.050 73.050 ;
        RECT 277.950 71.400 355.050 72.600 ;
        RECT 277.950 70.950 280.050 71.400 ;
        RECT 352.950 70.950 355.050 71.400 ;
        RECT 520.950 72.600 523.050 73.050 ;
        RECT 553.950 72.600 556.050 73.050 ;
        RECT 520.950 71.400 556.050 72.600 ;
        RECT 520.950 70.950 523.050 71.400 ;
        RECT 553.950 70.950 556.050 71.400 ;
        RECT 646.950 72.600 649.050 73.050 ;
        RECT 745.950 72.600 748.050 73.050 ;
        RECT 646.950 71.400 748.050 72.600 ;
        RECT 646.950 70.950 649.050 71.400 ;
        RECT 745.950 70.950 748.050 71.400 ;
        RECT 838.950 72.600 841.050 73.050 ;
        RECT 868.950 72.600 871.050 73.050 ;
        RECT 838.950 71.400 871.050 72.600 ;
        RECT 838.950 70.950 841.050 71.400 ;
        RECT 868.950 70.950 871.050 71.400 ;
        RECT 127.950 69.600 130.050 70.050 ;
        RECT 133.950 69.600 136.050 70.050 ;
        RECT 139.950 69.600 142.050 70.050 ;
        RECT 127.950 68.400 142.050 69.600 ;
        RECT 127.950 67.950 130.050 68.400 ;
        RECT 133.950 67.950 136.050 68.400 ;
        RECT 139.950 67.950 142.050 68.400 ;
        RECT 175.950 69.600 178.050 70.050 ;
        RECT 190.950 69.600 193.050 70.050 ;
        RECT 211.950 69.600 214.050 70.050 ;
        RECT 175.950 68.400 214.050 69.600 ;
        RECT 175.950 67.950 178.050 68.400 ;
        RECT 190.950 67.950 193.050 68.400 ;
        RECT 211.950 67.950 214.050 68.400 ;
        RECT 256.950 69.600 259.050 70.050 ;
        RECT 271.950 69.600 274.050 70.050 ;
        RECT 256.950 68.400 274.050 69.600 ;
        RECT 256.950 67.950 259.050 68.400 ;
        RECT 271.950 67.950 274.050 68.400 ;
        RECT 412.950 69.600 415.050 70.050 ;
        RECT 478.950 69.600 481.050 70.050 ;
        RECT 412.950 68.400 481.050 69.600 ;
        RECT 412.950 67.950 415.050 68.400 ;
        RECT 478.950 67.950 481.050 68.400 ;
        RECT 490.950 69.600 493.050 70.050 ;
        RECT 535.950 69.600 538.050 70.050 ;
        RECT 490.950 68.400 538.050 69.600 ;
        RECT 490.950 67.950 493.050 68.400 ;
        RECT 535.950 67.950 538.050 68.400 ;
        RECT 565.950 69.600 568.050 70.050 ;
        RECT 652.950 69.600 655.050 70.050 ;
        RECT 565.950 68.400 655.050 69.600 ;
        RECT 565.950 67.950 568.050 68.400 ;
        RECT 652.950 67.950 655.050 68.400 ;
        RECT 832.950 69.600 835.050 70.050 ;
        RECT 859.950 69.600 862.050 70.050 ;
        RECT 832.950 68.400 862.050 69.600 ;
        RECT 832.950 67.950 835.050 68.400 ;
        RECT 859.950 67.950 862.050 68.400 ;
        RECT 73.950 66.600 76.050 67.050 ;
        RECT 91.950 66.600 94.050 67.050 ;
        RECT 73.950 65.400 94.050 66.600 ;
        RECT 73.950 64.950 76.050 65.400 ;
        RECT 91.950 64.950 94.050 65.400 ;
        RECT 235.950 66.600 238.050 67.050 ;
        RECT 295.950 66.600 298.050 67.050 ;
        RECT 235.950 65.400 298.050 66.600 ;
        RECT 235.950 64.950 238.050 65.400 ;
        RECT 295.950 64.950 298.050 65.400 ;
        RECT 355.950 66.600 358.050 67.050 ;
        RECT 367.950 66.600 370.050 67.050 ;
        RECT 355.950 65.400 370.050 66.600 ;
        RECT 355.950 64.950 358.050 65.400 ;
        RECT 367.950 64.950 370.050 65.400 ;
        RECT 391.950 66.600 394.050 67.050 ;
        RECT 424.950 66.600 427.050 67.050 ;
        RECT 427.950 66.600 430.050 67.050 ;
        RECT 451.950 66.600 454.050 67.050 ;
        RECT 391.950 65.400 454.050 66.600 ;
        RECT 391.950 64.950 394.050 65.400 ;
        RECT 424.950 64.950 427.050 65.400 ;
        RECT 427.950 64.950 430.050 65.400 ;
        RECT 451.950 64.950 454.050 65.400 ;
        RECT 460.950 66.600 463.050 67.050 ;
        RECT 481.950 66.600 484.050 67.050 ;
        RECT 460.950 65.400 484.050 66.600 ;
        RECT 460.950 64.950 463.050 65.400 ;
        RECT 481.950 64.950 484.050 65.400 ;
        RECT 571.950 66.600 574.050 67.050 ;
        RECT 595.950 66.600 598.050 67.050 ;
        RECT 622.950 66.600 625.050 67.050 ;
        RECT 571.950 65.400 625.050 66.600 ;
        RECT 571.950 64.950 574.050 65.400 ;
        RECT 595.950 64.950 598.050 65.400 ;
        RECT 622.950 64.950 625.050 65.400 ;
        RECT 757.950 66.600 760.050 67.050 ;
        RECT 772.950 66.600 775.050 67.050 ;
        RECT 757.950 65.400 775.050 66.600 ;
        RECT 757.950 64.950 760.050 65.400 ;
        RECT 772.950 64.950 775.050 65.400 ;
        RECT 889.950 66.600 892.050 67.050 ;
        RECT 910.950 66.600 913.050 67.050 ;
        RECT 889.950 65.400 913.050 66.600 ;
        RECT 889.950 64.950 892.050 65.400 ;
        RECT 910.950 64.950 913.050 65.400 ;
        RECT 22.950 63.600 25.050 64.050 ;
        RECT 31.950 63.600 34.050 64.050 ;
        RECT 46.950 63.600 49.050 64.050 ;
        RECT 208.950 63.600 211.050 64.050 ;
        RECT 22.950 62.400 49.050 63.600 ;
        RECT 22.950 61.950 25.050 62.400 ;
        RECT 31.950 61.950 34.050 62.400 ;
        RECT 46.950 61.950 49.050 62.400 ;
        RECT 176.400 62.400 211.050 63.600 ;
        RECT 28.950 60.600 31.050 61.050 ;
        RECT 76.950 60.600 79.050 61.200 ;
        RECT 23.400 59.400 31.050 60.600 ;
        RECT 19.950 54.600 22.050 54.900 ;
        RECT 23.400 54.600 24.600 59.400 ;
        RECT 28.950 58.950 31.050 59.400 ;
        RECT 65.400 59.400 79.050 60.600 ;
        RECT 65.400 54.900 66.600 59.400 ;
        RECT 76.950 59.100 79.050 59.400 ;
        RECT 94.950 60.750 97.050 61.200 ;
        RECT 103.950 60.750 106.050 61.200 ;
        RECT 94.950 59.550 106.050 60.750 ;
        RECT 94.950 59.100 97.050 59.550 ;
        RECT 103.950 59.100 106.050 59.550 ;
        RECT 109.950 59.100 112.050 61.200 ;
        RECT 19.950 53.400 24.600 54.600 ;
        RECT 19.950 52.800 22.050 53.400 ;
        RECT 64.950 52.800 67.050 54.900 ;
        RECT 85.950 54.600 88.050 54.900 ;
        RECT 94.950 54.600 97.050 55.050 ;
        RECT 85.950 53.400 97.050 54.600 ;
        RECT 85.950 52.800 88.050 53.400 ;
        RECT 94.950 52.950 97.050 53.400 ;
        RECT 100.950 54.600 103.050 55.050 ;
        RECT 110.400 54.600 111.600 59.100 ;
        RECT 166.950 58.950 169.050 61.050 ;
        RECT 167.400 55.050 168.600 58.950 ;
        RECT 176.400 57.600 177.600 62.400 ;
        RECT 208.950 61.950 211.050 62.400 ;
        RECT 180.000 60.600 184.050 61.050 ;
        RECT 173.400 56.400 177.600 57.600 ;
        RECT 179.400 58.950 184.050 60.600 ;
        RECT 196.950 60.750 199.050 61.200 ;
        RECT 220.950 60.750 223.050 61.200 ;
        RECT 196.950 59.550 223.050 60.750 ;
        RECT 247.950 60.600 250.050 61.200 ;
        RECT 196.950 59.100 199.050 59.550 ;
        RECT 220.950 59.100 223.050 59.550 ;
        RECT 233.400 59.400 250.050 60.600 ;
        RECT 100.950 53.400 111.600 54.600 ;
        RECT 118.950 54.600 121.050 55.050 ;
        RECT 124.950 54.600 127.050 54.900 ;
        RECT 118.950 53.400 127.050 54.600 ;
        RECT 100.950 52.950 103.050 53.400 ;
        RECT 118.950 52.950 121.050 53.400 ;
        RECT 124.950 52.800 127.050 53.400 ;
        RECT 142.950 54.600 145.050 55.050 ;
        RECT 151.950 54.600 154.050 54.900 ;
        RECT 142.950 53.400 154.050 54.600 ;
        RECT 142.950 52.950 145.050 53.400 ;
        RECT 151.950 52.800 154.050 53.400 ;
        RECT 166.950 52.950 169.050 55.050 ;
        RECT 173.400 54.900 174.600 56.400 ;
        RECT 179.400 54.900 180.600 58.950 ;
        RECT 211.950 57.600 214.050 58.050 ;
        RECT 233.400 57.600 234.600 59.400 ;
        RECT 247.950 59.100 250.050 59.400 ;
        RECT 259.950 60.750 262.050 61.200 ;
        RECT 265.950 60.750 268.050 61.200 ;
        RECT 259.950 59.550 268.050 60.750 ;
        RECT 259.950 59.100 262.050 59.550 ;
        RECT 265.950 59.100 268.050 59.550 ;
        RECT 277.950 60.600 280.050 61.200 ;
        RECT 289.950 60.600 292.050 61.200 ;
        RECT 277.950 59.400 292.050 60.600 ;
        RECT 277.950 59.100 280.050 59.400 ;
        RECT 289.950 59.100 292.050 59.400 ;
        RECT 307.950 60.750 310.050 61.200 ;
        RECT 331.950 60.750 334.050 64.050 ;
        RECT 368.400 63.600 369.600 64.950 ;
        RECT 457.950 63.600 460.050 64.050 ;
        RECT 472.950 63.600 475.050 64.050 ;
        RECT 368.400 62.400 475.050 63.600 ;
        RECT 457.950 61.950 460.050 62.400 ;
        RECT 472.950 61.950 475.050 62.400 ;
        RECT 487.950 63.600 490.050 64.050 ;
        RECT 493.950 63.600 496.050 64.050 ;
        RECT 487.950 62.400 496.050 63.600 ;
        RECT 487.950 61.950 490.050 62.400 ;
        RECT 493.950 61.950 496.050 62.400 ;
        RECT 529.950 63.600 532.050 64.050 ;
        RECT 544.950 63.600 547.050 64.050 ;
        RECT 556.950 63.600 559.050 64.050 ;
        RECT 529.950 62.400 559.050 63.600 ;
        RECT 529.950 61.950 532.050 62.400 ;
        RECT 544.950 61.950 547.050 62.400 ;
        RECT 556.950 61.950 559.050 62.400 ;
        RECT 658.950 63.600 661.050 64.050 ;
        RECT 706.950 63.600 709.050 64.050 ;
        RECT 658.950 62.400 709.050 63.600 ;
        RECT 658.950 61.950 661.050 62.400 ;
        RECT 706.950 61.950 709.050 62.400 ;
        RECT 754.950 61.950 757.050 64.050 ;
        RECT 814.950 63.600 817.050 64.050 ;
        RECT 823.950 63.600 826.050 64.050 ;
        RECT 841.950 63.600 844.050 64.050 ;
        RECT 814.950 62.400 844.050 63.600 ;
        RECT 814.950 61.950 817.050 62.400 ;
        RECT 823.950 61.950 826.050 62.400 ;
        RECT 841.950 61.950 844.050 62.400 ;
        RECT 871.950 63.600 874.050 64.050 ;
        RECT 880.950 63.600 883.050 64.050 ;
        RECT 871.950 62.400 883.050 63.600 ;
        RECT 871.950 61.950 874.050 62.400 ;
        RECT 880.950 61.950 883.050 62.400 ;
        RECT 334.950 60.750 337.050 61.200 ;
        RECT 307.950 59.550 337.050 60.750 ;
        RECT 307.950 59.100 310.050 59.550 ;
        RECT 332.400 59.400 333.600 59.550 ;
        RECT 334.950 59.100 337.050 59.550 ;
        RECT 361.950 59.100 364.050 61.200 ;
        RECT 385.950 60.600 388.050 61.200 ;
        RECT 412.950 60.600 415.050 61.200 ;
        RECT 385.950 59.400 415.050 60.600 ;
        RECT 385.950 59.100 388.050 59.400 ;
        RECT 412.950 59.100 415.050 59.400 ;
        RECT 484.950 60.750 487.050 61.200 ;
        RECT 511.950 60.750 514.050 61.200 ;
        RECT 484.950 59.550 514.050 60.750 ;
        RECT 484.950 59.100 487.050 59.550 ;
        RECT 511.950 59.100 514.050 59.550 ;
        RECT 562.950 60.750 565.050 61.200 ;
        RECT 577.950 60.750 580.050 61.200 ;
        RECT 562.950 60.600 580.050 60.750 ;
        RECT 589.950 60.600 592.050 61.200 ;
        RECT 562.950 59.550 592.050 60.600 ;
        RECT 562.950 59.100 565.050 59.550 ;
        RECT 577.950 59.400 592.050 59.550 ;
        RECT 577.950 59.100 580.050 59.400 ;
        RECT 589.950 59.100 592.050 59.400 ;
        RECT 604.950 60.600 607.050 61.050 ;
        RECT 616.950 60.600 619.050 61.200 ;
        RECT 631.950 60.600 634.050 61.200 ;
        RECT 604.950 59.400 634.050 60.600 ;
        RECT 211.950 56.400 234.600 57.600 ;
        RECT 290.400 57.600 291.600 59.100 ;
        RECT 362.400 57.600 363.600 59.100 ;
        RECT 604.950 58.950 607.050 59.400 ;
        RECT 616.950 59.100 619.050 59.400 ;
        RECT 631.950 59.100 634.050 59.400 ;
        RECT 664.950 60.600 667.050 61.200 ;
        RECT 679.950 60.600 682.050 61.200 ;
        RECT 664.950 59.400 682.050 60.600 ;
        RECT 715.950 61.050 718.050 61.500 ;
        RECT 727.950 61.050 730.050 61.500 ;
        RECT 715.950 59.850 730.050 61.050 ;
        RECT 715.950 59.400 718.050 59.850 ;
        RECT 727.950 59.400 730.050 59.850 ;
        RECT 664.950 59.100 667.050 59.400 ;
        RECT 679.950 59.100 682.050 59.400 ;
        RECT 418.950 57.600 421.050 58.050 ;
        RECT 445.950 57.600 448.050 58.050 ;
        RECT 290.400 56.400 411.600 57.600 ;
        RECT 211.950 55.950 214.050 56.400 ;
        RECT 172.950 52.800 175.050 54.900 ;
        RECT 178.950 54.600 181.050 54.900 ;
        RECT 187.950 54.600 190.050 54.900 ;
        RECT 178.950 53.400 190.050 54.600 ;
        RECT 178.950 52.800 181.050 53.400 ;
        RECT 187.950 52.800 190.050 53.400 ;
        RECT 274.950 54.600 277.050 54.900 ;
        RECT 292.950 54.600 295.050 54.900 ;
        RECT 274.950 53.400 295.050 54.600 ;
        RECT 296.400 54.600 297.600 56.400 ;
        RECT 313.950 54.600 316.050 54.900 ;
        RECT 296.400 53.400 316.050 54.600 ;
        RECT 274.950 52.800 277.050 53.400 ;
        RECT 292.950 52.800 295.050 53.400 ;
        RECT 313.950 52.800 316.050 53.400 ;
        RECT 319.950 54.450 322.050 54.900 ;
        RECT 325.800 54.450 327.900 54.900 ;
        RECT 319.950 53.250 327.900 54.450 ;
        RECT 319.950 52.800 322.050 53.250 ;
        RECT 325.800 52.800 327.900 53.250 ;
        RECT 328.950 54.450 331.050 54.900 ;
        RECT 337.950 54.450 340.050 54.900 ;
        RECT 328.950 53.250 340.050 54.450 ;
        RECT 328.950 52.800 331.050 53.250 ;
        RECT 337.950 52.800 340.050 53.250 ;
        RECT 343.950 54.600 346.050 54.900 ;
        RECT 355.950 54.600 358.050 55.050 ;
        RECT 343.950 53.400 358.050 54.600 ;
        RECT 343.950 52.800 346.050 53.400 ;
        RECT 355.950 52.950 358.050 53.400 ;
        RECT 370.950 54.600 373.050 54.900 ;
        RECT 382.950 54.600 385.050 54.900 ;
        RECT 391.950 54.600 394.050 55.050 ;
        RECT 370.950 53.400 394.050 54.600 ;
        RECT 370.950 52.800 373.050 53.400 ;
        RECT 382.950 52.800 385.050 53.400 ;
        RECT 391.950 52.950 394.050 53.400 ;
        RECT 397.950 54.600 400.050 55.050 ;
        RECT 410.400 54.900 411.600 56.400 ;
        RECT 418.950 56.400 448.050 57.600 ;
        RECT 418.950 55.950 421.050 56.400 ;
        RECT 445.950 55.950 448.050 56.400 ;
        RECT 403.950 54.600 406.050 54.900 ;
        RECT 397.950 53.400 406.050 54.600 ;
        RECT 397.950 52.950 400.050 53.400 ;
        RECT 403.950 52.800 406.050 53.400 ;
        RECT 409.950 54.600 412.050 54.900 ;
        RECT 427.950 54.600 430.050 54.900 ;
        RECT 409.950 53.400 430.050 54.600 ;
        RECT 409.950 52.800 412.050 53.400 ;
        RECT 427.950 52.800 430.050 53.400 ;
        RECT 454.950 54.600 457.050 54.900 ;
        RECT 484.950 54.600 487.050 55.050 ;
        RECT 454.950 53.400 487.050 54.600 ;
        RECT 454.950 52.800 457.050 53.400 ;
        RECT 484.950 52.950 487.050 53.400 ;
        RECT 508.950 54.450 511.050 54.900 ;
        RECT 520.950 54.450 523.050 54.900 ;
        RECT 508.950 53.250 523.050 54.450 ;
        RECT 508.950 52.800 511.050 53.250 ;
        RECT 520.950 52.800 523.050 53.250 ;
        RECT 544.950 54.450 547.050 54.900 ;
        RECT 550.950 54.450 553.050 54.900 ;
        RECT 544.950 53.250 553.050 54.450 ;
        RECT 544.950 52.800 547.050 53.250 ;
        RECT 550.950 52.800 553.050 53.250 ;
        RECT 598.950 54.600 601.050 54.900 ;
        RECT 628.950 54.600 631.050 54.900 ;
        RECT 598.950 53.400 631.050 54.600 ;
        RECT 598.950 52.800 601.050 53.400 ;
        RECT 628.950 52.800 631.050 53.400 ;
        RECT 634.950 54.600 637.050 54.900 ;
        RECT 646.950 54.600 649.050 55.050 ;
        RECT 755.400 54.900 756.600 61.950 ;
        RECT 763.950 60.600 766.050 61.200 ;
        RECT 778.950 60.600 781.050 61.200 ;
        RECT 852.000 60.600 856.050 61.050 ;
        RECT 763.950 59.400 781.050 60.600 ;
        RECT 763.950 59.100 766.050 59.400 ;
        RECT 778.950 59.100 781.050 59.400 ;
        RECT 851.400 58.950 856.050 60.600 ;
        RECT 895.950 60.750 898.050 61.200 ;
        RECT 913.950 60.750 916.050 61.200 ;
        RECT 895.950 59.550 916.050 60.750 ;
        RECT 895.950 59.100 898.050 59.550 ;
        RECT 913.950 59.100 916.050 59.550 ;
        RECT 838.950 57.600 841.050 58.050 ;
        RECT 788.400 56.400 841.050 57.600 ;
        RECT 634.950 53.400 649.050 54.600 ;
        RECT 634.950 52.800 637.050 53.400 ;
        RECT 646.950 52.950 649.050 53.400 ;
        RECT 682.950 54.600 685.050 54.900 ;
        RECT 682.950 53.400 691.050 54.600 ;
        RECT 682.950 52.800 685.050 53.400 ;
        RECT 688.950 52.500 691.050 53.400 ;
        RECT 754.950 52.800 757.050 54.900 ;
        RECT 788.400 54.600 789.600 56.400 ;
        RECT 838.950 55.950 841.050 56.400 ;
        RECT 851.400 54.600 852.600 58.950 ;
        RECT 787.950 52.500 790.050 54.600 ;
        RECT 850.950 52.500 853.050 54.600 ;
        RECT 865.950 54.450 868.050 54.900 ;
        RECT 880.950 54.450 883.050 54.900 ;
        RECT 865.950 53.250 883.050 54.450 ;
        RECT 865.950 52.800 868.050 53.250 ;
        RECT 880.950 52.800 883.050 53.250 ;
        RECT 886.950 54.450 889.050 54.900 ;
        RECT 904.950 54.450 907.050 54.900 ;
        RECT 886.950 53.250 907.050 54.450 ;
        RECT 886.950 52.800 889.050 53.250 ;
        RECT 904.950 52.800 907.050 53.250 ;
        RECT 97.950 51.600 100.050 52.050 ;
        RECT 106.950 51.600 109.050 52.050 ;
        RECT 97.950 50.400 109.050 51.600 ;
        RECT 97.950 49.950 100.050 50.400 ;
        RECT 106.950 49.950 109.050 50.400 ;
        RECT 208.950 51.600 211.050 52.050 ;
        RECT 259.950 51.600 262.050 52.050 ;
        RECT 208.950 50.400 262.050 51.600 ;
        RECT 208.950 49.950 211.050 50.400 ;
        RECT 259.950 49.950 262.050 50.400 ;
        RECT 292.950 51.600 295.050 52.050 ;
        RECT 304.950 51.600 307.050 52.050 ;
        RECT 292.950 50.400 307.050 51.600 ;
        RECT 292.950 49.950 295.050 50.400 ;
        RECT 304.950 49.950 307.050 50.400 ;
        RECT 412.950 51.600 415.050 52.050 ;
        RECT 418.950 51.600 421.050 52.050 ;
        RECT 412.950 50.400 421.050 51.600 ;
        RECT 412.950 49.950 415.050 50.400 ;
        RECT 418.950 49.950 421.050 50.400 ;
        RECT 460.950 51.600 463.050 52.050 ;
        RECT 469.950 51.600 472.050 52.050 ;
        RECT 481.950 51.600 484.050 52.050 ;
        RECT 460.950 50.400 484.050 51.600 ;
        RECT 460.950 49.950 463.050 50.400 ;
        RECT 469.950 49.950 472.050 50.400 ;
        RECT 481.950 49.950 484.050 50.400 ;
        RECT 553.950 51.600 556.050 52.050 ;
        RECT 574.950 51.600 577.050 52.050 ;
        RECT 592.950 51.600 595.050 52.050 ;
        RECT 553.950 50.400 595.050 51.600 ;
        RECT 553.950 49.950 556.050 50.400 ;
        RECT 574.950 49.950 577.050 50.400 ;
        RECT 592.950 49.950 595.050 50.400 ;
        RECT 661.950 51.600 664.050 52.050 ;
        RECT 721.950 51.600 724.050 52.050 ;
        RECT 760.950 51.600 763.050 52.050 ;
        RECT 769.950 51.600 772.050 52.050 ;
        RECT 661.950 50.400 772.050 51.600 ;
        RECT 661.950 49.950 664.050 50.400 ;
        RECT 721.950 49.950 724.050 50.400 ;
        RECT 760.950 49.950 763.050 50.400 ;
        RECT 769.950 49.950 772.050 50.400 ;
        RECT 34.950 48.600 37.050 49.050 ;
        RECT 46.950 48.600 49.050 49.050 ;
        RECT 34.950 47.400 49.050 48.600 ;
        RECT 34.950 46.950 37.050 47.400 ;
        RECT 46.950 46.950 49.050 47.400 ;
        RECT 58.950 48.600 61.050 49.050 ;
        RECT 100.950 48.600 103.050 49.050 ;
        RECT 121.950 48.600 124.050 49.050 ;
        RECT 58.950 47.400 124.050 48.600 ;
        RECT 58.950 46.950 61.050 47.400 ;
        RECT 100.950 46.950 103.050 47.400 ;
        RECT 121.950 46.950 124.050 47.400 ;
        RECT 139.950 48.600 142.050 49.050 ;
        RECT 166.950 48.600 169.050 49.050 ;
        RECT 139.950 47.400 169.050 48.600 ;
        RECT 139.950 46.950 142.050 47.400 ;
        RECT 166.950 46.950 169.050 47.400 ;
        RECT 190.950 48.600 193.050 49.050 ;
        RECT 205.950 48.600 208.050 49.050 ;
        RECT 190.950 47.400 208.050 48.600 ;
        RECT 190.950 46.950 193.050 47.400 ;
        RECT 205.950 46.950 208.050 47.400 ;
        RECT 310.950 48.600 313.050 49.050 ;
        RECT 424.950 48.600 427.050 49.050 ;
        RECT 310.950 47.400 427.050 48.600 ;
        RECT 310.950 46.950 313.050 47.400 ;
        RECT 424.950 46.950 427.050 47.400 ;
        RECT 475.950 48.600 478.050 49.050 ;
        RECT 484.950 48.600 487.050 49.050 ;
        RECT 475.950 47.400 487.050 48.600 ;
        RECT 475.950 46.950 478.050 47.400 ;
        RECT 484.950 46.950 487.050 47.400 ;
        RECT 496.950 48.600 499.050 49.050 ;
        RECT 502.950 48.600 505.050 49.050 ;
        RECT 514.950 48.600 517.050 49.050 ;
        RECT 547.950 48.600 550.050 49.050 ;
        RECT 562.950 48.600 565.050 49.050 ;
        RECT 496.950 47.400 565.050 48.600 ;
        RECT 496.950 46.950 499.050 47.400 ;
        RECT 502.950 46.950 505.050 47.400 ;
        RECT 514.950 46.950 517.050 47.400 ;
        RECT 547.950 46.950 550.050 47.400 ;
        RECT 562.950 46.950 565.050 47.400 ;
        RECT 589.950 48.600 592.050 49.050 ;
        RECT 607.950 48.600 610.050 49.050 ;
        RECT 589.950 47.400 610.050 48.600 ;
        RECT 589.950 46.950 592.050 47.400 ;
        RECT 607.950 46.950 610.050 47.400 ;
        RECT 655.950 48.600 658.050 49.050 ;
        RECT 700.950 48.600 703.050 49.050 ;
        RECT 655.950 47.400 703.050 48.600 ;
        RECT 655.950 46.950 658.050 47.400 ;
        RECT 700.950 46.950 703.050 47.400 ;
        RECT 892.950 48.600 895.050 49.050 ;
        RECT 901.950 48.600 904.050 49.050 ;
        RECT 892.950 47.400 904.050 48.600 ;
        RECT 892.950 46.950 895.050 47.400 ;
        RECT 901.950 46.950 904.050 47.400 ;
        RECT 79.950 45.600 82.050 46.050 ;
        RECT 91.950 45.600 94.050 46.050 ;
        RECT 79.950 44.400 94.050 45.600 ;
        RECT 79.950 43.950 82.050 44.400 ;
        RECT 91.950 43.950 94.050 44.400 ;
        RECT 223.950 45.600 226.050 46.050 ;
        RECT 259.950 45.600 262.050 46.050 ;
        RECT 223.950 44.400 262.050 45.600 ;
        RECT 223.950 43.950 226.050 44.400 ;
        RECT 259.950 43.950 262.050 44.400 ;
        RECT 265.950 45.600 268.050 46.050 ;
        RECT 406.950 45.600 409.050 46.050 ;
        RECT 265.950 44.400 409.050 45.600 ;
        RECT 265.950 43.950 268.050 44.400 ;
        RECT 406.950 43.950 409.050 44.400 ;
        RECT 454.950 45.600 457.050 46.050 ;
        RECT 487.950 45.600 490.050 46.050 ;
        RECT 454.950 44.400 490.050 45.600 ;
        RECT 454.950 43.950 457.050 44.400 ;
        RECT 487.950 43.950 490.050 44.400 ;
        RECT 526.950 45.600 529.050 46.050 ;
        RECT 535.950 45.600 538.050 46.050 ;
        RECT 526.950 44.400 538.050 45.600 ;
        RECT 526.950 43.950 529.050 44.400 ;
        RECT 535.950 43.950 538.050 44.400 ;
        RECT 856.950 45.600 859.050 46.050 ;
        RECT 865.950 45.600 868.050 46.050 ;
        RECT 856.950 44.400 868.050 45.600 ;
        RECT 856.950 43.950 859.050 44.400 ;
        RECT 865.950 43.950 868.050 44.400 ;
        RECT 871.950 45.600 874.050 46.050 ;
        RECT 919.950 45.600 922.050 46.050 ;
        RECT 871.950 44.400 922.050 45.600 ;
        RECT 871.950 43.950 874.050 44.400 ;
        RECT 919.950 43.950 922.050 44.400 ;
        RECT 13.950 42.600 16.050 43.050 ;
        RECT 19.950 42.600 22.050 43.050 ;
        RECT 73.950 42.600 76.050 43.050 ;
        RECT 97.950 42.600 100.050 43.050 ;
        RECT 13.950 41.400 100.050 42.600 ;
        RECT 13.950 40.950 16.050 41.400 ;
        RECT 19.950 40.950 22.050 41.400 ;
        RECT 73.950 40.950 76.050 41.400 ;
        RECT 97.950 40.950 100.050 41.400 ;
        RECT 136.950 42.600 139.050 43.050 ;
        RECT 184.950 42.600 187.050 43.050 ;
        RECT 136.950 41.400 187.050 42.600 ;
        RECT 136.950 40.950 139.050 41.400 ;
        RECT 184.950 40.950 187.050 41.400 ;
        RECT 229.950 42.600 232.050 43.050 ;
        RECT 256.950 42.600 259.050 43.050 ;
        RECT 298.950 42.600 301.050 43.050 ;
        RECT 229.950 41.400 301.050 42.600 ;
        RECT 229.950 40.950 232.050 41.400 ;
        RECT 256.950 40.950 259.050 41.400 ;
        RECT 298.950 40.950 301.050 41.400 ;
        RECT 388.950 42.600 391.050 43.050 ;
        RECT 421.950 42.600 424.050 43.050 ;
        RECT 388.950 41.400 424.050 42.600 ;
        RECT 388.950 40.950 391.050 41.400 ;
        RECT 421.950 40.950 424.050 41.400 ;
        RECT 433.950 42.600 436.050 43.050 ;
        RECT 484.950 42.600 487.050 43.050 ;
        RECT 433.950 41.400 487.050 42.600 ;
        RECT 433.950 40.950 436.050 41.400 ;
        RECT 484.950 40.950 487.050 41.400 ;
        RECT 490.950 42.600 493.050 43.050 ;
        RECT 532.950 42.600 535.050 43.050 ;
        RECT 490.950 41.400 535.050 42.600 ;
        RECT 490.950 40.950 493.050 41.400 ;
        RECT 532.950 40.950 535.050 41.400 ;
        RECT 895.950 42.600 898.050 43.050 ;
        RECT 907.950 42.600 910.050 43.050 ;
        RECT 895.950 41.400 910.050 42.600 ;
        RECT 895.950 40.950 898.050 41.400 ;
        RECT 907.950 40.950 910.050 41.400 ;
        RECT 79.950 39.600 82.050 40.050 ;
        RECT 109.950 39.600 112.050 40.050 ;
        RECT 79.950 38.400 112.050 39.600 ;
        RECT 79.950 37.950 82.050 38.400 ;
        RECT 109.950 37.950 112.050 38.400 ;
        RECT 124.950 39.600 127.050 40.050 ;
        RECT 133.950 39.600 136.050 40.050 ;
        RECT 124.950 38.400 136.050 39.600 ;
        RECT 124.950 37.950 127.050 38.400 ;
        RECT 133.950 37.950 136.050 38.400 ;
        RECT 148.950 39.600 151.050 40.050 ;
        RECT 157.950 39.600 160.050 40.050 ;
        RECT 220.950 39.600 223.050 40.050 ;
        RECT 301.950 39.600 304.050 40.050 ;
        RECT 316.950 39.600 319.050 40.050 ;
        RECT 148.950 38.400 223.050 39.600 ;
        RECT 148.950 37.950 151.050 38.400 ;
        RECT 157.950 37.950 160.050 38.400 ;
        RECT 220.950 37.950 223.050 38.400 ;
        RECT 227.400 38.400 319.050 39.600 ;
        RECT 227.400 37.050 228.600 38.400 ;
        RECT 301.950 37.950 304.050 38.400 ;
        RECT 316.950 37.950 319.050 38.400 ;
        RECT 382.950 39.600 385.050 40.050 ;
        RECT 481.950 39.600 484.050 40.050 ;
        RECT 382.950 38.400 484.050 39.600 ;
        RECT 382.950 37.950 385.050 38.400 ;
        RECT 481.950 37.950 484.050 38.400 ;
        RECT 487.950 39.600 490.050 40.050 ;
        RECT 568.950 39.600 571.050 40.050 ;
        RECT 613.950 39.600 616.050 40.050 ;
        RECT 652.950 39.600 655.050 40.050 ;
        RECT 487.950 38.400 655.050 39.600 ;
        RECT 487.950 37.950 490.050 38.400 ;
        RECT 568.950 37.950 571.050 38.400 ;
        RECT 613.950 37.950 616.050 38.400 ;
        RECT 652.950 37.950 655.050 38.400 ;
        RECT 736.950 39.600 739.050 40.050 ;
        RECT 751.950 39.600 754.050 40.050 ;
        RECT 736.950 38.400 754.050 39.600 ;
        RECT 736.950 37.950 739.050 38.400 ;
        RECT 751.950 37.950 754.050 38.400 ;
        RECT 772.950 39.600 775.050 40.050 ;
        RECT 778.950 39.600 781.050 40.050 ;
        RECT 772.950 38.400 781.050 39.600 ;
        RECT 772.950 37.950 775.050 38.400 ;
        RECT 778.950 37.950 781.050 38.400 ;
        RECT 1.950 36.600 4.050 37.050 ;
        RECT 13.950 36.600 16.050 37.050 ;
        RECT 1.950 35.400 16.050 36.600 ;
        RECT 1.950 34.950 4.050 35.400 ;
        RECT 13.950 34.950 16.050 35.400 ;
        RECT 40.950 36.600 43.050 37.050 ;
        RECT 61.950 36.600 64.050 37.050 ;
        RECT 40.950 35.400 64.050 36.600 ;
        RECT 40.950 34.950 43.050 35.400 ;
        RECT 61.950 34.950 64.050 35.400 ;
        RECT 163.950 36.600 166.050 37.050 ;
        RECT 175.950 36.600 178.050 37.050 ;
        RECT 163.950 35.400 178.050 36.600 ;
        RECT 163.950 34.950 166.050 35.400 ;
        RECT 175.950 34.950 178.050 35.400 ;
        RECT 193.950 36.600 196.050 37.050 ;
        RECT 226.950 36.600 229.050 37.050 ;
        RECT 193.950 35.400 229.050 36.600 ;
        RECT 193.950 34.950 196.050 35.400 ;
        RECT 226.950 34.950 229.050 35.400 ;
        RECT 337.950 36.600 340.050 37.050 ;
        RECT 364.950 36.600 367.050 37.050 ;
        RECT 511.950 36.600 514.050 37.050 ;
        RECT 529.950 36.600 532.050 37.050 ;
        RECT 337.950 35.400 367.050 36.600 ;
        RECT 337.950 34.950 340.050 35.400 ;
        RECT 364.950 34.950 367.050 35.400 ;
        RECT 392.400 35.400 532.050 36.600 ;
        RECT 37.950 33.600 40.050 34.050 ;
        RECT 88.950 33.600 91.050 34.050 ;
        RECT 112.950 33.600 115.050 34.050 ;
        RECT 130.950 33.600 133.050 34.050 ;
        RECT 244.950 33.600 247.050 34.050 ;
        RECT 37.950 32.400 247.050 33.600 ;
        RECT 37.950 31.950 40.050 32.400 ;
        RECT 88.950 31.950 91.050 32.400 ;
        RECT 112.950 31.950 115.050 32.400 ;
        RECT 130.950 31.950 133.050 32.400 ;
        RECT 244.950 31.950 247.050 32.400 ;
        RECT 253.950 33.600 256.050 34.050 ;
        RECT 268.950 33.600 271.050 34.050 ;
        RECT 253.950 32.400 271.050 33.600 ;
        RECT 253.950 31.950 256.050 32.400 ;
        RECT 268.950 31.950 271.050 32.400 ;
        RECT 298.950 33.600 301.050 34.050 ;
        RECT 313.950 33.600 316.050 34.050 ;
        RECT 298.950 32.400 316.050 33.600 ;
        RECT 298.950 31.950 301.050 32.400 ;
        RECT 313.950 31.950 316.050 32.400 ;
        RECT 331.950 33.600 334.050 34.050 ;
        RECT 361.950 33.600 364.050 34.050 ;
        RECT 331.950 32.400 364.050 33.600 ;
        RECT 331.950 31.950 334.050 32.400 ;
        RECT 361.950 31.950 364.050 32.400 ;
        RECT 367.950 33.600 370.050 34.050 ;
        RECT 392.400 33.600 393.600 35.400 ;
        RECT 511.950 34.950 514.050 35.400 ;
        RECT 529.950 34.950 532.050 35.400 ;
        RECT 367.950 32.400 393.600 33.600 ;
        RECT 400.950 33.600 403.050 34.050 ;
        RECT 505.950 33.600 508.050 34.050 ;
        RECT 400.950 32.400 508.050 33.600 ;
        RECT 367.950 31.950 370.050 32.400 ;
        RECT 400.950 31.950 403.050 32.400 ;
        RECT 505.950 31.950 508.050 32.400 ;
        RECT 532.950 33.600 535.050 34.050 ;
        RECT 559.950 33.600 562.050 34.050 ;
        RECT 574.950 33.600 577.050 34.050 ;
        RECT 532.950 32.400 577.050 33.600 ;
        RECT 532.950 31.950 535.050 32.400 ;
        RECT 559.950 31.950 562.050 32.400 ;
        RECT 574.950 31.950 577.050 32.400 ;
        RECT 604.950 33.600 607.050 34.050 ;
        RECT 724.950 33.600 727.050 34.050 ;
        RECT 742.950 33.600 745.050 34.050 ;
        RECT 604.950 32.400 636.600 33.600 ;
        RECT 604.950 31.950 607.050 32.400 ;
        RECT 58.950 28.950 61.050 31.050 ;
        RECT 121.950 28.950 124.050 31.050 ;
        RECT 247.950 30.600 250.050 31.050 ;
        RECT 292.950 30.600 295.050 31.050 ;
        RECT 325.950 30.600 328.050 31.050 ;
        RECT 247.950 29.400 328.050 30.600 ;
        RECT 247.950 28.950 250.050 29.400 ;
        RECT 292.950 28.950 295.050 29.400 ;
        RECT 325.950 28.950 328.050 29.400 ;
        RECT 364.950 30.600 367.050 31.050 ;
        RECT 394.950 30.600 397.050 31.050 ;
        RECT 438.000 30.600 442.050 31.050 ;
        RECT 364.950 29.400 397.050 30.600 ;
        RECT 437.400 29.400 459.600 30.600 ;
        RECT 364.950 28.950 367.050 29.400 ;
        RECT 394.950 28.950 397.050 29.400 ;
        RECT 438.000 28.950 442.050 29.400 ;
        RECT 40.950 27.600 43.050 28.050 ;
        RECT 17.400 26.400 43.050 27.600 ;
        RECT 17.400 21.900 18.600 26.400 ;
        RECT 40.950 25.950 43.050 26.400 ;
        RECT 46.950 27.600 49.050 28.050 ;
        RECT 55.950 27.600 58.050 28.200 ;
        RECT 46.950 26.400 58.050 27.600 ;
        RECT 46.950 25.950 49.050 26.400 ;
        RECT 55.950 26.100 58.050 26.400 ;
        RECT 59.400 21.900 60.600 28.950 ;
        RECT 61.950 27.600 64.050 28.200 ;
        RECT 118.950 27.600 121.050 28.200 ;
        RECT 61.950 26.400 121.050 27.600 ;
        RECT 61.950 26.100 64.050 26.400 ;
        RECT 118.950 26.100 121.050 26.400 ;
        RECT 122.400 21.900 123.600 28.950 ;
        RECT 129.000 27.600 133.050 28.050 ;
        RECT 128.400 25.950 133.050 27.600 ;
        RECT 148.950 27.600 151.050 28.200 ;
        RECT 166.950 27.600 169.050 28.200 ;
        RECT 172.950 27.600 175.050 28.050 ;
        RECT 148.950 26.400 162.600 27.600 ;
        RECT 148.950 26.100 151.050 26.400 ;
        RECT 128.400 21.900 129.600 25.950 ;
        RECT 136.950 24.600 139.050 25.050 ;
        RECT 161.400 24.600 162.600 26.400 ;
        RECT 166.950 26.400 175.050 27.600 ;
        RECT 166.950 26.100 169.050 26.400 ;
        RECT 172.950 25.950 175.050 26.400 ;
        RECT 199.950 27.750 202.050 28.200 ;
        RECT 208.950 27.750 211.050 28.200 ;
        RECT 199.950 26.550 211.050 27.750 ;
        RECT 199.950 26.100 202.050 26.550 ;
        RECT 208.950 26.100 211.050 26.550 ;
        RECT 214.950 27.600 217.050 28.200 ;
        RECT 241.950 27.600 244.050 28.050 ;
        RECT 214.950 26.400 244.050 27.600 ;
        RECT 214.950 26.100 217.050 26.400 ;
        RECT 241.950 25.950 244.050 26.400 ;
        RECT 259.950 27.600 262.050 28.200 ;
        RECT 277.950 27.600 280.050 28.200 ;
        RECT 259.950 26.400 280.050 27.600 ;
        RECT 259.950 26.100 262.050 26.400 ;
        RECT 277.950 26.100 280.050 26.400 ;
        RECT 283.950 27.600 286.050 28.200 ;
        RECT 289.950 27.600 292.050 28.050 ;
        RECT 307.950 27.600 310.050 28.200 ;
        RECT 283.950 26.400 292.050 27.600 ;
        RECT 283.950 26.100 286.050 26.400 ;
        RECT 289.950 25.950 292.050 26.400 ;
        RECT 293.400 26.400 310.050 27.600 ;
        RECT 293.400 24.600 294.600 26.400 ;
        RECT 307.950 26.100 310.050 26.400 ;
        RECT 343.950 27.750 346.050 28.200 ;
        RECT 352.950 27.750 355.050 28.200 ;
        RECT 343.950 26.550 355.050 27.750 ;
        RECT 343.950 26.100 346.050 26.550 ;
        RECT 352.950 26.100 355.050 26.550 ;
        RECT 370.950 27.750 373.050 28.200 ;
        RECT 379.950 27.750 382.050 28.200 ;
        RECT 370.950 26.550 382.050 27.750 ;
        RECT 433.950 27.600 436.050 28.200 ;
        RECT 370.950 26.100 373.050 26.550 ;
        RECT 379.950 26.100 382.050 26.550 ;
        RECT 413.400 26.400 436.050 27.600 ;
        RECT 413.400 24.600 414.600 26.400 ;
        RECT 433.950 26.100 436.050 26.400 ;
        RECT 445.950 27.600 448.050 28.050 ;
        RECT 454.950 27.600 457.050 28.200 ;
        RECT 445.950 26.400 457.050 27.600 ;
        RECT 445.950 25.950 448.050 26.400 ;
        RECT 454.950 26.100 457.050 26.400 ;
        RECT 136.950 23.400 159.600 24.600 ;
        RECT 161.400 23.400 165.600 24.600 ;
        RECT 136.950 22.950 139.050 23.400 ;
        RECT 16.950 19.800 19.050 21.900 ;
        RECT 22.950 21.600 25.050 21.900 ;
        RECT 34.950 21.600 37.050 21.900 ;
        RECT 52.950 21.600 55.050 21.900 ;
        RECT 22.950 20.400 55.050 21.600 ;
        RECT 22.950 19.800 25.050 20.400 ;
        RECT 34.950 19.800 37.050 20.400 ;
        RECT 52.950 19.800 55.050 20.400 ;
        RECT 58.950 19.800 61.050 21.900 ;
        RECT 88.950 21.450 91.050 21.900 ;
        RECT 94.950 21.450 97.050 21.900 ;
        RECT 88.950 20.250 97.050 21.450 ;
        RECT 88.950 19.800 91.050 20.250 ;
        RECT 94.950 19.800 97.050 20.250 ;
        RECT 121.950 19.800 124.050 21.900 ;
        RECT 127.950 19.800 130.050 21.900 ;
        RECT 139.950 21.600 142.050 22.050 ;
        RECT 158.400 21.900 159.600 23.400 ;
        RECT 145.950 21.600 148.050 21.900 ;
        RECT 139.950 20.400 148.050 21.600 ;
        RECT 139.950 19.950 142.050 20.400 ;
        RECT 145.950 19.800 148.050 20.400 ;
        RECT 157.950 19.800 160.050 21.900 ;
        RECT 164.400 21.600 165.600 23.400 ;
        RECT 281.400 23.400 453.600 24.600 ;
        RECT 281.400 21.900 282.600 23.400 ;
        RECT 452.400 21.900 453.600 23.400 ;
        RECT 458.400 21.900 459.600 29.400 ;
        RECT 460.950 27.600 463.050 28.200 ;
        RECT 469.950 27.600 472.050 28.050 ;
        RECT 460.950 26.400 472.050 27.600 ;
        RECT 460.950 26.100 463.050 26.400 ;
        RECT 469.950 25.950 472.050 26.400 ;
        RECT 505.950 27.600 508.050 28.050 ;
        RECT 532.950 27.600 535.050 28.050 ;
        RECT 505.950 26.400 535.050 27.600 ;
        RECT 505.950 25.950 508.050 26.400 ;
        RECT 532.950 25.950 535.050 26.400 ;
        RECT 541.950 26.100 544.050 28.200 ;
        RECT 546.000 27.600 550.050 28.050 ;
        RECT 472.950 24.600 475.050 25.050 ;
        RECT 472.950 23.400 486.600 24.600 ;
        RECT 472.950 22.950 475.050 23.400 ;
        RECT 485.400 21.900 486.600 23.400 ;
        RECT 181.950 21.600 184.050 21.900 ;
        RECT 164.400 20.400 184.050 21.600 ;
        RECT 181.950 19.800 184.050 20.400 ;
        RECT 211.950 21.450 214.050 21.900 ;
        RECT 220.950 21.450 223.050 21.900 ;
        RECT 211.950 20.250 223.050 21.450 ;
        RECT 211.950 19.800 214.050 20.250 ;
        RECT 220.950 19.800 223.050 20.250 ;
        RECT 226.950 21.450 229.050 21.900 ;
        RECT 232.950 21.450 235.050 21.900 ;
        RECT 226.950 20.250 235.050 21.450 ;
        RECT 226.950 19.800 229.050 20.250 ;
        RECT 232.950 19.800 235.050 20.250 ;
        RECT 256.950 21.600 259.050 21.900 ;
        RECT 274.950 21.600 277.050 21.900 ;
        RECT 256.950 20.400 277.050 21.600 ;
        RECT 256.950 19.800 259.050 20.400 ;
        RECT 274.950 19.800 277.050 20.400 ;
        RECT 280.950 19.800 283.050 21.900 ;
        RECT 292.950 21.450 295.050 21.900 ;
        RECT 298.950 21.450 301.050 21.900 ;
        RECT 292.950 20.250 301.050 21.450 ;
        RECT 292.950 19.800 295.050 20.250 ;
        RECT 298.950 19.800 301.050 20.250 ;
        RECT 304.950 21.450 307.050 21.900 ;
        RECT 310.950 21.450 313.050 21.900 ;
        RECT 304.950 20.250 313.050 21.450 ;
        RECT 304.950 19.800 307.050 20.250 ;
        RECT 310.950 19.800 313.050 20.250 ;
        RECT 316.950 21.450 319.050 21.900 ;
        RECT 322.950 21.450 325.050 21.900 ;
        RECT 316.950 20.250 325.050 21.450 ;
        RECT 316.950 19.800 319.050 20.250 ;
        RECT 322.950 19.800 325.050 20.250 ;
        RECT 328.950 21.450 331.050 21.900 ;
        RECT 337.950 21.450 340.050 21.900 ;
        RECT 328.950 20.250 340.050 21.450 ;
        RECT 328.950 19.800 331.050 20.250 ;
        RECT 337.950 19.800 340.050 20.250 ;
        RECT 346.950 21.600 349.050 21.900 ;
        RECT 391.950 21.600 394.050 21.900 ;
        RECT 346.950 20.400 394.050 21.600 ;
        RECT 346.950 19.800 349.050 20.400 ;
        RECT 391.950 19.800 394.050 20.400 ;
        RECT 400.950 21.450 403.050 21.900 ;
        RECT 409.950 21.450 412.050 21.900 ;
        RECT 400.950 20.250 412.050 21.450 ;
        RECT 400.950 19.800 403.050 20.250 ;
        RECT 409.950 19.800 412.050 20.250 ;
        RECT 424.950 21.450 427.050 21.900 ;
        RECT 430.950 21.450 433.050 21.900 ;
        RECT 424.950 20.250 433.050 21.450 ;
        RECT 424.950 19.800 427.050 20.250 ;
        RECT 430.950 19.800 433.050 20.250 ;
        RECT 436.950 21.450 439.050 21.900 ;
        RECT 445.950 21.450 448.050 21.900 ;
        RECT 436.950 20.250 448.050 21.450 ;
        RECT 436.950 19.800 439.050 20.250 ;
        RECT 445.950 19.800 448.050 20.250 ;
        RECT 451.950 19.800 454.050 21.900 ;
        RECT 457.950 19.800 460.050 21.900 ;
        RECT 469.950 21.450 472.050 21.900 ;
        RECT 478.950 21.450 481.050 21.900 ;
        RECT 469.950 20.250 481.050 21.450 ;
        RECT 469.950 19.800 472.050 20.250 ;
        RECT 478.950 19.800 481.050 20.250 ;
        RECT 484.950 19.800 487.050 21.900 ;
        RECT 508.950 21.600 511.050 22.050 ;
        RECT 526.950 21.600 529.050 22.050 ;
        RECT 508.950 20.400 529.050 21.600 ;
        RECT 508.950 19.950 511.050 20.400 ;
        RECT 526.950 19.950 529.050 20.400 ;
        RECT 52.950 18.600 55.050 19.050 ;
        RECT 70.950 18.600 73.050 19.050 ;
        RECT 52.950 17.400 73.050 18.600 ;
        RECT 52.950 16.950 55.050 17.400 ;
        RECT 70.950 16.950 73.050 17.400 ;
        RECT 76.950 18.600 79.050 19.050 ;
        RECT 85.950 18.600 88.050 19.050 ;
        RECT 76.950 17.400 88.050 18.600 ;
        RECT 76.950 16.950 79.050 17.400 ;
        RECT 85.950 16.950 88.050 17.400 ;
        RECT 190.950 18.600 193.050 19.050 ;
        RECT 205.950 18.600 208.050 19.050 ;
        RECT 190.950 17.400 208.050 18.600 ;
        RECT 190.950 16.950 193.050 17.400 ;
        RECT 205.950 16.950 208.050 17.400 ;
        RECT 262.950 18.600 265.050 19.050 ;
        RECT 280.950 18.600 283.050 19.050 ;
        RECT 262.950 17.400 283.050 18.600 ;
        RECT 262.950 16.950 265.050 17.400 ;
        RECT 280.950 16.950 283.050 17.400 ;
        RECT 361.950 18.600 364.050 19.050 ;
        RECT 379.950 18.600 382.050 19.050 ;
        RECT 385.950 18.600 388.050 19.050 ;
        RECT 361.950 17.400 388.050 18.600 ;
        RECT 361.950 16.950 364.050 17.400 ;
        RECT 379.950 16.950 382.050 17.400 ;
        RECT 385.950 16.950 388.050 17.400 ;
        RECT 391.950 18.600 394.050 19.050 ;
        RECT 415.950 18.600 418.050 19.050 ;
        RECT 391.950 17.400 418.050 18.600 ;
        RECT 391.950 16.950 394.050 17.400 ;
        RECT 415.950 16.950 418.050 17.400 ;
        RECT 529.950 18.600 532.050 19.050 ;
        RECT 538.950 18.600 541.050 19.050 ;
        RECT 529.950 17.400 541.050 18.600 ;
        RECT 542.400 18.600 543.600 26.100 ;
        RECT 545.400 25.950 550.050 27.600 ;
        RECT 565.950 26.100 568.050 28.200 ;
        RECT 613.950 27.600 616.050 28.200 ;
        RECT 619.950 27.600 622.050 31.050 ;
        RECT 613.950 27.000 622.050 27.600 ;
        RECT 622.950 27.750 625.050 28.200 ;
        RECT 631.950 27.750 634.050 28.200 ;
        RECT 613.950 26.400 621.600 27.000 ;
        RECT 622.950 26.550 634.050 27.750 ;
        RECT 613.950 26.100 616.050 26.400 ;
        RECT 622.950 26.100 625.050 26.550 ;
        RECT 631.950 26.100 634.050 26.550 ;
        RECT 545.400 21.900 546.600 25.950 ;
        RECT 553.950 24.600 556.050 25.050 ;
        RECT 566.400 24.600 567.600 26.100 ;
        RECT 553.950 23.400 567.600 24.600 ;
        RECT 553.950 22.950 556.050 23.400 ;
        RECT 635.400 21.900 636.600 32.400 ;
        RECT 724.950 32.400 745.050 33.600 ;
        RECT 724.950 31.950 727.050 32.400 ;
        RECT 742.950 31.950 745.050 32.400 ;
        RECT 781.950 33.600 784.050 34.050 ;
        RECT 805.950 33.600 808.050 34.050 ;
        RECT 781.950 32.400 808.050 33.600 ;
        RECT 781.950 31.950 784.050 32.400 ;
        RECT 805.950 31.950 808.050 32.400 ;
        RECT 637.950 27.600 640.050 28.200 ;
        RECT 646.950 27.600 649.050 28.050 ;
        RECT 637.950 26.400 649.050 27.600 ;
        RECT 637.950 26.100 640.050 26.400 ;
        RECT 646.950 25.950 649.050 26.400 ;
        RECT 658.950 27.750 661.050 28.200 ;
        RECT 664.950 27.750 667.050 28.200 ;
        RECT 658.950 26.550 667.050 27.750 ;
        RECT 658.950 26.100 661.050 26.550 ;
        RECT 664.950 26.100 667.050 26.550 ;
        RECT 682.950 27.750 685.050 28.200 ;
        RECT 694.950 27.750 697.050 28.200 ;
        RECT 682.950 26.550 697.050 27.750 ;
        RECT 682.950 26.100 685.050 26.550 ;
        RECT 694.950 26.100 697.050 26.550 ;
        RECT 736.950 27.600 739.050 28.500 ;
        RECT 751.950 27.600 754.050 28.200 ;
        RECT 736.950 26.400 754.050 27.600 ;
        RECT 793.950 27.600 796.050 28.500 ;
        RECT 805.950 27.600 808.050 28.200 ;
        RECT 793.950 26.400 808.050 27.600 ;
        RECT 751.950 26.100 754.050 26.400 ;
        RECT 805.950 26.100 808.050 26.400 ;
        RECT 826.950 27.750 829.050 28.200 ;
        RECT 838.950 27.750 841.050 28.200 ;
        RECT 826.950 26.550 841.050 27.750 ;
        RECT 826.950 26.100 829.050 26.550 ;
        RECT 838.950 26.100 841.050 26.550 ;
        RECT 710.400 23.400 729.600 24.600 ;
        RECT 544.950 19.800 547.050 21.900 ;
        RECT 568.950 21.450 571.050 21.900 ;
        RECT 604.950 21.450 607.050 21.900 ;
        RECT 568.950 20.250 607.050 21.450 ;
        RECT 568.950 19.800 571.050 20.250 ;
        RECT 604.950 19.800 607.050 20.250 ;
        RECT 610.950 21.600 613.050 21.900 ;
        RECT 628.950 21.600 631.050 21.900 ;
        RECT 610.950 20.400 631.050 21.600 ;
        RECT 610.950 19.800 613.050 20.400 ;
        RECT 628.950 19.800 631.050 20.400 ;
        RECT 634.950 19.800 637.050 21.900 ;
        RECT 655.950 21.600 658.050 21.900 ;
        RECT 673.950 21.600 676.050 21.900 ;
        RECT 710.400 21.600 711.600 23.400 ;
        RECT 728.400 21.600 729.600 23.400 ;
        RECT 655.950 20.400 676.050 21.600 ;
        RECT 655.950 19.800 658.050 20.400 ;
        RECT 673.950 19.800 676.050 20.400 ;
        RECT 709.950 19.500 712.050 21.600 ;
        RECT 718.950 21.150 721.050 21.600 ;
        RECT 724.800 21.150 726.900 21.600 ;
        RECT 718.950 19.950 726.900 21.150 ;
        RECT 718.950 19.500 721.050 19.950 ;
        RECT 724.800 19.500 726.900 19.950 ;
        RECT 727.950 21.150 730.050 21.600 ;
        RECT 766.950 21.150 769.050 21.600 ;
        RECT 727.950 19.950 769.050 21.150 ;
        RECT 727.950 19.500 730.050 19.950 ;
        RECT 766.950 19.500 769.050 19.950 ;
        RECT 775.950 21.150 778.050 21.600 ;
        RECT 781.950 21.150 784.050 21.600 ;
        RECT 775.950 19.950 784.050 21.150 ;
        RECT 775.950 19.500 778.050 19.950 ;
        RECT 781.950 19.500 784.050 19.950 ;
        RECT 877.950 21.450 880.050 21.900 ;
        RECT 889.950 21.450 892.050 21.900 ;
        RECT 877.950 20.250 892.050 21.450 ;
        RECT 877.950 19.800 880.050 20.250 ;
        RECT 889.950 19.800 892.050 20.250 ;
        RECT 646.950 18.600 649.050 19.050 ;
        RECT 661.950 18.600 664.050 19.050 ;
        RECT 542.400 17.400 552.600 18.600 ;
        RECT 529.950 16.950 532.050 17.400 ;
        RECT 538.950 16.950 541.050 17.400 ;
        RECT 133.950 15.600 136.050 16.050 ;
        RECT 181.950 15.600 184.050 16.050 ;
        RECT 133.950 14.400 184.050 15.600 ;
        RECT 133.950 13.950 136.050 14.400 ;
        RECT 181.950 13.950 184.050 14.400 ;
        RECT 187.950 15.600 190.050 15.900 ;
        RECT 238.950 15.600 241.050 16.050 ;
        RECT 247.950 15.600 250.050 16.050 ;
        RECT 187.950 14.400 250.050 15.600 ;
        RECT 187.950 13.800 190.050 14.400 ;
        RECT 238.950 13.950 241.050 14.400 ;
        RECT 247.950 13.950 250.050 14.400 ;
        RECT 289.950 15.600 292.050 16.050 ;
        RECT 352.950 15.600 355.050 16.050 ;
        RECT 367.950 15.600 370.050 16.050 ;
        RECT 289.950 14.400 370.050 15.600 ;
        RECT 289.950 13.950 292.050 14.400 ;
        RECT 352.950 13.950 355.050 14.400 ;
        RECT 367.950 13.950 370.050 14.400 ;
        RECT 448.950 15.600 451.050 16.050 ;
        RECT 472.950 15.600 475.050 16.050 ;
        RECT 448.950 14.400 475.050 15.600 ;
        RECT 551.400 15.600 552.600 17.400 ;
        RECT 646.950 17.400 664.050 18.600 ;
        RECT 646.950 16.950 649.050 17.400 ;
        RECT 661.950 16.950 664.050 17.400 ;
        RECT 553.950 15.600 556.050 16.050 ;
        RECT 616.950 15.600 619.050 16.050 ;
        RECT 622.950 15.600 625.050 16.050 ;
        RECT 551.400 14.400 625.050 15.600 ;
        RECT 448.950 13.950 451.050 14.400 ;
        RECT 472.950 13.950 475.050 14.400 ;
        RECT 553.950 13.950 556.050 14.400 ;
        RECT 616.950 13.950 619.050 14.400 ;
        RECT 622.950 13.950 625.050 14.400 ;
        RECT 631.950 15.600 634.050 16.050 ;
        RECT 664.950 15.600 667.050 16.050 ;
        RECT 631.950 14.400 667.050 15.600 ;
        RECT 631.950 13.950 634.050 14.400 ;
        RECT 664.950 13.950 667.050 14.400 ;
        RECT 109.950 12.600 112.050 13.050 ;
        RECT 223.950 12.600 226.050 13.050 ;
        RECT 109.950 11.400 226.050 12.600 ;
        RECT 109.950 10.950 112.050 11.400 ;
        RECT 223.950 10.950 226.050 11.400 ;
        RECT 268.950 12.600 271.050 13.050 ;
        RECT 478.950 12.600 481.050 13.050 ;
        RECT 610.950 12.600 613.050 13.050 ;
        RECT 268.950 11.400 351.600 12.600 ;
        RECT 268.950 10.950 271.050 11.400 ;
        RECT 46.950 9.600 49.050 10.050 ;
        RECT 256.950 9.600 259.050 10.050 ;
        RECT 46.950 8.400 259.050 9.600 ;
        RECT 350.400 9.600 351.600 11.400 ;
        RECT 478.950 11.400 613.050 12.600 ;
        RECT 478.950 10.950 481.050 11.400 ;
        RECT 610.950 10.950 613.050 11.400 ;
        RECT 361.950 9.600 364.050 10.050 ;
        RECT 350.400 8.400 364.050 9.600 ;
        RECT 46.950 7.950 49.050 8.400 ;
        RECT 256.950 7.950 259.050 8.400 ;
        RECT 361.950 7.950 364.050 8.400 ;
        RECT 421.950 9.600 424.050 10.050 ;
        RECT 601.950 9.600 604.050 10.050 ;
        RECT 421.950 8.400 604.050 9.600 ;
        RECT 421.950 7.950 424.050 8.400 ;
        RECT 601.950 7.950 604.050 8.400 ;
        RECT 112.950 6.600 115.050 7.050 ;
        RECT 199.950 6.600 202.050 7.050 ;
        RECT 112.950 5.400 202.050 6.600 ;
        RECT 112.950 4.950 115.050 5.400 ;
        RECT 199.950 4.950 202.050 5.400 ;
        RECT 319.950 6.600 322.050 7.050 ;
        RECT 415.950 6.600 418.050 7.050 ;
        RECT 319.950 5.400 418.050 6.600 ;
        RECT 319.950 4.950 322.050 5.400 ;
        RECT 415.950 4.950 418.050 5.400 ;
        RECT 427.950 6.600 430.050 7.050 ;
        RECT 508.950 6.600 511.050 7.050 ;
        RECT 427.950 5.400 511.050 6.600 ;
        RECT 427.950 4.950 430.050 5.400 ;
        RECT 508.950 4.950 511.050 5.400 ;
        RECT 517.950 6.600 520.050 7.050 ;
        RECT 562.950 6.600 565.050 7.050 ;
        RECT 517.950 5.400 565.050 6.600 ;
        RECT 517.950 4.950 520.050 5.400 ;
        RECT 562.950 4.950 565.050 5.400 ;
  END
END ALU_wrapper
END LIBRARY

