magic
tech scmos
magscale 1 30
timestamp 1719895877
<< checkpaint >>
rect 47800 171700 61200 180850
rect 18300 145440 61200 171700
rect 18300 145200 44800 145440
rect 47800 145200 61200 145440
rect 61300 145200 74700 180850
rect 74800 145200 88200 180850
rect 88300 146970 101700 180850
rect 101900 146970 115100 180850
rect 88300 145200 115100 146970
rect 115300 145200 128700 180850
rect 128800 171700 142200 180850
rect 128800 145440 171700 171700
rect 128800 145200 142200 145440
rect 145200 145200 171700 145440
rect 18300 142200 44650 145200
rect 9150 128800 44800 142200
rect 101100 140200 103040 145200
rect 145440 142200 171700 145200
rect 145200 128800 180850 142200
rect 9150 115300 44800 128700
rect 145200 115300 180850 128700
rect 9150 101800 44800 115200
rect 145200 101800 180850 115200
rect 9150 88300 44800 101700
rect 145200 88300 180850 101700
rect 9150 74900 44800 88100
rect 45930 85530 47165 85855
rect 45055 77480 47165 85530
rect 145200 74800 180850 88200
rect 9150 61300 44800 74700
rect 145200 61300 180850 74700
rect 9150 47800 44800 61200
rect 145200 47800 180850 61200
rect 18300 44800 44560 47800
rect 97740 45875 100710 47165
rect 99000 45640 100610 45875
rect 145440 44800 171700 47800
rect 18300 44560 44800 44800
rect 47800 44560 61200 44800
rect 18300 18300 61200 44560
rect 47800 9150 61200 18300
rect 61300 9150 74700 44800
rect 74800 9150 88200 44800
rect 88300 9150 101700 44800
rect 101800 9150 115200 44800
rect 115300 9150 128700 44800
rect 128800 44560 142200 44800
rect 145200 44560 171700 44800
rect 128800 18300 171700 44560
rect 128800 9150 142200 18300
<< metal1 >>
rect 103800 143060 104500 144200
rect 106100 143700 144145 144500
rect 143245 140000 144145 143700
rect 143650 114035 143860 114460
rect 143650 113320 144075 113530
rect 145400 87120 145650 103000
rect 145395 86800 145910 87120
rect 45955 75940 46235 76360
rect 143690 59375 143900 59815
rect 143740 57040 144260 57255
rect 145400 56820 145650 86800
rect 143740 56440 144260 56655
rect 98400 46240 99600 46475
rect 98400 45900 98700 46240
rect 60120 45600 98700 45900
rect 99000 45600 106555 45900
rect 99000 45300 99300 45600
rect 73620 45000 99300 45300
rect 73300 44135 73620 45000
<< metal2 >>
rect 49000 145510 49320 145940
rect 62500 144205 62820 145940
rect 76000 142900 76320 145940
rect 76000 142100 79780 142900
rect 79235 140900 79780 142100
rect 89500 141350 89820 145940
rect 101700 140800 102440 142970
rect 103800 140800 104500 143060
rect 116500 141800 116820 145940
rect 130000 143100 130320 145940
rect 130000 142400 135745 143100
rect 116500 141100 133045 141800
rect 135300 141000 135745 142400
rect 44060 129880 45500 130200
rect 44060 116380 44900 116700
rect 44500 105415 44900 116380
rect 45100 106015 45500 129880
rect 144900 130000 145940 130320
rect 143650 113530 143860 114035
rect 44900 105040 45720 105160
rect 44500 103200 44900 104185
rect 44060 102880 44900 103200
rect 45500 103840 45996 103960
rect 45100 102500 45500 103585
rect 44500 102100 45500 102500
rect 44500 89699 44900 102100
rect 44060 89379 44900 89699
rect 42300 78080 45655 84930
rect 44500 75940 45955 76360
rect 44500 62700 44900 75940
rect 44060 62380 44900 62700
rect 144400 59585 144650 116360
rect 143900 59375 144650 59585
rect 144900 57255 145150 130000
rect 144260 57040 145150 57255
rect 144260 56440 145400 56655
rect 44060 48880 45100 49200
rect 59800 44060 60120 45445
rect 67540 45000 67645 46265
rect 94240 45600 94505 46345
rect 94840 46200 94945 46365
rect 106840 45900 106945 46350
rect 107440 45300 107545 46285
rect 73300 44135 73620 45000
rect 99600 45000 107545 45300
rect 99600 44400 99900 45000
rect 108640 44400 108745 46465
rect 86800 44100 99900 44400
rect 100300 44100 108745 44400
rect 113800 44060 114120 44535
rect 127300 44060 127620 45200
rect 140800 44060 141120 45775
<< metal3 >>
rect 50845 144700 104500 145500
rect 103800 144200 104500 144700
rect 64455 143400 101700 144200
rect 78750 140900 88400 141350
rect 144650 116500 145440 116820
rect 144105 113740 145900 113950
rect 144075 113320 145400 113530
rect 143695 112240 144900 112360
rect 143840 111640 144400 111760
rect 45500 105640 46315 105760
rect 44900 105040 46590 105160
rect 44900 104440 46785 104560
rect 45500 103840 46530 103960
rect 45100 101440 47970 101561
rect 45100 49415 45500 101440
rect 143690 59815 143900 60460
rect 144150 60120 144400 111640
rect 144650 73620 144900 112240
rect 145150 87120 145400 113320
rect 145650 100905 145900 113740
rect 145150 86800 145395 87120
rect 144650 73300 145360 73620
rect 144150 59800 145545 60120
rect 95325 45900 140800 46200
rect 94725 45300 127300 45600
rect 68070 44700 113800 45000
<< m2contact >>
rect 106100 144500 113245 146000
rect 143440 115960 143860 116260
rect 145400 103000 145940 103320
rect 45655 78080 46530 84930
rect 145400 56440 145650 56820
rect 99600 46240 100050 46475
rect 59800 45445 60120 45900
rect 106555 45600 106945 45900
rect 73300 45000 73620 45300
<< m3contact >>
rect 49000 144700 50845 145510
rect 62500 143400 64455 144205
rect 77850 140900 78750 141350
rect 88400 140900 89820 141350
rect 101700 142970 102440 144200
rect 103800 143060 104500 144200
rect 144400 116360 144650 116820
rect 143440 115540 143860 115960
rect 143650 114035 143860 114460
rect 143650 113320 144075 113530
rect 45100 105640 45500 106015
rect 44500 105040 44900 105415
rect 44500 104185 44900 104560
rect 45100 103585 45500 103960
rect 45955 75940 46360 76360
rect 143690 59375 143900 59815
rect 145440 116500 145940 116820
rect 145650 100300 145940 100905
rect 145395 86800 145940 87120
rect 145360 73300 145940 73620
rect 145545 59800 145940 60120
rect 143740 57040 144260 57255
rect 143740 56440 144260 56655
rect 45100 48880 45500 49415
rect 94840 45900 95325 46200
rect 94240 45300 94725 45600
rect 67540 44700 68070 45000
rect 140800 45775 141120 46200
rect 127300 45200 127620 45600
rect 113800 44535 114120 45000
<< end >>