magic
tech scmos
magscale 1 2
timestamp 1726538409
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
<< ptransistor >>
rect 22 166 26 246
rect 36 166 40 246
rect 56 206 60 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 42 40 54
rect 24 14 26 42
rect 38 14 40 42
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
<< pdiffusion >>
rect 20 166 22 246
rect 26 166 36 246
rect 40 206 42 246
rect 54 206 56 246
rect 60 206 62 246
rect 40 166 51 206
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 42
rect 46 14 58 54
rect 66 14 78 54
<< pdcontact >>
rect 8 166 20 246
rect 42 206 54 246
rect 62 206 74 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 22 246 26 250
rect 36 246 40 250
rect 56 246 60 250
rect 22 162 26 166
rect 12 157 26 162
rect 36 162 40 166
rect 56 162 60 206
rect 36 157 44 162
rect 56 157 66 162
rect 12 129 16 157
rect 12 66 16 117
rect 40 103 44 157
rect 36 91 44 103
rect 12 59 24 66
rect 20 54 24 59
rect 40 54 44 91
rect 60 103 66 157
rect 60 54 64 103
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
<< polycontact >>
rect 4 117 16 129
rect 24 91 36 103
rect 64 91 76 103
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 8 246 20 252
rect 62 246 74 252
rect 43 117 51 206
rect 49 75 57 103
rect 49 68 74 75
rect 6 54 58 57
rect 18 48 46 54
rect 66 54 74 68
rect 26 8 38 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 3 103 17 117
rect 23 103 37 117
rect 43 103 57 117
rect 63 103 77 117
<< metal2 >>
rect 26 117 34 134
rect 66 117 74 134
rect 6 86 14 103
rect 46 86 54 103
<< m1p >>
rect -6 252 106 268
rect -6 -8 106 8
<< m2p >>
rect 26 119 34 134
rect 66 119 74 134
rect 6 86 14 101
rect 46 86 54 101
<< labels >>
rlabel metal1 -6 252 86 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal2 10 90 10 90 5 A
port 1 n signal input
rlabel metal2 30 130 30 130 5 B
port 2 n signal input
rlabel metal2 50 90 50 90 1 Y
port 4 n signal output
rlabel metal2 70 132 70 132 1 C
port 3 n signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
