magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -56 -56 84 204
<< diffusion >>
rect 5 5 23 143
<< genericcontact >>
rect 11 127 17 133
rect 11 99 17 105
rect 11 71 17 77
rect 11 43 17 49
rect 11 15 17 21
<< metal1 >>
rect 4 4 24 144
<< end >>
