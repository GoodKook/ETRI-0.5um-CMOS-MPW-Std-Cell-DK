magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -52 -52 1092 88
use p2res_CDNS_7230122529124  p2res_CDNS_7230122529124_0
timestamp 1555596690
transform 1 0 0 0 1 0
box 8 8 1032 28
<< end >>
