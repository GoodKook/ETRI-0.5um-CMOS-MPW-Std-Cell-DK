/* Verilog module written by vlog2Verilog (qflow) */

module cpu(
    output [15:0] AB,
    input [7:0] DI,
    output [7:0] DO,
    input IRQ,
    input NMI,
    input RDY,
    output WE,
    input clk,
    input reset
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire C ;
wire D ;
wire I ;
wire N ;
wire V ;
wire Z ;
wire _1677_ ;
wire _1257_ ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _1295_ ;
wire _703_ ;
wire _1389_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _1198_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _929_ ;
wire _509_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire _16_ ;
wire _1195_ ;
wire _54_ ;
wire _603_ ;
wire _1289_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _1098_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _926_ ;
wire _506_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire IRQ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _1727_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1__bF$buf10 ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire WE ;
wire _1383_ ;
wire _294_ ;
wire _13_ ;
wire _1439_ ;
wire _1019_ ;
wire php ;
wire _1192_ ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _1095_ ;
wire _7_ ;
wire RDY ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire adc_sbc ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _1724_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _10_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _1283_ ;
wire _194_ ;
wire _1339_ ;
wire _1092_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire write_back ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _1721_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _902__bF$buf0 ;
wire _902__bF$buf1 ;
wire _902__bF$buf2 ;
wire _902__bF$buf3 ;
wire _1718_ ;
wire _629_ ;
wire _209_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _1374_ ;
wire _285_ ;
wire _1_ ;
wire index_y ;
wire _1183_ ;
wire _1659_ ;
wire _1239_ ;
wire _42_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire clc ;
wire cld ;
wire cli ;
wire clk ;
wire clv ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _1715_ ;
wire _626_ ;
wire _206_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1371_ ;
wire _282_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _1319__bF$buf0 ;
wire _1319__bF$buf1 ;
wire _1319__bF$buf2 ;
wire _1319__bF$buf3 ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _1083_ ;
wire _1559_ ;
wire _1139_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _1027__bF$buf0 ;
wire _1027__bF$buf1 ;
wire _1027__bF$buf2 ;
wire _1027__bF$buf3 ;
wire _1027__bF$buf4 ;
wire _1712_ ;
wire _623_ ;
wire _203_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _1709_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire HC ;
wire _33_ ;
wire _1459_ ;
wire _1039_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire [6:0] ADD ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _1706_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _1609_ ;
wire _1362_ ;
wire RDY_bF$buf0 ;
wire RDY_bF$buf1 ;
wire RDY_bF$buf2 ;
wire RDY_bF$buf3 ;
wire RDY_bF$buf4 ;
wire RDY_bF$buf5 ;
wire RDY_bF$buf6 ;
wire RDY_bF$buf7 ;
wire RDY_bF$buf8 ;
wire RDY_bF$buf9 ;
wire _693_ ;
wire _273_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _1456_ ;
wire _1036_ ;
wire res ;
wire _787_ ;
wire _367_ ;
wire rotate ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire [3:0] alu_op ;
wire _1359_ ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire [1:0] dst_reg ;
wire \u_ALU8.BI7  ;
wire [7:0] DIHOLD ;
wire _805_ ;
wire _65_ ;
wire _1703_ ;
wire _614_ ;
wire _903__bF$buf0 ;
wire _903__bF$buf1 ;
wire _903__bF$buf2 ;
wire _903__bF$buf3 ;
wire [5:0] _1512_ ;
wire _843_ ;
wire _423_ ;
wire [15:0] _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _1738_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _24_ ;
wire _1679_ ;
wire _1259_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _1700_ ;
wire _611_ ;
wire _1714__bF$buf0 ;
wire _1714__bF$buf1 ;
wire _1714__bF$buf2 ;
wire _1714__bF$buf3 ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire \u_ALU8.BCD  ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _21_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire [7:0] \AXYS[1]  ;
wire _1579_ ;
wire _1159_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _928_ ;
wire _508_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _1729_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _1194_ ;
wire _53_ ;
wire _1479_ ;
wire _1059_ ;
wire store ;
wire _602_ ;
wire _1288_ ;
wire _199_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire IRHOLD_valid ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _1726_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _12_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _1285_ ;
wire _196_ ;
wire _1094_ ;
wire _1379_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire _1188_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _1723_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _1__bF$buf0 ;
wire _1__bF$buf1 ;
wire _1__bF$buf2 ;
wire _1__bF$buf3 ;
wire _1__bF$buf4 ;
wire _1__bF$buf5 ;
wire _1__bF$buf6 ;
wire _1__bF$buf7 ;
wire _1__bF$buf8 ;
wire _1__bF$buf9 ;
wire _919_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire backwards ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _44_ ;
wire _1699_ ;
wire _1279_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1720_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire [15:0] PC ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _1717_ ;
wire _628_ ;
wire _208_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _1373_ ;
wire _284_ ;
wire _0_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire adj_bcd ;
wire _41_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire _913_ ;
wire [7:0] \AXYS[3]  ;
wire _1599_ ;
wire _1179_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire compare ;
wire _816_ ;
wire _76_ ;
wire _1714_ ;
wire _625_ ;
wire _205_ ;
wire load_only ;
wire clk_bF$buf10 ;
wire shift ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1370_ ;
wire _281_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire [1:0] src_reg ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _1329_ ;
wire _1082_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire _35_ ;
wire _1149__bF$buf0 ;
wire _1149__bF$buf1 ;
wire _1149__bF$buf2 ;
wire _1149__bF$buf3 ;
wire _1149__bF$buf4 ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _1711_ ;
wire _622_ ;
wire _202_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _1708_ ;
wire _619_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _1593_ ;
wire _1173_ ;
wire _1649_ ;
wire _1229_ ;
wire _32_ ;
wire _1458_ ;
wire _1038_ ;
wire [2:0] cond_code ;
wire _789_ ;
wire _369_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _904_ ;
wire _713_ ;
wire _1399_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _1705_ ;
wire _616_ ;
wire [5:0] state ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire bit_ins ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire [7:0] DI ;
wire [7:0] DO ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _1493_ ;
wire _1073_ ;
wire _1549_ ;
wire _1129_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _1702_ ;
wire _613_ ;
wire _1299_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire [15:0] AB ;
wire [7:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _1737_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _1393_ ;
wire _23_ ;
wire _1449_ ;
wire _1029_ ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire _886__bF$buf0 ;
wire _886__bF$buf1 ;
wire _886__bF$buf2 ;
wire _886__bF$buf3 ;
wire _886__bF$buf4 ;
wire _886__bF$buf5 ;
wire _886__bF$buf6 ;
wire _704_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _1199_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire NMI ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _20_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _1293_ ;
wire _1349_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire plp ;
wire _1196_ ;
wire _55_ ;
wire _604_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _1099_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _1728_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire _295_ ;
wire _14_ ;
wire _1193_ ;
wire _1669_ ;
wire _1249_ ;
wire _52_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _1096_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _1725_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _11_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _1093_ ;
wire [7:0] \AXYS[0]  ;
wire _1569_ ;
wire _1149_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _1722_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _1719_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _1528_ ;
wire _1108_ ;
wire shift_right ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _914__bF$buf0 ;
wire _914__bF$buf1 ;
wire _914__bF$buf2 ;
wire _914__bF$buf3 ;
wire _914__bF$buf4 ;
wire _43_ ;
wire _1469_ ;
wire _1049_ ;
wire [7:0] DIMUX ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _1150__bF$buf0 ;
wire _1150__bF$buf1 ;
wire _1150__bF$buf2 ;
wire _1150__bF$buf3 ;
wire _1150__bF$buf4 ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire [3:0] op ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _1716_ ;
wire _627_ ;
wire _207_ ;
wire _720__bF$buf0 ;
wire _720__bF$buf1 ;
wire _720__bF$buf2 ;
wire _720__bF$buf3 ;
wire _380_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _1619_ ;
wire _1372_ ;
wire _283_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire sec ;
wire sed ;
wire sei ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire [7:0] IRHOLD ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire alu_shift_right ;
wire _1084_ ;
wire _1369_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _1713_ ;
wire _624_ ;
wire _204_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _1519_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire _34_ ;
wire _1689_ ;
wire _1269_ ;
wire NMI_1 ;
wire _812_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _1710_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire adc_bcd ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _1707_ ;
wire _618_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _931__bF$buf0 ;
wire _931__bF$buf1 ;
wire _931__bF$buf2 ;
wire _931__bF$buf3 ;
wire _931__bF$buf4 ;
wire _903_ ;
wire [7:0] \AXYS[2]  ;
wire _1589_ ;
wire _1169_ ;
wire _712_ ;
wire [7:0] ABH ;
wire [7:0] ABL ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire NMI_edge ;
wire _806_ ;
wire _66_ ;
wire _1704_ ;
wire _615_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire [7:0] _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire load_reg ;
wire _709_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire CI ;
wire CO ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _1739_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire inc ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _1701_ ;
wire _612_ ;
wire _1298_ ;
wire reset ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _22_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

FILL FILL_2__2620_ (
);

FILL FILL_2__2200_ (
);

FILL FILL_4__2966_ (
);

FILL FILL_4__2546_ (
);

FILL FILL_4__2126_ (
);

FILL FILL_0__2866_ (
);

FILL FILL_0__2446_ (
);

FILL FILL_0__2026_ (
);

FILL FILL_5__1830_ (
);

FILL FILL_7__1848_ (
);

FILL FILL_1__1822_ (
);

FILL FILL_3__1748_ (
);

FILL FILL_5__2615_ (
);

FILL FILL_1__2607_ (
);

FILL FILL_4__3084_ (
);

FILL FILL_4__1817_ (
);

DFFSR _3403_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_72_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[0] [3])
);

FILL FILL_1__2780_ (
);

FILL FILL_1__2360_ (
);

FILL FILL_3__2286_ (
);

FILL FILL_5__3573_ (
);

FILL FILL_5__3153_ (
);

FILL FILL_1__3565_ (
);

FILL FILL_1__3145_ (
);

FILL FILL_4__1990_ (
);

FILL FILL_0__1890_ (
);

FILL FILL_4__2775_ (
);

FILL FILL_4__2355_ (
);

FILL FILL_0__2675_ (
);

FILL FILL_6__3642_ (
);

FILL FILL_0__2255_ (
);

FILL FILL_6__3222_ (
);

FILL FILL_2__3634_ (
);

FILL FILL_2__3214_ (
);

FILL FILL_3__1977_ (
);

FILL FILL_5__2844_ (
);

FILL FILL_5__2424_ (
);

FILL FILL_5__2004_ (
);

FILL FILL_1__2836_ (
);

FILL FILL_1__2416_ (
);

FILL FILL_3__3703_ (
);

FILL FILL_5__3629_ (
);

FILL FILL_5__3209_ (
);

FILL FILL169050x64950 (
);

FILL FILL_7__2195_ (
);

FILL FILL_0__1946_ (
);

FILL FILL_6__2913_ (
);

NAND2X1 _3632_ (
    .A(_1602_),
    .B(_1604_),
    .Y(_1662_)
);

AOI21X1 _3212_ (
    .A(_744_),
    .B(_798_),
    .C(_801_),
    .Y(_87_)
);

FILL FILL_3__2095_ (
);

FILL FILL_2__2905_ (
);

FILL FILL_4__2584_ (
);

FILL FILL_4__2164_ (
);

FILL FILL_0__2484_ (
);

FILL FILL_6__3451_ (
);

FILL FILL_0__2064_ (
);

FILL FILL_6__3031_ (
);

FILL FILL_2__3023_ (
);

NOR2X1 _2903_ (
    .A(_1185_),
    .B(_1187_),
    .Y(_550_)
);

FILL FILL_1__1860_ (
);

FILL FILL_3__1786_ (
);

FILL FILL_0__3269_ (
);

FILL FILL_5__2653_ (
);

FILL FILL_5__2233_ (
);

FILL FILL_1__2645_ (
);

FILL FILL_7__3612_ (
);

FILL FILL_1__2225_ (
);

FILL FILL_3__3512_ (
);

FILL FILL_5__3018_ (
);

FILL FILL_4__1855_ (
);

FILL FILL_0__1755_ (
);

FILL FILL_6__2722_ (
);

DFFSR _3441_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(_109_),
    .CLK(clk_bF$buf2),
    .Q(ABH[0])
);

FILL FILL_6__2302_ (
);

OAI21X1 _3021_ (
    .A(_950_),
    .B(_1063_),
    .C(RDY_bF$buf2),
    .Y(_645_)
);

FILL FILL_2__2714_ (
);

FILL FILL_5__3191_ (
);

FILL FILL_6__3507_ (
);

FILL FILL_1__3183_ (
);

FILL FILL_5__1924_ (
);

FILL FILL_1__1916_ (
);

FILL FILL_4__2393_ (
);

FILL FILL_5__2709_ (
);

FILL FILL_0__2293_ (
);

FILL FILL_6__3260_ (
);

FILL FILL_2__3672_ (
);

FILL FILL_2__3252_ (
);

FILL FILL_4__3598_ (
);

FILL FILL_4__3178_ (
);

NOR2X1 _2712_ (
    .A(_377_),
    .B(_381_),
    .Y(_382_)
);

FILL FILL_0__3498_ (
);

FILL FILL_0__3078_ (
);

FILL FILL_5__2882_ (
);

FILL FILL_5__2462_ (
);

FILL FILL_5__2042_ (
);

FILL FILL_1__2874_ (
);

FILL FILL_1__2454_ (
);

FILL FILL_1__2034_ (
);

FILL FILL_7__3001_ (
);

FILL FILL_5__3667_ (
);

FILL FILL_5__3247_ (
);

FILL FILL_1__3659_ (
);

FILL FILL_1__3239_ (
);

FILL FILL_0__1984_ (
);

FILL FILL_6__2951_ (
);

OAI21X1 _3670_ (
    .A(_1693_),
    .B(_1692_),
    .C(_1691_),
    .Y(_1521_)
);

FILL FILL_6__2531_ (
);

NAND3X1 _3250_ (
    .A(_130_),
    .B(_825_),
    .C(_822_),
    .Y(_826_)
);

FILL FILL_6__2111_ (
);

FILL FILL_2__2943_ (
);

FILL FILL_2__2523_ (
);

FILL FILL_2__2103_ (
);

FILL FILL_4__2869_ (
);

FILL FILL_4__2449_ (
);

FILL FILL_4__2029_ (
);

FILL FILL_0__2769_ (
);

FILL FILL_0__2349_ (
);

FILL FILL_6__3316_ (
);

FILL FILL_0__3710_ (
);

FILL FILL_2__3308_ (
);

FILL FILL_5__2938_ (
);

FILL FILL_5__2518_ (
);

FILL FILL_0_BUFX2_insert20 (
);

FILL FILL_0_BUFX2_insert21 (
);

FILL FILL_2__3481_ (
);

FILL FILL_0_BUFX2_insert22 (
);

FILL FILL_0_BUFX2_insert23 (
);

FILL FILL_2__3061_ (
);

FILL FILL_0_BUFX2_insert24 (
);

FILL FILL_0_BUFX2_insert25 (
);

FILL FILL_6__1802_ (
);

AND2X2 _2941_ (
    .A(_583_),
    .B(_575_),
    .Y(_584_)
);

OAI21X1 _2521_ (
    .A(state[5]),
    .B(_996_),
    .C(_215_),
    .Y(_216_)
);

INVX1 _2101_ (
    .A(_1209_),
    .Y(_1210_)
);

FILL FILL_5__2691_ (
);

FILL FILL_5__2271_ (
);

NAND2X1 _3306_ (
    .A(_1741_[10]),
    .B(_869_),
    .Y(_872_)
);

FILL FILL_1__2683_ (
);

FILL FILL_7__3650_ (
);

FILL FILL_1__2263_ (
);

FILL FILL_7__3230_ (
);

FILL FILL_3__2189_ (
);

FILL FILL_3__3550_ (
);

FILL FILL_3__3130_ (
);

FILL FILL_5__3476_ (
);

FILL FILL_5__3056_ (
);

FILL FILL_1__3468_ (
);

FILL FILL_1__3048_ (
);

FILL FILL_4__1893_ (
);

FILL FILL_0__1793_ (
);

FILL FILL_6__2760_ (
);

FILL FILL_6__2340_ (
);

FILL FILL_2__2752_ (
);

FILL FILL_2__2332_ (
);

FILL FILL_4__2678_ (
);

FILL FILL_4__2258_ (
);

FILL FILL_0__2998_ (
);

FILL FILL_0__2578_ (
);

FILL FILL_6__3545_ (
);

FILL FILL_0__2158_ (
);

FILL FILL_6__3125_ (
);

FILL FILL_2__3537_ (
);

FILL FILL_2__3117_ (
);

FILL FILL_5__1962_ (
);

FILL FILL_1__1954_ (
);

FILL FILL_7__2501_ (
);

FILL FILL_3__2821_ (
);

FILL FILL_3__2401_ (
);

FILL FILL_5__2747_ (
);

FILL FILL_5__2327_ (
);

FILL FILL_1__2739_ (
);

FILL FILL_1__2319_ (
);

FILL FILL_2__3290_ (
);

FILL FILL_3__3606_ (
);

NAND3X1 _2750_ (
    .A(_392_),
    .B(_399_),
    .C(_415_),
    .Y(_416_)
);

OAI21X1 _2330_ (
    .A(RDY_bF$buf8),
    .B(_1027__bF$buf1),
    .C(_1436_),
    .Y(_1437_)
);

FILL FILL_4__1949_ (
);

FILL FILL_5__2080_ (
);

FILL FILL_7__2098_ (
);

FILL FILL_0__1849_ (
);

FILL FILL_6__2816_ (
);

INVX1 _3535_ (
    .A(BI[1]),
    .Y(_1565_)
);

NAND2X1 _3115_ (
    .A(_966_),
    .B(_1319__bF$buf3),
    .Y(_723_)
);

FILL FILL_1__2492_ (
);

FILL FILL_1__2072_ (
);

FILL FILL_2__2808_ (
);

FILL FILL_5__3285_ (
);

FILL FILL_1__3697_ (
);

FILL FILL_1__3277_ (
);

FILL FILL_2__2981_ (
);

FILL FILL_2__2561_ (
);

FILL FILL_2__2141_ (
);

FILL FILL_4__2487_ (
);

FILL FILL_4__2067_ (
);

FILL FILL_0__2387_ (
);

FILL FILL_5__1771_ (
);

NAND2X1 _2806_ (
    .A(_392_),
    .B(_399_),
    .Y(_469_)
);

FILL FILL_1__1763_ (
);

FILL FILL_7__2730_ (
);

FILL FILL_3__2630_ (
);

FILL FILL_3__2210_ (
);

FILL FILL_5__2976_ (
);

FILL FILL_5__2556_ (
);

FILL FILL_5__2136_ (
);

FILL FILL_1__2968_ (
);

FILL FILL_1__2548_ (
);

FILL FILL_1__2128_ (
);

FILL FILL_6__1840_ (
);

FILL FILL_2__1832_ (
);

FILL FILL_4__1758_ (
);

FILL FILL_6__2625_ (
);

DFFSR _3344_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_21_),
    .CLK(clk_bF$buf1),
    .Q(cond_code[2])
);

FILL FILL_6__2205_ (
);

FILL FILL_2__2617_ (
);

FILL FILL_5__3094_ (
);

FILL FILL_1__3086_ (
);

FILL FILL_3__1901_ (
);

FILL FILL_5__1827_ (
);

FILL FILL_1__1819_ (
);

FILL FILL_2__2790_ (
);

FILL FILL_2__2370_ (
);

FILL FILL_4__2296_ (
);

NAND2X1 _1830_ (
    .A(_903__bF$buf2),
    .B(_955_),
    .Y(_956_)
);

FILL FILL_6__3583_ (
);

FILL FILL_0__2196_ (
);

FILL FILL_6__3163_ (
);

FILL FILL_2__3575_ (
);

FILL FILL_2__3155_ (
);

AOI22X1 _2615_ (
    .A(ABH[5]),
    .B(_925_),
    .C(_198_),
    .D(ADD[5]),
    .Y(_297_)
);

FILL FILL_1__1992_ (
);

FILL FILL_5__2785_ (
);

FILL FILL_5__2365_ (
);

FILL FILL_1__2777_ (
);

FILL FILL_1__2357_ (
);

BUFX2 BUFX2_insert37 (
    .A(_720_),
    .Y(_720__bF$buf3)
);

BUFX2 BUFX2_insert38 (
    .A(_720_),
    .Y(_720__bF$buf2)
);

FILL FILL_3__3644_ (
);

BUFX2 BUFX2_insert39 (
    .A(_720_),
    .Y(_720__bF$buf1)
);

FILL FILL_3__3224_ (
);

FILL FILL169950x3750 (
);

FILL FILL_4__1987_ (
);

FILL FILL_0__1887_ (
);

FILL FILL_6__2854_ (
);

OAI21X1 _3573_ (
    .A(_1562_),
    .B(_1600_),
    .C(_1602_),
    .Y(_1603_)
);

FILL FILL_6__2434_ (
);

FILL FILL_6__2014_ (
);

OAI21X1 _3153_ (
    .A(DIMUX[4]),
    .B(_1018_),
    .C(_756_),
    .Y(_757_)
);

FILL FILL_2__2846_ (
);

FILL FILL_2__2426_ (
);

FILL FILL_2__2006_ (
);

FILL FILL_4__3713_ (
);

FILL FILL_6__3639_ (
);

FILL FILL_6__3219_ (
);

FILL FILL_0__3613_ (
);

FILL FILL_3__2915_ (
);

OAI21X1 _2844_ (
    .A(_1015_),
    .B(_351_),
    .C(_504_),
    .Y(_505_)
);

OAI21X1 _2424_ (
    .A(_128_),
    .B(_129_),
    .C(_131_),
    .Y(alu_op[0])
);

INVX1 _2004_ (
    .A(_1116_),
    .Y(_1117_)
);

FILL FILL_5__2594_ (
);

FILL FILL_5__2174_ (
);

NAND2X1 _3629_ (
    .A(_1657_),
    .B(_1656_),
    .Y(_1659_)
);

NOR2X1 _3209_ (
    .A(\AXYS[2] [1]),
    .B(_798_),
    .Y(_800_)
);

FILL FILL_1__2586_ (
);

FILL FILL_7__3553_ (
);

FILL FILL_1__2166_ (
);

FILL FILL_7__3133_ (
);

FILL FILL_3__3453_ (
);

FILL FILL_3__3033_ (
);

FILL FILL_2__1870_ (
);

FILL FILL_4__1796_ (
);

FILL FILL_6__2663_ (
);

DFFSR _3382_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(DIMUX[7]),
    .CLK(clk_bF$buf3),
    .Q(DIHOLD[7])
);

FILL FILL_6__2243_ (
);

FILL FILL_2__2655_ (
);

FILL FILL_2__2235_ (
);

FILL FILL_4__3522_ (
);

FILL FILL_4__3102_ (
);

FILL FILL_6__3028_ (
);

FILL FILL_0__3002_ (
);

FILL FILL_5__1865_ (
);

FILL FILL_1__1857_ (
);

FILL FILL_7__2824_ (
);

FILL FILL_7__2404_ (
);

FILL FILL_3__2724_ (
);

FILL FILL_3__2304_ (
);

FILL FILL_7__3609_ (
);

FILL FILL_2__3193_ (
);

FILL FILL_3__3509_ (
);

FILL FILL_6__1934_ (
);

AOI21X1 _2653_ (
    .A(_929_),
    .B(_935_),
    .C(_327_),
    .Y(_328_)
);

AND2X2 _2233_ (
    .A(_1340_),
    .B(_1336_),
    .Y(_1341_)
);

FILL FILL_2__1926_ (
);

FILL FILL169950x111750 (
);

FILL FILL_6__2719_ (
);

DFFSR _3438_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_106_),
    .CLK(clk_bF$buf1),
    .Q(ABL[5])
);

NOR2X1 _3018_ (
    .A(_643_),
    .B(_620_),
    .Y(_644_)
);

FILL FILL_1__2395_ (
);

FILL FILL169350x39750 (
);

FILL FILL_3__3262_ (
);

FILL FILL_5__3188_ (
);

FILL FILL_6__2892_ (
);

FILL FILL_6__2472_ (
);

OAI21X1 _3191_ (
    .A(_724_),
    .B(_789_),
    .C(_790_),
    .Y(_77_)
);

FILL FILL_6__2052_ (
);

FILL FILL_2__2884_ (
);

FILL FILL_2__2464_ (
);

FILL FILL_2__2044_ (
);

OAI21X1 _1924_ (
    .A(_1029_),
    .B(_1033_),
    .C(index_y),
    .Y(_1041_)
);

FILL FILL_6__3677_ (
);

FILL FILL_6__3257_ (
);

FILL FILL_2__3669_ (
);

FILL FILL_0__3651_ (
);

FILL FILL_0__3231_ (
);

FILL FILL_2__3249_ (
);

OAI21X1 _2709_ (
    .A(_251_),
    .B(_378_),
    .C(_148_),
    .Y(_379_)
);

FILL FILL_7__2633_ (
);

FILL FILL_7__2213_ (
);

FILL FILL_3__2953_ (
);

FILL FILL_3__2533_ (
);

FILL FILL_3__2113_ (
);

FILL FILL_5__2879_ (
);

FILL FILL_5__2459_ (
);

FILL FILL_5__2039_ (
);

OAI22X1 _2882_ (
    .A(_147_),
    .B(_1150__bF$buf1),
    .C(_535_),
    .D(_533_),
    .Y(_23_)
);

INVX1 _2462_ (
    .A(_162_),
    .Y(_163_)
);

INVX1 _2042_ (
    .A(IRHOLD[1]),
    .Y(_1151_)
);

FILL FILL_4__2602_ (
);

FILL FILL_6__2948_ (
);

NAND2X1 _3667_ (
    .A(ADD[4]),
    .B(_1714__bF$buf0),
    .Y(_1691_)
);

FILL FILL_6__2528_ (
);

INVX1 _3247_ (
    .A(_1030_),
    .Y(_823_)
);

FILL FILL_6__2108_ (
);

FILL FILL_0__2922_ (
);

FILL FILL_0__2502_ (
);

FILL FILL_3__3491_ (
);

FILL FILL_3__3071_ (
);

FILL FILL_0__3707_ (
);

FILL FILL_3__1804_ (
);

FILL FILL_6__2281_ (
);

FILL FILL_2__2693_ (
);

FILL FILL_2__2273_ (
);

FILL FILL_4__2199_ (
);

FILL FILL_4__3560_ (
);

FILL FILL_4__3140_ (
);

FILL FILL_6__3486_ (
);

FILL FILL_0__2099_ (
);

FILL FILL_6__3066_ (
);

FILL FILL_2__3478_ (
);

FILL FILL_0__3460_ (
);

FILL FILL_0__3040_ (
);

FILL FILL_2__3058_ (
);

NAND2X1 _2938_ (
    .A(_550_),
    .B(_1182_),
    .Y(_581_)
);

OAI22X1 _2518_ (
    .A(_914__bF$buf3),
    .B(_974_),
    .C(_931__bF$buf3),
    .D(_984_),
    .Y(_213_)
);

FILL FILL_1__1895_ (
);

FILL FILL_7__2862_ (
);

FILL FILL_7__2442_ (
);

FILL FILL_7__2022_ (
);

FILL FILL_3__2762_ (
);

FILL FILL_3__2342_ (
);

FILL FILL_5__2688_ (
);

FILL FILL_5__2268_ (
);

FILL FILL_7__3227_ (
);

FILL FILL_1__3621_ (
);

FILL FILL_1__3201_ (
);

FILL FILL_3__3547_ (
);

FILL FILL_3__3127_ (
);

FILL FILL_6__1972_ (
);

OAI21X1 _2691_ (
    .A(_362_),
    .B(_340_),
    .C(RDY_bF$buf3),
    .Y(_363_)
);

OAI21X1 _2271_ (
    .A(cond_code[2]),
    .B(_1377_),
    .C(_1378_),
    .Y(_1379_)
);

FILL FILL_2__1964_ (
);

FILL FILL_4__2831_ (
);

FILL FILL_4__2411_ (
);

FILL FILL_6__2757_ (
);

INVX2 _3476_ (
    .A(alu_shift_right),
    .Y(_1722_)
);

FILL FILL_6__2337_ (
);

NOR2X1 _3056_ (
    .A(plp),
    .B(cld),
    .Y(_670_)
);

FILL FILL_2__2749_ (
);

FILL FILL_0__2731_ (
);

FILL FILL_2__2329_ (
);

FILL FILL_0__2311_ (
);

FILL FILL_4__3616_ (
);

FILL FILL_0__3516_ (
);

FILL FILL_5__1959_ (
);

FILL FILL_6__2090_ (
);

FILL FILL_5__2900_ (
);

FILL FILL_2__2082_ (
);

FILL FILL_3__2818_ (
);

NAND2X1 _1962_ (
    .A(_969_),
    .B(_1078_),
    .Y(_1079_)
);

FILL FILL_6__3295_ (
);

FILL FILL_2__3287_ (
);

OAI21X1 _2747_ (
    .A(_329_),
    .B(_365_),
    .C(PC[5]),
    .Y(_413_)
);

OAI21X1 _2327_ (
    .A(_886__bF$buf0),
    .B(_1079_),
    .C(_1433_),
    .Y(_1434_)
);

FILL FILL_7__2251_ (
);

FILL FILL_3__2991_ (
);

FILL FILL_3__2571_ (
);

FILL FILL_3__2151_ (
);

FILL FILL_5__2497_ (
);

FILL FILL_5__2077_ (
);

FILL FILL_1__2489_ (
);

FILL FILL_7__3456_ (
);

FILL FILL_1__2069_ (
);

FILL FILL_7__3036_ (
);

FILL FILL_1__3010_ (
);

FILL FILL_6__1781_ (
);

INVX1 _2080_ (
    .A(_1188_),
    .Y(_1189_)
);

FILL FILL_5_BUFX2_insert40 (
);

FILL FILL_5_BUFX2_insert41 (
);

FILL FILL_5_BUFX2_insert42 (
);

FILL FILL_5_BUFX2_insert43 (
);

FILL FILL_5_BUFX2_insert44 (
);

FILL FILL_5_BUFX2_insert45 (
);

FILL FILL_2__1773_ (
);

FILL FILL_5_BUFX2_insert46 (
);

FILL FILL_5_BUFX2_insert47 (
);

FILL FILL_5_BUFX2_insert48 (
);

FILL FILL_5_BUFX2_insert49 (
);

FILL FILL_4__2640_ (
);

FILL FILL_4__2220_ (
);

FILL FILL_6__2986_ (
);

FILL FILL_6__2566_ (
);

NAND2X1 _3285_ (
    .A(ABL[0]),
    .B(_860_),
    .Y(_861_)
);

FILL FILL_6__2146_ (
);

FILL FILL_0__2960_ (
);

FILL FILL_2__2978_ (
);

FILL FILL_2__2558_ (
);

FILL FILL_0__2540_ (
);

FILL FILL_0__2120_ (
);

FILL FILL_2__2138_ (
);

FILL FILL_7__1942_ (
);

FILL FILL_4__3005_ (
);

FILL FILL_3__1842_ (
);

FILL FILL_5__1768_ (
);

FILL FILL_7__2727_ (
);

FILL FILL_1__2701_ (
);

FILL FILL_3__2627_ (
);

FILL FILL_3__2207_ (
);

INVX1 _1771_ (
    .A(state[3]),
    .Y(_897_)
);

FILL FILL_2__3096_ (
);

FILL FILL_4__1911_ (
);

FILL FILL_6__1837_ (
);

AOI21X1 _2976_ (
    .A(_596_),
    .B(_606_),
    .C(_1326_),
    .Y(_607_)
);

AND2X2 _2556_ (
    .A(_243_),
    .B(_246_),
    .Y(_247_)
);

AOI22X1 _2136_ (
    .A(_1193_),
    .B(_1244_),
    .C(_1243_),
    .D(_1242_),
    .Y(_1245_)
);

FILL FILL_7__2480_ (
);

FILL FILL_2__1829_ (
);

FILL FILL_0__1811_ (
);

FILL FILL_3__2380_ (
);

FILL FILL_1__2298_ (
);

FILL FILL_7__3265_ (
);

FILL FILL_3__3585_ (
);

FILL FILL_3__3165_ (
);

FILL FILL_6__2795_ (
);

FILL FILL_6__2375_ (
);

NAND2X1 _3094_ (
    .A(_895_),
    .B(_703_),
    .Y(_704_)
);

FILL FILL_2__2787_ (
);

FILL FILL_2__2367_ (
);

NAND2X1 _1827_ (
    .A(_903__bF$buf3),
    .B(_952_),
    .Y(_953_)
);

FILL FILL_7__1751_ (
);

FILL FILL_4__3654_ (
);

FILL FILL_4__3234_ (
);

FILL FILL_0__3554_ (
);

FILL FILL_0__3134_ (
);

FILL FILL_5__1997_ (
);

FILL FILL_1__1989_ (
);

FILL FILL_7__2956_ (
);

FILL FILL_7__2116_ (
);

FILL FILL_1__2930_ (
);

FILL FILL_1__2510_ (
);

FILL FILL_3__2856_ (
);

FILL FILL_3__2436_ (
);

FILL FILL_3__2016_ (
);

FILL FILL_5__3303_ (
);

FILL FILL_1__3715_ (
);

MUX2X1 _2785_ (
    .A(_448_),
    .B(_285_),
    .S(_1154_),
    .Y(_449_)
);

NOR2X1 _2365_ (
    .A(RDY_bF$buf1),
    .B(_1470_),
    .Y(_1471_)
);

FILL FILL_4__2925_ (
);

FILL FILL_4__2505_ (
);

FILL FILL_7__3074_ (
);

FILL FILL_0__2825_ (
);

FILL FILL_0__2405_ (
);

FILL FILL_6__2184_ (
);

FILL FILL_2__2596_ (
);

FILL FILL_2__2176_ (
);

FILL FILL_7__1980_ (
);

FILL FILL_4__3463_ (
);

FILL FILL_4__3043_ (
);

FILL FILL_3__1880_ (
);

FILL FILL_2_CLKBUF1_insert26 (
);

FILL FILL_2_CLKBUF1_insert27 (
);

FILL FILL_2_CLKBUF1_insert28 (
);

FILL FILL_2_CLKBUF1_insert29 (
);

FILL FILL_1__1798_ (
);

FILL FILL_7__2345_ (
);

FILL FILL_3__2665_ (
);

FILL FILL_3__2245_ (
);

FILL FILL_5__3532_ (
);

FILL FILL_5__3112_ (
);

FILL FILL_1__3524_ (
);

FILL FILL_1__3104_ (
);

FILL FILL_6__1875_ (
);

OAI21X1 _2594_ (
    .A(_276_),
    .B(_218_),
    .C(_279_),
    .Y(_1741_[9])
);

NOR2X1 _2174_ (
    .A(_1172_),
    .B(_1212_),
    .Y(_1283_)
);

FILL FILL_2__1867_ (
);

FILL FILL_4__2734_ (
);

FILL FILL_4__2314_ (
);

DFFSR _3379_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(DIMUX[4]),
    .CLK(clk_bF$buf5),
    .Q(DIHOLD[4])
);

FILL FILL_0__2634_ (
);

FILL FILL_6__3601_ (
);

FILL FILL_0__2214_ (
);

FILL FILL_4__3519_ (
);

FILL FILL_3__1936_ (
);

FILL FILL_5__2803_ (
);

NOR2X1 _1865_ (
    .A(_931__bF$buf4),
    .B(_989_),
    .Y(_990_)
);

FILL FILL_4__3692_ (
);

FILL FILL_4__3272_ (
);

FILL FILL_6__3198_ (
);

FILL FILL_0__3592_ (
);

FILL FILL_0__3172_ (
);

FILL FILL_7__2574_ (
);

FILL FILL_0__1905_ (
);

FILL FILL_3__2894_ (
);

FILL FILL_3__2474_ (
);

FILL FILL_3__2054_ (
);

FILL FILL_3__3259_ (
);

FILL FILL_4__2963_ (
);

FILL FILL_4__2543_ (
);

FILL FILL_4__2123_ (
);

FILL FILL_6__2889_ (
);

FILL FILL_6__2469_ (
);

OAI21X1 _3188_ (
    .A(_722_),
    .B(_787_),
    .C(_788_),
    .Y(_76_)
);

FILL FILL_6__2049_ (
);

FILL FILL_0__2863_ (
);

FILL FILL_0__2443_ (
);

FILL FILL_0__2023_ (
);

FILL FILL_7__1845_ (
);

FILL FILL_3__1745_ (
);

FILL FILL_0__3648_ (
);

FILL FILL_0__3228_ (
);

FILL FILL_5__2612_ (
);

FILL FILL_1__2604_ (
);

FILL FILL_4__3081_ (
);

FILL FILL_4__1814_ (
);

INVX1 _2879_ (
    .A(_531_),
    .Y(_533_)
);

OAI21X1 _2459_ (
    .A(_1319__bF$buf2),
    .B(_1263_),
    .C(PC[10]),
    .Y(_160_)
);

OAI21X1 _2039_ (
    .A(_1074_),
    .B(_1143_),
    .C(_1148_),
    .Y(AI[7])
);

FILL FILL_7__2383_ (
);

DFFSR _3400_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_69_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[0] [0])
);

FILL FILL_3__2283_ (
);

FILL FILL_7__3588_ (
);

FILL FILL_5__3570_ (
);

FILL FILL_5__3150_ (
);

FILL FILL_0__2919_ (
);

FILL FILL_1__3562_ (
);

FILL FILL_1__3142_ (
);

FILL FILL_3__3488_ (
);

FILL FILL_3__3068_ (
);

FILL FILL_4__2772_ (
);

FILL FILL_4__2352_ (
);

FILL FILL_6__2698_ (
);

FILL FILL_6__2278_ (
);

FILL FILL_0__2672_ (
);

FILL FILL_0__2252_ (
);

FILL FILL_2__3631_ (
);

FILL FILL_2__3211_ (
);

FILL FILL_4__3557_ (
);

FILL FILL_4__3137_ (
);

FILL FILL_3__1974_ (
);

FILL FILL_0__3457_ (
);

FILL FILL_0__3037_ (
);

FILL FILL_7__2859_ (
);

FILL FILL_5__2841_ (
);

FILL FILL_5__2421_ (
);

FILL FILL_7__2019_ (
);

FILL FILL_5__2001_ (
);

FILL FILL_1__2833_ (
);

FILL FILL_1__2413_ (
);

FILL FILL_3__2759_ (
);

FILL FILL_3__2339_ (
);

FILL FILL_3__3700_ (
);

FILL FILL_5__3626_ (
);

FILL FILL_5__3206_ (
);

FILL FILL_1__3618_ (
);

FILL FILL_6__1969_ (
);

AOI21X1 _2688_ (
    .A(_342_),
    .B(_347_),
    .C(_359_),
    .Y(_360_)
);

OAI21X1 _2268_ (
    .A(cond_code[2]),
    .B(_1374_),
    .C(_1375_),
    .Y(_1376_)
);

FILL FILL_7__2192_ (
);

FILL FILL_0__1943_ (
);

FILL FILL_6__2910_ (
);

FILL FILL_3__2092_ (
);

FILL FILL_2__2902_ (
);

FILL FILL_4__2828_ (
);

FILL FILL_4__2408_ (
);

FILL FILL_0__2728_ (
);

FILL FILL_0__2308_ (
);

FILL FILL_3__3297_ (
);

FILL FILL_4__2581_ (
);

FILL FILL_4__2161_ (
);

FILL FILL_6__2087_ (
);

FILL FILL_0__2481_ (
);

FILL FILL_2__2499_ (
);

FILL FILL_0__2061_ (
);

FILL FILL_2__2079_ (
);

FILL FILL_2__3020_ (
);

OAI21X1 _1959_ (
    .A(_914__bF$buf4),
    .B(_1075_),
    .C(_953_),
    .Y(_1076_)
);

INVX1 _2900_ (
    .A(sei),
    .Y(_548_)
);

FILL FILL_3__1783_ (
);

FILL FILL_0__3266_ (
);

FILL FILL_5__2650_ (
);

FILL FILL_5__2230_ (
);

FILL FILL_7__2248_ (
);

FILL FILL_1__2642_ (
);

FILL FILL_1__2222_ (
);

FILL FILL_3__2988_ (
);

FILL FILL_3__2568_ (
);

FILL FILL_3__2148_ (
);

FILL FILL_5__3015_ (
);

FILL FILL_1__3007_ (
);

FILL FILL_4__1852_ (
);

FILL FILL_6__1778_ (
);

OAI21X1 _2497_ (
    .A(_143_),
    .B(_1143_),
    .C(_192_),
    .Y(_1742_[7])
);

MUX2X1 _2077_ (
    .A(DIMUX[6]),
    .B(IRHOLD[6]),
    .S(_1168_),
    .Y(_1186_)
);

FILL FILL_0__1752_ (
);

FILL FILL_2__2711_ (
);

FILL FILL_4__2637_ (
);

FILL FILL_4__2217_ (
);

FILL FILL_0__2957_ (
);

FILL FILL_0__2537_ (
);

FILL FILL_6__3504_ (
);

FILL FILL_0__2117_ (
);

FILL FILL_1__3180_ (
);

FILL FILL_5__1921_ (
);

FILL FILL_1__1913_ (
);

FILL FILL_3__1839_ (
);

FILL FILL_4__2390_ (
);

FILL FILL_5__2706_ (
);

FILL FILL_0__2290_ (
);

INVX1 _1768_ (
    .A(C),
    .Y(_894_)
);

FILL FILL_4__3595_ (
);

FILL FILL_4__3175_ (
);

FILL FILL_0__3495_ (
);

FILL FILL_0__3075_ (
);

FILL FILL_4__1908_ (
);

FILL FILL_7__2477_ (
);

FILL FILL_0__1808_ (
);

FILL FILL_1__2871_ (
);

FILL FILL_1__2451_ (
);

FILL FILL_1__2031_ (
);

FILL FILL_3__2797_ (
);

FILL FILL_3__2377_ (
);

FILL FILL_5__3664_ (
);

FILL FILL_5__3244_ (
);

FILL FILL_1__3656_ (
);

FILL FILL_1__3236_ (
);

FILL FILL_0__1981_ (
);

FILL FILL_2__1999_ (
);

FILL FILL_2__2940_ (
);

FILL FILL_2__2520_ (
);

FILL FILL_2__2100_ (
);

FILL FILL_4__2866_ (
);

FILL FILL_4__2446_ (
);

FILL FILL_4__2026_ (
);

FILL FILL_0__2766_ (
);

FILL FILL_0__2346_ (
);

FILL FILL_6__3313_ (
);

FILL FILL_2__3305_ (
);

FILL FILL_7__1748_ (
);

FILL FILL_1_CLKBUF1_insert30 (
);

FILL FILL_1_CLKBUF1_insert31 (
);

FILL FILL_1_CLKBUF1_insert32 (
);

FILL FILL_1_CLKBUF1_insert33 (
);

FILL FILL_1_CLKBUF1_insert34 (
);

FILL FILL_1_CLKBUF1_insert35 (
);

FILL FILL_1_CLKBUF1_insert36 (
);

FILL FILL_5__2935_ (
);

FILL FILL_5__2515_ (
);

FILL FILL_1__2927_ (
);

FILL FILL_1__2507_ (
);

OAI21X1 _1997_ (
    .A(_1010_),
    .B(_983_),
    .C(_1110_),
    .Y(_1111_)
);

OAI21X1 _3303_ (
    .A(_269_),
    .B(_869_),
    .C(_870_),
    .Y(_109_)
);

FILL FILL_1__2680_ (
);

FILL FILL_1__2260_ (
);

FILL FILL_3__2186_ (
);

FILL FILL_5__3473_ (
);

FILL FILL_5__3053_ (
);

FILL FILL_1__3465_ (
);

FILL FILL_1__3045_ (
);

FILL FILL_4__1890_ (
);

FILL FILL_0__1790_ (
);

FILL FILL_4__2675_ (
);

FILL FILL_4__2255_ (
);

FILL FILL_0__2995_ (
);

FILL FILL_0__2575_ (
);

FILL FILL_6__3542_ (
);

FILL FILL_0__2155_ (
);

FILL FILL_6__3122_ (
);

FILL FILL_2__3534_ (
);

FILL FILL_2__3114_ (
);

FILL FILL_7__1977_ (
);

FILL FILL_1__1951_ (
);

FILL FILL_3__1877_ (
);

FILL FILL_5__2744_ (
);

FILL FILL_5__2324_ (
);

FILL FILL_1__2736_ (
);

FILL FILL_1__2316_ (
);

FILL FILL_7__3703_ (
);

FILL FILL_3__3603_ (
);

FILL FILL_5__3529_ (
);

FILL FILL_5__3109_ (
);

FILL FILL_4__1946_ (
);

FILL FILL_7__2095_ (
);

FILL FILL_0__1846_ (
);

FILL FILL_6__2813_ (
);

INVX1 _3532_ (
    .A(_1561_),
    .Y(_1562_)
);

OAI21X1 _3112_ (
    .A(_719_),
    .B(_718_),
    .C(RDY_bF$buf2),
    .Y(_720_)
);

FILL FILL_2__2805_ (
);

FILL FILL_5__3282_ (
);

FILL FILL_1__3694_ (
);

FILL FILL_1__3274_ (
);

FILL FILL_4__2484_ (
);

FILL FILL_4__2064_ (
);

FILL FILL_0__2384_ (
);

FILL FILL_4__3269_ (
);

NOR3X1 _2803_ (
    .A(_456_),
    .B(_416_),
    .C(_370_),
    .Y(_466_)
);

FILL FILL_1__1760_ (
);

FILL FILL_0__3589_ (
);

FILL FILL_0__3169_ (
);

FILL FILL_5__2973_ (
);

FILL FILL_5__2553_ (
);

FILL FILL_5__2133_ (
);

FILL FILL_1__2965_ (
);

FILL FILL_1__2545_ (
);

FILL FILL_1__2125_ (
);

FILL FILL_4__1755_ (
);

FILL FILL_6__2622_ (
);

DFFSR _3341_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_18_),
    .CLK(clk_bF$buf1),
    .Q(NMI_edge)
);

FILL FILL_6__2202_ (
);

FILL FILL_2__2614_ (
);

FILL FILL_5__3091_ (
);

FILL FILL_1__3083_ (
);

FILL FILL_5__1824_ (
);

FILL FILL_1__1816_ (
);

FILL FILL_4__2293_ (
);

FILL FILL_5__2609_ (
);

FILL FILL_6__3580_ (
);

FILL FILL_0__2193_ (
);

FILL FILL_6__3160_ (
);

FILL FILL_2__3572_ (
);

FILL FILL_2__3152_ (
);

FILL FILL_4__3498_ (
);

FILL FILL_4__3078_ (
);

OAI21X1 _2612_ (
    .A(_290_),
    .B(_218_),
    .C(_294_),
    .Y(_1741_[12])
);

FILL FILL_5__2782_ (
);

FILL FILL_5__2362_ (
);

FILL FILL_1__2774_ (
);

FILL FILL_1__2354_ (
);

FILL FILL_3__3641_ (
);

FILL FILL_3__3221_ (
);

FILL FILL_5__3567_ (
);

FILL FILL_5__3147_ (
);

FILL FILL_1__3559_ (
);

FILL FILL_1__3139_ (
);

FILL FILL_4__1984_ (
);

FILL FILL_0__1884_ (
);

FILL FILL_6__2851_ (
);

AND2X2 _3570_ (
    .A(_1595_),
    .B(_1599_),
    .Y(_1600_)
);

FILL FILL_6__2431_ (
);

FILL FILL_6__2011_ (
);

NAND2X1 _3150_ (
    .A(\AXYS[0] [3]),
    .B(_722_),
    .Y(_755_)
);

FILL FILL_2__2843_ (
);

FILL FILL_2__2423_ (
);

FILL FILL_2__2003_ (
);

FILL FILL_4__2769_ (
);

FILL FILL_4__2349_ (
);

FILL FILL_4__3710_ (
);

FILL FILL_0__2669_ (
);

FILL FILL_6__3636_ (
);

FILL FILL_0__2249_ (
);

FILL FILL_6__3216_ (
);

FILL FILL_0__3610_ (
);

FILL FILL_2__3628_ (
);

FILL FILL_2__3208_ (
);

FILL FILL_3__2912_ (
);

FILL FILL_5__2838_ (
);

FILL FILL_5__2418_ (
);

NOR2X1 _2841_ (
    .A(_1334_),
    .B(_1135_),
    .Y(_502_)
);

INVX2 _2421_ (
    .A(_915_),
    .Y(_129_)
);

AOI22X1 _2001_ (
    .A(_1049_),
    .B(\AXYS[3] [4]),
    .C(\AXYS[2] [4]),
    .D(_1057_),
    .Y(_1114_)
);

FILL FILL_5__2591_ (
);

FILL FILL_5__2171_ (
);

FILL FILL_6__2907_ (
);

OAI21X1 _3626_ (
    .A(_1655_),
    .B(_1636_),
    .C(_1650_),
    .Y(_1656_)
);

AND2X2 _3206_ (
    .A(_1057_),
    .B(_721_),
    .Y(_798_)
);

FILL FILL_1__2583_ (
);

FILL FILL_7__3550_ (
);

FILL FILL_1__2163_ (
);

FILL FILL_7__3130_ (
);

FILL FILL_3__2089_ (
);

FILL FILL_3__3450_ (
);

FILL FILL_3__3030_ (
);

FILL FILL_4__1793_ (
);

FILL FILL_6__2660_ (
);

FILL FILL_6__2240_ (
);

FILL FILL_2__2652_ (
);

FILL FILL_2__2232_ (
);

FILL FILL_4__2998_ (
);

FILL FILL_4__2578_ (
);

FILL FILL_4__2158_ (
);

FILL FILL_0__2898_ (
);

FILL FILL_0__2478_ (
);

FILL FILL_0__2058_ (
);

FILL FILL_6__3025_ (
);

FILL FILL_2__3017_ (
);

FILL FILL_5__1862_ (
);

FILL FILL_1__1854_ (
);

FILL FILL_7__2401_ (
);

FILL FILL_3__2721_ (
);

FILL FILL_3__2301_ (
);

FILL FILL_5__2647_ (
);

FILL FILL_5__2227_ (
);

FILL FILL_1__2639_ (
);

FILL FILL_7__3606_ (
);

FILL FILL_1__2219_ (
);

FILL FILL_2__3190_ (
);

FILL FILL_3__3506_ (
);

FILL FILL_6__1931_ (
);

AOI22X1 _2650_ (
    .A(_902__bF$buf0),
    .B(_931__bF$buf2),
    .C(_984_),
    .D(_912_),
    .Y(_325_)
);

NAND2X1 _2230_ (
    .A(RDY_bF$buf2),
    .B(_1063_),
    .Y(_1338_)
);

FILL FILL_2__1923_ (
);

FILL FILL_4__1849_ (
);

FILL FILL_0__1749_ (
);

FILL FILL_6__2716_ (
);

DFFSR _3435_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_103_),
    .CLK(clk_bF$buf1),
    .Q(ABL[2])
);

NAND3X1 _3015_ (
    .A(_1159_),
    .B(_1178_),
    .C(_640_),
    .Y(_641_)
);

FILL FILL_1__2392_ (
);

FILL FILL_2__2708_ (
);

FILL FILL_1_BUFX2_insert60 (
);

FILL FILL_1_BUFX2_insert61 (
);

FILL FILL_1_BUFX2_insert62 (
);

FILL FILL_1_BUFX2_insert63 (
);

FILL FILL_5__3185_ (
);

FILL FILL_1_BUFX2_insert64 (
);

FILL FILL_1_BUFX2_insert65 (
);

FILL FILL_1_BUFX2_insert66 (
);

FILL FILL_1_BUFX2_insert67 (
);

FILL FILL_1_BUFX2_insert68 (
);

FILL FILL_1_BUFX2_insert69 (
);

FILL FILL_1__3597_ (
);

FILL FILL_1__3177_ (
);

FILL FILL_5__1918_ (
);

FILL FILL_2__2881_ (
);

FILL FILL_2__2461_ (
);

FILL FILL_2__2041_ (
);

FILL FILL_4__2387_ (
);

INVX1 _1921_ (
    .A(_1034_),
    .Y(_1038_)
);

FILL FILL_6__3674_ (
);

FILL FILL_0__2287_ (
);

FILL FILL_6__3254_ (
);

FILL FILL_2__3666_ (
);

FILL FILL_2__3246_ (
);

OAI22X1 _2706_ (
    .A(RDY_bF$buf3),
    .B(_1011_),
    .C(_376_),
    .D(_375_),
    .Y(_6_)
);

FILL FILL_7__2630_ (
);

FILL FILL_3__2950_ (
);

FILL FILL_3__2530_ (
);

FILL FILL_3__2110_ (
);

FILL FILL_5__2876_ (
);

FILL FILL_5__2456_ (
);

FILL FILL_5__2036_ (
);

FILL FILL_1__2868_ (
);

FILL FILL_1__2448_ (
);

FILL FILL_1__2028_ (
);

FILL FILL_3__3315_ (
);

FILL FILL_0__1978_ (
);

FILL FILL_6__2945_ (
);

OAI21X1 _3664_ (
    .A(_1714__bF$buf1),
    .B(_1620_),
    .C(_1689_),
    .Y(_1519_)
);

FILL FILL_6__2525_ (
);

OAI21X1 _3244_ (
    .A(_902__bF$buf1),
    .B(_928_),
    .C(_1272_),
    .Y(_820_)
);

FILL FILL_6__2105_ (
);

FILL FILL_2__2937_ (
);

FILL FILL_2__2517_ (
);

FILL FILL_7__1901_ (
);

FILL FILL168150x75750 (
);

FILL FILL_3__1801_ (
);

FILL FILL_0__3704_ (
);

FILL FILL_2__2690_ (
);

FILL FILL_2__2270_ (
);

FILL FILL_4__2196_ (
);

FILL FILL_6__3483_ (
);

FILL FILL_0__2096_ (
);

FILL FILL_6__3063_ (
);

FILL FILL_2__3475_ (
);

FILL FILL_2__3055_ (
);

INVX2 _2935_ (
    .A(_1397_),
    .Y(_578_)
);

NAND2X1 _2515_ (
    .A(_903__bF$buf1),
    .B(_1427_),
    .Y(_210_)
);

FILL FILL_1__1892_ (
);

FILL FILL_5__2685_ (
);

FILL FILL_5__2265_ (
);

FILL FILL_1__2677_ (
);

FILL FILL_1__2257_ (
);

FILL FILL_7__3224_ (
);

FILL FILL_3__3544_ (
);

FILL FILL_3__3124_ (
);

FILL FILL_2__1961_ (
);

FILL FILL_4__1887_ (
);

FILL FILL_0__1787_ (
);

FILL FILL_6__2754_ (
);

AND2X2 _3473_ (
    .A(_1718_),
    .B(BI[7]),
    .Y(_1719_)
);

FILL FILL_6__2334_ (
);

AND2X2 _3053_ (
    .A(_663_),
    .B(AV),
    .Y(_668_)
);

FILL FILL_2__2746_ (
);

FILL FILL_2__2326_ (
);

FILL FILL_4__3613_ (
);

FILL FILL_6__3539_ (
);

FILL FILL_6__3119_ (
);

FILL FILL_0__3513_ (
);

FILL FILL_5__1956_ (
);

FILL FILL_1__1948_ (
);

FILL FILL_3__2815_ (
);

FILL FILL_6__3292_ (
);

FILL FILL_2__3284_ (
);

AND2X2 _2744_ (
    .A(_401_),
    .B(_410_),
    .Y(_411_)
);

NOR2X1 _2324_ (
    .A(_1383_),
    .B(_1430_),
    .Y(_1431_)
);

FILL FILL_5__2494_ (
);

FILL FILL_5__2074_ (
);

AOI21X1 _3529_ (
    .A(_1725_),
    .B(_1553_),
    .C(_1740_),
    .Y(_1559_)
);

OAI21X1 _3109_ (
    .A(_935_),
    .B(_992_),
    .C(_969_),
    .Y(_717_)
);

FILL FILL_1__2486_ (
);

FILL FILL_7__3453_ (
);

FILL FILL_1__2066_ (
);

FILL FILL_7__3033_ (
);

FILL FILL_5__3699_ (
);

FILL FILL_5__3279_ (
);

FILL FILL_5_BUFX2_insert10 (
);

FILL FILL_5_BUFX2_insert11 (
);

FILL FILL_5_BUFX2_insert12 (
);

FILL FILL_5_BUFX2_insert13 (
);

FILL FILL_5_BUFX2_insert14 (
);

FILL FILL_5_BUFX2_insert15 (
);

FILL FILL_2__1770_ (
);

FILL FILL_5_BUFX2_insert16 (
);

FILL FILL_5_BUFX2_insert17 (
);

FILL FILL_5_BUFX2_insert18 (
);

FILL FILL_5_BUFX2_insert19 (
);

FILL FILL_6__2983_ (
);

FILL FILL_6__2563_ (
);

NOR2X1 _3282_ (
    .A(_857_),
    .B(_1000_),
    .Y(_858_)
);

FILL FILL_6__2143_ (
);

FILL FILL_2__2975_ (
);

FILL FILL_2__2555_ (
);

FILL FILL_2__2135_ (
);

FILL FILL_4__3002_ (
);

FILL FILL_5__1765_ (
);

FILL FILL_1__1757_ (
);

FILL FILL_7__2724_ (
);

FILL FILL_7__2304_ (
);

FILL FILL_3__2624_ (
);

FILL FILL_3__2204_ (
);

FILL FILL_7__3509_ (
);

FILL FILL_2__3093_ (
);

FILL FILL_6__1834_ (
);

OAI21X1 _2973_ (
    .A(_601_),
    .B(_604_),
    .C(_602_),
    .Y(_45_)
);

INVX1 _2553_ (
    .A(ABL[4]),
    .Y(_244_)
);

NOR2X1 _2133_ (
    .A(write_back),
    .B(_1241_),
    .Y(_1242_)
);

FILL FILL_2__1826_ (
);

FILL FILL_6__2619_ (
);

DFFSR _3338_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_16_),
    .CLK(clk_bF$buf0),
    .Q(PC[14])
);

FILL FILL_1__2295_ (
);

FILL FILL_7__3262_ (
);

FILL FILL_3__3582_ (
);

FILL FILL_3__3162_ (
);

FILL FILL_5__3088_ (
);

FILL FILL_6__2792_ (
);

FILL FILL_6__2372_ (
);

MUX2X1 _3091_ (
    .A(_701_),
    .B(_697_),
    .S(_698_),
    .Y(_66_)
);

FILL FILL_2__2784_ (
);

FILL FILL_2__2364_ (
);

NOR2X1 _1824_ (
    .A(_931__bF$buf2),
    .B(_949_),
    .Y(_950_)
);

FILL FILL_4__3651_ (
);

FILL FILL_4__3231_ (
);

FILL FILL_6__3577_ (
);

FILL FILL_6__3157_ (
);

FILL FILL_2__3569_ (
);

FILL FILL_0__3551_ (
);

FILL FILL_2__3149_ (
);

FILL FILL_0__3131_ (
);

FILL FILL_5__1994_ (
);

AOI22X1 _2609_ (
    .A(ABH[4]),
    .B(_925_),
    .C(_198_),
    .D(ADD[4]),
    .Y(_292_)
);

FILL FILL_1__1986_ (
);

FILL FILL_7__2953_ (
);

FILL FILL_7__2533_ (
);

FILL FILL_7__2113_ (
);

FILL FILL_3__2853_ (
);

FILL FILL_3__2433_ (
);

FILL FILL_3__2013_ (
);

FILL FILL_5__2779_ (
);

FILL FILL_5__2359_ (
);

FILL FILL_5__3300_ (
);

FILL FILL_1__3712_ (
);

FILL FILL_3__3638_ (
);

FILL FILL_3__3218_ (
);

AOI21X1 _2782_ (
    .A(ADD[3]),
    .B(_1299_),
    .C(_1334_),
    .Y(_446_)
);

NAND2X1 _2362_ (
    .A(RDY_bF$buf6),
    .B(_1020_),
    .Y(_1468_)
);

FILL FILL_4__2922_ (
);

FILL FILL_4__2502_ (
);

FILL FILL_6__2848_ (
);

INVX1 _3567_ (
    .A(_1596_),
    .Y(_1597_)
);

FILL FILL_6__2428_ (
);

FILL FILL_6__2008_ (
);

NOR2X1 _3147_ (
    .A(_750_),
    .B(_747_),
    .Y(_752_)
);

FILL FILL_0__2822_ (
);

FILL FILL_0__2402_ (
);

FILL FILL_4__3707_ (
);

FILL FILL_0__3607_ (
);

FILL FILL_6__2181_ (
);

FILL FILL_2__2593_ (
);

FILL FILL_2__2173_ (
);

FILL FILL_4__2099_ (
);

FILL FILL_3__2909_ (
);

FILL FILL_4__3460_ (
);

FILL FILL_4__3040_ (
);

FILL FILL_6_BUFX2_insert60 (
);

FILL FILL_6_BUFX2_insert61 (
);

FILL FILL_6_BUFX2_insert62 (
);

FILL FILL_6_BUFX2_insert63 (
);

FILL FILL_6_BUFX2_insert64 (
);

FILL FILL_6_BUFX2_insert65 (
);

FILL FILL_6_BUFX2_insert66 (
);

FILL FILL_6_BUFX2_insert67 (
);

FILL FILL_6_BUFX2_insert68 (
);

FILL FILL_6_BUFX2_insert69 (
);

OAI21X1 _2838_ (
    .A(RDY_bF$buf4),
    .B(_295_),
    .C(_499_),
    .Y(_15_)
);

NOR2X1 _2418_ (
    .A(_1445_),
    .B(_126_),
    .Y(_127_)
);

FILL FILL_1__1795_ (
);

FILL FILL_7__2762_ (
);

FILL FILL_7__2342_ (
);

FILL FILL_3__2662_ (
);

FILL FILL_3__2242_ (
);

FILL FILL_5__2588_ (
);

FILL FILL_5__2168_ (
);

FILL FILL_7__3127_ (
);

FILL FILL_1__3521_ (
);

FILL FILL_1__3101_ (
);

FILL FILL_3__3027_ (
);

FILL FILL_6__1872_ (
);

AOI21X1 _2591_ (
    .A(_198_),
    .B(ADD[1]),
    .C(_1093_),
    .Y(_277_)
);

NAND3X1 _2171_ (
    .A(_1256_),
    .B(_1279_),
    .C(_1254_),
    .Y(_1280_)
);

FILL FILL_2__1864_ (
);

FILL FILL_4__2731_ (
);

FILL FILL_4__2311_ (
);

FILL FILL_6__2657_ (
);

DFFSR _3376_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(DIMUX[1]),
    .CLK(clk_bF$buf5),
    .Q(DIHOLD[1])
);

FILL FILL_6__2237_ (
);

FILL FILL_2__2649_ (
);

FILL FILL_0__2631_ (
);

FILL FILL_2__2229_ (
);

FILL FILL_0__2211_ (
);

FILL FILL_4__3516_ (
);

FILL FILL_3__1933_ (
);

FILL FILL_5__1859_ (
);

FILL FILL_5__2800_ (
);

FILL FILL_3__2718_ (
);

NAND2X1 _1862_ (
    .A(_913_),
    .B(_935_),
    .Y(_987_)
);

FILL FILL_6__3195_ (
);

FILL FILL_2__3187_ (
);

FILL FILL_6__1928_ (
);

NAND3X1 _2647_ (
    .A(_1092_),
    .B(_321_),
    .C(_211_),
    .Y(_322_)
);

OAI21X1 _2227_ (
    .A(_914__bF$buf0),
    .B(_984_),
    .C(RDY_bF$buf6),
    .Y(_1335_)
);

FILL FILL_7__2991_ (
);

FILL FILL_7__2151_ (
);

FILL FILL_0__1902_ (
);

FILL FILL_3__2891_ (
);

FILL FILL_3__2471_ (
);

FILL FILL_3__2051_ (
);

FILL FILL_5__2397_ (
);

FILL FILL_1__2389_ (
);

FILL FILL_3__3676_ (
);

FILL FILL_3__3256_ (
);

FILL FILL_4__2960_ (
);

FILL FILL_4__2540_ (
);

FILL FILL_4__2120_ (
);

FILL FILL_6__2886_ (
);

FILL FILL_6__2466_ (
);

AOI21X1 _3185_ (
    .A(_780_),
    .B(_784_),
    .C(_785_),
    .Y(_786_)
);

FILL FILL_6__2046_ (
);

FILL FILL_0__2860_ (
);

FILL FILL_2__2878_ (
);

FILL FILL_2__2458_ (
);

FILL FILL_0__2440_ (
);

FILL FILL_2__2038_ (
);

FILL FILL_0__2020_ (
);

AND2X2 _1918_ (
    .A(_1034_),
    .B(_1027__bF$buf0),
    .Y(_1035_)
);

FILL FILL_7__1842_ (
);

FILL FILL_0__3645_ (
);

FILL FILL_0__3225_ (
);

FILL FILL_7__2627_ (
);

FILL FILL_1__2601_ (
);

FILL FILL_3__2947_ (
);

FILL FILL_3__2527_ (
);

FILL FILL_3__2107_ (
);

FILL FILL_4__1811_ (
);

NOR2X1 _2876_ (
    .A(_1149__bF$buf0),
    .B(_530_),
    .Y(_531_)
);

INVX1 _2456_ (
    .A(_157_),
    .Y(_158_)
);

INVX1 _2036_ (
    .A(_1145_),
    .Y(_1146_)
);

FILL FILL_7__2380_ (
);

FILL FILL_3__2280_ (
);

FILL FILL_7__3585_ (
);

FILL FILL_1__2198_ (
);

FILL FILL_7__3165_ (
);

FILL FILL_0__2916_ (
);

FILL FILL_3__3485_ (
);

FILL FILL_3__3065_ (
);

FILL FILL_6__2695_ (
);

FILL FILL_6__2275_ (
);

FILL FILL_2__2687_ (
);

FILL FILL_2__2267_ (
);

FILL FILL_4__3554_ (
);

FILL FILL_4__3134_ (
);

FILL FILL_3__1971_ (
);

FILL FILL_0__3454_ (
);

FILL FILL_0__3034_ (
);

FILL FILL_5__1897_ (
);

FILL FILL_1__1889_ (
);

FILL FILL_7__2856_ (
);

FILL FILL_7__2016_ (
);

FILL FILL_1__2830_ (
);

FILL FILL_1__2410_ (
);

FILL FILL_3__2756_ (
);

FILL FILL_3__2336_ (
);

FILL FILL_5__3623_ (
);

FILL FILL_5__3203_ (
);

FILL FILL_1__3615_ (
);

FILL FILL_6__1966_ (
);

OAI21X1 _2685_ (
    .A(_355_),
    .B(_326_),
    .C(_356_),
    .Y(_357_)
);

INVX1 _2265_ (
    .A(cond_code[0]),
    .Y(_1373_)
);

FILL FILL_0__1940_ (
);

FILL FILL_2__1958_ (
);

FILL FILL_4__2825_ (
);

FILL FILL_4__2405_ (
);

FILL FILL_0__2725_ (
);

FILL FILL_0__2305_ (
);

FILL FILL_3__3294_ (
);

FILL FILL_6__2084_ (
);

FILL FILL_2__2496_ (
);

FILL FILL_2__2076_ (
);

NAND3X1 _1956_ (
    .A(_1071_),
    .B(_1072_),
    .C(_1066_),
    .Y(_1073_)
);

FILL FILL_7__1880_ (
);

FILL FILL_6__3289_ (
);

FILL FILL_3__1780_ (
);

FILL FILL_0__3263_ (
);

FILL FILL_7__2245_ (
);

FILL FILL_3__2985_ (
);

FILL FILL_3__2565_ (
);

FILL FILL_3__2145_ (
);

FILL FILL_5__3012_ (
);

FILL FILL_1__3004_ (
);

FILL FILL_6__1775_ (
);

AOI21X1 _2494_ (
    .A(AN),
    .B(_144_),
    .C(_189_),
    .Y(_190_)
);

NAND2X1 _2074_ (
    .A(IRHOLD_valid),
    .B(IRHOLD[7]),
    .Y(_1183_)
);

FILL FILL_2__1767_ (
);

FILL FILL_4__2634_ (
);

FILL FILL_4__2214_ (
);

BUFX2 _3699_ (
    .A(_1741_[2]),
    .Y(AB[2])
);

OAI21X1 _3279_ (
    .A(_850_),
    .B(_854_),
    .C(_843_),
    .Y(_855_)
);

FILL FILL_0__2954_ (
);

FILL FILL_0__2534_ (
);

FILL FILL_6__3501_ (
);

FILL FILL_0__2114_ (
);

FILL FILL_1__1910_ (
);

FILL FILL_3__1836_ (
);

FILL FILL_5__2703_ (
);

OAI21X1 _1765_ (
    .A(RDY_bF$buf3),
    .B(_891_),
    .C(_892_),
    .Y(DIMUX[6])
);

FILL FILL_4__3592_ (
);

FILL FILL_4__3172_ (
);

FILL FILL_6__3098_ (
);

FILL FILL_0__3492_ (
);

FILL FILL_0__3072_ (
);

FILL FILL_4__1905_ (
);

FILL FILL_7__2474_ (
);

FILL FILL_0__1805_ (
);

FILL FILL_3__2794_ (
);

FILL FILL_3__2374_ (
);

FILL FILL_5__3661_ (
);

FILL FILL_7__3259_ (
);

FILL FILL_5__3241_ (
);

FILL FILL_1__3653_ (
);

FILL FILL_1__3233_ (
);

FILL FILL_3__3579_ (
);

FILL FILL_3__3159_ (
);

FILL FILL_2__1996_ (
);

FILL FILL_4__2863_ (
);

FILL FILL_4__2443_ (
);

FILL FILL_4__2023_ (
);

FILL FILL_6__2789_ (
);

FILL FILL_6__2369_ (
);

MUX2X1 _3088_ (
    .A(ADD[1]),
    .B(AZ),
    .S(plp),
    .Y(_699_)
);

FILL FILL_0__2763_ (
);

FILL FILL_0__2343_ (
);

FILL FILL_6__3310_ (
);

FILL FILL_2__3302_ (
);

FILL FILL_7__1745_ (
);

FILL FILL_4__3648_ (
);

FILL FILL_4__3228_ (
);

FILL FILL_0__3548_ (
);

FILL FILL_0__3128_ (
);

FILL FILL_5__2932_ (
);

FILL FILL_5__2512_ (
);

FILL FILL_1__2924_ (
);

FILL FILL_1__2504_ (
);

NAND3X1 _1994_ (
    .A(_1107_),
    .B(_1105_),
    .C(_1106_),
    .Y(_1108_)
);

FILL FILL_1__3709_ (
);

OAI21X1 _2779_ (
    .A(_443_),
    .B(_440_),
    .C(RDY_bF$buf4),
    .Y(_444_)
);

MUX2X1 _2359_ (
    .A(_1464_),
    .B(_998_),
    .S(_886__bF$buf1),
    .Y(_1465_)
);

FILL FILL_7__2283_ (
);

OAI21X1 _3300_ (
    .A(_267_),
    .B(_860_),
    .C(_868_),
    .Y(_108_)
);

FILL FILL_3__2183_ (
);

FILL FILL_4__2919_ (
);

FILL FILL_7__3488_ (
);

FILL FILL_5__3470_ (
);

FILL FILL_5__3050_ (
);

FILL FILL_0__2819_ (
);

FILL FILL_1__3462_ (
);

FILL FILL_1__3042_ (
);

FILL FILL169950x21750 (
);

FILL FILL_4__2672_ (
);

FILL FILL_4__2252_ (
);

FILL FILL_6__2598_ (
);

FILL FILL_6__2178_ (
);

FILL FILL_0__2992_ (
);

FILL FILL_0__2572_ (
);

FILL FILL_0__2152_ (
);

FILL FILL_2__3531_ (
);

FILL FILL_2__3111_ (
);

FILL FILL_7__1974_ (
);

FILL FILL_4__3457_ (
);

FILL FILL_4__3037_ (
);

FILL FILL_3__1874_ (
);

FILL FILL_5__2741_ (
);

FILL FILL_7__2759_ (
);

FILL FILL_5__2321_ (
);

FILL FILL_1__2733_ (
);

FILL FILL_1__2313_ (
);

FILL FILL_7__3700_ (
);

FILL FILL_3__2659_ (
);

FILL FILL_3__2239_ (
);

FILL FILL_3__3600_ (
);

FILL FILL_5__3526_ (
);

FILL FILL_5__3106_ (
);

FILL FILL_1__3518_ (
);

FILL FILL_4__1943_ (
);

FILL FILL_6__1869_ (
);

NOR2X1 _2588_ (
    .A(_271_),
    .B(_274_),
    .Y(_275_)
);

OAI21X1 _2168_ (
    .A(RDY_bF$buf1),
    .B(_1275_),
    .C(_1276_),
    .Y(_1277_)
);

FILL FILL_7__2092_ (
);

FILL FILL_0__1843_ (
);

FILL FILL_6__2810_ (
);

FILL FILL_2__2802_ (
);

FILL FILL_4__2728_ (
);

FILL FILL_4__2308_ (
);

FILL FILL_0__2628_ (
);

FILL FILL_0__2208_ (
);

FILL FILL_1__3691_ (
);

FILL FILL_1__3271_ (
);

FILL FILL_3__3197_ (
);

FILL FILL_4__2481_ (
);

FILL FILL_4__2061_ (
);

FILL FILL_0__2381_ (
);

FILL FILL_2__2399_ (
);

NAND2X1 _1859_ (
    .A(_911_),
    .B(_957_),
    .Y(_984_)
);

FILL FILL_4__3266_ (
);

OAI21X1 _2800_ (
    .A(_888_),
    .B(_351_),
    .C(_462_),
    .Y(_463_)
);

FILL FILL_0__3586_ (
);

FILL FILL_0__3166_ (
);

FILL FILL_5__2970_ (
);

FILL FILL_7__2988_ (
);

FILL FILL_5__2550_ (
);

FILL FILL_7__2148_ (
);

FILL FILL_5__2130_ (
);

FILL FILL_1__2962_ (
);

FILL FILL_1__2542_ (
);

FILL FILL_1__2122_ (
);

FILL FILL_3__2888_ (
);

FILL FILL_3__2468_ (
);

FILL FILL_3__2048_ (
);

FILL FILL_4__1752_ (
);

NAND3X1 _2397_ (
    .A(_1448_),
    .B(_1496_),
    .C(_1501_),
    .Y(_1502_)
);

FILL FILL_2__2611_ (
);

FILL FILL_4__2957_ (
);

FILL FILL_4__2537_ (
);

FILL FILL_4__2117_ (
);

FILL FILL_0__2857_ (
);

FILL FILL_0__2437_ (
);

FILL FILL_0__2017_ (
);

FILL FILL_1__3080_ (
);

FILL FILL_5__1821_ (
);

FILL FILL_1__1813_ (
);

FILL FILL_4__2290_ (
);

FILL FILL_5__2606_ (
);

FILL FILL_0__2190_ (
);

FILL FILL_4__3495_ (
);

FILL FILL_4__3075_ (
);

FILL FILL_4__1808_ (
);

FILL FILL_7__2377_ (
);

FILL FILL_1__2771_ (
);

FILL FILL_1__2351_ (
);

FILL FILL_3__2697_ (
);

FILL FILL_3__2277_ (
);

FILL FILL_5__3564_ (
);

FILL FILL_5__3144_ (
);

FILL FILL_1__3556_ (
);

FILL FILL_1__3136_ (
);

FILL FILL_4__1981_ (
);

FILL FILL_0__1881_ (
);

FILL FILL_2__1899_ (
);

FILL FILL_2__2840_ (
);

FILL FILL_2__2420_ (
);

FILL FILL_2__2000_ (
);

FILL FILL_4__2766_ (
);

FILL FILL_4__2346_ (
);

FILL FILL_0__2666_ (
);

FILL FILL_6__3633_ (
);

FILL FILL_0__2246_ (
);

FILL FILL_6__3213_ (
);

FILL FILL_2__3625_ (
);

FILL FILL_2__3205_ (
);

FILL FILL_3__1968_ (
);

FILL FILL_5__2835_ (
);

FILL FILL_5__2415_ (
);

FILL FILL_1__2827_ (
);

FILL FILL_1__2407_ (
);

OAI22X1 _1897_ (
    .A(_1014_),
    .B(_968_),
    .C(_1015_),
    .D(_1004_),
    .Y(BI[6])
);

FILL FILL_0__1937_ (
);

FILL FILL_6__2904_ (
);

OAI21X1 _3623_ (
    .A(_1645_),
    .B(_1652_),
    .C(_1648_),
    .Y(_1653_)
);

OAI21X1 _3203_ (
    .A(_778_),
    .B(_789_),
    .C(_796_),
    .Y(_83_)
);

FILL FILL_1__2580_ (
);

FILL FILL_1__2160_ (
);

FILL FILL_3__2086_ (
);

FILL FILL_4__1790_ (
);

FILL FILL_4__2995_ (
);

FILL FILL_4__2575_ (
);

FILL FILL_4__2155_ (
);

FILL FILL_0__2895_ (
);

FILL FILL_0__2475_ (
);

FILL FILL_0__2055_ (
);

FILL FILL_6__3022_ (
);

FILL FILL_2__3014_ (
);

FILL FILL_7__1877_ (
);

FILL FILL_1__1851_ (
);

FILL FILL_3__1777_ (
);

FILL FILL_5__2644_ (
);

FILL FILL_5__2224_ (
);

FILL FILL_1__2636_ (
);

FILL FILL_7__3603_ (
);

FILL FILL_1__2216_ (
);

FILL FILL_3__3503_ (
);

FILL FILL_5__3009_ (
);

FILL FILL_2__1920_ (
);

FILL FILL_4__1846_ (
);

FILL FILL_0__1746_ (
);

FILL FILL_6__2713_ (
);

DFFSR _3432_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_100_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[3] [7])
);

NOR2X1 _3012_ (
    .A(_1214_),
    .B(_1213_),
    .Y(_638_)
);

FILL FILL_2__2705_ (
);

FILL FILL_5__3182_ (
);

FILL FILL_1_BUFX2_insert37 (
);

FILL FILL_1_BUFX2_insert38 (
);

FILL FILL_1_BUFX2_insert39 (
);

FILL FILL_1__3594_ (
);

FILL FILL_1__3174_ (
);

FILL FILL_5__1915_ (
);

FILL FILL_1__1907_ (
);

FILL FILL_4__2384_ (
);

FILL FILL_6__3671_ (
);

FILL FILL_0__2284_ (
);

FILL FILL_6__3251_ (
);

FILL FILL_2__3663_ (
);

FILL FILL_2__3243_ (
);

FILL FILL_4__3589_ (
);

FILL FILL_4__3169_ (
);

AOI21X1 _2703_ (
    .A(PC[4]),
    .B(_371_),
    .C(_373_),
    .Y(_374_)
);

FILL FILL_0__3489_ (
);

FILL FILL_0__3069_ (
);

FILL FILL_5__2873_ (
);

FILL FILL_5__2453_ (
);

FILL FILL_5__2033_ (
);

FILL FILL_1__2865_ (
);

FILL FILL_1__2445_ (
);

FILL FILL_1__2025_ (
);

FILL FILL_3__3312_ (
);

FILL FILL_5__3658_ (
);

FILL FILL_5__3238_ (
);

FILL FILL_0__1975_ (
);

FILL FILL_6__2942_ (
);

NAND2X1 _3661_ (
    .A(ADD[1]),
    .B(_1714__bF$buf1),
    .Y(_1688_)
);

FILL FILL_6__2522_ (
);

FILL FILL_6__2102_ (
);

OAI21X1 _3241_ (
    .A(_931__bF$buf3),
    .B(_1069_),
    .C(_1202_),
    .Y(_817_)
);

FILL FILL_2__2934_ (
);

FILL FILL_2__2514_ (
);

FILL FILL_6__3307_ (
);

FILL FILL_0__3701_ (
);

FILL FILL_4__2193_ (
);

FILL FILL_5__2929_ (
);

FILL FILL_5__2509_ (
);

FILL FILL_6__3480_ (
);

FILL FILL_0__2093_ (
);

FILL FILL_6__3060_ (
);

FILL FILL_2__3472_ (
);

FILL FILL_2__3052_ (
);

AOI22X1 _2932_ (
    .A(_543_),
    .B(_574_),
    .C(_572_),
    .D(_1351_),
    .Y(_575_)
);

NAND3X1 _2512_ (
    .A(_940_),
    .B(_1028_),
    .C(_1267_),
    .Y(_207_)
);

FILL FILL_0__3298_ (
);

FILL FILL_5__2682_ (
);

FILL FILL_5__2262_ (
);

FILL FILL_1__2674_ (
);

FILL FILL_1__2254_ (
);

FILL FILL_3__3541_ (
);

FILL FILL_3__3121_ (
);

FILL FILL_5__3467_ (
);

FILL FILL_5__3047_ (
);

FILL FILL_1__3459_ (
);

FILL FILL_1__3039_ (
);

FILL FILL_4__1884_ (
);

FILL FILL_0__1784_ (
);

FILL FILL_6__2751_ (
);

INVX2 _3470_ (
    .A(alu_op[1]),
    .Y(_1716_)
);

FILL FILL_6__2331_ (
);

OAI21X1 _3050_ (
    .A(_914__bF$buf4),
    .B(_989_),
    .C(DIMUX[6]),
    .Y(_665_)
);

FILL FILL_2__2743_ (
);

FILL FILL_2__2323_ (
);

FILL FILL_4__2669_ (
);

FILL FILL_4__2249_ (
);

FILL FILL_4__3610_ (
);

FILL FILL_0__2989_ (
);

FILL FILL_0__2569_ (
);

FILL FILL_6__3536_ (
);

FILL FILL_0__2149_ (
);

FILL FILL_6__3116_ (
);

FILL FILL_2__3528_ (
);

FILL FILL_0__3510_ (
);

FILL FILL_2__3108_ (
);

FILL FILL_5__1953_ (
);

FILL FILL_1__1945_ (
);

FILL FILL_7__2912_ (
);

FILL FILL_3__2812_ (
);

FILL FILL_5__2738_ (
);

FILL FILL_5__2318_ (
);

FILL FILL_2_BUFX2_insert80 (
);

FILL FILL_2_BUFX2_insert81 (
);

FILL FILL_2_BUFX2_insert82 (
);

FILL FILL_2_BUFX2_insert83 (
);

FILL FILL_2__3281_ (
);

NOR3X1 _2741_ (
    .A(_403_),
    .B(_404_),
    .C(_407_),
    .Y(_408_)
);

OAI21X1 _2321_ (
    .A(_941_),
    .B(_1427_),
    .C(_903__bF$buf0),
    .Y(_1428_)
);

FILL FILL_5__2491_ (
);

FILL FILL_5__2071_ (
);

FILL FILL_6__2807_ (
);

NAND2X1 _3526_ (
    .A(_1722_),
    .B(_1555_),
    .Y(_1556_)
);

INVX1 _3106_ (
    .A(backwards),
    .Y(_715_)
);

FILL FILL_1__2483_ (
);

FILL FILL_7__3450_ (
);

FILL FILL_1__2063_ (
);

FILL FILL_7__3030_ (
);

FILL FILL_5__3696_ (
);

FILL FILL_5__3276_ (
);

FILL FILL_1__3268_ (
);

FILL FILL_6__2980_ (
);

FILL FILL_6__2560_ (
);

FILL FILL_6__2140_ (
);

FILL FILL_2__2972_ (
);

FILL FILL_2__2552_ (
);

FILL FILL_2__2132_ (
);

FILL FILL_4__2898_ (
);

FILL FILL_4__2478_ (
);

FILL FILL_4__2058_ (
);

FILL FILL_0__2798_ (
);

FILL FILL_0__2378_ (
);

FILL FILL_5__1762_ (
);

FILL FILL_1__1754_ (
);

FILL FILL_7__2301_ (
);

FILL FILL_3__2621_ (
);

FILL FILL_3__2201_ (
);

FILL FILL_5__2967_ (
);

FILL FILL_5__2547_ (
);

FILL FILL_5__2127_ (
);

FILL FILL_1__2959_ (
);

FILL FILL_1__2539_ (
);

FILL FILL_7__3506_ (
);

FILL FILL_1__2119_ (
);

FILL FILL_2__3090_ (
);

OAI21X1 _2970_ (
    .A(_886__bF$buf5),
    .B(_1027__bF$buf0),
    .C(store),
    .Y(_602_)
);

FILL FILL_6__1831_ (
);

AOI21X1 _2550_ (
    .A(_1108_),
    .B(_195_),
    .C(_241_),
    .Y(_242_)
);

OAI21X1 _2130_ (
    .A(RDY_bF$buf8),
    .B(_1222_),
    .C(_1238_),
    .Y(_1239_)
);

FILL FILL_2__1823_ (
);

FILL FILL_4__1749_ (
);

FILL FILL_6__2616_ (
);

DFFSR _3335_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_13_),
    .CLK(clk_bF$buf2),
    .Q(PC[11])
);

FILL FILL_1__2292_ (
);

FILL FILL_2__2608_ (
);

FILL FILL_5__3085_ (
);

FILL FILL_1__3497_ (
);

FILL FILL_1__3077_ (
);

FILL FILL_5__1818_ (
);

FILL FILL_2__2781_ (
);

FILL FILL_2__2361_ (
);

FILL FILL_4__2287_ (
);

NOR2X1 _1821_ (
    .A(_902__bF$buf1),
    .B(_946_),
    .Y(_947_)
);

FILL FILL_6__3574_ (
);

FILL FILL_0__2187_ (
);

FILL FILL_6__3154_ (
);

FILL FILL_2__3566_ (
);

FILL FILL_2__3146_ (
);

FILL FILL_5__1991_ (
);

OAI21X1 _2606_ (
    .A(_285_),
    .B(_218_),
    .C(_289_),
    .Y(_1741_[11])
);

FILL FILL_1__1983_ (
);

FILL FILL_7__2530_ (
);

FILL FILL_3__2850_ (
);

FILL FILL_3__2430_ (
);

FILL FILL_3__2010_ (
);

FILL FILL_5__2776_ (
);

FILL FILL_5__2356_ (
);

FILL FILL_1__2768_ (
);

FILL FILL_1__2348_ (
);

FILL FILL_7__3315_ (
);

FILL FILL_3__3635_ (
);

FILL FILL_3__3215_ (
);

FILL FILL_4__1978_ (
);

FILL FILL_0__1878_ (
);

FILL FILL_6__2845_ (
);

NOR2X1 _3564_ (
    .A(_1570_),
    .B(_1568_),
    .Y(_1594_)
);

FILL FILL_6__2425_ (
);

FILL FILL_6__2005_ (
);

NAND2X1 _3144_ (
    .A(ADD[3]),
    .B(_731_),
    .Y(_749_)
);

FILL FILL_2__2837_ (
);

FILL FILL_2__2417_ (
);

FILL FILL_7__1801_ (
);

FILL FILL_4__3704_ (
);

FILL FILL_0__3604_ (
);

FILL FILL_2__2590_ (
);

FILL FILL_2__2170_ (
);

FILL FILL_4__2096_ (
);

FILL FILL_3__2906_ (
);

FILL FILL_6_BUFX2_insert37 (
);

FILL FILL_6_BUFX2_insert38 (
);

FILL FILL_6_BUFX2_insert39 (
);

INVX1 _2835_ (
    .A(_495_),
    .Y(_497_)
);

NAND3X1 _2415_ (
    .A(_1259_),
    .B(_1318_),
    .C(_123_),
    .Y(_124_)
);

FILL FILL_1__1792_ (
);

FILL FILL_5__2585_ (
);

FILL FILL_5__2165_ (
);

FILL FILL_1__2997_ (
);

FILL FILL_1__2577_ (
);

FILL FILL_1__2157_ (
);

FILL FILL_7__3124_ (
);

FILL FILL_3__3024_ (
);

FILL FILL_2__1861_ (
);

FILL FILL_4__1787_ (
);

FILL FILL_6__2654_ (
);

DFFSR _3373_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_50_),
    .CLK(clk_bF$buf10),
    .Q(dst_reg[1])
);

FILL FILL_6__2234_ (
);

FILL FILL_2__2646_ (
);

FILL FILL_2__2226_ (
);

FILL FILL_4__3513_ (
);

FILL FILL_6__3019_ (
);

FILL FILL_3__1930_ (
);

FILL FILL_5__1856_ (
);

FILL FILL_1__1848_ (
);

FILL FILL_3__2715_ (
);

FILL FILL_6__3192_ (
);

FILL FILL_2__3184_ (
);

FILL FILL_6__1925_ (
);

AND2X2 _2644_ (
    .A(_317_),
    .B(_318_),
    .Y(_319_)
);

NOR2X1 _2224_ (
    .A(_1173_),
    .B(_1215_),
    .Y(_1332_)
);

FILL FILL_2__1917_ (
);

FILL FILL_5__2394_ (
);

DFFSR _3429_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_97_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[3] [4])
);

NAND2X1 _3009_ (
    .A(_603_),
    .B(_552_),
    .Y(_635_)
);

FILL FILL168150x61350 (
);

FILL FILL_1__2386_ (
);

FILL FILL_3__3673_ (
);

FILL FILL_3__3253_ (
);

FILL FILL_5__3599_ (
);

FILL FILL_5__3179_ (
);

FILL FILL_6__2883_ (
);

FILL FILL_6__2463_ (
);

FILL FILL_6__2043_ (
);

NAND2X1 _3182_ (
    .A(_781_),
    .B(_782_),
    .Y(_783_)
);

FILL FILL_2__2875_ (
);

FILL FILL_2__2455_ (
);

FILL FILL_2__2035_ (
);

NAND2X1 _1915_ (
    .A(_1030_),
    .B(_1031_),
    .Y(_1032_)
);

FILL FILL_1_BUFX2_insert0 (
);

FILL FILL_6__3668_ (
);

FILL FILL_6__3248_ (
);

FILL FILL_1_BUFX2_insert1 (
);

FILL FILL_1_BUFX2_insert2 (
);

FILL FILL_1_BUFX2_insert3 (
);

FILL FILL_1_BUFX2_insert4 (
);

FILL FILL_1_BUFX2_insert5 (
);

FILL FILL_1_BUFX2_insert6 (
);

FILL FILL_1_BUFX2_insert7 (
);

FILL FILL_1_BUFX2_insert8 (
);

FILL FILL_1_BUFX2_insert9 (
);

FILL FILL_0__3642_ (
);

FILL FILL_0__3222_ (
);

FILL FILL_7__2624_ (
);

FILL FILL_7__2204_ (
);

FILL FILL_3__2944_ (
);

FILL FILL_3__2524_ (
);

FILL FILL_3__2104_ (
);

FILL FILL_3__3309_ (
);

OAI21X1 _2873_ (
    .A(_886__bF$buf5),
    .B(_1185_),
    .C(_528_),
    .Y(_21_)
);

OAI21X1 _2453_ (
    .A(_1334_),
    .B(_154_),
    .C(Z),
    .Y(_155_)
);

INVX1 _2033_ (
    .A(_1142_),
    .Y(_1143_)
);

FILL FILL_6__2939_ (
);

OAI21X1 _3658_ (
    .A(_1580_),
    .B(_1610_),
    .C(_1611_),
    .Y(_1686_)
);

FILL FILL_6__2519_ (
);

OAI21X1 _3238_ (
    .A(_778_),
    .B(_807_),
    .C(_815_),
    .Y(_99_)
);

FILL FILL_7__3582_ (
);

FILL FILL_1__2195_ (
);

FILL FILL_7__3162_ (
);

FILL FILL_0__2913_ (
);

FILL FILL_3__3482_ (
);

FILL FILL_3__3062_ (
);

FILL FILL_6__2692_ (
);

FILL FILL_6__2272_ (
);

FILL FILL_2__2684_ (
);

FILL FILL_2__2264_ (
);

FILL FILL_4__3551_ (
);

FILL FILL_4__3131_ (
);

FILL FILL_6__3477_ (
);

FILL FILL_6__3057_ (
);

FILL FILL_0__3451_ (
);

FILL FILL_2__3469_ (
);

FILL FILL_2__3049_ (
);

FILL FILL_0__3031_ (
);

FILL FILL_5__1894_ (
);

AND2X2 _2929_ (
    .A(_543_),
    .B(_1178_),
    .Y(_572_)
);

OAI21X1 _2509_ (
    .A(_993_),
    .B(_992_),
    .C(_903__bF$buf3),
    .Y(_204_)
);

FILL FILL_1__1886_ (
);

FILL FILL_7__2853_ (
);

FILL FILL_7__2433_ (
);

FILL FILL_7__2013_ (
);

FILL FILL_3__2753_ (
);

FILL FILL_3__2333_ (
);

FILL FILL_5__2679_ (
);

FILL FILL_5__2259_ (
);

FILL FILL_7__3638_ (
);

FILL FILL_5__3620_ (
);

FILL FILL_5__3200_ (
);

FILL FILL_1__3612_ (
);

FILL FILL_3__3538_ (
);

FILL FILL_3__3118_ (
);

FILL FILL_6__1963_ (
);

AOI21X1 _2682_ (
    .A(_352_),
    .B(_353_),
    .C(_1009_),
    .Y(_354_)
);

NOR2X1 _2262_ (
    .A(_1188_),
    .B(_1355_),
    .Y(_1370_)
);

FILL FILL_2__1955_ (
);

FILL FILL_4__2822_ (
);

FILL FILL_4__2402_ (
);

FILL FILL_6__2748_ (
);

INVX4 _3467_ (
    .A(reset),
    .Y(_1513_)
);

FILL FILL_6__2328_ (
);

INVX1 _3047_ (
    .A(_661_),
    .Y(_662_)
);

FILL FILL_0__2722_ (
);

FILL FILL_0__2302_ (
);

FILL FILL_3__3291_ (
);

FILL FILL_4__3607_ (
);

FILL FILL_0__3507_ (
);

FILL FILL_6__2081_ (
);

FILL FILL_7__2909_ (
);

FILL FILL_2__2493_ (
);

FILL FILL_2__2073_ (
);

FILL FILL_3__2809_ (
);

OAI21X1 _1953_ (
    .A(_914__bF$buf2),
    .B(_1069_),
    .C(_1032_),
    .Y(_1070_)
);

FILL FILL_6__3286_ (
);

FILL FILL_2__3698_ (
);

FILL FILL_0__3260_ (
);

FILL FILL_2__3278_ (
);

NAND2X1 _2738_ (
    .A(ADD[0]),
    .B(_1299_),
    .Y(_405_)
);

NOR2X1 _2318_ (
    .A(_1424_),
    .B(_916_),
    .Y(_1425_)
);

FILL FILL_7__2662_ (
);

FILL FILL_7__2242_ (
);

FILL FILL_3__2982_ (
);

FILL FILL_3__2562_ (
);

FILL FILL_3__2142_ (
);

FILL FILL_5__2488_ (
);

FILL FILL_5__2068_ (
);

FILL FILL_7__3027_ (
);

FILL FILL_1__3001_ (
);

FILL FILL_6__1772_ (
);

OAI21X1 _2491_ (
    .A(_143_),
    .B(_1133_),
    .C(_187_),
    .Y(_1742_[6])
);

OAI21X1 _2071_ (
    .A(_1168_),
    .B(IRHOLD[5]),
    .C(_1167_),
    .Y(_1180_)
);

FILL FILL_2__1764_ (
);

FILL FILL_4__2631_ (
);

FILL FILL_4__2211_ (
);

FILL FILL_6__2977_ (
);

BUFX2 _3696_ (
    .A(_1741_[13]),
    .Y(AB[13])
);

FILL FILL_6__2557_ (
);

NOR2X1 _3276_ (
    .A(_975_),
    .B(_851_),
    .Y(_852_)
);

FILL FILL_6__2137_ (
);

FILL FILL_0__2951_ (
);

FILL FILL_2__2969_ (
);

FILL FILL_2__2549_ (
);

FILL FILL_0__2531_ (
);

FILL FILL_2__2129_ (
);

FILL FILL_0__2111_ (
);

FILL FILL_3__1833_ (
);

FILL FILL_0__3316_ (
);

FILL FILL_5__1759_ (
);

FILL FILL_5__2700_ (
);

FILL FILL_3__2618_ (
);

OAI21X1 _1762_ (
    .A(RDY_bF$buf4),
    .B(_889_),
    .C(_890_),
    .Y(DIMUX[5])
);

FILL FILL_6__3095_ (
);

FILL FILL_2__3087_ (
);

FILL FILL_4__1902_ (
);

FILL FILL_6__1828_ (
);

NAND2X1 _2967_ (
    .A(_1150__bF$buf0),
    .B(_596_),
    .Y(_600_)
);

OAI22X1 _2547_ (
    .A(_1010_),
    .B(_201_),
    .C(_238_),
    .D(_199_),
    .Y(_239_)
);

NAND2X1 _2127_ (
    .A(_886__bF$buf0),
    .B(_1235_),
    .Y(_1236_)
);

FILL FILL_7__2891_ (
);

FILL FILL_7__2471_ (
);

FILL FILL_7__2051_ (
);

FILL FILL_0__1802_ (
);

FILL FILL_3__2791_ (
);

FILL FILL_3__2371_ (
);

FILL FILL_5__2297_ (
);

FILL FILL_1__2289_ (
);

FILL FILL_7__3256_ (
);

FILL FILL_1__3650_ (
);

FILL FILL_1__3230_ (
);

FILL FILL_3__3576_ (
);

FILL FILL_3__3156_ (
);

FILL FILL_2__1993_ (
);

FILL FILL_4__2860_ (
);

FILL FILL_4__2440_ (
);

FILL FILL_4__2020_ (
);

FILL FILL_6__2786_ (
);

FILL FILL_6__2366_ (
);

OAI21X1 _3085_ (
    .A(_1377_),
    .B(_690_),
    .C(_696_),
    .Y(_65_)
);

FILL FILL_2__2778_ (
);

FILL FILL_0__2760_ (
);

FILL FILL_2__2358_ (
);

FILL FILL_0__2340_ (
);

INVX1 _1818_ (
    .A(_943_),
    .Y(_944_)
);

FILL FILL_4__3645_ (
);

FILL FILL_4__3225_ (
);

FILL FILL_0__3545_ (
);

FILL FILL_0__3125_ (
);

FILL FILL_5__1988_ (
);

FILL FILL_3_BUFX2_insert0 (
);

FILL FILL_3_BUFX2_insert1 (
);

FILL FILL_3_BUFX2_insert2 (
);

FILL FILL_3_BUFX2_insert3 (
);

FILL FILL_3_BUFX2_insert4 (
);

FILL FILL_3_BUFX2_insert5 (
);

FILL FILL_7__2527_ (
);

FILL FILL_3_BUFX2_insert6 (
);

FILL FILL_3_BUFX2_insert7 (
);

FILL FILL_3_BUFX2_insert8 (
);

FILL FILL_3_BUFX2_insert9 (
);

FILL FILL_1__2921_ (
);

FILL FILL_1__2501_ (
);

FILL FILL_3__2847_ (
);

FILL FILL_3__2427_ (
);

FILL FILL_3__2007_ (
);

NAND2X1 _1991_ (
    .A(\AXYS[1] [3]),
    .B(_1047_),
    .Y(_1105_)
);

FILL FILL_5__3714_ (
);

FILL FILL_1__3706_ (
);

NAND2X1 _2776_ (
    .A(_280_),
    .B(_365_),
    .Y(_441_)
);

NAND3X1 _2356_ (
    .A(_1441_),
    .B(_1451_),
    .C(_1461_),
    .Y(_1462_)
);

FILL FILL_7__2280_ (
);

FILL FILL_3__2180_ (
);

FILL FILL_4__2916_ (
);

FILL FILL_7__3485_ (
);

FILL FILL_1__2098_ (
);

FILL FILL_7__3065_ (
);

FILL FILL_0__2816_ (
);

FILL FILL_6__2595_ (
);

FILL FILL_6__2175_ (
);

FILL FILL_2__2587_ (
);

FILL FILL_2__2167_ (
);

FILL FILL_7__1971_ (
);

FILL FILL_4__3454_ (
);

FILL FILL_4__3034_ (
);

FILL FILL_3__1871_ (
);

FILL FILL_5__1797_ (
);

FILL FILL_1__1789_ (
);

FILL FILL_7__2756_ (
);

FILL FILL_1__2730_ (
);

FILL FILL_1__2310_ (
);

FILL FILL_3__2656_ (
);

FILL FILL_3__2236_ (
);

FILL FILL_5__3523_ (
);

FILL FILL_5__3103_ (
);

FILL FILL_1__3515_ (
);

FILL FILL_4__1940_ (
);

FILL FILL_6__1866_ (
);

INVX2 _2585_ (
    .A(_215_),
    .Y(_272_)
);

AOI21X1 _2165_ (
    .A(_1271_),
    .B(_1273_),
    .C(_1270_),
    .Y(_1274_)
);

FILL FILL_0__1840_ (
);

FILL FILL_2__1858_ (
);

FILL FILL_4__2725_ (
);

FILL FILL_4__2305_ (
);

FILL FILL_7__3294_ (
);

FILL FILL_0__2625_ (
);

FILL FILL_0__2205_ (
);

FILL FILL169050x133350 (
);

FILL FILL_3__3194_ (
);

FILL FILL_3__1927_ (
);

FILL FILL_2__2396_ (
);

INVX1 _1856_ (
    .A(_900_),
    .Y(_981_)
);

FILL FILL_7__1780_ (
);

FILL FILL_4__3263_ (
);

FILL FILL_6__3189_ (
);

FILL FILL_0__3583_ (
);

FILL FILL_0__3163_ (
);

FILL FILL_7__2985_ (
);

FILL FILL_7__2145_ (
);

FILL FILL_3__2885_ (
);

FILL FILL_3__2465_ (
);

FILL FILL_3__2045_ (
);

NAND3X1 _2394_ (
    .A(_1197_),
    .B(_1497_),
    .C(_1498_),
    .Y(_1499_)
);

FILL FILL169350x3750 (
);

FILL FILL_4__2954_ (
);

FILL FILL_4__2534_ (
);

FILL FILL_4__2114_ (
);

OAI21X1 _3599_ (
    .A(_1533_),
    .B(_1628_),
    .C(_1536_),
    .Y(_1629_)
);

OAI21X1 _3179_ (
    .A(_769_),
    .B(_759_),
    .C(_773_),
    .Y(_780_)
);

FILL FILL_0__2854_ (
);

FILL FILL_0__2434_ (
);

FILL FILL_0__2014_ (
);

FILL FILL_1__1810_ (
);

FILL FILL_0__3639_ (
);

FILL FILL_0__3219_ (
);

FILL FILL_5__2603_ (
);

FILL FILL_4__3492_ (
);

FILL FILL_4__3072_ (
);

FILL FILL_4__1805_ (
);

FILL FILL_7__2374_ (
);

FILL FILL_3__2694_ (
);

FILL FILL_3__2274_ (
);

FILL FILL_7__3579_ (
);

FILL FILL_5__3561_ (
);

FILL FILL_7__3159_ (
);

FILL FILL_5__3141_ (
);

FILL FILL_1__3553_ (
);

FILL FILL_1__3133_ (
);

FILL FILL_3__3479_ (
);

FILL FILL_3__3059_ (
);

FILL FILL_2__1896_ (
);

FILL FILL_4__2763_ (
);

FILL FILL_4__2343_ (
);

FILL FILL_6__2689_ (
);

FILL FILL_6__2269_ (
);

FILL FILL_0__2663_ (
);

FILL FILL_6__3630_ (
);

FILL FILL_0__2243_ (
);

FILL FILL_6__3210_ (
);

FILL FILL_2__3622_ (
);

FILL FILL_2__3202_ (
);

FILL FILL_4__3548_ (
);

FILL FILL_4__3128_ (
);

FILL FILL_3__1965_ (
);

FILL FILL_0__3028_ (
);

FILL FILL_5__2832_ (
);

FILL FILL_5__2412_ (
);

FILL FILL_1__2824_ (
);

FILL FILL_1__2404_ (
);

OAI22X1 _1894_ (
    .A(_1012_),
    .B(_968_),
    .C(_1013_),
    .D(_1004_),
    .Y(BI[5])
);

FILL FILL_5__3617_ (
);

FILL FILL_1__3609_ (
);

NOR2X1 _2679_ (
    .A(_1291_),
    .B(_325_),
    .Y(_351_)
);

NOR2X1 _2259_ (
    .A(_1366_),
    .B(_1355_),
    .Y(_1367_)
);

FILL FILL_0__1934_ (
);

FILL FILL_6__2901_ (
);

AOI22X1 _3620_ (
    .A(_1724_),
    .B(_1729_),
    .C(_1639_),
    .D(_1649_),
    .Y(_1650_)
);

OAI21X1 _3200_ (
    .A(_720__bF$buf1),
    .B(_687_),
    .C(\AXYS[1] [5]),
    .Y(_795_)
);

FILL FILL_3__2083_ (
);

FILL FILL_4__2819_ (
);

FILL FILL_0__2719_ (
);

FILL FILL_3__3288_ (
);

FILL FILL_4__2992_ (
);

FILL FILL_4__2572_ (
);

FILL FILL_4__2152_ (
);

FILL FILL_6__2498_ (
);

FILL FILL_6__2078_ (
);

FILL FILL_0__2892_ (
);

FILL FILL_0__2472_ (
);

FILL FILL_0__2052_ (
);

FILL FILL_2__3011_ (
);

FILL FILL_7__1874_ (
);

FILL FILL_0__3677_ (
);

FILL FILL_3__1774_ (
);

FILL FILL_0__3257_ (
);

FILL FILL_7__2659_ (
);

FILL FILL_5__2641_ (
);

FILL FILL_5__2221_ (
);

FILL FILL_1__2633_ (
);

FILL FILL_7__3600_ (
);

FILL FILL_1__2213_ (
);

FILL FILL_3__2979_ (
);

FILL FILL_3__2559_ (
);

FILL FILL_3__2139_ (
);

FILL FILL_3__3500_ (
);

FILL FILL_5__3006_ (
);

FILL FILL_4__1843_ (
);

FILL FILL_6__1769_ (
);

AOI21X1 _2488_ (
    .A(ADD[6]),
    .B(_144_),
    .C(_184_),
    .Y(_185_)
);

OAI21X1 _2068_ (
    .A(IRHOLD_valid),
    .B(_888_),
    .C(_1176_),
    .Y(_1177_)
);

FILL FILL_6__2710_ (
);

FILL FILL_2__2702_ (
);

FILL FILL_4__2628_ (
);

FILL FILL_4__2208_ (
);

FILL FILL_0__2948_ (
);

FILL FILL_0__2528_ (
);

FILL FILL_0__2108_ (
);

FILL FILL_1__3591_ (
);

FILL FILL_1__3171_ (
);

FILL FILL_3__3097_ (
);

FILL FILL_5__1912_ (
);

FILL FILL_1__1904_ (
);

FILL FILL_4__2381_ (
);

FILL FILL_0__2281_ (
);

FILL FILL_2__2299_ (
);

FILL FILL_2__3660_ (
);

FILL FILL_2__3240_ (
);

INVX1 _1759_ (
    .A(_888_),
    .Y(DIMUX[4])
);

FILL FILL_4__3586_ (
);

FILL FILL_4__3166_ (
);

OAI21X1 _2700_ (
    .A(_364_),
    .B(_322_),
    .C(_353_),
    .Y(_371_)
);

FILL FILL_0__3486_ (
);

FILL FILL_0__3066_ (
);

FILL FILL_5__2870_ (
);

FILL FILL_7__2888_ (
);

FILL FILL_5__2450_ (
);

FILL FILL_5__2030_ (
);

FILL FILL_7__2048_ (
);

FILL FILL_1__2862_ (
);

FILL FILL_1__2442_ (
);

FILL FILL_1__2022_ (
);

FILL FILL_3__2788_ (
);

FILL FILL_3__2368_ (
);

FILL FILL_5__3655_ (
);

FILL FILL_5__3235_ (
);

FILL FILL_1__3647_ (
);

FILL FILL_1__3227_ (
);

FILL FILL_6__1998_ (
);

INVX1 _2297_ (
    .A(_1156_),
    .Y(_1404_)
);

FILL FILL_0__1972_ (
);

FILL FILL_2__2931_ (
);

FILL FILL_2__2511_ (
);

FILL FILL_4__2857_ (
);

FILL FILL_4__2437_ (
);

FILL FILL_4__2017_ (
);

FILL FILL_0__2757_ (
);

FILL FILL_0__2337_ (
);

FILL FILL_6__3304_ (
);

FILL FILL_4__2190_ (
);

FILL FILL_5__2926_ (
);

FILL FILL_5__2506_ (
);

FILL FILL_0__2090_ (
);

FILL FILL_1__2918_ (
);

OAI22X1 _1988_ (
    .A(_1102_),
    .B(_1092_),
    .C(_1008_),
    .D(_983_),
    .Y(_1103_)
);

FILL FILL_0__3295_ (
);

FILL FILL_7__2277_ (
);

BUFX2 _3714_ (
    .A(_1742_[7]),
    .Y(DO[7])
);

FILL FILL_1__2671_ (
);

FILL FILL_1__2251_ (
);

FILL FILL_3__2597_ (
);

FILL FILL_3__2177_ (
);

FILL FILL_5__3464_ (
);

FILL FILL_5__3044_ (
);

FILL FILL_1__3456_ (
);

FILL FILL_1__3036_ (
);

FILL FILL_4__1881_ (
);

FILL FILL_2__1799_ (
);

FILL FILL_0__1781_ (
);

FILL FILL_2__2740_ (
);

FILL FILL_2__2320_ (
);

FILL FILL_4__2666_ (
);

FILL FILL_4__2246_ (
);

FILL FILL_0__2986_ (
);

FILL FILL_0__2566_ (
);

FILL FILL_6__3533_ (
);

FILL FILL_0__2146_ (
);

FILL FILL_6__3113_ (
);

FILL FILL_2__3525_ (
);

FILL FILL_2__3105_ (
);

FILL FILL_5__1950_ (
);

FILL FILL_1__1942_ (
);

FILL FILL_3__1868_ (
);

FILL FILL_5__2735_ (
);

FILL FILL_5__2315_ (
);

FILL FILL_2_BUFX2_insert50 (
);

FILL FILL_2_BUFX2_insert51 (
);

FILL FILL_2_BUFX2_insert52 (
);

FILL FILL_2_BUFX2_insert53 (
);

FILL FILL_2_BUFX2_insert54 (
);

FILL FILL_2_BUFX2_insert55 (
);

FILL FILL_2_BUFX2_insert56 (
);

FILL FILL_1__2727_ (
);

FILL FILL_2_BUFX2_insert57 (
);

FILL FILL_2_BUFX2_insert58 (
);

FILL FILL_1__2307_ (
);

FILL FILL_2_BUFX2_insert59 (
);

OAI22X1 _1797_ (
    .A(_909_),
    .B(_922_),
    .C(_921_),
    .D(_917_),
    .Y(_923_)
);

FILL FILL_4__1937_ (
);

FILL FILL_0__1837_ (
);

FILL FILL_6__2804_ (
);

INVX1 _3523_ (
    .A(BI[2]),
    .Y(_1553_)
);

OAI21X1 _3103_ (
    .A(_704_),
    .B(_711_),
    .C(_712_),
    .Y(_713_)
);

FILL FILL_1__2480_ (
);

FILL FILL_1__2060_ (
);

FILL FILL_5__3693_ (
);

FILL FILL_5__3273_ (
);

FILL FILL_1__3265_ (
);

FILL FILL_4__2895_ (
);

FILL FILL_4__2475_ (
);

FILL FILL_4__2055_ (
);

FILL FILL_0__2795_ (
);

FILL FILL_0__2375_ (
);

FILL FILL_7__1777_ (
);

FILL FILL_1__1751_ (
);

FILL FILL_5__2964_ (
);

FILL FILL_5__2544_ (
);

FILL FILL_5__2124_ (
);

FILL FILL_1__2956_ (
);

FILL FILL_1__2536_ (
);

FILL FILL_7__3503_ (
);

FILL FILL_1__2116_ (
);

FILL FILL_2__1820_ (
);

FILL FILL_4__1746_ (
);

FILL FILL_6__2613_ (
);

DFFSR _3332_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(_10_),
    .CLK(clk_bF$buf2),
    .Q(PC[8])
);

FILL FILL_2__2605_ (
);

FILL FILL_5__3082_ (
);

FILL FILL_1__3494_ (
);

FILL FILL_1__3074_ (
);

FILL FILL_5__1815_ (
);

FILL FILL_1__1807_ (
);

FILL FILL_4__2284_ (
);

FILL FILL_6__3571_ (
);

FILL FILL_0__2184_ (
);

FILL FILL_6__3151_ (
);

FILL FILL_2__3563_ (
);

FILL FILL_2__3143_ (
);

FILL FILL_4__3489_ (
);

FILL FILL_4__3069_ (
);

OAI21X1 _2603_ (
    .A(_925_),
    .B(_196_),
    .C(ABH[3]),
    .Y(_287_)
);

FILL FILL_1__1980_ (
);

FILL FILL_5__2773_ (
);

FILL FILL_5__2353_ (
);

FILL FILL_1__2765_ (
);

FILL FILL_1__2345_ (
);

FILL FILL_7__3312_ (
);

FILL FILL_3__3632_ (
);

FILL FILL_3__3212_ (
);

FILL FILL_5__3558_ (
);

FILL FILL_5__3138_ (
);

FILL FILL_4__1975_ (
);

FILL FILL_0__1875_ (
);

FILL FILL_6__2842_ (
);

NAND2X1 _3561_ (
    .A(_1590_),
    .B(_1589_),
    .Y(_1591_)
);

FILL FILL_6__2422_ (
);

FILL FILL_6__2002_ (
);

NOR2X1 _3141_ (
    .A(_732_),
    .B(_741_),
    .Y(_746_)
);

FILL FILL_2__2834_ (
);

FILL FILL_2__2414_ (
);

FILL FILL_4__3701_ (
);

FILL FILL_6__3627_ (
);

FILL FILL_6__3207_ (
);

FILL FILL_0__3601_ (
);

FILL FILL_2__3619_ (
);

FILL FILL_4__2093_ (
);

FILL FILL_3__2903_ (
);

FILL FILL_5__2829_ (
);

FILL FILL_5__2409_ (
);

FILL FILL_4__3298_ (
);

NOR2X1 _2832_ (
    .A(_295_),
    .B(_352_),
    .Y(_494_)
);

NAND2X1 _2412_ (
    .A(_119_),
    .B(_120_),
    .Y(_121_)
);

FILL FILL_0__3198_ (
);

FILL FILL_5__2582_ (
);

FILL FILL_5__2162_ (
);

OAI21X1 _3617_ (
    .A(BI[6]),
    .B(_1739_),
    .C(_1646_),
    .Y(_1647_)
);

FILL FILL_1__2994_ (
);

FILL FILL_1__2574_ (
);

FILL FILL_1__2154_ (
);

FILL FILL_3__3021_ (
);

FILL FILL_4__1784_ (
);

FILL FILL_6__2651_ (
);

FILL FILL_6__2231_ (
);

DFFSR _3370_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_47_),
    .CLK(clk_bF$buf10),
    .Q(src_reg[0])
);

FILL FILL_2__2643_ (
);

FILL FILL_2__2223_ (
);

FILL FILL_4__2989_ (
);

FILL FILL_4__2569_ (
);

FILL FILL_4__2149_ (
);

FILL FILL_4__3510_ (
);

FILL FILL_0__2889_ (
);

FILL FILL_0__2469_ (
);

FILL FILL_0__2049_ (
);

FILL FILL_6__3016_ (
);

FILL FILL_2__3008_ (
);

FILL FILL_5__1853_ (
);

FILL FILL_1__1845_ (
);

FILL FILL_7__2812_ (
);

FILL FILL_3__2712_ (
);

FILL FILL_5__2638_ (
);

FILL FILL_5__2218_ (
);

FILL FILL_2__3181_ (
);

FILL FILL_6__1922_ (
);

NOR2X1 _2641_ (
    .A(_311_),
    .B(_315_),
    .Y(_316_)
);

INVX1 _2221_ (
    .A(_1328_),
    .Y(_1329_)
);

FILL FILL_2__1914_ (
);

FILL FILL_5__2391_ (
);

FILL FILL_6__2707_ (
);

DFFSR _3426_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_94_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[3] [1])
);

NAND2X1 _3006_ (
    .A(_632_),
    .B(_630_),
    .Y(_50_)
);

FILL FILL_1__2383_ (
);

FILL FILL_3__3670_ (
);

FILL FILL_3__3250_ (
);

FILL FILL_5__3596_ (
);

FILL FILL_5__3176_ (
);

FILL FILL_1__3588_ (
);

FILL FILL_1__3168_ (
);

FILL FILL_5__1909_ (
);

FILL FILL_6__2880_ (
);

FILL FILL_6__2460_ (
);

FILL FILL_6__2040_ (
);

FILL FILL_2__2872_ (
);

FILL FILL_2__2452_ (
);

FILL FILL_2__2032_ (
);

FILL FILL_4__2798_ (
);

FILL FILL_4__2378_ (
);

OAI21X1 _1912_ (
    .A(_914__bF$buf0),
    .B(_949_),
    .C(_1028_),
    .Y(_1029_)
);

FILL FILL_0__2698_ (
);

FILL FILL_6__3665_ (
);

FILL FILL_0__2278_ (
);

FILL FILL_6__3245_ (
);

FILL FILL_2__3657_ (
);

FILL FILL_2__3237_ (
);

FILL FILL_7__2201_ (
);

FILL FILL_3__2941_ (
);

FILL FILL_3__2521_ (
);

FILL FILL_3__2101_ (
);

FILL FILL_5__2867_ (
);

FILL FILL_5__2447_ (
);

FILL FILL_5__2027_ (
);

FILL FILL_1__2859_ (
);

FILL FILL_1__2439_ (
);

FILL FILL_1__2019_ (
);

FILL FILL_3__3306_ (
);

NAND2X1 _2870_ (
    .A(cond_code[1]),
    .B(_886__bF$buf5),
    .Y(_527_)
);

OAI21X1 _2450_ (
    .A(_143_),
    .B(_1060_),
    .C(_152_),
    .Y(_1742_[0])
);

AOI22X1 _2030_ (
    .A(_1049_),
    .B(\AXYS[3] [7]),
    .C(\AXYS[2] [7]),
    .D(_1057_),
    .Y(_1140_)
);

FILL FILL_0__1969_ (
);

FILL FILL_6__2936_ (
);

OAI21X1 _3655_ (
    .A(_1714__bF$buf3),
    .B(_1626_),
    .C(_1683_),
    .Y(_1516_)
);

FILL FILL_6__2516_ (
);

OAI21X1 _3235_ (
    .A(_720__bF$buf3),
    .B(_808_),
    .C(\AXYS[3] [5]),
    .Y(_814_)
);

FILL FILL_1__2192_ (
);

FILL FILL_2__2928_ (
);

FILL FILL_0__2910_ (
);

FILL FILL_2__2508_ (
);

FILL FILL_2__2681_ (
);

FILL FILL_2__2261_ (
);

FILL FILL_4__2187_ (
);

FILL FILL_6__3474_ (
);

FILL FILL_0__2087_ (
);

FILL FILL_6__3054_ (
);

FILL FILL167850x64950 (
);

FILL FILL_2__3466_ (
);

FILL FILL_2__3046_ (
);

FILL FILL_5__1891_ (
);

OAI21X1 _2926_ (
    .A(_1395_),
    .B(_569_),
    .C(_1185_),
    .Y(_570_)
);

NOR2X1 _2506_ (
    .A(_1201_),
    .B(_943_),
    .Y(_201_)
);

FILL FILL_1__1883_ (
);

FILL FILL_7__2430_ (
);

FILL FILL_3__2750_ (
);

FILL FILL_3__2330_ (
);

FILL FILL_5__2676_ (
);

FILL FILL_5__2256_ (
);

FILL FILL_1__2668_ (
);

FILL FILL_7__3635_ (
);

FILL FILL_1__2248_ (
);

FILL FILL_7__3215_ (
);

FILL FILL_3__3535_ (
);

FILL FILL_3__3115_ (
);

FILL FILL_6__1960_ (
);

FILL FILL_2__1952_ (
);

FILL FILL_4__1878_ (
);

FILL FILL_0__1778_ (
);

FILL FILL_6__2745_ (
);

NOR2X1 _3464_ (
    .A(_1708_),
    .B(_1710_),
    .Y(_1712_)
);

FILL FILL_6__2325_ (
);

OAI21X1 _3044_ (
    .A(_656_),
    .B(_917_),
    .C(_658_),
    .Y(_659_)
);

FILL FILL_2__2737_ (
);

FILL FILL_2__2317_ (
);

FILL FILL_4__3604_ (
);

FILL FILL_0__3504_ (
);

FILL FILL_5__1947_ (
);

FILL FILL_1__1939_ (
);

FILL FILL_7__2906_ (
);

FILL FILL_2__2490_ (
);

FILL FILL_2__2070_ (
);

FILL FILL_3__2806_ (
);

OAI21X1 _1950_ (
    .A(_903__bF$buf2),
    .B(_969_),
    .C(_935_),
    .Y(_1067_)
);

FILL FILL_6__3283_ (
);

FILL FILL_2__3695_ (
);

FILL FILL_2__3275_ (
);

OAI22X1 _2735_ (
    .A(RDY_bF$buf0),
    .B(_1016_),
    .C(_400_),
    .D(_402_),
    .Y(_9_)
);

NAND3X1 _2315_ (
    .A(_1408_),
    .B(_1415_),
    .C(_1421_),
    .Y(_1422_)
);

FILL FILL_5__2485_ (
);

FILL FILL_5__2065_ (
);

FILL FILL_1__2897_ (
);

FILL FILL_1__2477_ (
);

FILL FILL_1__2057_ (
);

FILL FILL_7__3024_ (
);

FILL FILL_2__1761_ (
);

FILL FILL_6__2974_ (
);

BUFX2 _3693_ (
    .A(_1741_[10]),
    .Y(AB[10])
);

FILL FILL_6__2554_ (
);

NAND3X1 _3273_ (
    .A(_848_),
    .B(_839_),
    .C(_847_),
    .Y(_849_)
);

FILL FILL_6__2134_ (
);

FILL FILL_2__2966_ (
);

FILL FILL_2__2546_ (
);

FILL FILL_2__2126_ (
);

FILL FILL_7__1930_ (
);

FILL FILL_3__1830_ (
);

FILL FILL_0__3313_ (
);

FILL FILL_5__1756_ (
);

FILL FILL_1__1748_ (
);

FILL FILL_3__2615_ (
);

FILL FILL_6__3092_ (
);

FILL FILL_2__3084_ (
);

FILL FILL_6__1825_ (
);

OAI21X1 _2964_ (
    .A(_1149__bF$buf4),
    .B(_597_),
    .C(_598_),
    .Y(_42_)
);

INVX1 _2544_ (
    .A(_236_),
    .Y(_1741_[2])
);

NOR2X1 _2124_ (
    .A(_902__bF$buf3),
    .B(_989_),
    .Y(_1233_)
);

FILL FILL_2__1817_ (
);

FILL FILL_5__2294_ (
);

DFFSR _3329_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(_7_),
    .CLK(clk_bF$buf5),
    .Q(PC[5])
);

FILL FILL_1__2286_ (
);

FILL FILL_7__3253_ (
);

FILL FILL_7_BUFX2_insert71 (
);

FILL FILL_7_BUFX2_insert72 (
);

FILL FILL_3__3573_ (
);

FILL FILL_3__3153_ (
);

FILL FILL_7_BUFX2_insert74 (
);

FILL FILL_7_BUFX2_insert75 (
);

FILL FILL_7_BUFX2_insert77 (
);

FILL FILL_5__3499_ (
);

FILL FILL_5__3079_ (
);

FILL FILL_7_BUFX2_insert79 (
);

FILL FILL_2__1990_ (
);

FILL FILL_6__2783_ (
);

FILL FILL_6__2363_ (
);

AOI21X1 _3082_ (
    .A(DIMUX[7]),
    .B(_1027__bF$buf3),
    .C(_693_),
    .Y(_694_)
);

FILL FILL_2__2775_ (
);

FILL FILL_2__2355_ (
);

NOR2X1 _1815_ (
    .A(_924_),
    .B(_898_),
    .Y(_941_)
);

FILL FILL_4__3642_ (
);

FILL FILL_4__3222_ (
);

FILL FILL_6__3568_ (
);

FILL FILL_6__3148_ (
);

FILL FILL_0__3542_ (
);

FILL FILL_0__3122_ (
);

FILL FILL_5__1985_ (
);

FILL FILL_1__1977_ (
);

FILL FILL_7__2524_ (
);

FILL FILL_3__2844_ (
);

FILL FILL_3__2424_ (
);

FILL FILL_3__2004_ (
);

FILL FILL_5__3711_ (
);

FILL FILL_7__3309_ (
);

FILL FILL_1__3703_ (
);

FILL FILL_3__3629_ (
);

FILL FILL_3__3209_ (
);

MUX2X1 _2773_ (
    .A(_437_),
    .B(_280_),
    .S(_352_),
    .Y(_438_)
);

NAND2X1 _2353_ (
    .A(_1420_),
    .B(_1419_),
    .Y(_1459_)
);

FILL FILL_4__2913_ (
);

FILL FILL_6__2839_ (
);

NAND2X1 _3558_ (
    .A(BI[0]),
    .B(_1573_),
    .Y(_1588_)
);

FILL FILL_6__2419_ (
);

AOI21X1 _3138_ (
    .A(DIMUX[2]),
    .B(_1319__bF$buf3),
    .C(_743_),
    .Y(_744_)
);

FILL FILL_7__3482_ (
);

FILL FILL_1__2095_ (
);

FILL FILL_7__3062_ (
);

FILL FILL_0__2813_ (
);

FILL FILL169350x32550 (
);

FILL FILL_6__2592_ (
);

FILL FILL_6__2172_ (
);

FILL FILL_2__2584_ (
);

FILL FILL_2__2164_ (
);

FILL FILL_4__3451_ (
);

FILL FILL_4__3031_ (
);

FILL FILL_5__1794_ (
);

OAI21X1 _2829_ (
    .A(_296_),
    .B(_378_),
    .C(_490_),
    .Y(_491_)
);

AND2X2 _2409_ (
    .A(_117_),
    .B(_1254_),
    .Y(_118_)
);

FILL FILL_1__1786_ (
);

FILL FILL_7__2753_ (
);

FILL FILL_7__2333_ (
);

FILL FILL_3__2653_ (
);

FILL FILL_3__2233_ (
);

FILL FILL_5__2999_ (
);

FILL FILL_5__2579_ (
);

FILL FILL_5__2159_ (
);

FILL FILL_5__3520_ (
);

FILL FILL_7__3538_ (
);

FILL FILL_5__3100_ (
);

FILL FILL_1__3512_ (
);

FILL FILL_3__3018_ (
);

FILL FILL_6__1863_ (
);

INVX1 _2582_ (
    .A(ABH[0]),
    .Y(_269_)
);

OAI21X1 _2162_ (
    .A(_931__bF$buf4),
    .B(_974_),
    .C(_886__bF$buf2),
    .Y(_1271_)
);

FILL FILL_2__1855_ (
);

FILL FILL_4__2722_ (
);

FILL FILL_4__2302_ (
);

FILL FILL_6__2648_ (
);

FILL FILL_6__2228_ (
);

DFFSR _3367_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_44_),
    .CLK(clk_bF$buf6),
    .Q(write_back)
);

FILL FILL_7__3291_ (
);

FILL FILL_0__2622_ (
);

FILL FILL_0__2202_ (
);

FILL FILL_3__3191_ (
);

FILL FILL_4__3507_ (
);

FILL FILL_3__1924_ (
);

FILL FILL_7__2809_ (
);

FILL FILL_2__2393_ (
);

FILL FILL_3__2709_ (
);

NAND2X1 _1853_ (
    .A(_903__bF$buf1),
    .B(_977_),
    .Y(_978_)
);

FILL FILL_4__3260_ (
);

FILL FILL_6__3186_ (
);

FILL FILL_2__3598_ (
);

FILL FILL_0__3580_ (
);

FILL FILL_0__3160_ (
);

FILL FILL_2__3178_ (
);

FILL FILL_6__1919_ (
);

INVX1 _2638_ (
    .A(_312_),
    .Y(_313_)
);

NOR2X1 _2218_ (
    .A(_1213_),
    .B(_1215_),
    .Y(_1326_)
);

FILL FILL_7__2982_ (
);

FILL FILL_7__2562_ (
);

FILL FILL_7__2142_ (
);

FILL FILL_3__2882_ (
);

FILL FILL_3__2462_ (
);

FILL FILL_3__2042_ (
);

FILL FILL_5__2388_ (
);

FILL FILL_3__3667_ (
);

FILL FILL_3__3247_ (
);

NOR2X1 _2391_ (
    .A(_1239_),
    .B(_1434_),
    .Y(_1496_)
);

FILL FILL_4__2951_ (
);

FILL FILL_4__2531_ (
);

FILL FILL_4__2111_ (
);

FILL FILL_6__2877_ (
);

AOI22X1 _3596_ (
    .A(_1550_),
    .B(_1625_),
    .C(_1607_),
    .D(_1624_),
    .Y(_1626_)
);

FILL FILL_6__2457_ (
);

FILL FILL_6__2037_ (
);

INVX1 _3176_ (
    .A(_777_),
    .Y(_778_)
);

FILL FILL_0__2851_ (
);

FILL FILL_2__2869_ (
);

FILL FILL_2__2449_ (
);

FILL FILL_0__2431_ (
);

FILL FILL_0__2011_ (
);

FILL FILL_2__2029_ (
);

NOR2X1 _1909_ (
    .A(_1023_),
    .B(_1025_),
    .Y(_1026_)
);

FILL FILL_4__3316_ (
);

FILL FILL_0__3636_ (
);

FILL FILL_0__3216_ (
);

FILL FILL_5__2600_ (
);

FILL FILL_3__2938_ (
);

FILL FILL_3__2518_ (
);

FILL FILL_4__1802_ (
);

OAI21X1 _2867_ (
    .A(_1153_),
    .B(_1021_),
    .C(_525_),
    .Y(_18_)
);

AOI22X1 _2447_ (
    .A(PC[0]),
    .B(_1080_),
    .C(_149_),
    .D(C),
    .Y(_150_)
);

AOI21X1 _2027_ (
    .A(_1082_),
    .B(ADD[6]),
    .C(_1137_),
    .Y(_1138_)
);

FILL FILL_7__2791_ (
);

FILL FILL_7__2371_ (
);

FILL FILL167250x144150 (
);

FILL FILL_3__2691_ (
);

FILL FILL_3__2271_ (
);

FILL FILL_5__2197_ (
);

FILL FILL_1__2189_ (
);

FILL FILL_7__3156_ (
);

FILL FILL_0__2907_ (
);

FILL FILL_1__3550_ (
);

FILL FILL_1__3130_ (
);

FILL FILL_3__3476_ (
);

FILL FILL_3__3056_ (
);

FILL FILL169650x75750 (
);

FILL FILL_2__1893_ (
);

FILL FILL_4__2760_ (
);

FILL FILL_4__2340_ (
);

FILL FILL_6__2686_ (
);

FILL FILL_6__2266_ (
);

FILL FILL_2__2678_ (
);

FILL FILL_0__2660_ (
);

FILL FILL_2__2258_ (
);

FILL FILL_0__2240_ (
);

FILL FILL_4__3545_ (
);

FILL FILL_4__3125_ (
);

FILL FILL_3__1962_ (
);

FILL FILL_0__3025_ (
);

FILL FILL_5__1888_ (
);

FILL FILL_7__2427_ (
);

FILL FILL_1__2821_ (
);

FILL FILL_1__2401_ (
);

FILL FILL_3__2747_ (
);

FILL FILL_3__2327_ (
);

OAI22X1 _1891_ (
    .A(_1011_),
    .B(_968_),
    .C(_888_),
    .D(_1004_),
    .Y(BI[4])
);

FILL FILL_5__3614_ (
);

FILL FILL_1__3606_ (
);

FILL FILL168450x57750 (
);

FILL FILL_6__1957_ (
);

INVX1 _2676_ (
    .A(_347_),
    .Y(_349_)
);

NOR2X1 _2256_ (
    .A(_1363_),
    .B(_1358_),
    .Y(_1364_)
);

FILL FILL_7__2180_ (
);

FILL FILL_2__1949_ (
);

FILL FILL_0__1931_ (
);

FILL FILL_3__2080_ (
);

FILL FILL_4__2816_ (
);

FILL FILL_0__2716_ (
);

FILL FILL_3__3285_ (
);

FILL FILL_6__2495_ (
);

FILL FILL_6__2075_ (
);

FILL FILL_2__2487_ (
);

FILL FILL_2__2067_ (
);

NOR2X1 _1947_ (
    .A(_990_),
    .B(_1063_),
    .Y(_1064_)
);

FILL FILL_7__1871_ (
);

FILL FILL169350x133350 (
);

FILL FILL_0__3674_ (
);

FILL FILL_3__1771_ (
);

FILL FILL_0__3254_ (
);

FILL FILL_7__2656_ (
);

FILL FILL_1__2630_ (
);

FILL FILL_1__2210_ (
);

FILL FILL_3__2976_ (
);

FILL FILL_3__2556_ (
);

FILL FILL_3__2136_ (
);

FILL FILL169950x126150 (
);

FILL FILL_5__3003_ (
);

FILL FILL_4__1840_ (
);

FILL FILL_6__1766_ (
);

OAI21X1 _2485_ (
    .A(_143_),
    .B(_1125_),
    .C(_182_),
    .Y(_1742_[5])
);

INVX1 _2065_ (
    .A(_1173_),
    .Y(_1174_)
);

FILL FILL_2__1758_ (
);

FILL FILL_4__2625_ (
);

FILL FILL_4__2205_ (
);

FILL FILL_7__3194_ (
);

FILL FILL_0__2945_ (
);

FILL FILL_0__2525_ (
);

FILL FILL_0__2105_ (
);

FILL FILL_3__3094_ (
);

FILL FILL_7__1927_ (
);

FILL FILL_1__1901_ (
);

FILL FILL_3__1827_ (
);

FILL FILL_2__2296_ (
);

INVX8 _1756_ (
    .A(RDY_bF$buf5),
    .Y(_886_)
);

FILL FILL_4__3583_ (
);

FILL FILL_4__3163_ (
);

FILL FILL_6__3089_ (
);

FILL FILL_0__3483_ (
);

FILL FILL_0__3063_ (
);

FILL FILL_7__2885_ (
);

FILL FILL_7__2045_ (
);

FILL FILL_3__2785_ (
);

FILL FILL_3__2365_ (
);

FILL FILL_5__3652_ (
);

FILL FILL_5__3232_ (
);

FILL FILL_1__3644_ (
);

FILL FILL_1__3224_ (
);

FILL FILL_6__1995_ (
);

NAND2X1 _2294_ (
    .A(_1400_),
    .B(_1398_),
    .Y(_1401_)
);

FILL FILL_2__1987_ (
);

FILL FILL_4__2854_ (
);

FILL FILL_4__2434_ (
);

FILL FILL_4__2014_ (
);

AND2X2 _3499_ (
    .A(_1718_),
    .B(BI[4]),
    .Y(_1529_)
);

AOI21X1 _3079_ (
    .A(_662_),
    .B(_1227_),
    .C(AN),
    .Y(_691_)
);

FILL FILL_0__2754_ (
);

FILL FILL_0__2334_ (
);

FILL FILL_6__3301_ (
);

FILL FILL_2__3713_ (
);

FILL FILL_4__3639_ (
);

FILL FILL_4__3219_ (
);

FILL FILL_0__3539_ (
);

FILL FILL_0__3119_ (
);

FILL FILL_5__2923_ (
);

FILL FILL_5__2503_ (
);

FILL FILL_1__2915_ (
);

NAND3X1 _1985_ (
    .A(_1099_),
    .B(_1097_),
    .C(_1098_),
    .Y(_1100_)
);

FILL FILL_5__3708_ (
);

FILL FILL_0__3292_ (
);

FILL FILL_7__2274_ (
);

BUFX2 _3711_ (
    .A(_1742_[4]),
    .Y(DO[4])
);

FILL FILL_3__2594_ (
);

FILL FILL_3__2174_ (
);

FILL FILL_7__3479_ (
);

FILL FILL_5__3461_ (
);

FILL FILL_7__3059_ (
);

FILL FILL_5__3041_ (
);

FILL FILL_1__3453_ (
);

FILL FILL_1__3033_ (
);

FILL FILL_2__1796_ (
);

FILL FILL_4__2663_ (
);

FILL FILL_4__2243_ (
);

FILL FILL_6__2589_ (
);

FILL FILL_6__2169_ (
);

FILL FILL_0__2983_ (
);

FILL FILL_0__2563_ (
);

FILL FILL_6__3530_ (
);

FILL FILL_0__2143_ (
);

FILL FILL_6__3110_ (
);

FILL FILL_2__3522_ (
);

FILL FILL_2__3102_ (
);

FILL FILL_4__3028_ (
);

FILL FILL_3__1865_ (
);

FILL FILL_5__2732_ (
);

FILL FILL_5__2312_ (
);

FILL FILL_2_BUFX2_insert20 (
);

FILL FILL_2_BUFX2_insert21 (
);

FILL FILL_2_BUFX2_insert22 (
);

FILL FILL_2_BUFX2_insert23 (
);

FILL FILL_2_BUFX2_insert24 (
);

FILL FILL_2_BUFX2_insert25 (
);

FILL FILL_1__2724_ (
);

FILL FILL_1__2304_ (
);

INVX1 _1794_ (
    .A(rotate),
    .Y(_920_)
);

FILL FILL_5__3517_ (
);

FILL FILL_1__3509_ (
);

FILL FILL_4__1934_ (
);

OAI21X1 _2999_ (
    .A(_612_),
    .B(_578_),
    .C(_1252_),
    .Y(_627_)
);

AOI21X1 _2579_ (
    .A(_1142_),
    .B(_195_),
    .C(_266_),
    .Y(_267_)
);

INVX1 _2159_ (
    .A(_1032_),
    .Y(_1268_)
);

FILL FILL_0__1834_ (
);

FILL FILL_6__2801_ (
);

OR2X2 _3520_ (
    .A(_1545_),
    .B(_1549_),
    .Y(_1550_)
);

NAND2X1 _3100_ (
    .A(C),
    .B(_709_),
    .Y(_710_)
);

FILL FILL_4__2719_ (
);

FILL FILL_7__3288_ (
);

FILL FILL_5__3270_ (
);

FILL FILL_0__2619_ (
);

FILL FILL_1__3262_ (
);

FILL FILL_3__3188_ (
);

FILL FILL_4__2892_ (
);

FILL FILL_4__2472_ (
);

FILL FILL_4__2052_ (
);

FILL FILL_6__2398_ (
);

FILL FILL_0__2792_ (
);

FILL FILL_0__2372_ (
);

FILL FILL_4__3677_ (
);

FILL FILL_7__1774_ (
);

FILL FILL_4__3257_ (
);

FILL FILL_0__3577_ (
);

FILL FILL_0__3157_ (
);

FILL FILL_5__2961_ (
);

FILL FILL_5__2541_ (
);

FILL FILL_7__2559_ (
);

FILL FILL_5__2121_ (
);

FILL FILL_1__2953_ (
);

FILL FILL_1__2533_ (
);

FILL FILL_7__3500_ (
);

FILL FILL_1__2113_ (
);

FILL FILL_3__2879_ (
);

FILL FILL_3__2459_ (
);

FILL FILL_3__2039_ (
);

OAI21X1 _2388_ (
    .A(_1462_),
    .B(_1484_),
    .C(_1493_),
    .Y(_1512_[3])
);

FILL FILL_6__2610_ (
);

FILL FILL_2__2602_ (
);

FILL FILL_4__2948_ (
);

FILL FILL_4__2528_ (
);

FILL FILL_4__2108_ (
);

FILL FILL_0__2848_ (
);

FILL FILL_0__2428_ (
);

FILL FILL_0__2008_ (
);

FILL FILL_1__3491_ (
);

FILL FILL_1__3071_ (
);

FILL FILL_5__1812_ (
);

FILL FILL_1__1804_ (
);

FILL FILL_4__2281_ (
);

FILL FILL_0__2181_ (
);

FILL FILL_2__2199_ (
);

FILL FILL_2__3560_ (
);

FILL FILL_2__3140_ (
);

FILL FILL_4__3486_ (
);

FILL FILL_4__3066_ (
);

OAI21X1 _2600_ (
    .A(_280_),
    .B(_218_),
    .C(_284_),
    .Y(_1741_[10])
);

FILL FILL_7__2788_ (
);

FILL FILL_5__2770_ (
);

FILL FILL_5__2350_ (
);

FILL FILL_1__2762_ (
);

FILL FILL_1__2342_ (
);

FILL FILL_3__2688_ (
);

FILL FILL_3__2268_ (
);

FILL FILL_5__3555_ (
);

FILL FILL_5__3135_ (
);

FILL FILL_1__3547_ (
);

FILL FILL_1__3127_ (
);

FILL FILL_4__1972_ (
);

FILL FILL_6__1898_ (
);

OAI21X1 _2197_ (
    .A(_886__bF$buf2),
    .B(_1304_),
    .C(_1305_),
    .Y(_1306_)
);

FILL FILL_0__1872_ (
);

FILL FILL_2__2831_ (
);

FILL FILL_2__2411_ (
);

FILL FILL_4__2757_ (
);

FILL FILL_4__2337_ (
);

FILL FILL_0__2657_ (
);

FILL FILL_6__3624_ (
);

FILL FILL_0__2237_ (
);

FILL FILL_6__3204_ (
);

FILL FILL_2__3616_ (
);

FILL FILL_3__1959_ (
);

FILL FILL_4__2090_ (
);

FILL FILL_3__2900_ (
);

FILL FILL_5__2826_ (
);

FILL FILL_5__2406_ (
);

FILL FILL_1__2818_ (
);

INVX2 _1888_ (
    .A(DIMUX[3]),
    .Y(_1010_)
);

FILL FILL_4__3295_ (
);

FILL FILL_0__3195_ (
);

FILL FILL_7__2177_ (
);

FILL FILL_0__1928_ (
);

OAI21X1 _3614_ (
    .A(AI[6]),
    .B(_1641_),
    .C(_1722_),
    .Y(_1644_)
);

FILL FILL_1__2991_ (
);

FILL FILL_1__2571_ (
);

FILL FILL_1__2151_ (
);

FILL FILL_3__2497_ (
);

FILL FILL_3__2077_ (
);

FILL FILL_4__1781_ (
);

FILL FILL_2__2640_ (
);

FILL FILL_2__2220_ (
);

FILL FILL_4__2986_ (
);

FILL FILL_4__2566_ (
);

FILL FILL_4__2146_ (
);

FILL FILL_0__2886_ (
);

FILL FILL_0__2466_ (
);

FILL FILL_0__2046_ (
);

FILL FILL_6__3013_ (
);

FILL FILL_2__3005_ (
);

FILL FILL_5__1850_ (
);

FILL FILL_1__1842_ (
);

FILL FILL_3__1768_ (
);

FILL FILL_5__2635_ (
);

FILL FILL_5__2215_ (
);

FILL FILL_1__2627_ (
);

FILL FILL_1__2207_ (
);

FILL FILL_2__1911_ (
);

FILL FILL_4__1837_ (
);

FILL FILL_6__2704_ (
);

DFFSR _3423_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_92_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[2] [7])
);

OAI21X1 _3003_ (
    .A(_626_),
    .B(_629_),
    .C(_1150__bF$buf4),
    .Y(_630_)
);

FILL FILL_1__2380_ (
);

FILL FILL_5__3593_ (
);

FILL FILL_5__3173_ (
);

FILL FILL_1__3585_ (
);

FILL FILL_1__3165_ (
);

FILL FILL_5__1906_ (
);

FILL FILL_4__2795_ (
);

FILL FILL_4__2375_ (
);

FILL FILL_0__2695_ (
);

FILL FILL_6__3662_ (
);

FILL FILL_0__2275_ (
);

FILL FILL_6__3242_ (
);

FILL FILL_2__3654_ (
);

FILL FILL_2__3234_ (
);

FILL FILL_3__1997_ (
);

FILL FILL_5__2864_ (
);

FILL FILL_5__2444_ (
);

FILL FILL_5__2024_ (
);

FILL FILL_1__2856_ (
);

FILL FILL_1__2436_ (
);

FILL FILL_1__2016_ (
);

FILL FILL_3__3303_ (
);

FILL FILL_5__3649_ (
);

FILL FILL_5__3229_ (
);

FILL FILL_0__1966_ (
);

FILL FILL_6__2933_ (
);

AOI22X1 _3652_ (
    .A(_1658_),
    .B(_1659_),
    .C(_1675_),
    .D(_1681_),
    .Y(_1682_)
);

FILL FILL_6__2513_ (
);

OAI21X1 _3232_ (
    .A(_754_),
    .B(_807_),
    .C(_812_),
    .Y(_96_)
);

FILL FILL_2__2925_ (
);

FILL FILL_2__2505_ (
);

FILL FILL_4__2184_ (
);

FILL FILL_6__3471_ (
);

FILL FILL_0__2084_ (
);

FILL FILL_6__3051_ (
);

FILL FILL_2__3463_ (
);

FILL FILL_2__3043_ (
);

AOI22X1 _2923_ (
    .A(_128_),
    .B(_1149__bF$buf2),
    .C(_567_),
    .D(_563_),
    .Y(_32_)
);

NAND3X1 _2503_ (
    .A(_1202_),
    .B(_197_),
    .C(_1224_),
    .Y(_198_)
);

FILL FILL_1__1880_ (
);

FILL FILL_0__3289_ (
);

FILL FILL_5__2673_ (
);

FILL FILL_5__2253_ (
);

BUFX2 _3708_ (
    .A(_1742_[1]),
    .Y(DO[1])
);

FILL FILL_1__2665_ (
);

FILL FILL_7__3632_ (
);

FILL FILL_1__2245_ (
);

FILL FILL_7__3212_ (
);

FILL FILL_3__3532_ (
);

FILL FILL_3__3112_ (
);

FILL FILL_5__3458_ (
);

FILL FILL_5__3038_ (
);

FILL FILL_4__1875_ (
);

FILL FILL_0__1775_ (
);

FILL FILL_6__2742_ (
);

NAND2X1 _3461_ (
    .A(\u_ALU8.BI7 ),
    .B(_1707_),
    .Y(_1709_)
);

FILL FILL_6__2322_ (
);

INVX1 _3041_ (
    .A(bit_ins),
    .Y(_656_)
);

FILL FILL_2__2734_ (
);

FILL FILL_2__2314_ (
);

FILL FILL_4__3601_ (
);

FILL FILL_6__3527_ (
);

FILL FILL_6__3107_ (
);

FILL FILL_2__3519_ (
);

FILL FILL_0__3501_ (
);

FILL FILL_5__1944_ (
);

FILL FILL_1__1936_ (
);

FILL FILL_7__2903_ (
);

FILL FILL_3__2803_ (
);

FILL FILL_5__2729_ (
);

FILL FILL_5__2309_ (
);

FILL FILL_6__3280_ (
);

FILL FILL_2__3692_ (
);

FILL FILL_2__3272_ (
);

FILL FILL_4__3198_ (
);

AOI21X1 _2732_ (
    .A(_386_),
    .B(_392_),
    .C(_399_),
    .Y(_400_)
);

AND2X2 _2312_ (
    .A(_1416_),
    .B(_1418_),
    .Y(_1419_)
);

FILL FILL_0__3098_ (
);

FILL FILL_5__2482_ (
);

FILL FILL_5__2062_ (
);

OAI21X1 _3517_ (
    .A(alu_op[3]),
    .B(BI[3]),
    .C(_1740_),
    .Y(_1547_)
);

FILL FILL_1__2894_ (
);

FILL FILL_1__2474_ (
);

FILL FILL_1__2054_ (
);

FILL FILL_5__3267_ (
);

FILL FILL_1__3259_ (
);

FILL FILL_6__2971_ (
);

DFFSR _3690_ (
    .R(_1513_),
    .S(vdd),
    .D(_1525_),
    .CLK(clk_bF$buf3),
    .Q(\u_ALU8.AI7 )
);

FILL FILL_6__2551_ (
);

NAND3X1 _3270_ (
    .A(_840_),
    .B(_844_),
    .C(_845_),
    .Y(_846_)
);

FILL FILL_6__2131_ (
);

FILL FILL_2__2963_ (
);

FILL FILL_2__2543_ (
);

FILL FILL_2__2123_ (
);

FILL FILL_4__2889_ (
);

FILL FILL_4__2469_ (
);

FILL FILL_4__2049_ (
);

FILL FILL_0__2789_ (
);

FILL FILL_0__2369_ (
);

FILL FILL_0__3310_ (
);

FILL FILL_5__1753_ (
);

FILL FILL_1__1745_ (
);

FILL FILL_7__2712_ (
);

FILL FILL_3__2612_ (
);

FILL FILL_5__2958_ (
);

FILL FILL_5__2538_ (
);

FILL FILL_5__2118_ (
);

FILL FILL_2__3081_ (
);

FILL FILL_6__1822_ (
);

INVX1 _2961_ (
    .A(_576_),
    .Y(_596_)
);

AND2X2 _2541_ (
    .A(_232_),
    .B(_233_),
    .Y(_234_)
);

INVX1 _2121_ (
    .A(_1229_),
    .Y(_1230_)
);

FILL FILL_2__1814_ (
);

FILL FILL_5__2291_ (
);

FILL FILL_6__2607_ (
);

DFFSR _3326_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(_4_),
    .CLK(clk_bF$buf3),
    .Q(PC[2])
);

FILL FILL_1__2283_ (
);

FILL FILL_7_BUFX2_insert40 (
);

FILL FILL_7_BUFX2_insert42 (
);

FILL FILL_3__3570_ (
);

FILL FILL_7_BUFX2_insert43 (
);

FILL FILL_3__3150_ (
);

FILL FILL_7_BUFX2_insert45 (
);

FILL FILL_7_BUFX2_insert46 (
);

FILL FILL_5__3496_ (
);

FILL FILL_7_BUFX2_insert48 (
);

FILL FILL_5__3076_ (
);

FILL FILL_1__3488_ (
);

FILL FILL_1__3068_ (
);

FILL FILL_5__1809_ (
);

FILL FILL_6__2780_ (
);

FILL FILL_6__2360_ (
);

FILL FILL_2__2772_ (
);

FILL FILL_2__2352_ (
);

FILL FILL_4__2698_ (
);

FILL FILL_4__2278_ (
);

NAND2X1 _1812_ (
    .A(_937_),
    .B(_910_),
    .Y(_938_)
);

FILL FILL_0__2598_ (
);

FILL FILL_6__3565_ (
);

FILL FILL_0__2178_ (
);

FILL FILL_6__3145_ (
);

FILL FILL_2__3557_ (
);

FILL FILL_2__3137_ (
);

FILL FILL_5__1982_ (
);

FILL FILL_1__1974_ (
);

FILL FILL_7__2941_ (
);

FILL FILL_7__2521_ (
);

FILL FILL_7__2101_ (
);

FILL FILL_3__2841_ (
);

FILL FILL_3__2421_ (
);

FILL FILL_3__2001_ (
);

FILL FILL_5__2767_ (
);

FILL FILL_5__2347_ (
);

FILL FILL_1__2759_ (
);

FILL FILL_1__2339_ (
);

FILL FILL_7__3306_ (
);

FILL FILL_1__3700_ (
);

FILL FILL_3__3626_ (
);

FILL FILL_3__3206_ (
);

AOI22X1 _2770_ (
    .A(_925_),
    .B(ABH[2]),
    .C(PC[10]),
    .D(_312_),
    .Y(_435_)
);

NAND3X1 _2350_ (
    .A(_1451_),
    .B(_1443_),
    .C(_1456_),
    .Y(_1512_[2])
);

FILL FILL_4__1969_ (
);

FILL FILL_4__2910_ (
);

FILL FILL_0__1869_ (
);

FILL FILL_6__2836_ (
);

OAI21X1 _3555_ (
    .A(_1725_),
    .B(_1740_),
    .C(CI),
    .Y(_1585_)
);

FILL FILL_6__2416_ (
);

OR2X2 _3135_ (
    .A(_740_),
    .B(_739_),
    .Y(_741_)
);

FILL FILL_1__2092_ (
);

FILL FILL_0__2810_ (
);

FILL FILL_2__2828_ (
);

FILL FILL_2__2408_ (
);

FILL FILL_1__3297_ (
);

FILL FILL_2__2581_ (
);

FILL FILL_2__2161_ (
);

FILL FILL_4__2087_ (
);

FILL FILL_5__1791_ (
);

INVX1 _2826_ (
    .A(_465_),
    .Y(_488_)
);

AND2X2 _2406_ (
    .A(_1509_),
    .B(_1436_),
    .Y(_1510_)
);

FILL FILL_1__1783_ (
);

FILL FILL_7__2330_ (
);

FILL FILL_3__2650_ (
);

FILL FILL_3__2230_ (
);

FILL FILL_5__2996_ (
);

FILL FILL_5__2576_ (
);

FILL FILL_5__2156_ (
);

FILL FILL_1__2988_ (
);

FILL FILL_1__2568_ (
);

FILL FILL_7__3535_ (
);

FILL FILL_1__2148_ (
);

FILL FILL_7__3115_ (
);

FILL FILL_3__3015_ (
);

FILL FILL168150x133350 (
);

FILL FILL_6__1860_ (
);

FILL FILL_2__1852_ (
);

FILL FILL_4__1778_ (
);

FILL FILL_6__2645_ (
);

DFFSR _3364_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_41_),
    .CLK(clk_bF$buf4),
    .Q(adc_sbc)
);

FILL FILL_6__2225_ (
);

FILL FILL_2__2637_ (
);

FILL FILL_2__2217_ (
);

FILL FILL_4__3504_ (
);

FILL FILL_3__1921_ (
);

FILL FILL_5__1847_ (
);

FILL FILL_1__1839_ (
);

FILL FILL_7__2806_ (
);

FILL FILL_2__2390_ (
);

FILL FILL_3__2706_ (
);

OAI21X1 _1850_ (
    .A(_914__bF$buf2),
    .B(_974_),
    .C(_972_),
    .Y(_975_)
);

FILL FILL_6__3183_ (
);

FILL FILL_2__3595_ (
);

FILL FILL_2__3175_ (
);

FILL FILL_6__1916_ (
);

INVX8 _2635_ (
    .A(reset),
    .Y(_1_)
);

NAND3X1 _2215_ (
    .A(_1323_),
    .B(_1282_),
    .C(_1302_),
    .Y(_1324_)
);

FILL FILL_2__1908_ (
);

FILL FILL_5__2385_ (
);

FILL FILL_1__2797_ (
);

FILL FILL_1__2377_ (
);

FILL FILL_3__3664_ (
);

FILL FILL_3__3244_ (
);

FILL FILL_6__2874_ (
);

NAND2X1 _3593_ (
    .A(_1622_),
    .B(_1618_),
    .Y(_1623_)
);

FILL FILL_6__2454_ (
);

FILL FILL_6__2034_ (
);

NOR2X1 _3173_ (
    .A(_1319__bF$buf1),
    .B(_774_),
    .Y(_775_)
);

FILL FILL_2__2866_ (
);

FILL FILL_2__2446_ (
);

FILL FILL_2__2026_ (
);

NAND3X1 _1906_ (
    .A(_1018_),
    .B(_1019_),
    .C(_1022_),
    .Y(_1023_)
);

FILL FILL_7__1830_ (
);

FILL FILL_4__3313_ (
);

FILL FILL_6__3659_ (
);

FILL FILL_6__3239_ (
);

FILL FILL_0__3633_ (
);

FILL FILL_0__3213_ (
);

FILL FILL_3__2935_ (
);

FILL FILL_3__2515_ (
);

AOI22X1 _2864_ (
    .A(_886__bF$buf3),
    .B(_304_),
    .C(_520_),
    .D(_523_),
    .Y(_17_)
);

INVX1 _2444_ (
    .A(php),
    .Y(_147_)
);

NOR2X1 _2024_ (
    .A(_1134_),
    .B(_1092_),
    .Y(_1135_)
);

FILL FILL_5__2194_ (
);

NAND2X1 _3649_ (
    .A(_1653_),
    .B(_1636_),
    .Y(_1679_)
);

OAI21X1 _3229_ (
    .A(_720__bF$buf0),
    .B(_808_),
    .C(\AXYS[3] [2]),
    .Y(_811_)
);

FILL FILL_1__2186_ (
);

FILL FILL_7__3153_ (
);

FILL FILL_0__2904_ (
);

FILL FILL_3__3473_ (
);

FILL FILL_3__3053_ (
);

FILL FILL_2__1890_ (
);

FILL FILL_6__2683_ (
);

FILL FILL_6__2263_ (
);

FILL FILL_2__2675_ (
);

FILL FILL_2__2255_ (
);

FILL FILL_4__3542_ (
);

FILL FILL_4__3122_ (
);

FILL FILL_6__3468_ (
);

FILL FILL_6__3048_ (
);

FILL FILL_0__3022_ (
);

FILL FILL_5__1885_ (
);

FILL FILL_1__1877_ (
);

FILL FILL_7__2424_ (
);

FILL FILL_3__2744_ (
);

FILL FILL_3__2324_ (
);

FILL FILL_5__3611_ (
);

FILL FILL_7__3629_ (
);

FILL FILL_7__3209_ (
);

FILL FILL_1__3603_ (
);

FILL FILL_3__3529_ (
);

FILL FILL_3__3109_ (
);

FILL FILL_6__1954_ (
);

INVX1 _2673_ (
    .A(_345_),
    .Y(_346_)
);

NAND2X1 _2253_ (
    .A(_886__bF$buf6),
    .B(_1360_),
    .Y(_1361_)
);

FILL FILL_2__1946_ (
);

FILL FILL_4__2813_ (
);

FILL FILL_6__2739_ (
);

NOR2X1 _3458_ (
    .A(_1705_),
    .B(_1704_),
    .Y(_1706_)
);

FILL FILL_6__2319_ (
);

OAI21X1 _3038_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[7]),
    .Y(_655_)
);

FILL FILL_0__2713_ (
);

FILL FILL_3__3282_ (
);

FILL FILL_6__2492_ (
);

FILL FILL_6__2072_ (
);

FILL FILL_2__2484_ (
);

FILL FILL_2__2064_ (
);

AOI21X1 _1944_ (
    .A(_901_),
    .B(_941_),
    .C(_988_),
    .Y(_1061_)
);

FILL FILL_6__3697_ (
);

FILL FILL_6__3277_ (
);

FILL FILL_0__3671_ (
);

FILL FILL_2__3269_ (
);

FILL FILL_0__3251_ (
);

OAI21X1 _2729_ (
    .A(_396_),
    .B(_378_),
    .C(_148_),
    .Y(_397_)
);

NAND2X1 _2309_ (
    .A(_1365_),
    .B(_1350_),
    .Y(_1416_)
);

FILL FILL_7__2653_ (
);

FILL FILL_3__2973_ (
);

FILL FILL_3__2553_ (
);

FILL FILL_3__2133_ (
);

FILL FILL_5__2899_ (
);

FILL FILL_5__2479_ (
);

FILL FILL_5__2059_ (
);

FILL FILL_5__3000_ (
);

FILL FILL_6__1763_ (
);

OAI21X1 _2482_ (
    .A(_1319__bF$buf0),
    .B(_1263_),
    .C(PC[13]),
    .Y(_180_)
);

OAI21X1 _2062_ (
    .A(_1168_),
    .B(_1169_),
    .C(_1170_),
    .Y(_1171_)
);

FILL FILL_2__1755_ (
);

FILL FILL_4__2622_ (
);

FILL FILL_4__2202_ (
);

FILL FILL_6__2968_ (
);

DFFSR _3687_ (
    .R(_1513_),
    .S(vdd),
    .D(_1522_),
    .CLK(clk_bF$buf3),
    .Q(ADD[5])
);

FILL FILL_6__2548_ (
);

NAND2X1 _3267_ (
    .A(_842_),
    .B(_835_),
    .Y(_843_)
);

FILL FILL_6__2128_ (
);

FILL FILL_7__3191_ (
);

FILL FILL_0__2942_ (
);

FILL FILL_0__2522_ (
);

FILL FILL_0__2102_ (
);

FILL FILL_3__3091_ (
);

FILL FILL_7__1924_ (
);

FILL FILL_3__1824_ (
);

FILL FILL_0__3307_ (
);

FILL FILL_7__2709_ (
);

FILL FILL169950x147750 (
);

FILL FILL_2__2293_ (
);

FILL FILL_3__2609_ (
);

INVX1 _1753_ (
    .A(DIHOLD[3]),
    .Y(_884_)
);

FILL FILL_4__3580_ (
);

FILL FILL_4__3160_ (
);

FILL FILL_6__3086_ (
);

FILL FILL_2__3498_ (
);

FILL FILL_0__3480_ (
);

FILL FILL_2__3078_ (
);

FILL FILL_0__3060_ (
);

FILL FILL_6__1819_ (
);

NAND3X1 _2958_ (
    .A(_559_),
    .B(_1405_),
    .C(_593_),
    .Y(_595_)
);

INVX1 _2538_ (
    .A(_231_),
    .Y(_1741_[1])
);

NAND2X1 _2118_ (
    .A(_903__bF$buf1),
    .B(_971_),
    .Y(_1227_)
);

FILL FILL_7__2882_ (
);

FILL FILL_7__2462_ (
);

FILL FILL_7__2042_ (
);

FILL FILL_3__2782_ (
);

FILL FILL_3__2362_ (
);

FILL FILL_5__2288_ (
);

FILL FILL_7__3667_ (
);

FILL FILL_1__3641_ (
);

FILL FILL_1__3221_ (
);

FILL FILL_3__3567_ (
);

FILL FILL_3__3147_ (
);

FILL FILL_6__1992_ (
);

AOI21X1 _2291_ (
    .A(_1394_),
    .B(_1251_),
    .C(_1397_),
    .Y(_1398_)
);

FILL FILL_2__1984_ (
);

FILL FILL_4__2851_ (
);

FILL FILL167550x144150 (
);

FILL FILL_4__2431_ (
);

FILL FILL_4__2011_ (
);

FILL FILL_6__2777_ (
);

OAI21X1 _3496_ (
    .A(alu_op[3]),
    .B(BI[5]),
    .C(_1740_),
    .Y(_1526_)
);

FILL FILL_6__2357_ (
);

NAND2X1 _3076_ (
    .A(_921_),
    .B(_661_),
    .Y(_688_)
);

FILL FILL_0__2751_ (
);

FILL FILL_2__2769_ (
);

FILL FILL_0__2331_ (
);

FILL FILL_2__2349_ (
);

FILL FILL_2__3710_ (
);

NOR2X1 _1809_ (
    .A(_924_),
    .B(_934_),
    .Y(_935_)
);

FILL FILL_4__3636_ (
);

FILL FILL_4__3216_ (
);

FILL FILL_0__3536_ (
);

FILL FILL_0__3116_ (
);

FILL FILL_5__1979_ (
);

FILL FILL_5__2920_ (
);

FILL FILL_7__2938_ (
);

FILL FILL_5__2500_ (
);

FILL FILL_1__2912_ (
);

FILL FILL_3__2838_ (
);

FILL FILL_3__2418_ (
);

NAND2X1 _1982_ (
    .A(\AXYS[1] [2]),
    .B(_1047_),
    .Y(_1097_)
);

FILL FILL_5__3705_ (
);

OAI21X1 _2767_ (
    .A(_431_),
    .B(_197_),
    .C(_148_),
    .Y(_432_)
);

NAND2X1 _2347_ (
    .A(_1354_),
    .B(_1453_),
    .Y(_1454_)
);

FILL FILL_7__2691_ (
);

FILL FILL_7__2271_ (
);

FILL FILL_3__2591_ (
);

FILL FILL_3__2171_ (
);

FILL FILL_5__2097_ (
);

FILL FILL_4__2907_ (
);

FILL FILL_1__2089_ (
);

FILL FILL_7__3056_ (
);

FILL FILL_0__2807_ (
);

FILL FILL_1__3450_ (
);

FILL FILL_1__3030_ (
);

FILL FILL_2__1793_ (
);

FILL FILL_4__2660_ (
);

FILL FILL_4__2240_ (
);

FILL FILL_6__2586_ (
);

FILL FILL_6__2166_ (
);

FILL FILL_2__2998_ (
);

FILL FILL_0__2980_ (
);

FILL FILL_0__2560_ (
);

FILL FILL_2__2578_ (
);

FILL FILL_2__2158_ (
);

FILL FILL_0__2140_ (
);

FILL FILL_4__3025_ (
);

FILL FILL_3__1862_ (
);

FILL FILL_5__1788_ (
);

FILL FILL_7__2327_ (
);

FILL FILL_1__2721_ (
);

FILL FILL_1__2301_ (
);

FILL FILL_3__2647_ (
);

FILL FILL_3__2227_ (
);

INVX1 _1791_ (
    .A(_916_),
    .Y(_917_)
);

FILL FILL_5__3514_ (
);

FILL FILL169650x133350 (
);

FILL FILL_1__3506_ (
);

FILL FILL_4__1931_ (
);

FILL FILL_6__1857_ (
);

AOI22X1 _2996_ (
    .A(_1017_),
    .B(_1149__bF$buf0),
    .C(_617_),
    .D(_624_),
    .Y(_48_)
);

AOI22X1 _2576_ (
    .A(DIMUX[7]),
    .B(_227_),
    .C(_200_),
    .D(ABL[7]),
    .Y(_264_)
);

OAI21X1 _2156_ (
    .A(_886__bF$buf2),
    .B(_1263_),
    .C(_1264_),
    .Y(_1265_)
);

FILL FILL_7__2080_ (
);

FILL FILL_2__1849_ (
);

FILL FILL_0__1831_ (
);

FILL FILL_4__2716_ (
);

FILL FILL_7__3285_ (
);

FILL FILL_0__2616_ (
);

FILL FILL_3__3185_ (
);

FILL FILL_3__1918_ (
);

FILL FILL_6__2395_ (
);

FILL FILL_2__2387_ (
);

NAND2X1 _1847_ (
    .A(_969_),
    .B(_971_),
    .Y(_972_)
);

FILL FILL_4__3674_ (
);

FILL FILL_7__1771_ (
);

FILL FILL_4__3254_ (
);

FILL FILL_0__3574_ (
);

FILL FILL_0__3154_ (
);

FILL FILL_7__2556_ (
);

FILL FILL_1__2950_ (
);

FILL FILL_1__2530_ (
);

FILL FILL_1__2110_ (
);

FILL FILL_3__2876_ (
);

FILL FILL_3__2456_ (
);

FILL FILL_3__2036_ (
);

FILL FILL169650x61350 (
);

FILL FILL_1__3315_ (
);

AND2X2 _2385_ (
    .A(_1490_),
    .B(_1487_),
    .Y(_1491_)
);

FILL FILL_4__2945_ (
);

FILL FILL_4__2525_ (
);

FILL FILL_4__2105_ (
);

FILL FILL_0__2845_ (
);

FILL FILL_0__2425_ (
);

FILL FILL_0__2005_ (
);

FILL FILL_7__1827_ (
);

FILL FILL_1__1801_ (
);

FILL FILL_2__2196_ (
);

FILL FILL_4__3483_ (
);

FILL FILL_4__3063_ (
);

FILL FILL_7__2785_ (
);

FILL FILL_3__2685_ (
);

FILL FILL_3__2265_ (
);

FILL FILL_5__3552_ (
);

FILL FILL_5__3132_ (
);

FILL FILL_1__3544_ (
);

FILL FILL_1__3124_ (
);

FILL FILL_6__1895_ (
);

NAND2X1 _2194_ (
    .A(_929_),
    .B(_941_),
    .Y(_1303_)
);

FILL FILL_2__1887_ (
);

FILL FILL_4__2754_ (
);

FILL FILL_4__2334_ (
);

DFFSR _3399_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(_68_),
    .CLK(clk_bF$buf5),
    .Q(backwards)
);

FILL FILL_0__2654_ (
);

FILL FILL_6__3621_ (
);

FILL FILL_0__2234_ (
);

FILL FILL_6__3201_ (
);

FILL FILL_2__3613_ (
);

FILL FILL_4__3539_ (
);

FILL FILL_4__3119_ (
);

FILL FILL_3__1956_ (
);

FILL FILL_0__3019_ (
);

FILL FILL_5__2823_ (
);

FILL FILL_5__2403_ (
);

FILL FILL_1__2815_ (
);

INVX1 _1885_ (
    .A(DIMUX[2]),
    .Y(_1008_)
);

FILL FILL_4__3292_ (
);

FILL FILL_5__3608_ (
);

FILL FILL_0__3192_ (
);

FILL FILL_7__2174_ (
);

FILL FILL_0__1925_ (
);

AND2X2 _3611_ (
    .A(_1718_),
    .B(BI[6]),
    .Y(_1641_)
);

FILL FILL_3__2494_ (
);

FILL FILL_3__2074_ (
);

FILL FILL_3__3699_ (
);

FILL FILL_3__3279_ (
);

FILL FILL_4__2983_ (
);

FILL FILL_4__2563_ (
);

FILL FILL_4__2143_ (
);

FILL FILL_6__2489_ (
);

FILL FILL_6__2069_ (
);

FILL FILL_0__2883_ (
);

FILL FILL_0__2463_ (
);

FILL FILL_0__2043_ (
);

FILL FILL_6__3010_ (
);

FILL FILL_2__3002_ (
);

FILL FILL_3__1765_ (
);

FILL FILL_0__3668_ (
);

FILL FILL_0__3248_ (
);

FILL FILL_5__2632_ (
);

FILL FILL_5__2212_ (
);

FILL FILL_1__2624_ (
);

FILL FILL_1__2204_ (
);

FILL FILL_4__1834_ (
);

OAI21X1 _2899_ (
    .A(_537_),
    .B(_547_),
    .C(_546_),
    .Y(_28_)
);

OAI21X1 _2479_ (
    .A(_143_),
    .B(_1117_),
    .C(_177_),
    .Y(_1742_[4])
);

INVX2 _2059_ (
    .A(IRHOLD_valid),
    .Y(_1168_)
);

FILL FILL_6__2701_ (
);

DFFSR _3420_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_89_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[2] [4])
);

OAI21X1 _3000_ (
    .A(_627_),
    .B(_626_),
    .C(_1150__bF$buf4),
    .Y(_628_)
);

FILL FILL_4__2619_ (
);

FILL FILL_5__3590_ (
);

FILL FILL_5__3170_ (
);

FILL FILL_7__3188_ (
);

FILL FILL_0__2939_ (
);

FILL FILL_0__2519_ (
);

FILL FILL_1__3582_ (
);

FILL FILL_1__3162_ (
);

FILL FILL_3__3088_ (
);

FILL FILL_5__1903_ (
);

FILL FILL_4__2792_ (
);

FILL FILL_4__2372_ (
);

FILL FILL_6__2298_ (
);

FILL FILL_0__2692_ (
);

FILL FILL_0__2272_ (
);

FILL FILL_2__3651_ (
);

FILL FILL_2__3231_ (
);

FILL FILL_4__3577_ (
);

FILL FILL_4__3157_ (
);

FILL FILL_3__1994_ (
);

FILL FILL_0__3477_ (
);

FILL FILL_0__3057_ (
);

FILL FILL_5__2861_ (
);

FILL FILL_7__2459_ (
);

FILL FILL_5__2441_ (
);

FILL FILL_5__2021_ (
);

FILL FILL_1__2853_ (
);

FILL FILL_1__2433_ (
);

FILL FILL_1__2013_ (
);

FILL FILL_3__2779_ (
);

FILL FILL_3__2359_ (
);

FILL FILL_3__3300_ (
);

FILL FILL_5__3646_ (
);

FILL FILL_5__3226_ (
);

FILL FILL_1__3638_ (
);

FILL FILL_1__3218_ (
);

FILL FILL_6__1989_ (
);

NOR2X1 _2288_ (
    .A(_1156_),
    .B(_1214_),
    .Y(_1395_)
);

FILL FILL_0__1963_ (
);

FILL FILL_6__2930_ (
);

FILL FILL_6__2510_ (
);

FILL FILL_3_BUFX2_insert60 (
);

FILL FILL_3_BUFX2_insert61 (
);

FILL FILL_3_BUFX2_insert62 (
);

FILL FILL_3_BUFX2_insert63 (
);

FILL FILL_2__2922_ (
);

FILL FILL_2__2502_ (
);

FILL FILL_3_BUFX2_insert64 (
);

FILL FILL_3_BUFX2_insert65 (
);

FILL FILL_3_BUFX2_insert66 (
);

FILL FILL_3_BUFX2_insert67 (
);

FILL FILL_4__2848_ (
);

FILL FILL_3_BUFX2_insert68 (
);

FILL FILL_4__2428_ (
);

FILL FILL_3_BUFX2_insert69 (
);

FILL FILL_4__2008_ (
);

FILL FILL_0__2748_ (
);

FILL FILL_6__3715_ (
);

FILL FILL_0__2328_ (
);

FILL FILL_2__3707_ (
);

FILL FILL_4__2181_ (
);

FILL FILL_5__2917_ (
);

FILL FILL_0__2081_ (
);

FILL FILL_2__2099_ (
);

FILL FILL_1__2909_ (
);

FILL FILL_2__3460_ (
);

OAI21X1 _1979_ (
    .A(_1006_),
    .B(_983_),
    .C(_1094_),
    .Y(_1095_)
);

FILL FILL_2__3040_ (
);

INVX1 _2920_ (
    .A(_564_),
    .Y(_565_)
);

INVX2 _2500_ (
    .A(_194_),
    .Y(_195_)
);

FILL FILL_0__3286_ (
);

FILL FILL_7__2688_ (
);

FILL FILL_5__2670_ (
);

FILL FILL_5__2250_ (
);

BUFX2 _3705_ (
    .A(_1741_[8]),
    .Y(AB[8])
);

FILL FILL_1__2662_ (
);

FILL FILL_1__2242_ (
);

FILL FILL_3__2588_ (
);

FILL FILL_3__2168_ (
);

FILL FILL_5__3455_ (
);

FILL FILL_5__3035_ (
);

FILL FILL_1__3027_ (
);

FILL FILL_4__1872_ (
);

FILL FILL_6__1798_ (
);

INVX1 _2097_ (
    .A(_1205_),
    .Y(_1206_)
);

FILL FILL_0__1772_ (
);

FILL FILL_2__2731_ (
);

FILL FILL_2__2311_ (
);

FILL FILL_4__2657_ (
);

FILL FILL_4__2237_ (
);

FILL FILL_0__2977_ (
);

FILL FILL_0__2557_ (
);

FILL FILL_6__3524_ (
);

FILL FILL_0__2137_ (
);

FILL FILL_6__3104_ (
);

FILL FILL_2__3516_ (
);

FILL FILL_5__1941_ (
);

FILL FILL_7__1959_ (
);

FILL FILL_1__1933_ (
);

FILL FILL_3__1859_ (
);

FILL FILL_3__2800_ (
);

FILL FILL_5__2726_ (
);

FILL FILL_5__2306_ (
);

FILL FILL_1__2718_ (
);

NAND2X1 _1788_ (
    .A(_913_),
    .B(_901_),
    .Y(_914_)
);

FILL FILL_4__3195_ (
);

FILL FILL_0__3095_ (
);

FILL FILL_4__1928_ (
);

FILL FILL_7__2077_ (
);

FILL FILL_0__1828_ (
);

NAND2X1 _3514_ (
    .A(_1543_),
    .B(_1542_),
    .Y(_1544_)
);

FILL FILL_1__2891_ (
);

FILL FILL_1__2471_ (
);

FILL FILL_1__2051_ (
);

FILL FILL_3__2397_ (
);

FILL FILL_5__3264_ (
);

FILL FILL_1__3676_ (
);

FILL FILL_1__3256_ (
);

FILL FILL_2__2960_ (
);

FILL FILL_2__2540_ (
);

FILL FILL_2__2120_ (
);

FILL FILL_4__2886_ (
);

FILL FILL_4__2466_ (
);

FILL FILL_4__2046_ (
);

FILL FILL_0__2786_ (
);

FILL FILL_0__2366_ (
);

FILL FILL_5__1750_ (
);

FILL FILL_7__1768_ (
);

FILL FILL_5__2955_ (
);

FILL FILL_5__2535_ (
);

FILL FILL_5__2115_ (
);

FILL FILL_1__2947_ (
);

FILL FILL_1__2527_ (
);

FILL FILL_1__2107_ (
);

FILL FILL_2__1811_ (
);

FILL FILL_6__2604_ (
);

DFFSR _3323_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_1512_[5]),
    .CLK(clk_bF$buf6),
    .Q(state[5])
);

FILL FILL_1__2280_ (
);

FILL FILL_7_BUFX2_insert11 (
);

FILL FILL_7_BUFX2_insert13 (
);

FILL FILL_7_BUFX2_insert14 (
);

FILL FILL_7_BUFX2_insert16 (
);

FILL FILL_7_BUFX2_insert17 (
);

FILL FILL_5__3493_ (
);

FILL FILL_7_BUFX2_insert19 (
);

FILL FILL_5__3073_ (
);

FILL FILL_1__3485_ (
);

FILL FILL_1__3065_ (
);

FILL FILL_5__1806_ (
);

FILL FILL_4__2695_ (
);

FILL FILL_4__2275_ (
);

FILL FILL_0__2595_ (
);

FILL FILL_6__3562_ (
);

FILL FILL_0__2175_ (
);

FILL FILL_6__3142_ (
);

FILL FILL_2__3554_ (
);

FILL FILL_2__3134_ (
);

FILL FILL_1__1971_ (
);

FILL FILL_3__1897_ (
);

FILL FILL_5__2764_ (
);

FILL FILL_5__2344_ (
);

FILL FILL_1__2756_ (
);

FILL FILL_1__2336_ (
);

FILL FILL_7__3303_ (
);

FILL FILL_3__3623_ (
);

FILL FILL_3__3203_ (
);

FILL FILL_5__3549_ (
);

FILL FILL_5__3129_ (
);

FILL FILL_4__1966_ (
);

FILL FILL_0__1866_ (
);

FILL FILL_6__2833_ (
);

INVX1 _3552_ (
    .A(_1581_),
    .Y(_1582_)
);

FILL FILL_6__2413_ (
);

OAI21X1 _3132_ (
    .A(_722_),
    .B(_737_),
    .C(_738_),
    .Y(_70_)
);

FILL FILL169950x36150 (
);

FILL FILL_2__2825_ (
);

FILL FILL_2__2405_ (
);

FILL FILL_6__3618_ (
);

FILL FILL_1__3294_ (
);

FILL FILL_4__2084_ (
);

FILL FILL_4__3289_ (
);

OAI21X1 _2823_ (
    .A(_463_),
    .B(_464_),
    .C(_485_),
    .Y(_486_)
);

NOR2X1 _2403_ (
    .A(_1372_),
    .B(_1506_),
    .Y(_1507_)
);

FILL FILL_1__1780_ (
);

FILL FILL_0__3189_ (
);

FILL FILL168750x18150 (
);

FILL FILL_5__2993_ (
);

FILL FILL_5__2573_ (
);

FILL FILL_5__2153_ (
);

OAI21X1 _3608_ (
    .A(_1724_),
    .B(_1727_),
    .C(_1637_),
    .Y(_1638_)
);

FILL FILL_1__2985_ (
);

FILL FILL_1__2565_ (
);

FILL FILL_7__3532_ (
);

FILL FILL_1__2145_ (
);

FILL FILL_7__3112_ (
);

FILL FILL_3__3012_ (
);

FILL FILL_4__1775_ (
);

FILL FILL_6__2642_ (
);

DFFSR _3361_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_38_),
    .CLK(clk_bF$buf9),
    .Q(compare)
);

FILL FILL_6__2222_ (
);

FILL FILL_2__2634_ (
);

FILL FILL_2__2214_ (
);

FILL FILL_4__3501_ (
);

FILL FILL_6__3007_ (
);

FILL FILL_5__1844_ (
);

FILL FILL_1__1836_ (
);

FILL FILL_7__2803_ (
);

FILL FILL_3__2703_ (
);

FILL FILL_5__2629_ (
);

FILL FILL_5__2209_ (
);

FILL FILL_6__3180_ (
);

FILL FILL_2__3592_ (
);

FILL FILL_2__3172_ (
);

FILL FILL_4__3098_ (
);

FILL FILL_6__1913_ (
);

NOR2X1 _2632_ (
    .A(_309_),
    .B(_917_),
    .Y(\u_ALU8.BCD )
);

OAI21X1 _2212_ (
    .A(_886__bF$buf2),
    .B(_1319__bF$buf3),
    .C(_1320_),
    .Y(_1321_)
);

FILL FILL_2__1905_ (
);

FILL FILL_5__2382_ (
);

DFFSR _3417_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_86_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[2] [1])
);

FILL FILL_1__2794_ (
);

FILL FILL_1__2374_ (
);

FILL FILL_3__3661_ (
);

FILL FILL_3__3241_ (
);

FILL FILL_5__3587_ (
);

FILL FILL_5__3167_ (
);

FILL FILL_1__3579_ (
);

FILL FILL_1__3159_ (
);

FILL FILL_6__2871_ (
);

NAND2X1 _3590_ (
    .A(_1609_),
    .B(_1619_),
    .Y(_1620_)
);

FILL FILL_6__2451_ (
);

NOR2X1 _3170_ (
    .A(_770_),
    .B(_771_),
    .Y(_772_)
);

FILL FILL_6__2031_ (
);

FILL FILL_2__2863_ (
);

FILL FILL_2__2443_ (
);

FILL FILL_2__2023_ (
);

FILL FILL_4__2789_ (
);

FILL FILL_4__2369_ (
);

NOR2X1 _1903_ (
    .A(_931__bF$buf0),
    .B(_938_),
    .Y(_1020_)
);

FILL FILL_4__3310_ (
);

FILL FILL_0__2689_ (
);

FILL FILL_6__3656_ (
);

FILL FILL_0__2269_ (
);

FILL FILL_6__3236_ (
);

FILL FILL_2__3648_ (
);

FILL FILL_0__3630_ (
);

FILL FILL_2__3228_ (
);

FILL FILL_0__3210_ (
);

FILL FILL_7__2612_ (
);

FILL FILL_3__2932_ (
);

FILL FILL_3__2512_ (
);

FILL FILL_5__2858_ (
);

FILL FILL_5__2438_ (
);

FILL FILL_5__2018_ (
);

INVX1 _2861_ (
    .A(_519_),
    .Y(_521_)
);

OAI21X1 _2441_ (
    .A(php),
    .B(_1337_),
    .C(_1227_),
    .Y(_144_)
);

NAND3X1 _2021_ (
    .A(_1131_),
    .B(_1129_),
    .C(_1130_),
    .Y(_1132_)
);

FILL FILL_5__2191_ (
);

FILL FILL_6__2927_ (
);

NAND2X1 _3646_ (
    .A(_1635_),
    .B(_1630_),
    .Y(_1676_)
);

FILL FILL_6__2507_ (
);

OAI21X1 _3226_ (
    .A(_724_),
    .B(_807_),
    .C(_809_),
    .Y(_93_)
);

FILL FILL_1__2183_ (
);

FILL FILL_2__2919_ (
);

FILL FILL_0__2901_ (
);

FILL FILL_3__3470_ (
);

FILL FILL_3__3050_ (
);

FILL FILL_6__2680_ (
);

FILL FILL_6__2260_ (
);

FILL FILL_2__2672_ (
);

FILL FILL_2__2252_ (
);

FILL FILL_4__2598_ (
);

FILL FILL_4__2178_ (
);

FILL FILL_0__2498_ (
);

FILL FILL_6__3465_ (
);

FILL FILL_0__2078_ (
);

FILL FILL_6__3045_ (
);

FILL FILL_2__3457_ (
);

FILL FILL_2__3037_ (
);

FILL FILL_5__1882_ (
);

OAI21X1 _2917_ (
    .A(_1217_),
    .B(_1396_),
    .C(_557_),
    .Y(_562_)
);

FILL FILL_1__1874_ (
);

FILL FILL_7__2841_ (
);

FILL FILL_7__2421_ (
);

FILL FILL_7__2001_ (
);

FILL FILL_3__2741_ (
);

FILL FILL_3__2321_ (
);

FILL FILL_5__2667_ (
);

FILL FILL_5__2247_ (
);

FILL FILL_1__2659_ (
);

FILL FILL_1__2239_ (
);

FILL FILL_7__3206_ (
);

FILL FILL_1__3600_ (
);

FILL FILL_3__3526_ (
);

FILL FILL_3__3106_ (
);

FILL FILL_6__1951_ (
);

OAI21X1 _2670_ (
    .A(_1153_),
    .B(res),
    .C(_1334_),
    .Y(_343_)
);

OAI22X1 _2250_ (
    .A(RDY_bF$buf5),
    .B(_972_),
    .C(_1149__bF$buf3),
    .D(_1357_),
    .Y(_1358_)
);

FILL FILL_2__1943_ (
);

FILL FILL_4__1869_ (
);

FILL FILL_4__2810_ (
);

FILL FILL_0__1769_ (
);

FILL FILL_6__2736_ (
);

INVX1 _3455_ (
    .A(\u_ALU8.AI7 ),
    .Y(_1703_)
);

FILL FILL_6__2316_ (
);

OAI21X1 _3035_ (
    .A(_1013_),
    .B(_647_),
    .C(_653_),
    .Y(_58_)
);

FILL FILL_0__2710_ (
);

FILL FILL_2__2728_ (
);

FILL FILL_2__2308_ (
);

FILL FILL_1__3197_ (
);

FILL FILL168450x133350 (
);

FILL FILL_5__1938_ (
);

FILL FILL_2__2481_ (
);

FILL FILL_2__2061_ (
);

NAND2X1 _1941_ (
    .A(\AXYS[2] [0]),
    .B(_1057_),
    .Y(_1058_)
);

FILL FILL_6__3694_ (
);

FILL FILL_6__3274_ (
);

FILL FILL_2__3266_ (
);

OAI21X1 _2726_ (
    .A(_394_),
    .B(_387_),
    .C(RDY_bF$buf0),
    .Y(_395_)
);

OAI21X1 _2306_ (
    .A(_1181_),
    .B(_1412_),
    .C(_1393_),
    .Y(_1413_)
);

FILL FILL_7__2650_ (
);

FILL FILL_7__2230_ (
);

FILL FILL_3__2970_ (
);

FILL FILL_3__2550_ (
);

FILL FILL_3__2130_ (
);

FILL FILL_5__2896_ (
);

FILL FILL_5__2476_ (
);

FILL FILL_5__2056_ (
);

FILL FILL_1__2888_ (
);

FILL FILL_1__2468_ (
);

FILL FILL_1__2048_ (
);

FILL FILL_6__1760_ (
);

FILL FILL_2__1752_ (
);

FILL FILL_0__1998_ (
);

FILL FILL_6__2965_ (
);

DFFSR _3684_ (
    .R(_1513_),
    .S(vdd),
    .D(_1519_),
    .CLK(clk_bF$buf3),
    .Q(ADD[2])
);

FILL FILL_6__2545_ (
);

NOR2X1 _3264_ (
    .A(_1201_),
    .B(_1309_),
    .Y(_840_)
);

FILL FILL_6__2125_ (
);

FILL FILL_2__2957_ (
);

FILL FILL_2__2537_ (
);

FILL FILL_2__2117_ (
);

FILL FILL_7__1921_ (
);

FILL FILL_3__1821_ (
);

FILL FILL_0__3304_ (
);

FILL FILL_5__1747_ (
);

FILL FILL_7__2706_ (
);

FILL FILL_2__2290_ (
);

FILL FILL_3__2606_ (
);

INVX1 _1750_ (
    .A(DIHOLD[2]),
    .Y(_882_)
);

FILL FILL_6__3083_ (
);

FILL FILL_2__3495_ (
);

FILL FILL_2__3075_ (
);

FILL FILL_6__1816_ (
);

OAI21X1 _2955_ (
    .A(_1037_),
    .B(_1263_),
    .C(RDY_bF$buf2),
    .Y(_592_)
);

AND2X2 _2535_ (
    .A(_226_),
    .B(_228_),
    .Y(_229_)
);

INVX1 _2115_ (
    .A(_1196_),
    .Y(_1224_)
);

FILL FILL_2__1808_ (
);

FILL FILL_5__2285_ (
);

FILL FILL_1__2697_ (
);

FILL FILL_7__3664_ (
);

FILL FILL_1__2277_ (
);

FILL FILL_7__3244_ (
);

FILL FILL_3__3564_ (
);

FILL FILL_3__3144_ (
);

FILL FILL_2__1981_ (
);

FILL FILL_6__2774_ (
);

OAI21X1 _3493_ (
    .A(_1737_),
    .B(_1736_),
    .C(_1733_),
    .Y(_1738_)
);

FILL FILL_6__2354_ (
);

OAI21X1 _3073_ (
    .A(_680_),
    .B(_684_),
    .C(_685_),
    .Y(_64_)
);

FILL FILL_2__2766_ (
);

FILL FILL_2__2346_ (
);

OAI21X1 _1806_ (
    .A(_928_),
    .B(_931__bF$buf3),
    .C(_930_),
    .Y(_932_)
);

FILL FILL_4__3633_ (
);

FILL FILL_4__3213_ (
);

FILL FILL_6__3559_ (
);

FILL FILL_6__3139_ (
);

FILL FILL_0__3533_ (
);

FILL FILL_0__3113_ (
);

FILL FILL_5__1976_ (
);

FILL FILL_1__1968_ (
);

FILL FILL_7__2935_ (
);

FILL FILL_3__2835_ (
);

FILL FILL_3__2415_ (
);

FILL FILL_5__3702_ (
);

OAI22X1 _2764_ (
    .A(RDY_bF$buf4),
    .B(_276_),
    .C(_424_),
    .D(_429_),
    .Y(_11_)
);

NOR2X1 _2344_ (
    .A(_1450_),
    .B(_1445_),
    .Y(_1451_)
);

FILL FILL_5__2094_ (
);

FILL FILL_4__2904_ (
);

NAND2X1 _3549_ (
    .A(alu_shift_right),
    .B(AI[1]),
    .Y(_1579_)
);

OAI21X1 _3129_ (
    .A(_1006_),
    .B(_1018_),
    .C(_735_),
    .Y(_736_)
);

FILL FILL_1__2086_ (
);

FILL FILL_7__3053_ (
);

FILL FILL_0__2804_ (
);

FILL FILL_5__3299_ (
);

FILL FILL_2__1790_ (
);

FILL FILL_6__2583_ (
);

FILL FILL_6__2163_ (
);

FILL FILL_2__2995_ (
);

FILL FILL_2__2575_ (
);

FILL FILL_2__2155_ (
);

FILL FILL_4__3022_ (
);

FILL FILL_5__1785_ (
);

FILL FILL_1__1777_ (
);

FILL FILL_7__2324_ (
);

FILL FILL_3__2644_ (
);

FILL FILL_3__2224_ (
);

FILL FILL_7__3529_ (
);

FILL FILL_5__3511_ (
);

FILL FILL_7__3109_ (
);

FILL FILL_1__3503_ (
);

FILL FILL_3__3009_ (
);

FILL FILL_6__1854_ (
);

OAI21X1 _2993_ (
    .A(_596_),
    .B(_1397_),
    .C(_609_),
    .Y(_622_)
);

AOI21X1 _2573_ (
    .A(_1132_),
    .B(_195_),
    .C(_261_),
    .Y(_262_)
);

OAI21X1 _2153_ (
    .A(_886__bF$buf6),
    .B(_1260_),
    .C(_1261_),
    .Y(_1262_)
);

FILL FILL_2__1846_ (
);

FILL FILL_4__2713_ (
);

FILL FILL_6__2639_ (
);

DFFSR _3358_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_35_),
    .CLK(clk_bF$buf4),
    .Q(op[3])
);

FILL FILL_6__2219_ (
);

FILL FILL_7__3282_ (
);

FILL FILL_0__2613_ (
);

FILL FILL_3__3182_ (
);

FILL FILL_3__1915_ (
);

FILL FILL169050x18150 (
);

FILL FILL_6__2392_ (
);

FILL FILL_2__2384_ (
);

INVX4 _1844_ (
    .A(_931__bF$buf3),
    .Y(_969_)
);

FILL FILL_4__3671_ (
);

FILL FILL_4__3251_ (
);

FILL FILL_6__3597_ (
);

FILL FILL_6__3177_ (
);

FILL FILL_2__3589_ (
);

FILL FILL_0__3571_ (
);

FILL FILL_2__3169_ (
);

FILL FILL_0__3151_ (
);

FILL FILL_7_CLKBUF1_insert30 (
);

FILL FILL_7_CLKBUF1_insert32 (
);

FILL FILL_7_CLKBUF1_insert34 (
);

FILL FILL_7_CLKBUF1_insert35 (
);

INVX1 _2629_ (
    .A(adc_sbc),
    .Y(_308_)
);

INVX1 _2209_ (
    .A(_1317_),
    .Y(_1318_)
);

FILL FILL_7__2553_ (
);

FILL FILL_3__2873_ (
);

FILL FILL_3__2453_ (
);

FILL FILL_3__2033_ (
);

FILL FILL_5__2799_ (
);

FILL FILL_5__2379_ (
);

FILL FILL_1__3312_ (
);

FILL FILL_3__3658_ (
);

FILL FILL_3__3238_ (
);

INVX1 _2382_ (
    .A(_1266_),
    .Y(_1488_)
);

FILL FILL_4__2942_ (
);

FILL FILL_4__2522_ (
);

FILL FILL_4__2102_ (
);

FILL FILL_6__2868_ (
);

MUX2X1 _3587_ (
    .A(_1616_),
    .B(_1615_),
    .S(_1568_),
    .Y(_1617_)
);

FILL FILL_6__2448_ (
);

FILL FILL_6__2028_ (
);

INVX1 _3167_ (
    .A(ADD[6]),
    .Y(_769_)
);

FILL FILL_7__3091_ (
);

FILL FILL_0__2842_ (
);

FILL FILL_0__2422_ (
);

FILL FILL_0__2002_ (
);

FILL FILL_7__1824_ (
);

FILL FILL_4__3307_ (
);

FILL FILL_0__3627_ (
);

FILL FILL_0__3207_ (
);

FILL FILL_7__2609_ (
);

FILL FILL169650x82950 (
);

FILL FILL167850x144150 (
);

FILL FILL_2__2193_ (
);

FILL FILL_3__2929_ (
);

FILL FILL_3__2509_ (
);

FILL FILL_4__3480_ (
);

FILL FILL_4__3060_ (
);

OAI21X1 _2858_ (
    .A(_893_),
    .B(_351_),
    .C(_517_),
    .Y(_518_)
);

OAI21X1 _2438_ (
    .A(_1199_),
    .B(_141_),
    .C(store),
    .Y(_142_)
);

NAND2X1 _2018_ (
    .A(\AXYS[1] [6]),
    .B(_1047_),
    .Y(_1129_)
);

FILL FILL_7__2782_ (
);

FILL FILL_7__2362_ (
);

FILL FILL_3__2682_ (
);

FILL FILL_3__2262_ (
);

FILL FILL_5__2188_ (
);

FILL FILL_7__3567_ (
);

FILL FILL_1__3541_ (
);

FILL FILL_1__3121_ (
);

FILL FILL_3__3467_ (
);

FILL FILL_3__3047_ (
);

FILL FILL_6__1892_ (
);

OAI21X1 _2191_ (
    .A(RDY_bF$buf7),
    .B(_1299_),
    .C(_1298_),
    .Y(_1300_)
);

FILL FILL_2__1884_ (
);

FILL FILL168450x64950 (
);

FILL FILL_4__2751_ (
);

FILL FILL_4__2331_ (
);

FILL FILL_6__2677_ (
);

DFFSR _3396_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_65_),
    .CLK(clk_bF$buf1),
    .Q(N)
);

FILL FILL_6__2257_ (
);

FILL FILL_2__2669_ (
);

FILL FILL_0__2651_ (
);

FILL FILL_0__2231_ (
);

FILL FILL_2__2249_ (
);

FILL FILL_2__3610_ (
);

FILL FILL_4__3536_ (
);

FILL FILL_4__3116_ (
);

FILL FILL_3__1953_ (
);

FILL FILL_0__3016_ (
);

FILL FILL_5__1879_ (
);

FILL FILL_7__2838_ (
);

FILL FILL_5__2820_ (
);

FILL FILL_5__2400_ (
);

FILL FILL_1__2812_ (
);

FILL FILL_3__2738_ (
);

FILL FILL_3__2318_ (
);

INVX2 _1882_ (
    .A(DIMUX[1]),
    .Y(_1006_)
);

FILL FILL_5__3605_ (
);

FILL FILL_6__1948_ (
);

NAND2X1 _2667_ (
    .A(RDY_bF$buf3),
    .B(_340_),
    .Y(_341_)
);

NAND2X1 _2247_ (
    .A(_1178_),
    .B(_1181_),
    .Y(_1355_)
);

FILL FILL_7__2591_ (
);

FILL FILL_7__2171_ (
);

FILL FILL_0__1922_ (
);

FILL FILL_3__2491_ (
);

FILL FILL_3__2071_ (
);

FILL FILL_4__2807_ (
);

FILL FILL_0__2707_ (
);

FILL FILL_3__3696_ (
);

FILL FILL_3__3276_ (
);

FILL FILL169950x133350 (
);

FILL FILL_4__2980_ (
);

FILL FILL_4__2560_ (
);

FILL FILL_4__2140_ (
);

FILL FILL_6__2486_ (
);

FILL FILL_6__2066_ (
);

FILL FILL_0__2880_ (
);

FILL FILL_2__2898_ (
);

FILL FILL_2__2478_ (
);

FILL FILL_0__2460_ (
);

FILL FILL_2__2058_ (
);

FILL FILL_0__2040_ (
);

INVX1 _1938_ (
    .A(src_reg[0]),
    .Y(_1055_)
);

FILL FILL_3__1762_ (
);

FILL FILL_0__3665_ (
);

FILL FILL_0__3245_ (
);

FILL FILL_7__2227_ (
);

FILL FILL_1__2621_ (
);

FILL FILL_1__2201_ (
);

FILL FILL_3__2967_ (
);

FILL FILL_3__2547_ (
);

FILL FILL_3__2127_ (
);

FILL FILL_4__1831_ (
);

FILL FILL_6__1757_ (
);

OAI22X1 _2896_ (
    .A(_545_),
    .B(_1150__bF$buf2),
    .C(_541_),
    .D(_544_),
    .Y(_27_)
);

OAI21X1 _2476_ (
    .A(_1319__bF$buf0),
    .B(_1263_),
    .C(PC[12]),
    .Y(_175_)
);

INVX1 _2056_ (
    .A(I),
    .Y(_1165_)
);

FILL FILL_2__1749_ (
);

FILL FILL_4__2616_ (
);

FILL FILL_7__3185_ (
);

FILL FILL_0__2936_ (
);

FILL FILL_0__2516_ (
);

FILL FILL_3__3085_ (
);

FILL FILL_5__1900_ (
);

FILL FILL_3__1818_ (
);

FILL FILL_6__2295_ (
);

FILL FILL_2__2287_ (
);

INVX1 _1747_ (
    .A(DIHOLD[1]),
    .Y(_880_)
);

FILL FILL_4__3574_ (
);

FILL FILL_4__3154_ (
);

FILL FILL_3__1991_ (
);

FILL FILL_0__3474_ (
);

FILL FILL_0__3054_ (
);

FILL FILL_7__2456_ (
);

FILL FILL_1__2850_ (
);

FILL FILL_1__2430_ (
);

FILL FILL_1__2010_ (
);

FILL FILL_3__2776_ (
);

FILL FILL_3__2356_ (
);

FILL FILL_5__3643_ (
);

FILL FILL_5__3223_ (
);

FILL FILL_1__3635_ (
);

FILL FILL_1__3215_ (
);

FILL FILL_6__1986_ (
);

NAND2X1 _2285_ (
    .A(_1343_),
    .B(_1392_),
    .Y(_1512_[1])
);

FILL FILL_2__1978_ (
);

FILL FILL_0__1960_ (
);

FILL FILL_3_BUFX2_insert37 (
);

FILL FILL_4__2845_ (
);

FILL FILL_3_BUFX2_insert38 (
);

FILL FILL_3_BUFX2_insert39 (
);

FILL FILL_4__2425_ (
);

FILL FILL_4__2005_ (
);

FILL FILL_0__2745_ (
);

FILL FILL_6__3712_ (
);

FILL FILL_0__2325_ (
);

FILL FILL_2__3704_ (
);

FILL FILL_5__2914_ (
);

FILL FILL_2__2096_ (
);

FILL FILL_1__2906_ (
);

NAND2X1 _1976_ (
    .A(_929_),
    .B(_952_),
    .Y(_1092_)
);

FILL FILL_0__3283_ (
);

FILL FILL_7__2685_ (
);

BUFX2 _3702_ (
    .A(_1741_[5]),
    .Y(AB[5])
);

FILL FILL_3__2585_ (
);

FILL FILL_3__2165_ (
);

FILL FILL_5__3452_ (
);

FILL FILL_5__3032_ (
);

FILL FILL_1__3024_ (
);

FILL FILL_6__1795_ (
);

OAI21X1 _2094_ (
    .A(_914__bF$buf3),
    .B(_974_),
    .C(_1202_),
    .Y(_1203_)
);

FILL FILL_2__1787_ (
);

FILL FILL_4__2654_ (
);

FILL FILL_4__2234_ (
);

NAND2X1 _3299_ (
    .A(ABL[7]),
    .B(_860_),
    .Y(_868_)
);

FILL FILL_0__2974_ (
);

FILL FILL_0__2554_ (
);

FILL FILL_6__3521_ (
);

FILL FILL_0__2134_ (
);

FILL FILL_6__3101_ (
);

FILL FILL_2__3513_ (
);

FILL FILL_7__1956_ (
);

FILL FILL_4__3019_ (
);

FILL FILL_1__1930_ (
);

FILL FILL_3__1856_ (
);

FILL FILL_5__2723_ (
);

FILL FILL_5__2303_ (
);

FILL FILL_1__2715_ (
);

NOR2X1 _1785_ (
    .A(state[1]),
    .B(_906_),
    .Y(_911_)
);

FILL FILL_4__3192_ (
);

FILL FILL169650x14550 (
);

FILL FILL_5__3508_ (
);

FILL FILL_0__3092_ (
);

FILL FILL_4__1925_ (
);

FILL FILL_7__2074_ (
);

FILL FILL_0__1825_ (
);

OAI21X1 _3511_ (
    .A(_1539_),
    .B(_1540_),
    .C(_1717_),
    .Y(_1541_)
);

FILL FILL_3__2394_ (
);

FILL FILL_7__3699_ (
);

FILL FILL_5__3261_ (
);

FILL FILL_1__3673_ (
);

FILL FILL_1__3253_ (
);

FILL FILL_3__3599_ (
);

FILL FILL_3__3179_ (
);

FILL FILL_4__2883_ (
);

FILL FILL_4__2463_ (
);

FILL FILL_4__2043_ (
);

FILL FILL_6__2389_ (
);

FILL FILL_0__2783_ (
);

FILL FILL_0__2363_ (
);

FILL FILL_4__3668_ (
);

FILL FILL_4__3248_ (
);

FILL FILL_0__3568_ (
);

FILL FILL_0__3148_ (
);

FILL FILL_4_BUFX2_insert80 (
);

FILL FILL_4_BUFX2_insert81 (
);

FILL FILL_4_BUFX2_insert82 (
);

FILL FILL_4_BUFX2_insert83 (
);

FILL FILL_5__2952_ (
);

FILL FILL_5__2532_ (
);

FILL FILL_5__2112_ (
);

FILL FILL_1__2944_ (
);

FILL FILL_1__2524_ (
);

FILL FILL_1__2104_ (
);

FILL FILL_5__3317_ (
);

FILL FILL_1__3309_ (
);

NOR2X1 _2799_ (
    .A(_459_),
    .B(_461_),
    .Y(_462_)
);

INVX1 _2379_ (
    .A(_1248_),
    .Y(_1485_)
);

FILL FILL_6__2601_ (
);

DFFSR _3320_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_1512_[2]),
    .CLK(clk_bF$buf6),
    .Q(state[2])
);

FILL FILL_4__2939_ (
);

FILL FILL_4__2519_ (
);

FILL FILL_5__3490_ (
);

FILL FILL_7__3088_ (
);

FILL FILL_5__3070_ (
);

FILL FILL_0__2839_ (
);

FILL FILL_0__2419_ (
);

FILL FILL_1__3482_ (
);

FILL FILL_1__3062_ (
);

FILL FILL_5__1803_ (
);

FILL FILL_4__2692_ (
);

FILL FILL_4__2272_ (
);

FILL FILL_6__2198_ (
);

FILL FILL_0__2592_ (
);

FILL FILL_0__2172_ (
);

FILL FILL_2__3551_ (
);

FILL FILL_2__3131_ (
);

FILL FILL_4__3477_ (
);

FILL FILL_4__3057_ (
);

FILL FILL_3__1894_ (
);

FILL FILL_5__2761_ (
);

FILL FILL_7__2359_ (
);

FILL FILL_5__2341_ (
);

FILL FILL_1__2753_ (
);

FILL FILL_1__2333_ (
);

FILL FILL_3__2679_ (
);

FILL FILL_3__2259_ (
);

FILL FILL_3__3620_ (
);

FILL FILL_3__3200_ (
);

FILL FILL_5__3546_ (
);

FILL FILL_5__3126_ (
);

FILL FILL_1__3538_ (
);

FILL FILL_1__3118_ (
);

FILL FILL_4__1963_ (
);

FILL FILL_6__1889_ (
);

NAND2X1 _2188_ (
    .A(_1295_),
    .B(_1296_),
    .Y(_1297_)
);

FILL FILL_0__1863_ (
);

FILL FILL_6__2830_ (
);

FILL FILL_6__2410_ (
);

FILL FILL_2__2822_ (
);

FILL FILL_2__2402_ (
);

FILL FILL_4__2748_ (
);

FILL FILL_4__2328_ (
);

FILL FILL_0__2648_ (
);

FILL FILL_6__3615_ (
);

FILL FILL_0__2228_ (
);

FILL FILL_1__3291_ (
);

FILL FILL_2__3607_ (
);

FILL FILL_4__2081_ (
);

FILL FILL_5__2817_ (
);

FILL FILL169950x90150 (
);

FILL FILL_1__2809_ (
);

NAND3X1 _1879_ (
    .A(_980_),
    .B(_986_),
    .C(_1003_),
    .Y(_1004_)
);

FILL FILL_4__3286_ (
);

OAI22X1 _2820_ (
    .A(_481_),
    .B(_482_),
    .C(_427_),
    .D(_426_),
    .Y(_483_)
);

NOR2X1 _2400_ (
    .A(_1358_),
    .B(_1504_),
    .Y(_1505_)
);

FILL FILL_0__3186_ (
);

FILL FILL169950x57750 (
);

FILL FILL_5__2990_ (
);

FILL FILL_7__2588_ (
);

FILL FILL_5__2570_ (
);

FILL FILL_5__2150_ (
);

FILL FILL_0__1919_ (
);

INVX1 _3605_ (
    .A(_1634_),
    .Y(_1635_)
);

FILL FILL_1__2982_ (
);

FILL FILL_1__2562_ (
);

FILL FILL_1__2142_ (
);

FILL FILL_3__2488_ (
);

FILL FILL_3__2068_ (
);

FILL FILL_4__1772_ (
);

FILL FILL_2__2631_ (
);

FILL FILL_2__2211_ (
);

FILL FILL_4__2977_ (
);

FILL FILL_4__2557_ (
);

FILL FILL_4__2137_ (
);

FILL FILL_0__2877_ (
);

FILL FILL_0__2457_ (
);

FILL FILL_0__2037_ (
);

FILL FILL_6__3004_ (
);

FILL FILL_5__1841_ (
);

FILL FILL_7__1859_ (
);

FILL FILL168750x39750 (
);

FILL FILL_1__1833_ (
);

FILL FILL_3__1759_ (
);

FILL FILL_3__2700_ (
);

FILL FILL_5__2626_ (
);

FILL FILL_5__2206_ (
);

FILL FILL_1__2618_ (
);

FILL FILL_4__3095_ (
);

FILL FILL_6__1910_ (
);

FILL FILL_2__1902_ (
);

FILL FILL_4__1828_ (
);

DFFSR _3414_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_83_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[1] [6])
);

FILL FILL_1__2791_ (
);

FILL FILL_1__2371_ (
);

FILL FILL_3__2297_ (
);

FILL FILL_5__3584_ (
);

FILL FILL_5__3164_ (
);

FILL FILL_1__3576_ (
);

FILL FILL_1__3156_ (
);

FILL FILL_2__2860_ (
);

FILL FILL_2__2440_ (
);

FILL FILL_2__2020_ (
);

FILL FILL_4__2786_ (
);

FILL FILL_4__2366_ (
);

INVX1 _1900_ (
    .A(src_reg[1]),
    .Y(_1017_)
);

FILL FILL_0__2686_ (
);

FILL FILL_6__3653_ (
);

FILL FILL_0__2266_ (
);

FILL FILL_6__3233_ (
);

FILL FILL_2__3645_ (
);

FILL FILL_2__3225_ (
);

FILL FILL_3__1988_ (
);

FILL FILL_5__2855_ (
);

FILL FILL_5__2435_ (
);

FILL FILL_5__2015_ (
);

FILL FILL_1__2847_ (
);

FILL FILL_1__2427_ (
);

FILL FILL_1__2007_ (
);

FILL FILL_3__3714_ (
);

FILL FILL_0__1957_ (
);

FILL FILL_6__2924_ (
);

NAND2X1 _3643_ (
    .A(_1654_),
    .B(_1672_),
    .Y(_1673_)
);

FILL FILL_6__2504_ (
);

NAND2X1 _3223_ (
    .A(_721_),
    .B(_1049_),
    .Y(_807_)
);

FILL FILL_1__2180_ (
);

FILL FILL_2__2916_ (
);

FILL FILL_6__3709_ (
);

FILL FILL_4__2595_ (
);

FILL FILL_4__2175_ (
);

FILL FILL_0__2495_ (
);

FILL FILL_6__3462_ (
);

FILL FILL_0__2075_ (
);

FILL FILL_6__3042_ (
);

FILL FILL_2__3454_ (
);

FILL FILL_2__3034_ (
);

FILL FILL_7__1897_ (
);

NOR2X1 _2914_ (
    .A(_1412_),
    .B(_1348_),
    .Y(_559_)
);

FILL FILL_1__1871_ (
);

FILL FILL_3__1797_ (
);

FILL FILL_5__2664_ (
);

FILL FILL_5__2244_ (
);

FILL FILL_1__2656_ (
);

FILL FILL_1__2236_ (
);

FILL FILL_7__3203_ (
);

FILL FILL_3__3523_ (
);

FILL FILL_3__3103_ (
);

FILL FILL_5__3449_ (
);

FILL FILL_5__3029_ (
);

FILL FILL_2__1940_ (
);

FILL FILL_4__1866_ (
);

FILL FILL_0__1766_ (
);

FILL FILL_6__2733_ (
);

NOR2X1 _3452_ (
    .A(ADD[1]),
    .B(ADD[2]),
    .Y(_1701_)
);

FILL FILL_6__2313_ (
);

OAI21X1 _3032_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[4]),
    .Y(_652_)
);

FILL FILL_2__2725_ (
);

FILL FILL_2__2305_ (
);

FILL FILL_6__3518_ (
);

FILL FILL_1__3194_ (
);

FILL FILL_5__1935_ (
);

FILL FILL_1__1927_ (
);

FILL FILL_6__3691_ (
);

FILL FILL_6__3271_ (
);

FILL FILL_2__3263_ (
);

FILL FILL_4__3189_ (
);

OAI21X1 _2723_ (
    .A(_1014_),
    .B(_330_),
    .C(_391_),
    .Y(_392_)
);

OAI21X1 _2303_ (
    .A(_1190_),
    .B(_1409_),
    .C(_1252_),
    .Y(_1410_)
);

FILL FILL_0__3089_ (
);

FILL FILL_5__2893_ (
);

FILL FILL_5__2473_ (
);

FILL FILL_5__2053_ (
);

INVX1 _3508_ (
    .A(BI[3]),
    .Y(_1538_)
);

FILL FILL_1__2885_ (
);

FILL FILL_1__2465_ (
);

FILL FILL_1__2045_ (
);

FILL FILL_7__3012_ (
);

FILL FILL_5__3678_ (
);

FILL FILL_5__3258_ (
);

FILL FILL_0__1995_ (
);

FILL FILL_6__2962_ (
);

DFFSR _3681_ (
    .R(_1513_),
    .S(vdd),
    .D(_1516_),
    .CLK(clk_bF$buf3),
    .Q(HC)
);

FILL FILL_6__2542_ (
);

AND2X2 _3261_ (
    .A(_836_),
    .B(_1019_),
    .Y(_837_)
);

FILL FILL_6__2122_ (
);

FILL FILL_2__2954_ (
);

FILL FILL_2__2534_ (
);

FILL FILL_2__2114_ (
);

FILL FILL_0__3301_ (
);

FILL FILL_5__1744_ (
);

FILL FILL_7__2703_ (
);

FILL FILL_3__2603_ (
);

FILL FILL_5__2949_ (
);

FILL FILL_5__2529_ (
);

FILL FILL_5__2109_ (
);

FILL FILL_6__3080_ (
);

FILL FILL_2__3492_ (
);

FILL FILL_2__3072_ (
);

FILL FILL_6__1813_ (
);

OAI21X1 _2952_ (
    .A(_1149__bF$buf4),
    .B(_575_),
    .C(_590_),
    .Y(_38_)
);

OAI21X1 _2532_ (
    .A(_216_),
    .B(_209_),
    .C(ADD[1]),
    .Y(_226_)
);

NOR2X1 _2112_ (
    .A(_970_),
    .B(_976_),
    .Y(_1221_)
);

FILL FILL_2__1805_ (
);

FILL FILL_5__2282_ (
);

OAI21X1 _3317_ (
    .A(_1144_),
    .B(_869_),
    .C(_877_),
    .Y(_116_)
);

FILL FILL_1__2694_ (
);

FILL FILL_7__3661_ (
);

FILL FILL_1__2274_ (
);

FILL FILL_7__3241_ (
);

FILL FILL_3__3561_ (
);

FILL FILL_3__3141_ (
);

FILL FILL_5__3487_ (
);

FILL FILL_5__3067_ (
);

FILL FILL_1__3479_ (
);

FILL FILL_1__3059_ (
);

FILL FILL_6__2771_ (
);

NAND2X1 _3490_ (
    .A(AI[5]),
    .B(_1734_),
    .Y(_1735_)
);

FILL FILL_6__2351_ (
);

OAI21X1 _3070_ (
    .A(_1008_),
    .B(_956_),
    .C(_682_),
    .Y(_683_)
);

FILL FILL_2__2763_ (
);

FILL FILL_2__2343_ (
);

FILL FILL_4__2689_ (
);

FILL FILL_4__2269_ (
);

NOR2X1 _1803_ (
    .A(state[5]),
    .B(state[4]),
    .Y(_929_)
);

FILL FILL_4__3630_ (
);

FILL FILL_4__3210_ (
);

FILL FILL_0__2589_ (
);

FILL FILL_6__3556_ (
);

FILL FILL_0__2169_ (
);

FILL FILL_6__3136_ (
);

FILL FILL_0__3530_ (
);

FILL FILL_2__3548_ (
);

FILL FILL_2__3128_ (
);

FILL FILL_0__3110_ (
);

FILL FILL_5__1973_ (
);

FILL FILL_1__1965_ (
);

FILL FILL_7__2932_ (
);

FILL FILL_7__2512_ (
);

FILL FILL_3__2832_ (
);

FILL FILL_3__2412_ (
);

FILL FILL_5__2758_ (
);

FILL FILL_5__2338_ (
);

FILL FILL_3__3617_ (
);

NOR2X1 _2761_ (
    .A(_268_),
    .B(_352_),
    .Y(_427_)
);

OAI21X1 _2341_ (
    .A(_886__bF$buf0),
    .B(_1309_),
    .C(_1447_),
    .Y(_1448_)
);

FILL FILL_5__2091_ (
);

FILL FILL_4__2901_ (
);

FILL FILL_6__2827_ (
);

INVX1 _3546_ (
    .A(AI[0]),
    .Y(_1576_)
);

FILL FILL_6__2407_ (
);

INVX1 _3126_ (
    .A(_732_),
    .Y(_733_)
);

FILL FILL_1__2083_ (
);

FILL FILL_2__2819_ (
);

FILL FILL_0__2801_ (
);

FILL FILL_5__3296_ (
);

FILL FILL_1__3288_ (
);

FILL FILL_6__2580_ (
);

FILL FILL_6__2160_ (
);

FILL FILL_2__2992_ (
);

FILL FILL_2__2572_ (
);

FILL FILL_2__2152_ (
);

FILL FILL_4__2498_ (
);

FILL FILL_4__2078_ (
);

FILL FILL_0__2398_ (
);

FILL FILL_5__1782_ (
);

FILL FILL168750x133350 (
);

NAND2X1 _2817_ (
    .A(_1037_),
    .B(_449_),
    .Y(_480_)
);

FILL FILL_1__1774_ (
);

FILL FILL_7__2741_ (
);

FILL FILL_7__2321_ (
);

FILL FILL_3__2641_ (
);

FILL FILL_3__2221_ (
);

FILL FILL_5__2987_ (
);

FILL FILL_5__2567_ (
);

FILL FILL_5__2147_ (
);

FILL FILL_1__2979_ (
);

FILL FILL_1__2559_ (
);

FILL FILL_1__2139_ (
);

FILL FILL_7__3106_ (
);

FILL FILL_1__3500_ (
);

FILL FILL_3__3006_ (
);

FILL FILL_6__1851_ (
);

OAI21X1 _2990_ (
    .A(_1055_),
    .B(_1150__bF$buf4),
    .C(_619_),
    .Y(_47_)
);

AOI22X1 _2570_ (
    .A(DIMUX[6]),
    .B(_227_),
    .C(_200_),
    .D(ABL[6]),
    .Y(_259_)
);

OAI21X1 _2150_ (
    .A(_886__bF$buf6),
    .B(_1257_),
    .C(_1258_),
    .Y(_1259_)
);

FILL FILL_2__1843_ (
);

FILL FILL_4__1769_ (
);

FILL FILL_4__2710_ (
);

FILL FILL_6__2636_ (
);

DFFSR _3355_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_32_),
    .CLK(clk_bF$buf10),
    .Q(op[0])
);

FILL FILL_6__2216_ (
);

FILL FILL_0__2610_ (
);

FILL FILL_2__2628_ (
);

FILL FILL_2__2208_ (
);

FILL FILL_1__3097_ (
);

FILL FILL_3__1912_ (
);

FILL FILL_5__1838_ (
);

CLKBUF1 CLKBUF1_insert26 (
    .A(clk),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert27 (
    .A(clk),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert28 (
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert29 (
    .A(clk),
    .Y(clk_bF$buf7)
);

FILL FILL_2__2381_ (
);

INVX2 _1841_ (
    .A(DIMUX[0]),
    .Y(_966_)
);

FILL FILL_6__3594_ (
);

FILL FILL_6__3174_ (
);

FILL FILL_2__3586_ (
);

FILL FILL_2__3166_ (
);

FILL FILL_6__1907_ (
);

OAI21X1 _2626_ (
    .A(_1144_),
    .B(_270_),
    .C(_305_),
    .Y(_306_)
);

OAI21X1 _2206_ (
    .A(_902__bF$buf2),
    .B(_1075_),
    .C(RDY_bF$buf1),
    .Y(_1315_)
);

FILL FILL_7__2970_ (
);

FILL FILL_7__2550_ (
);

FILL FILL_7__2130_ (
);

FILL FILL_3__2870_ (
);

FILL FILL_3__2450_ (
);

FILL FILL_3__2030_ (
);

FILL FILL_5__2796_ (
);

FILL FILL_5__2376_ (
);

FILL FILL_1__2788_ (
);

FILL FILL_1__2368_ (
);

FILL FILL_3__3655_ (
);

FILL FILL_3__3235_ (
);

FILL FILL169050x39750 (
);

FILL FILL_4__1998_ (
);

FILL FILL_0__1898_ (
);

FILL FILL_6__2865_ (
);

OAI21X1 _3584_ (
    .A(_1612_),
    .B(_1613_),
    .C(_1611_),
    .Y(_1614_)
);

FILL FILL_6__2445_ (
);

FILL FILL_6__2025_ (
);

AOI22X1 _3164_ (
    .A(DIMUX[5]),
    .B(_1319__bF$buf1),
    .C(_766_),
    .D(_761_),
    .Y(_767_)
);

FILL FILL_2__2857_ (
);

FILL FILL_2__2437_ (
);

FILL FILL_2__2017_ (
);

FILL FILL_7__1821_ (
);

FILL FILL_4__3304_ (
);

FILL FILL_0__3624_ (
);

FILL FILL_0__3204_ (
);

FILL FILL_7__2606_ (
);

FILL FILL_2__2190_ (
);

FILL FILL_3__2926_ (
);

FILL FILL_3__2506_ (
);

NOR2X1 _2855_ (
    .A(_1334_),
    .B(_1145_),
    .Y(_515_)
);

INVX1 _2435_ (
    .A(op[3]),
    .Y(_140_)
);

OAI21X1 _2015_ (
    .A(_1013_),
    .B(_983_),
    .C(_1126_),
    .Y(_1127_)
);

FILL FILL_5__2185_ (
);

FILL FILL_1__2597_ (
);

FILL FILL_7__3564_ (
);

FILL FILL_1__2177_ (
);

FILL FILL_3__3464_ (
);

FILL FILL_3__3044_ (
);

FILL FILL_2__1881_ (
);

FILL FILL_6__2674_ (
);

DFFSR _3393_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_62_),
    .CLK(clk_bF$buf6),
    .Q(V)
);

FILL FILL_6__2254_ (
);

FILL FILL_2__2666_ (
);

FILL FILL_2__2246_ (
);

FILL FILL168750x3750 (
);

FILL FILL_4__3533_ (
);

FILL FILL_4__3113_ (
);

FILL FILL_6__3459_ (
);

FILL FILL_6__3039_ (
);

FILL FILL_3__1950_ (
);

FILL FILL_0__3013_ (
);

FILL FILL_5__1876_ (
);

FILL FILL_1__1868_ (
);

FILL FILL_7__2835_ (
);

FILL FILL_3__2735_ (
);

FILL FILL_3__2315_ (
);

FILL FILL_5__3602_ (
);

FILL FILL_6__1945_ (
);

OAI21X1 _2664_ (
    .A(_1005_),
    .B(_330_),
    .C(_337_),
    .Y(_338_)
);

NAND3X1 _2244_ (
    .A(_1150__bF$buf3),
    .B(_1351_),
    .C(_1350_),
    .Y(_1352_)
);

FILL FILL_2__1937_ (
);

FILL FILL_4__2804_ (
);

OR2X2 _3449_ (
    .A(ADD[0]),
    .B(ADD[3]),
    .Y(_1698_)
);

OAI21X1 _3029_ (
    .A(_1008_),
    .B(_647_),
    .C(_650_),
    .Y(_55_)
);

FILL FILL_0__2704_ (
);

FILL FILL_3__3693_ (
);

FILL FILL_3__3273_ (
);

FILL FILL_5__3199_ (
);

FILL FILL_6__2483_ (
);

FILL FILL_6__2063_ (
);

FILL FILL_2__2895_ (
);

FILL FILL_2__2475_ (
);

FILL FILL_2__2055_ (
);

NAND3X1 _1935_ (
    .A(_1041_),
    .B(_1044_),
    .C(_1036_),
    .Y(_1052_)
);

FILL FILL_6__3268_ (
);

FILL FILL_0__3662_ (
);

FILL FILL_0__3242_ (
);

FILL FILL_7__2224_ (
);

FILL FILL_3__2964_ (
);

FILL FILL_3__2544_ (
);

FILL FILL_3__2124_ (
);

FILL FILL_7__3009_ (
);

FILL FILL_6__1754_ (
);

NAND2X1 _2893_ (
    .A(_543_),
    .B(_1251_),
    .Y(_544_)
);

OAI21X1 _2473_ (
    .A(_148_),
    .B(_1166_),
    .C(_171_),
    .Y(_172_)
);

INVX1 _2053_ (
    .A(IRHOLD[3]),
    .Y(_1162_)
);

FILL FILL_2__1746_ (
);

FILL FILL_4__2613_ (
);

FILL FILL_6__2959_ (
);

FILL FILL_6__2539_ (
);

OAI21X1 _3678_ (
    .A(RDY_bF$buf7),
    .B(_1703_),
    .C(_1697_),
    .Y(_1525_)
);

FILL FILL_6__2119_ (
);

NAND3X1 _3258_ (
    .A(_148_),
    .B(_1067_),
    .C(_833_),
    .Y(_834_)
);

FILL FILL_7__3182_ (
);

FILL FILL_0__2933_ (
);

FILL FILL_0__2513_ (
);

FILL FILL_3__3082_ (
);

FILL FILL_3__1815_ (
);

FILL FILL_6__2292_ (
);

FILL FILL_2__2284_ (
);

INVX1 _1744_ (
    .A(DIHOLD[0]),
    .Y(_878_)
);

FILL FILL_4__3571_ (
);

FILL FILL_4__3151_ (
);

FILL FILL_6__3497_ (
);

FILL FILL_6__3077_ (
);

FILL FILL_2__3489_ (
);

FILL FILL_0__3471_ (
);

FILL FILL_0__3051_ (
);

FILL FILL_2__3069_ (
);

AOI21X1 _2949_ (
    .A(_310_),
    .B(_1149__bF$buf2),
    .C(_585_),
    .Y(_37_)
);

OAI21X1 _2529_ (
    .A(_965_),
    .B(_218_),
    .C(_223_),
    .Y(_224_)
);

NAND2X1 _2109_ (
    .A(_1172_),
    .B(_1217_),
    .Y(_1218_)
);

FILL FILL_7__2453_ (
);

FILL FILL_3__2773_ (
);

FILL FILL_3__2353_ (
);

FILL FILL_5__2699_ (
);

FILL FILL_5__2279_ (
);

FILL FILL_7__3658_ (
);

FILL FILL_5__3640_ (
);

FILL FILL_5__3220_ (
);

FILL FILL_7__3238_ (
);

FILL FILL_1__3632_ (
);

FILL FILL_1__3212_ (
);

FILL FILL_3__3558_ (
);

FILL FILL_3__3138_ (
);

FILL FILL_6__1983_ (
);

NOR3X1 _2282_ (
    .A(_1369_),
    .B(_1372_),
    .C(_1389_),
    .Y(_1390_)
);

FILL FILL_2__1975_ (
);

FILL FILL_4__2842_ (
);

FILL FILL_4__2422_ (
);

FILL FILL_4__2002_ (
);

FILL FILL_6__2768_ (
);

NAND2X1 _3487_ (
    .A(CO),
    .B(_1714__bF$buf2),
    .Y(_1732_)
);

FILL FILL_6__2348_ (
);

OAI21X1 _3067_ (
    .A(_988_),
    .B(_679_),
    .C(_678_),
    .Y(_680_)
);

FILL FILL_0__2742_ (
);

FILL FILL_0__2322_ (
);

FILL FILL_2__3701_ (
);

FILL FILL_4__3627_ (
);

FILL FILL_4__3207_ (
);

FILL FILL_0__3527_ (
);

FILL FILL_0__3107_ (
);

FILL FILL_5__2911_ (
);

FILL FILL_7__2509_ (
);

FILL FILL_2__2093_ (
);

FILL FILL_1__2903_ (
);

FILL FILL_3__2829_ (
);

FILL FILL_3__2409_ (
);

NAND3X1 _1973_ (
    .A(_1088_),
    .B(_1086_),
    .C(_1087_),
    .Y(_1089_)
);

FILL FILL_2__3298_ (
);

FILL FILL_0__3280_ (
);

AOI21X1 _2758_ (
    .A(_417_),
    .B(_409_),
    .C(_423_),
    .Y(_424_)
);

OAI22X1 _2338_ (
    .A(RDY_bF$buf5),
    .B(_1444_),
    .C(_1149__bF$buf3),
    .D(_1398_),
    .Y(_1445_)
);

FILL FILL_7__2682_ (
);

FILL FILL_3__2582_ (
);

FILL FILL_3__2162_ (
);

FILL FILL_5__2088_ (
);

FILL FILL_7__3467_ (
);

FILL FILL_1__3021_ (
);

FILL FILL_6__1792_ (
);

INVX1 _2091_ (
    .A(_1199_),
    .Y(_1200_)
);

FILL FILL_2__1784_ (
);

FILL FILL169650x140550 (
);

FILL FILL_4__2651_ (
);

FILL FILL_4__2231_ (
);

FILL FILL_6__2997_ (
);

FILL FILL_6__2577_ (
);

OAI21X1 _3296_ (
    .A(_860_),
    .B(_257_),
    .C(_866_),
    .Y(_106_)
);

FILL FILL_6__2157_ (
);

FILL FILL_2__2989_ (
);

FILL FILL_0__2971_ (
);

FILL FILL_2__2569_ (
);

FILL FILL_0__2551_ (
);

FILL FILL_0__2131_ (
);

FILL FILL_2__2149_ (
);

FILL FILL_2__3510_ (
);

FILL FILL_7__1953_ (
);

FILL FILL_4__3016_ (
);

FILL FILL_3__1853_ (
);

FILL FILL_5__1779_ (
);

FILL FILL_7__2738_ (
);

FILL FILL_5__2720_ (
);

FILL FILL_5__2300_ (
);

FILL FILL_1__2712_ (
);

FILL FILL_3__2638_ (
);

FILL FILL_3__2218_ (
);

NOR2X1 _1782_ (
    .A(_904_),
    .B(_907_),
    .Y(_908_)
);

FILL FILL_5__3505_ (
);

FILL FILL_4__1922_ (
);

FILL FILL_6__1848_ (
);

AOI21X1 _2987_ (
    .A(_1161_),
    .B(_611_),
    .C(_616_),
    .Y(_617_)
);

AOI21X1 _2567_ (
    .A(_1124_),
    .B(_195_),
    .C(_256_),
    .Y(_257_)
);

AOI22X1 _2147_ (
    .A(_886__bF$buf1),
    .B(_967_),
    .C(_1255_),
    .D(_1150__bF$buf3),
    .Y(_1256_)
);

FILL FILL_7__2491_ (
);

FILL FILL_7__2071_ (
);

FILL FILL_0__1822_ (
);

FILL FILL_3__2391_ (
);

FILL FILL_4__2707_ (
);

FILL FILL_0__2607_ (
);

FILL FILL_1__3670_ (
);

FILL FILL_1__3250_ (
);

FILL FILL_3__3596_ (
);

FILL FILL_3__3176_ (
);

FILL FILL_3__1909_ (
);

FILL FILL_4__2880_ (
);

FILL FILL_4__2460_ (
);

FILL FILL_4__2040_ (
);

FILL FILL_6__2386_ (
);

FILL FILL_0__2780_ (
);

FILL FILL_2__2798_ (
);

FILL FILL_0__2360_ (
);

FILL FILL_2__2378_ (
);

AOI21X1 _1838_ (
    .A(_920_),
    .B(_923_),
    .C(_963_),
    .Y(_964_)
);

FILL FILL_4__3665_ (
);

FILL FILL_4__3245_ (
);

FILL FILL_0__3565_ (
);

FILL FILL_0__3145_ (
);

FILL FILL_4_BUFX2_insert50 (
);

FILL FILL_4_BUFX2_insert51 (
);

FILL FILL_4_BUFX2_insert52 (
);

FILL FILL_4_BUFX2_insert53 (
);

FILL FILL_4_BUFX2_insert54 (
);

FILL FILL_4_BUFX2_insert55 (
);

FILL FILL_4_BUFX2_insert56 (
);

FILL FILL_4_BUFX2_insert57 (
);

FILL FILL_4_BUFX2_insert58 (
);

FILL FILL_4_BUFX2_insert59 (
);

FILL FILL_7__2967_ (
);

FILL FILL_7__2127_ (
);

FILL FILL_1__2941_ (
);

FILL FILL_1__2521_ (
);

FILL FILL_1__2101_ (
);

FILL FILL_3__2867_ (
);

FILL FILL_3__2447_ (
);

FILL FILL_3__2027_ (
);

FILL FILL_5__3314_ (
);

FILL FILL_1__3306_ (
);

OAI21X1 _2796_ (
    .A(_290_),
    .B(_313_),
    .C(_1118_),
    .Y(_459_)
);

NAND3X1 _2376_ (
    .A(_1474_),
    .B(_1480_),
    .C(_1481_),
    .Y(_1482_)
);

FILL FILL_4__2936_ (
);

FILL FILL_4__2516_ (
);

FILL FILL_7__3085_ (
);

FILL FILL_0__2836_ (
);

FILL FILL_0__2416_ (
);

FILL FILL_7__1818_ (
);

FILL FILL_5__1800_ (
);

FILL FILL_6__2195_ (
);

FILL FILL_2__2187_ (
);

FILL FILL_4__3474_ (
);

FILL FILL_4__3054_ (
);

FILL FILL_3__1891_ (
);

FILL FILL_7__2356_ (
);

FILL FILL_1__2750_ (
);

FILL FILL_1__2330_ (
);

FILL FILL_3__2676_ (
);

FILL FILL_3__2256_ (
);

FILL FILL_5__3543_ (
);

FILL FILL_5__3123_ (
);

FILL FILL_1__3535_ (
);

FILL FILL_1__3115_ (
);

FILL FILL_4__1960_ (
);

FILL FILL_6__1886_ (
);

NOR2X1 _2185_ (
    .A(_1289_),
    .B(_1293_),
    .Y(_1294_)
);

FILL FILL_0__1860_ (
);

FILL FILL_2__1878_ (
);

FILL FILL_4__2745_ (
);

FILL FILL_4__2325_ (
);

FILL FILL_0__2645_ (
);

FILL FILL_6__3612_ (
);

FILL FILL_0__2225_ (
);

FILL FILL_2__3604_ (
);

FILL FILL_6_CLKBUF1_insert30 (
);

FILL FILL_6_CLKBUF1_insert31 (
);

FILL FILL_6_CLKBUF1_insert32 (
);

FILL FILL_3__1947_ (
);

FILL FILL_6_CLKBUF1_insert33 (
);

FILL FILL_6_CLKBUF1_insert34 (
);

FILL FILL_6_CLKBUF1_insert35 (
);

FILL FILL_6_CLKBUF1_insert36 (
);

FILL FILL_5__2814_ (
);

FILL FILL_1__2806_ (
);

INVX1 _1876_ (
    .A(_1000_),
    .Y(_1001_)
);

FILL FILL_4__3283_ (
);

FILL FILL_0__3183_ (
);

FILL FILL_7__2585_ (
);

FILL FILL_0__1916_ (
);

OAI21X1 _3602_ (
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1527_),
    .Y(_1632_)
);

FILL FILL_3__2485_ (
);

FILL FILL_3__2065_ (
);

FILL FILL_4__2974_ (
);

FILL FILL_4__2554_ (
);

FILL FILL_4__2134_ (
);

OAI21X1 _3199_ (
    .A(_757_),
    .B(_789_),
    .C(_794_),
    .Y(_81_)
);

FILL FILL_0__2874_ (
);

FILL FILL_0__2454_ (
);

FILL FILL_0__2034_ (
);

FILL FILL_6__3001_ (
);

FILL FILL_7__1856_ (
);

FILL FILL_1__1830_ (
);

FILL FILL_0__3659_ (
);

FILL FILL_3__1756_ (
);

FILL FILL_0__3239_ (
);

FILL FILL_5__2623_ (
);

FILL FILL_5__2203_ (
);

FILL FILL_1__2615_ (
);

FILL FILL_4__3092_ (
);

FILL FILL_4__1825_ (
);

DFFSR _3411_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_80_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[1] [3])
);

FILL FILL_3__2294_ (
);

FILL FILL_5__3581_ (
);

FILL FILL_5__3161_ (
);

FILL FILL_1__3573_ (
);

FILL FILL_1__3153_ (
);

FILL FILL_3__3499_ (
);

FILL FILL_3__3079_ (
);

FILL FILL_4__2783_ (
);

FILL FILL_4__2363_ (
);

FILL FILL_6__2289_ (
);

FILL FILL_0__2683_ (
);

FILL FILL_6__3650_ (
);

FILL FILL_0__2263_ (
);

FILL FILL_6__3230_ (
);

FILL FILL_2__3642_ (
);

FILL FILL_2__3222_ (
);

FILL FILL_4__3568_ (
);

FILL FILL_4__3148_ (
);

FILL FILL_3__1985_ (
);

FILL FILL_0__3468_ (
);

FILL FILL_0__3048_ (
);

FILL FILL_5__2852_ (
);

FILL FILL_5__2432_ (
);

FILL FILL_5__2012_ (
);

FILL FILL_1__2844_ (
);

FILL FILL_1__2424_ (
);

FILL FILL_1__2004_ (
);

FILL FILL_3__3711_ (
);

FILL FILL_5__3637_ (
);

FILL FILL_5__3217_ (
);

FILL FILL_1__3629_ (
);

FILL FILL_1__3209_ (
);

NAND3X1 _2699_ (
    .A(_338_),
    .B(_369_),
    .C(_333_),
    .Y(_370_)
);

OAI21X1 _2279_ (
    .A(RDY_bF$buf2),
    .B(_953_),
    .C(_1386_),
    .Y(_1387_)
);

FILL FILL_0__1954_ (
);

FILL FILL_6__2921_ (
);

INVX1 _3640_ (
    .A(_1629_),
    .Y(_1670_)
);

FILL FILL_6__2501_ (
);

AOI21X1 _3220_ (
    .A(_778_),
    .B(_798_),
    .C(_805_),
    .Y(_91_)
);

FILL FILL_2__2913_ (
);

FILL FILL_4__2839_ (
);

FILL FILL_4__2419_ (
);

FILL FILL_0__2739_ (
);

FILL FILL_6__3706_ (
);

FILL FILL_0__2319_ (
);

FILL FILL_4__2592_ (
);

FILL FILL_4__2172_ (
);

FILL FILL_6__2098_ (
);

FILL FILL_5__2908_ (
);

FILL FILL_0__2492_ (
);

FILL FILL_0__2072_ (
);

FILL FILL_2__3451_ (
);

FILL FILL_2__3031_ (
);

INVX1 _2911_ (
    .A(_556_),
    .Y(_557_)
);

FILL FILL_0__3697_ (
);

FILL FILL_3__1794_ (
);

FILL FILL_0__3277_ (
);

FILL FILL_7__2679_ (
);

FILL FILL_5__2661_ (
);

FILL FILL_7__2259_ (
);

FILL FILL_5__2241_ (
);

FILL FILL_1__2653_ (
);

FILL FILL_1__2233_ (
);

FILL FILL_3__2999_ (
);

BUFX2 BUFX2_insert0 (
    .A(RDY),
    .Y(RDY_bF$buf9)
);

FILL FILL_3__2579_ (
);

FILL FILL_3__2159_ (
);

BUFX2 BUFX2_insert1 (
    .A(RDY),
    .Y(RDY_bF$buf8)
);

BUFX2 BUFX2_insert2 (
    .A(RDY),
    .Y(RDY_bF$buf7)
);

BUFX2 BUFX2_insert3 (
    .A(RDY),
    .Y(RDY_bF$buf6)
);

BUFX2 BUFX2_insert4 (
    .A(RDY),
    .Y(RDY_bF$buf5)
);

BUFX2 BUFX2_insert5 (
    .A(RDY),
    .Y(RDY_bF$buf4)
);

BUFX2 BUFX2_insert6 (
    .A(RDY),
    .Y(RDY_bF$buf3)
);

BUFX2 BUFX2_insert7 (
    .A(RDY),
    .Y(RDY_bF$buf2)
);

BUFX2 BUFX2_insert8 (
    .A(RDY),
    .Y(RDY_bF$buf1)
);

BUFX2 BUFX2_insert9 (
    .A(RDY),
    .Y(RDY_bF$buf0)
);

FILL FILL_3__3520_ (
);

FILL FILL_3__3100_ (
);

FILL FILL_5__3026_ (
);

FILL FILL_1__3018_ (
);

FILL FILL_4__1863_ (
);

FILL FILL_6__1789_ (
);

OAI21X1 _2088_ (
    .A(RDY_bF$buf8),
    .B(_1196_),
    .C(_1195_),
    .Y(_1197_)
);

FILL FILL_0__1763_ (
);

FILL FILL_6__2730_ (
);

FILL FILL_6__2310_ (
);

FILL FILL_2__2722_ (
);

FILL FILL_2__2302_ (
);

FILL FILL_4__2648_ (
);

FILL FILL_4__2228_ (
);

FILL FILL_0__2968_ (
);

FILL FILL_0__2548_ (
);

FILL FILL_6__3515_ (
);

FILL FILL_0__2128_ (
);

FILL FILL_1__3191_ (
);

FILL FILL_2__3507_ (
);

FILL FILL_5__1932_ (
);

FILL FILL_1__1924_ (
);

FILL FILL_5__2717_ (
);

FILL FILL_1__2709_ (
);

FILL FILL_2__3260_ (
);

INVX1 _1779_ (
    .A(state[1]),
    .Y(_905_)
);

FILL FILL_4__3186_ (
);

INVX1 _2720_ (
    .A(ABL[6]),
    .Y(_389_)
);

OAI21X1 _2300_ (
    .A(_1405_),
    .B(_1395_),
    .C(_1406_),
    .Y(_1407_)
);

FILL FILL_0__3086_ (
);

FILL FILL_4__1919_ (
);

FILL FILL_5__2890_ (
);

FILL FILL_7__2488_ (
);

FILL FILL_5__2470_ (
);

FILL FILL_5__2050_ (
);

FILL FILL_0__1819_ (
);

OAI21X1 _3505_ (
    .A(BI[4]),
    .B(_1739_),
    .C(_1534_),
    .Y(_1535_)
);

FILL FILL_1__2882_ (
);

FILL FILL_1__2462_ (
);

FILL FILL_1__2042_ (
);

FILL FILL_3__2388_ (
);

FILL FILL_5__3675_ (
);

FILL FILL_5__3255_ (
);

FILL FILL_1__3667_ (
);

FILL FILL_1__3247_ (
);

FILL FILL_0__1992_ (
);

FILL FILL_2__2951_ (
);

FILL FILL_2__2531_ (
);

FILL FILL_2__2111_ (
);

FILL FILL_4__2877_ (
);

FILL FILL_4__2457_ (
);

FILL FILL_4__2037_ (
);

FILL FILL_0__2777_ (
);

FILL FILL_0__2357_ (
);

FILL FILL_2__3316_ (
);

FILL FILL_7__1759_ (
);

FILL FILL_3__2600_ (
);

FILL FILL_5__2946_ (
);

FILL FILL_5__2526_ (
);

FILL FILL_5__2106_ (
);

FILL FILL_1__2938_ (
);

FILL FILL_1__2518_ (
);

FILL FILL_6__1810_ (
);

FILL FILL_2__1802_ (
);

NAND2X1 _3314_ (
    .A(_1741_[14]),
    .B(_869_),
    .Y(_876_)
);

FILL FILL_1__2691_ (
);

FILL FILL_1__2271_ (
);

FILL FILL_3__2197_ (
);

FILL FILL_5__3484_ (
);

FILL FILL_5__3064_ (
);

FILL FILL_1__3476_ (
);

FILL FILL_1__3056_ (
);

FILL FILL_2__2760_ (
);

FILL FILL_2__2340_ (
);

FILL FILL_4__2686_ (
);

FILL FILL_4__2266_ (
);

NOR2X1 _1800_ (
    .A(state[3]),
    .B(_896_),
    .Y(_926_)
);

FILL FILL_0__2586_ (
);

FILL FILL_6__3553_ (
);

FILL FILL_0__2166_ (
);

FILL FILL_6__3133_ (
);

FILL FILL169950x43350 (
);

FILL FILL_2__3545_ (
);

FILL FILL_2__3125_ (
);

FILL FILL_7__1988_ (
);

FILL FILL_5__1970_ (
);

FILL FILL_1__1962_ (
);

FILL FILL_3__1888_ (
);

FILL FILL_5__2755_ (
);

FILL FILL_5__2335_ (
);

FILL FILL_1__2747_ (
);

FILL FILL_1__2327_ (
);

FILL FILL_3__3614_ (
);

FILL FILL_4__1957_ (
);

FILL FILL_0__1857_ (
);

FILL FILL_6__2824_ (
);

NAND2X1 _3543_ (
    .A(alu_op[1]),
    .B(AI[0]),
    .Y(_1573_)
);

FILL FILL_6__2404_ (
);

INVX1 _3123_ (
    .A(_727_),
    .Y(_730_)
);

FILL FILL_1__2080_ (
);

FILL FILL_2__2816_ (
);

FILL FILL_5__3293_ (
);

FILL FILL_6__3609_ (
);

FILL FILL_1__3285_ (
);

FILL FILL_4__2495_ (
);

FILL FILL_4__2075_ (
);

FILL FILL_0__2395_ (
);

FILL FILL_7__1797_ (
);

NAND3X1 _2814_ (
    .A(_472_),
    .B(_476_),
    .C(_475_),
    .Y(_477_)
);

FILL FILL_1__1771_ (
);

FILL FILL_5__2984_ (
);

FILL FILL_5__2564_ (
);

FILL FILL_5__2144_ (
);

FILL FILL_1__2976_ (
);

FILL FILL_1__2556_ (
);

FILL FILL_1__2136_ (
);

FILL FILL_7__3103_ (
);

FILL FILL_3__3003_ (
);

FILL FILL_2__1840_ (
);

FILL FILL_4__1766_ (
);

FILL FILL_6__2633_ (
);

DFFSR _3352_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_29_),
    .CLK(clk_bF$buf9),
    .Q(sei)
);

FILL FILL_6__2213_ (
);

FILL FILL_2__2625_ (
);

FILL FILL_2__2205_ (
);

FILL FILL_1__3094_ (
);

FILL FILL_5__1835_ (
);

FILL FILL_1__1827_ (
);

FILL FILL_6__3591_ (
);

FILL FILL_6__3171_ (
);

FILL FILL_2__3583_ (
);

FILL FILL_2__3163_ (
);

FILL FILL_4__3089_ (
);

FILL FILL_6__1904_ (
);

OAI21X1 _2623_ (
    .A(_300_),
    .B(_218_),
    .C(_303_),
    .Y(_1741_[14])
);

NAND3X1 _2203_ (
    .A(_1308_),
    .B(_1306_),
    .C(_1311_),
    .Y(_1312_)
);

FILL FILL_5__2793_ (
);

FILL FILL_5__2373_ (
);

DFFSR _3408_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_77_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[1] [0])
);

FILL FILL_1__2785_ (
);

FILL FILL_1__2365_ (
);

FILL FILL_3__3652_ (
);

FILL FILL_3__3232_ (
);

FILL FILL_5__3578_ (
);

FILL FILL_5__3158_ (
);

FILL FILL_4__1995_ (
);

FILL FILL_0__1895_ (
);

FILL FILL_6__2862_ (
);

OAI21X1 _3581_ (
    .A(_1728_),
    .B(_1610_),
    .C(_1580_),
    .Y(_1611_)
);

FILL FILL_6__2442_ (
);

FILL FILL_6__2022_ (
);

OAI21X1 _3161_ (
    .A(_763_),
    .B(_762_),
    .C(ADD[5]),
    .Y(_764_)
);

FILL FILL_2__2854_ (
);

FILL FILL_2__2434_ (
);

FILL FILL_2__2014_ (
);

FILL FILL_4__3301_ (
);

FILL FILL_6__3647_ (
);

FILL FILL_6__3227_ (
);

FILL FILL_2__3639_ (
);

FILL FILL_0__3621_ (
);

FILL FILL_0__3201_ (
);

FILL FILL_2__3219_ (
);

FILL FILL_7__2603_ (
);

FILL FILL_3__2923_ (
);

FILL FILL_3__2503_ (
);

FILL FILL_5__2849_ (
);

FILL FILL_5__2429_ (
);

FILL FILL_5__2009_ (
);

FILL FILL_3__3708_ (
);

AND2X2 _2852_ (
    .A(_511_),
    .B(_512_),
    .Y(_16_)
);

NOR2X1 _2432_ (
    .A(_135_),
    .B(_137_),
    .Y(_138_)
);

NAND3X1 _2012_ (
    .A(_1123_),
    .B(_1121_),
    .C(_1122_),
    .Y(_1124_)
);

FILL FILL_5__2182_ (
);

FILL FILL_6__2918_ (
);

NAND2X1 _3637_ (
    .A(\u_ALU8.BCD ),
    .B(_1666_),
    .Y(_1667_)
);

NOR2X1 _3217_ (
    .A(\AXYS[2] [5]),
    .B(_798_),
    .Y(_804_)
);

FILL FILL_1__2594_ (
);

FILL FILL_7__3561_ (
);

FILL FILL_1__2174_ (
);

FILL FILL_7__3141_ (
);

FILL FILL_3__3461_ (
);

FILL FILL_3__3041_ (
);

FILL FILL_6__2671_ (
);

DFFPOSX1 _3390_ (
    .D(_59_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD[6])
);

FILL FILL_6__2251_ (
);

FILL FILL_2__2663_ (
);

FILL FILL_2__2243_ (
);

FILL FILL_4__2589_ (
);

FILL FILL_4__2169_ (
);

FILL FILL_4__3530_ (
);

FILL FILL_4__3110_ (
);

FILL FILL_0__2489_ (
);

FILL FILL_6__3456_ (
);

FILL FILL_0__2069_ (
);

FILL FILL_6__3036_ (
);

FILL FILL_2__3028_ (
);

FILL FILL_0__3010_ (
);

FILL FILL_5__1873_ (
);

NAND3X1 _2908_ (
    .A(_1327_),
    .B(_1178_),
    .C(_1161_),
    .Y(_554_)
);

FILL FILL_1__1865_ (
);

FILL FILL_7__2832_ (
);

FILL FILL_7__2412_ (
);

FILL FILL_3__2732_ (
);

FILL FILL_3__2312_ (
);

FILL FILL_5__2658_ (
);

FILL FILL_5__2238_ (
);

FILL FILL_7__3617_ (
);

FILL FILL_3__3517_ (
);

FILL FILL_6__1942_ (
);

NAND2X1 _2661_ (
    .A(ABL[1]),
    .B(_323_),
    .Y(_335_)
);

NAND2X1 _2241_ (
    .A(_1178_),
    .B(_1348_),
    .Y(_1349_)
);

FILL FILL_2__1934_ (
);

FILL FILL_4__2801_ (
);

FILL FILL_6__2727_ (
);

DFFSR _3446_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_114_),
    .CLK(clk_bF$buf0),
    .Q(ABH[5])
);

FILL FILL_6__2307_ (
);

OAI21X1 _3026_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[1]),
    .Y(_649_)
);

FILL FILL_2__2719_ (
);

FILL FILL_0__2701_ (
);

FILL FILL_3__3270_ (
);

FILL FILL_5__3196_ (
);

FILL FILL_1__3188_ (
);

FILL FILL_5__1929_ (
);

FILL FILL_6__2480_ (
);

FILL FILL_6__2060_ (
);

FILL FILL_2__2892_ (
);

FILL FILL_2__2472_ (
);

FILL FILL_2__2052_ (
);

FILL FILL_4__2398_ (
);

AOI22X1 _1932_ (
    .A(_1048_),
    .B(_1039_),
    .C(_1045_),
    .D(_1046_),
    .Y(_1049_)
);

FILL FILL_0__2298_ (
);

FILL FILL_6__3265_ (
);

FILL FILL_2__3677_ (
);

FILL FILL_2__3257_ (
);

INVX1 _2717_ (
    .A(_386_),
    .Y(_387_)
);

FILL FILL_7__2641_ (
);

FILL FILL_7__2221_ (
);

FILL FILL_3__2961_ (
);

FILL FILL_3__2541_ (
);

FILL FILL_3__2121_ (
);

FILL FILL_5__2887_ (
);

FILL FILL_5__2467_ (
);

FILL FILL_5__2047_ (
);

FILL FILL_1__2879_ (
);

FILL FILL_1__2459_ (
);

FILL FILL_1__2039_ (
);

FILL FILL_7__3006_ (
);

FILL FILL_6__1751_ (
);

OAI22X1 _2890_ (
    .A(_539_),
    .B(_1150__bF$buf2),
    .C(_541_),
    .D(_538_),
    .Y(_25_)
);

INVX1 _2470_ (
    .A(_169_),
    .Y(_170_)
);

OAI21X1 _2050_ (
    .A(IRHOLD_valid),
    .B(DIMUX[0]),
    .C(_1158_),
    .Y(_1159_)
);

FILL FILL_4__2610_ (
);

FILL FILL_0__1989_ (
);

FILL FILL_6__2956_ (
);

NAND2X1 _3675_ (
    .A(RDY_bF$buf7),
    .B(_1675_),
    .Y(_1696_)
);

FILL FILL_6__2536_ (
);

FILL FILL_6__2116_ (
);

AOI22X1 _3255_ (
    .A(_1303_),
    .B(_822_),
    .C(_828_),
    .D(_830_),
    .Y(_831_)
);

FILL FILL_2__2948_ (
);

FILL FILL_0__2930_ (
);

FILL FILL_2__2528_ (
);

FILL FILL_0__2510_ (
);

FILL FILL_2__2108_ (
);

FILL FILL_0__3715_ (
);

FILL FILL_3__1812_ (
);

FILL FILL_2__2281_ (
);

FILL FILL_6__3494_ (
);

FILL FILL_6__3074_ (
);

FILL FILL_0_BUFX2_insert70 (
);

FILL FILL_0_BUFX2_insert71 (
);

FILL FILL_2__3486_ (
);

FILL FILL_0_BUFX2_insert72 (
);

FILL FILL_2__3066_ (
);

FILL FILL_0_BUFX2_insert73 (
);

FILL FILL_0_BUFX2_insert74 (
);

FILL FILL_0_BUFX2_insert75 (
);

FILL FILL_0_BUFX2_insert76 (
);

FILL FILL_0_BUFX2_insert77 (
);

FILL FILL_0_BUFX2_insert78 (
);

FILL FILL_0_BUFX2_insert79 (
);

OAI21X1 _2946_ (
    .A(_140_),
    .B(_1150__bF$buf1),
    .C(_587_),
    .Y(_35_)
);

FILL FILL_6__1807_ (
);

OAI21X1 _2526_ (
    .A(_966_),
    .B(_201_),
    .C(_220_),
    .Y(_221_)
);

NAND2X1 _2106_ (
    .A(_1156_),
    .B(_1214_),
    .Y(_1215_)
);

FILL FILL_7__2870_ (
);

FILL FILL_7__2450_ (
);

FILL FILL_7__2030_ (
);

FILL FILL_3__2770_ (
);

FILL FILL_3__2350_ (
);

FILL FILL_5__2696_ (
);

FILL FILL_5__2276_ (
);

FILL FILL_1__2688_ (
);

FILL FILL_1__2268_ (
);

FILL FILL_7__3235_ (
);

FILL FILL_3__3555_ (
);

FILL FILL_3__3135_ (
);

FILL FILL_6__1980_ (
);

FILL FILL_2__1972_ (
);

FILL FILL_4__1898_ (
);

FILL FILL_0__1798_ (
);

FILL FILL_6__2765_ (
);

OAI21X1 _3484_ (
    .A(_1727_),
    .B(_1724_),
    .C(_1729_),
    .Y(_1730_)
);

FILL FILL_6__2345_ (
);

NOR2X1 _3064_ (
    .A(cli),
    .B(_1444_),
    .Y(_677_)
);

FILL FILL_2__2757_ (
);

FILL FILL_2__2337_ (
);

FILL FILL_4__3624_ (
);

FILL FILL_4__3204_ (
);

FILL FILL_0__3524_ (
);

FILL FILL_0__3104_ (
);

FILL FILL_5__1967_ (
);

FILL FILL_1__1959_ (
);

FILL FILL_7__2506_ (
);

FILL FILL_2__2090_ (
);

FILL FILL_1__2900_ (
);

FILL FILL_3__2826_ (
);

FILL FILL_3__2406_ (
);

NAND2X1 _1970_ (
    .A(\AXYS[1] [1]),
    .B(_1047_),
    .Y(_1086_)
);

FILL FILL_2__3295_ (
);

NAND3X1 _2755_ (
    .A(_148_),
    .B(_420_),
    .C(_1094_),
    .Y(_421_)
);

OAI21X1 _2335_ (
    .A(_1401_),
    .B(_1422_),
    .C(_1441_),
    .Y(_1442_)
);

FILL FILL_5__2085_ (
);

FILL FILL_1__2497_ (
);

FILL FILL_7__3464_ (
);

FILL FILL_1__2077_ (
);

FILL FILL_2__1781_ (
);

FILL FILL_6__2994_ (
);

FILL FILL_6__2574_ (
);

NAND2X1 _3293_ (
    .A(ABL[4]),
    .B(_860_),
    .Y(_865_)
);

FILL FILL_6__2154_ (
);

FILL FILL_2__2986_ (
);

FILL FILL_2__2566_ (
);

FILL FILL_2__2146_ (
);

FILL FILL_7__1950_ (
);

FILL FILL_4__3013_ (
);

FILL FILL_3__1850_ (
);

FILL FILL_5__1776_ (
);

FILL FILL_1__1768_ (
);

FILL FILL_7__2735_ (
);

FILL FILL_3__2635_ (
);

FILL FILL_3__2215_ (
);

FILL FILL_5__3502_ (
);

FILL FILL_6__1845_ (
);

NOR2X1 _2984_ (
    .A(_613_),
    .B(_530_),
    .Y(_614_)
);

NAND2X1 _2564_ (
    .A(_253_),
    .B(_250_),
    .Y(_254_)
);

INVX1 _2144_ (
    .A(_1252_),
    .Y(_1253_)
);

FILL FILL_2__1837_ (
);

FILL FILL_4__2704_ (
);

DFFSR _3349_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_26_),
    .CLK(clk_bF$buf9),
    .Q(cld)
);

FILL FILL_7__3273_ (
);

FILL FILL_0__2604_ (
);

FILL FILL_3__3593_ (
);

FILL FILL_3__3173_ (
);

FILL FILL_5__3099_ (
);

FILL FILL_3__1906_ (
);

FILL FILL_6__2383_ (
);

FILL FILL_2__2795_ (
);

FILL FILL_2__2375_ (
);

NAND3X1 _1835_ (
    .A(_953_),
    .B(_951_),
    .C(_960_),
    .Y(_961_)
);

FILL FILL_4__3662_ (
);

FILL FILL_4__3242_ (
);

FILL FILL_6__3588_ (
);

FILL FILL_6__3168_ (
);

FILL FILL_0__3562_ (
);

FILL FILL_0__3142_ (
);

FILL FILL_4_BUFX2_insert20 (
);

FILL FILL_4_BUFX2_insert21 (
);

FILL FILL_4_BUFX2_insert22 (
);

FILL FILL_4_BUFX2_insert23 (
);

FILL FILL_4_BUFX2_insert24 (
);

FILL FILL_4_BUFX2_insert25 (
);

FILL FILL_1__1997_ (
);

FILL FILL_7__2964_ (
);

FILL FILL_7__2124_ (
);

FILL FILL_3__2864_ (
);

FILL FILL_3__2444_ (
);

FILL FILL_3__2024_ (
);

FILL FILL_5__3311_ (
);

BUFX2 BUFX2_insert80 (
    .A(_1319_),
    .Y(_1319__bF$buf3)
);

BUFX2 BUFX2_insert81 (
    .A(_1319_),
    .Y(_1319__bF$buf2)
);

BUFX2 BUFX2_insert82 (
    .A(_1319_),
    .Y(_1319__bF$buf1)
);

BUFX2 BUFX2_insert83 (
    .A(_1319_),
    .Y(_1319__bF$buf0)
);

FILL FILL_1__3303_ (
);

FILL FILL_3__3649_ (
);

FILL FILL_3__3229_ (
);

OAI21X1 _2793_ (
    .A(_456_),
    .B(_401_),
    .C(RDY_bF$buf4),
    .Y(_457_)
);

NAND3X1 _2373_ (
    .A(_1475_),
    .B(_1478_),
    .C(_1476_),
    .Y(_1479_)
);

FILL FILL_4__2933_ (
);

FILL FILL_4__2513_ (
);

FILL FILL_6__2859_ (
);

INVX1 _3578_ (
    .A(\u_ALU8.BCD ),
    .Y(_1608_)
);

FILL FILL_6__2439_ (
);

OR2X2 _3158_ (
    .A(_760_),
    .B(ADD[5]),
    .Y(_761_)
);

FILL FILL_6__2019_ (
);

FILL FILL_7__3082_ (
);

FILL FILL_0__2833_ (
);

FILL FILL_0__2413_ (
);

FILL FILL_0__3618_ (
);

FILL FILL_6__2192_ (
);

FILL FILL_2__2184_ (
);

FILL FILL_4__3471_ (
);

FILL FILL_4__3051_ (
);

OAI21X1 _2849_ (
    .A(_508_),
    .B(_485_),
    .C(_509_),
    .Y(_510_)
);

INVX1 _2429_ (
    .A(_134_),
    .Y(_135_)
);

NAND2X1 _2009_ (
    .A(\AXYS[1] [5]),
    .B(_1047_),
    .Y(_1121_)
);

FILL FILL_7__2353_ (
);

FILL FILL_3__2673_ (
);

FILL FILL_3__2253_ (
);

FILL FILL_5__2599_ (
);

FILL FILL_5__2179_ (
);

FILL FILL_5__3540_ (
);

FILL FILL_7__3558_ (
);

FILL FILL_5__3120_ (
);

FILL FILL_7__3138_ (
);

FILL FILL_1__3532_ (
);

FILL FILL_1__3112_ (
);

FILL FILL_3__3458_ (
);

FILL FILL_3__3038_ (
);

FILL FILL_6__1883_ (
);

NOR2X1 _2182_ (
    .A(_931__bF$buf2),
    .B(_954_),
    .Y(_1291_)
);

FILL FILL_2__1875_ (
);

FILL FILL_4__2742_ (
);

FILL FILL_4__2322_ (
);

FILL FILL_6__2668_ (
);

DFFPOSX1 _3387_ (
    .D(_56_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD[3])
);

FILL FILL_6__2248_ (
);

FILL FILL_0__2642_ (
);

FILL FILL_0__2222_ (
);

FILL FILL_2__3601_ (
);

FILL FILL_4__3527_ (
);

FILL FILL_4__3107_ (
);

FILL FILL_3__1944_ (
);

FILL FILL_0__3007_ (
);

FILL FILL_5__2811_ (
);

FILL FILL_7__2409_ (
);

FILL FILL169950x140550 (
);

FILL FILL_1__2803_ (
);

FILL FILL_3__2729_ (
);

FILL FILL_3__2309_ (
);

INVX1 _1873_ (
    .A(_940_),
    .Y(_998_)
);

FILL FILL_4__3280_ (
);

FILL FILL_0__3180_ (
);

FILL FILL_2__3198_ (
);

FILL FILL_6__1939_ (
);

AND2X2 _2658_ (
    .A(_331_),
    .B(_320_),
    .Y(_333_)
);

NAND3X1 _2238_ (
    .A(_1229_),
    .B(_1345_),
    .C(_1231_),
    .Y(_1346_)
);

FILL FILL_7__2582_ (
);

FILL FILL_0__1913_ (
);

FILL FILL_3__2482_ (
);

FILL FILL_3__2062_ (
);

FILL FILL_3__3267_ (
);

FILL FILL_4__2971_ (
);

FILL FILL_4__2551_ (
);

FILL FILL_4__2131_ (
);

FILL FILL_6__2897_ (
);

FILL FILL_6__2477_ (
);

FILL FILL_6__2057_ (
);

OAI21X1 _3196_ (
    .A(_720__bF$buf2),
    .B(_687_),
    .C(\AXYS[1] [3]),
    .Y(_793_)
);

FILL FILL_0__2871_ (
);

FILL FILL_2__2889_ (
);

FILL FILL_0__2451_ (
);

FILL FILL_2__2469_ (
);

FILL FILL_0__2031_ (
);

FILL FILL_2__2049_ (
);

NAND3X1 _1929_ (
    .A(src_reg[0]),
    .B(_1035_),
    .C(_1026_),
    .Y(_1046_)
);

FILL FILL_7__1853_ (
);

FILL FILL_3__1753_ (
);

FILL FILL_0__3656_ (
);

FILL FILL_0__3236_ (
);

FILL FILL_7__2638_ (
);

FILL FILL_5__2620_ (
);

FILL FILL_5__2200_ (
);

FILL FILL_1__2612_ (
);

FILL FILL_3__2958_ (
);

FILL FILL_3__2538_ (
);

FILL FILL_3__2118_ (
);

FILL FILL_4__1822_ (
);

FILL FILL_6__1748_ (
);

INVX1 _2887_ (
    .A(sec),
    .Y(_539_)
);

OAI21X1 _2467_ (
    .A(_1009_),
    .B(_136_),
    .C(_166_),
    .Y(_167_)
);

OAI21X1 _2047_ (
    .A(IRHOLD_valid),
    .B(DIMUX[1]),
    .C(_1155_),
    .Y(_1156_)
);

FILL FILL_3__2291_ (
);

FILL FILL_4__2607_ (
);

FILL FILL_7__3596_ (
);

FILL FILL_0__2927_ (
);

FILL FILL_0__2507_ (
);

FILL FILL_1__3570_ (
);

FILL FILL_1__3150_ (
);

FILL FILL_3__3496_ (
);

FILL FILL_3__3076_ (
);

FILL FILL_7__1909_ (
);

FILL FILL_3__1809_ (
);

FILL FILL_4__2780_ (
);

FILL FILL_4__2360_ (
);

FILL FILL_6__2286_ (
);

FILL FILL_2__2698_ (
);

FILL FILL_0__2680_ (
);

FILL FILL_2__2278_ (
);

FILL FILL_0__2260_ (
);

FILL FILL_4__3565_ (
);

FILL FILL_4__3145_ (
);

FILL FILL_3__1982_ (
);

FILL FILL_0__3465_ (
);

FILL FILL_0__3045_ (
);

FILL FILL_7__2867_ (
);

FILL FILL_7__2027_ (
);

FILL FILL_1__2841_ (
);

FILL FILL_1__2421_ (
);

FILL FILL_1__2001_ (
);

FILL FILL_3__2767_ (
);

FILL FILL_3__2347_ (
);

FILL FILL_5__3634_ (
);

FILL FILL_5__3214_ (
);

FILL FILL_1__3626_ (
);

FILL FILL_1__3206_ (
);

FILL FILL_6__1977_ (
);

OAI21X1 _2696_ (
    .A(_329_),
    .B(_365_),
    .C(PC[3]),
    .Y(_367_)
);

NOR2X1 _2276_ (
    .A(_886__bF$buf4),
    .B(_968_),
    .Y(_1384_)
);

FILL FILL_2__1969_ (
);

FILL FILL_0__1951_ (
);

FILL FILL_2__2910_ (
);

FILL FILL_4__2836_ (
);

FILL FILL_4__2416_ (
);

FILL FILL_0__2736_ (
);

FILL FILL_0__2316_ (
);

FILL FILL_6__3703_ (
);

FILL FILL_6__2095_ (
);

FILL FILL_5__2905_ (
);

FILL FILL_2__2087_ (
);

OAI21X1 _1967_ (
    .A(_966_),
    .B(_983_),
    .C(_1083_),
    .Y(_1084_)
);

FILL FILL_0__3694_ (
);

FILL FILL_3__1791_ (
);

FILL FILL_0__3274_ (
);

FILL FILL_7__2256_ (
);

FILL FILL_1__2650_ (
);

FILL FILL_1__2230_ (
);

FILL FILL_3__2996_ (
);

FILL FILL_3__2576_ (
);

FILL FILL_3__2156_ (
);

FILL FILL_5__3023_ (
);

FILL FILL_1__3015_ (
);

FILL FILL_4__1860_ (
);

FILL FILL_6__1786_ (
);

OAI21X1 _2085_ (
    .A(CO),
    .B(store),
    .C(_1193_),
    .Y(_1194_)
);

FILL FILL_0__1760_ (
);

FILL FILL_2__1778_ (
);

FILL FILL_4__2645_ (
);

FILL FILL_4__2225_ (
);

FILL FILL_0__2965_ (
);

FILL FILL_0__2545_ (
);

FILL FILL_6__3512_ (
);

FILL FILL_0__2125_ (
);

FILL FILL_2__3504_ (
);

FILL FILL_7__1947_ (
);

FILL FILL_1__1921_ (
);

FILL FILL_3__1847_ (
);

FILL FILL_5__2714_ (
);

FILL FILL_1__2706_ (
);

NAND2X1 _1776_ (
    .A(state[5]),
    .B(_901_),
    .Y(_902_)
);

FILL FILL_4__3183_ (
);

FILL FILL_0__3083_ (
);

FILL FILL_4__1916_ (
);

FILL FILL_7__2485_ (
);

FILL FILL_0__1816_ (
);

OAI21X1 _3502_ (
    .A(AI[4]),
    .B(_1529_),
    .C(_1722_),
    .Y(_1532_)
);

FILL FILL_3__2385_ (
);

FILL FILL_5__3672_ (
);

FILL FILL_5__3252_ (
);

FILL FILL_1__3664_ (
);

FILL FILL_1__3244_ (
);

FILL FILL_4__2874_ (
);

FILL FILL_4__2454_ (
);

FILL FILL_4__2034_ (
);

AOI21X1 _3099_ (
    .A(_702_),
    .B(_707_),
    .C(_708_),
    .Y(_709_)
);

FILL FILL_0__2774_ (
);

FILL FILL_0__2354_ (
);

FILL FILL_2__3313_ (
);

FILL FILL_4__3659_ (
);

FILL FILL_7__1756_ (
);

FILL FILL_4__3239_ (
);

FILL FILL_0__3559_ (
);

FILL FILL_0__3139_ (
);

FILL FILL_5__2943_ (
);

FILL FILL_5__2523_ (
);

FILL FILL_5__2103_ (
);

FILL FILL_1__2935_ (
);

FILL FILL_1__2515_ (
);

FILL FILL_5__3308_ (
);

OAI21X1 _3311_ (
    .A(_291_),
    .B(_869_),
    .C(_874_),
    .Y(_113_)
);

FILL FILL_3__2194_ (
);

FILL FILL_5__3481_ (
);

FILL FILL_5__3061_ (
);

FILL FILL_1__3473_ (
);

FILL FILL_1__3053_ (
);

FILL FILL_4__2683_ (
);

FILL FILL_4__2263_ (
);

FILL FILL_6__2189_ (
);

FILL FILL_0__2583_ (
);

FILL FILL_6__3550_ (
);

FILL FILL_0__2163_ (
);

FILL FILL_6__3130_ (
);

FILL FILL_2__3542_ (
);

FILL FILL_2__3122_ (
);

FILL FILL_7__1985_ (
);

FILL FILL_4__3468_ (
);

FILL FILL_4__3048_ (
);

FILL FILL_3__1885_ (
);

FILL FILL_5__2752_ (
);

FILL FILL_5__2332_ (
);

FILL FILL_1__2744_ (
);

FILL FILL_1__2324_ (
);

FILL FILL_3__3611_ (
);

FILL FILL_5__3537_ (
);

FILL FILL_5__3117_ (
);

FILL FILL_1__3529_ (
);

FILL FILL_1__3109_ (
);

FILL FILL_4__1954_ (
);

INVX1 _2599_ (
    .A(_283_),
    .Y(_284_)
);

NAND2X1 _2179_ (
    .A(_1287_),
    .B(_1285_),
    .Y(_1288_)
);

FILL FILL_0__1854_ (
);

FILL FILL_6__2821_ (
);

AOI21X1 _3540_ (
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1569_),
    .Y(_1570_)
);

FILL FILL_6__2401_ (
);

NAND2X1 _3120_ (
    .A(HC),
    .B(_726_),
    .Y(_727_)
);

FILL FILL169950x64950 (
);

FILL FILL_2__2813_ (
);

FILL FILL_4__2739_ (
);

FILL FILL_4__2319_ (
);

FILL FILL_5__3290_ (
);

FILL FILL_0__2639_ (
);

FILL FILL_6__3606_ (
);

FILL FILL_0__2219_ (
);

FILL FILL_1__3282_ (
);

FILL FILL_4__2492_ (
);

FILL FILL_4__2072_ (
);

FILL FILL_5__2808_ (
);

FILL FILL_0__2392_ (
);

FILL FILL_4__3697_ (
);

FILL FILL_4__3277_ (
);

OAI21X1 _2811_ (
    .A(_473_),
    .B(_197_),
    .C(_148_),
    .Y(_474_)
);

FILL FILL_0__3597_ (
);

FILL FILL_0__3177_ (
);

FILL FILL_7__2999_ (
);

FILL FILL_5__2981_ (
);

FILL FILL_5__2561_ (
);

FILL FILL_7__2579_ (
);

FILL FILL_7__2159_ (
);

FILL FILL_5__2141_ (
);

FILL FILL_1__2973_ (
);

FILL FILL_1__2553_ (
);

FILL FILL_1__2133_ (
);

FILL FILL_3__2899_ (
);

FILL FILL_3__2479_ (
);

FILL FILL_3__2059_ (
);

FILL FILL_3__3000_ (
);

FILL FILL_4__1763_ (
);

FILL FILL_6__2630_ (
);

FILL FILL_6__2210_ (
);

FILL FILL_2__2622_ (
);

FILL FILL_2__2202_ (
);

FILL FILL_4__2968_ (
);

FILL FILL_4__2548_ (
);

FILL FILL_4__2128_ (
);

FILL FILL_0__2868_ (
);

FILL FILL_0__2448_ (
);

FILL FILL_0__2028_ (
);

FILL FILL_1__3091_ (
);

FILL FILL_5__1832_ (
);

FILL FILL_1__1824_ (
);

FILL FILL_5__2617_ (
);

FILL FILL_1__2609_ (
);

FILL FILL_2__3580_ (
);

FILL FILL_2__3160_ (
);

FILL FILL_4__3086_ (
);

FILL FILL_6__1901_ (
);

AOI21X1 _2620_ (
    .A(_198_),
    .B(ADD[6]),
    .C(_1135_),
    .Y(_301_)
);

INVX1 _2200_ (
    .A(_1028_),
    .Y(_1309_)
);

FILL FILL_4__1819_ (
);

FILL FILL_5__2790_ (
);

FILL FILL_5__2370_ (
);

FILL FILL_7__2388_ (
);

DFFSR _3405_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_74_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[0] [5])
);

FILL FILL_1__2782_ (
);

FILL FILL_1__2362_ (
);

FILL FILL_3__2288_ (
);

FILL FILL_5__3575_ (
);

FILL FILL_5__3155_ (
);

FILL FILL_1__3567_ (
);

FILL FILL_1__3147_ (
);

FILL FILL_4__1992_ (
);

FILL FILL_0__1892_ (
);

FILL FILL_2__2851_ (
);

FILL FILL_2__2431_ (
);

FILL FILL_2__2011_ (
);

FILL FILL_4__2777_ (
);

FILL FILL_4__2357_ (
);

FILL FILL_0__2677_ (
);

FILL FILL_6__3644_ (
);

FILL FILL_0__2257_ (
);

FILL FILL_6__3224_ (
);

FILL FILL_2__3636_ (
);

FILL FILL_2__3216_ (
);

FILL FILL_7__2600_ (
);

FILL FILL_3__1979_ (
);

FILL FILL_3__2920_ (
);

FILL FILL_3__2500_ (
);

FILL FILL_5__2846_ (
);

FILL FILL_5__2426_ (
);

FILL FILL_5__2006_ (
);

FILL FILL_1__2838_ (
);

FILL FILL_1__2418_ (
);

FILL FILL_3__3705_ (
);

FILL FILL_0__1948_ (
);

FILL FILL_6__2915_ (
);

NAND2X1 _3634_ (
    .A(_1662_),
    .B(_1663_),
    .Y(_1664_)
);

AOI21X1 _3214_ (
    .A(_754_),
    .B(_798_),
    .C(_802_),
    .Y(_88_)
);

FILL FILL_1__2591_ (
);

FILL FILL_1__2171_ (
);

FILL FILL_3__2097_ (
);

FILL FILL_2__2907_ (
);

FILL FILL_2__2660_ (
);

FILL FILL_2__2240_ (
);

FILL FILL_4__2586_ (
);

FILL FILL_4__2166_ (
);

FILL FILL_0__2486_ (
);

FILL FILL_6__3453_ (
);

FILL FILL_0__2066_ (
);

FILL FILL_6__3033_ (
);

FILL FILL_2__3025_ (
);

FILL FILL_7__1888_ (
);

FILL FILL_5__1870_ (
);

NOR2X1 _2905_ (
    .A(_1178_),
    .B(_551_),
    .Y(_552_)
);

FILL FILL_1__1862_ (
);

FILL FILL_3__1788_ (
);

FILL FILL_5__2655_ (
);

FILL FILL_5__2235_ (
);

FILL FILL_1__2647_ (
);

FILL FILL_7__3614_ (
);

FILL FILL_1__2227_ (
);

FILL FILL_3__3514_ (
);

FILL FILL_2__1931_ (
);

FILL FILL_4__1857_ (
);

FILL FILL_0__1757_ (
);

FILL FILL_6__2724_ (
);

DFFSR _3443_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(_111_),
    .CLK(clk_bF$buf2),
    .Q(ABH[2])
);

FILL FILL_6__2304_ (
);

INVX2 _3023_ (
    .A(_646_),
    .Y(_647_)
);

FILL FILL_2__2716_ (
);

FILL FILL_5__3193_ (
);

FILL FILL_6__3509_ (
);

FILL FILL_1__3185_ (
);

FILL FILL_5__1926_ (
);

FILL FILL_1__1918_ (
);

FILL FILL_4__2395_ (
);

FILL FILL_0__2295_ (
);

FILL FILL_6__3262_ (
);

FILL FILL_2__3674_ (
);

FILL FILL_2__3254_ (
);

AOI21X1 _2714_ (
    .A(_352_),
    .B(_353_),
    .C(_1011_),
    .Y(_384_)
);

FILL FILL_5__2884_ (
);

FILL FILL_5__2464_ (
);

FILL FILL_5__2044_ (
);

FILL FILL_1__2876_ (
);

FILL FILL_1__2456_ (
);

FILL FILL_1__2036_ (
);

FILL FILL_7__3003_ (
);

FILL FILL_5__3669_ (
);

FILL FILL_5__3249_ (
);

FILL FILL_4_CLKBUF1_insert26 (
);

FILL FILL_4_CLKBUF1_insert27 (
);

FILL FILL_4_CLKBUF1_insert28 (
);

FILL FILL_4_CLKBUF1_insert29 (
);

FILL FILL_0__1986_ (
);

FILL FILL_6__2953_ (
);

OAI21X1 _3672_ (
    .A(_1714__bF$buf0),
    .B(_1678_),
    .C(_1694_),
    .Y(_1522_)
);

FILL FILL_6__2533_ (
);

NOR2X1 _3252_ (
    .A(_817_),
    .B(_827_),
    .Y(_828_)
);

FILL FILL_6__2113_ (
);

FILL FILL_2__2945_ (
);

FILL FILL_2__2525_ (
);

FILL FILL_2__2105_ (
);

FILL FILL_0__3712_ (
);

FILL FILL_6__3491_ (
);

FILL FILL_6__3071_ (
);

FILL FILL_0_BUFX2_insert40 (
);

FILL FILL_0_BUFX2_insert41 (
);

FILL FILL_2__3483_ (
);

FILL FILL_0_BUFX2_insert42 (
);

FILL FILL_2__3063_ (
);

FILL FILL_0_BUFX2_insert43 (
);

FILL FILL_0_BUFX2_insert44 (
);

FILL FILL_0_BUFX2_insert45 (
);

FILL FILL_0_BUFX2_insert46 (
);

FILL FILL_0_BUFX2_insert47 (
);

FILL FILL_0_BUFX2_insert48 (
);

FILL FILL_0_BUFX2_insert49 (
);

FILL FILL_6__1804_ (
);

AND2X2 _2943_ (
    .A(_566_),
    .B(_585_),
    .Y(_586_)
);

NAND2X1 _2523_ (
    .A(_203_),
    .B(_217_),
    .Y(_218_)
);

AOI21X1 _2103_ (
    .A(_1168_),
    .B(_1010_),
    .C(_1211_),
    .Y(_1212_)
);

FILL FILL_5__2693_ (
);

FILL FILL_5__2273_ (
);

NAND2X1 _3308_ (
    .A(_1741_[11]),
    .B(_869_),
    .Y(_873_)
);

FILL FILL_1__2685_ (
);

FILL FILL_1__2265_ (
);

FILL FILL_7__3232_ (
);

FILL FILL_3__3552_ (
);

FILL FILL_3__3132_ (
);

FILL FILL_5__3478_ (
);

FILL FILL_5__3058_ (
);

FILL FILL_4__1895_ (
);

FILL FILL_0__1795_ (
);

FILL FILL_6__2762_ (
);

AOI21X1 _3481_ (
    .A(BI[7]),
    .B(alu_op[2]),
    .C(_1726_),
    .Y(_1727_)
);

FILL FILL_6__2342_ (
);

OAI21X1 _3061_ (
    .A(_529_),
    .B(_355_),
    .C(_674_),
    .Y(_675_)
);

FILL FILL_2__2754_ (
);

FILL FILL_2__2334_ (
);

FILL FILL_4__3621_ (
);

FILL FILL_4__3201_ (
);

FILL FILL_6__3547_ (
);

FILL FILL_6__3127_ (
);

FILL FILL_2__3539_ (
);

FILL FILL_0__3521_ (
);

FILL FILL_2__3119_ (
);

FILL FILL_0__3101_ (
);

FILL FILL_5__1964_ (
);

FILL FILL_1__1956_ (
);

FILL FILL_7__2503_ (
);

FILL FILL_3__2823_ (
);

FILL FILL_3__2403_ (
);

FILL FILL_5__2749_ (
);

FILL FILL_5__2329_ (
);

FILL FILL_7__3708_ (
);

FILL FILL_2__3292_ (
);

FILL FILL_3__3608_ (
);

NOR2X1 _2752_ (
    .A(_312_),
    .B(_365_),
    .Y(_418_)
);

OAI21X1 _2332_ (
    .A(_886__bF$buf2),
    .B(_1432_),
    .C(_1438_),
    .Y(_1439_)
);

FILL FILL_5__2082_ (
);

FILL FILL_6__2818_ (
);

OAI21X1 _3537_ (
    .A(AI[1]),
    .B(_1566_),
    .C(_1722_),
    .Y(_1567_)
);

NAND2X1 _3117_ (
    .A(\AXYS[0] [0]),
    .B(_722_),
    .Y(_725_)
);

FILL FILL_1__2494_ (
);

FILL FILL_7__3461_ (
);

FILL FILL_1__2074_ (
);

FILL FILL_7__3041_ (
);

FILL FILL_5__3287_ (
);

FILL FILL_1__3699_ (
);

FILL FILL_1__3279_ (
);

FILL FILL_6__2991_ (
);

FILL FILL_6__2571_ (
);

OAI21X1 _3290_ (
    .A(_860_),
    .B(_236_),
    .C(_863_),
    .Y(_103_)
);

FILL FILL_6__2151_ (
);

FILL FILL_2__2983_ (
);

FILL FILL_2__2563_ (
);

FILL FILL_2__2143_ (
);

FILL FILL_4__2489_ (
);

FILL FILL_4__2069_ (
);

FILL FILL_4__3010_ (
);

FILL FILL_0__2389_ (
);

FILL FILL_5__1773_ (
);

NAND2X1 _2808_ (
    .A(_276_),
    .B(_365_),
    .Y(_471_)
);

FILL FILL_1__1765_ (
);

FILL FILL_7__2732_ (
);

FILL FILL_3__2632_ (
);

FILL FILL_3__2212_ (
);

FILL FILL_5__2978_ (
);

FILL FILL_5__2558_ (
);

FILL FILL_5__2138_ (
);

FILL FILL_7__3517_ (
);

FILL FILL_6__1842_ (
);

OAI21X1 _2981_ (
    .A(_1172_),
    .B(_610_),
    .C(_579_),
    .Y(_611_)
);

INVX1 _2561_ (
    .A(ABL[5]),
    .Y(_251_)
);

INVX1 _2141_ (
    .A(_1249_),
    .Y(_1250_)
);

FILL FILL_2__1834_ (
);

FILL FILL_4__2701_ (
);

FILL FILL_6__2627_ (
);

DFFSR _3346_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_23_),
    .CLK(clk_bF$buf4),
    .Q(php)
);

FILL FILL_6__2207_ (
);

FILL FILL_7__3270_ (
);

FILL FILL_0__2601_ (
);

FILL FILL_2__2619_ (
);

FILL FILL_3__3590_ (
);

FILL FILL_3__3170_ (
);

FILL FILL_5__3096_ (
);

FILL FILL_1__3088_ (
);

FILL FILL_3__1903_ (
);

FILL FILL_5__1829_ (
);

FILL FILL_6__2380_ (
);

FILL FILL_2__2792_ (
);

FILL FILL_2__2372_ (
);

FILL FILL_4__2298_ (
);

NAND2X1 _1832_ (
    .A(_937_),
    .B(_957_),
    .Y(_958_)
);

FILL FILL_6__3585_ (
);

FILL FILL_0__2198_ (
);

FILL FILL_6__3165_ (
);

FILL FILL_2__3577_ (
);

FILL FILL_2__3157_ (
);

AOI21X1 _2617_ (
    .A(_272_),
    .B(DIMUX[5]),
    .C(_298_),
    .Y(_299_)
);

FILL FILL_1__1994_ (
);

FILL FILL_7__2961_ (
);

FILL FILL_7__2541_ (
);

FILL FILL_7__2121_ (
);

FILL FILL_3__2861_ (
);

FILL FILL_3__2441_ (
);

FILL FILL_3__2021_ (
);

FILL FILL_5__2787_ (
);

FILL FILL_5__2367_ (
);

FILL FILL_1__2779_ (
);

FILL FILL_1__2359_ (
);

BUFX2 BUFX2_insert50 (
    .A(_931_),
    .Y(_931__bF$buf4)
);

BUFX2 BUFX2_insert51 (
    .A(_931_),
    .Y(_931__bF$buf3)
);

BUFX2 BUFX2_insert52 (
    .A(_931_),
    .Y(_931__bF$buf2)
);

BUFX2 BUFX2_insert53 (
    .A(_931_),
    .Y(_931__bF$buf1)
);

BUFX2 BUFX2_insert54 (
    .A(_931_),
    .Y(_931__bF$buf0)
);

FILL FILL_1__3300_ (
);

BUFX2 BUFX2_insert55 (
    .A(_1150_),
    .Y(_1150__bF$buf4)
);

BUFX2 BUFX2_insert56 (
    .A(_1150_),
    .Y(_1150__bF$buf3)
);

BUFX2 BUFX2_insert57 (
    .A(_1150_),
    .Y(_1150__bF$buf2)
);

BUFX2 BUFX2_insert58 (
    .A(_1150_),
    .Y(_1150__bF$buf1)
);

FILL FILL_3__3646_ (
);

BUFX2 BUFX2_insert59 (
    .A(_1150_),
    .Y(_1150__bF$buf0)
);

FILL FILL_3__3226_ (
);

NAND2X1 _2790_ (
    .A(PC[11]),
    .B(_365_),
    .Y(_454_)
);

NAND3X1 _2370_ (
    .A(_1150__bF$buf3),
    .B(_1370_),
    .C(_1351_),
    .Y(_1476_)
);

FILL FILL_4__1989_ (
);

FILL FILL_4__2930_ (
);

FILL FILL_4__2510_ (
);

FILL FILL_0__1889_ (
);

FILL FILL_6__2856_ (
);

INVX1 _3575_ (
    .A(_1602_),
    .Y(_1605_)
);

FILL FILL_6__2436_ (
);

FILL FILL_6__2016_ (
);

OAI21X1 _3155_ (
    .A(_722_),
    .B(_757_),
    .C(_758_),
    .Y(_73_)
);

FILL FILL_2__2848_ (
);

FILL FILL_0__2830_ (
);

FILL FILL_2__2428_ (
);

FILL FILL_0__2410_ (
);

FILL FILL_2__2008_ (
);

FILL FILL_4__3715_ (
);

FILL FILL_0__3615_ (
);

FILL FILL_2__2181_ (
);

FILL FILL_3__2917_ (
);

NAND3X1 _2846_ (
    .A(_500_),
    .B(_506_),
    .C(_466_),
    .Y(_507_)
);

OAI21X1 _2426_ (
    .A(_132_),
    .B(_129_),
    .C(_131_),
    .Y(alu_op[1])
);

OAI21X1 _2006_ (
    .A(_888_),
    .B(_983_),
    .C(_1118_),
    .Y(_1119_)
);

FILL FILL_7__2770_ (
);

FILL FILL_7__2350_ (
);

FILL FILL_3__2670_ (
);

FILL FILL_3__2250_ (
);

FILL FILL_5__2596_ (
);

FILL FILL_5__2176_ (
);

FILL FILL_1__2588_ (
);

FILL FILL_1__2168_ (
);

FILL FILL_7__3135_ (
);

FILL FILL_3__3455_ (
);

FILL FILL_3__3035_ (
);

FILL FILL_6__1880_ (
);

FILL FILL_2__1872_ (
);

FILL FILL_4__1798_ (
);

FILL FILL_6__2665_ (
);

DFFPOSX1 _3384_ (
    .D(_53_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD[0])
);

FILL FILL_6__2245_ (
);

FILL FILL_2__2657_ (
);

FILL FILL_2__2237_ (
);

FILL FILL_4__3524_ (
);

FILL FILL_4__3104_ (
);

FILL FILL_3__1941_ (
);

FILL FILL_0__3004_ (
);

FILL FILL_5__1867_ (
);

FILL FILL_1__1859_ (
);

FILL FILL_7__2406_ (
);

FILL FILL_1__2800_ (
);

FILL FILL_3__2726_ (
);

FILL FILL_3__2306_ (
);

NAND3X1 _1870_ (
    .A(_987_),
    .B(_994_),
    .C(_991_),
    .Y(_995_)
);

FILL FILL_2__3195_ (
);

FILL FILL_6__1936_ (
);

AOI21X1 _2655_ (
    .A(_326_),
    .B(_328_),
    .C(_329_),
    .Y(_330_)
);

INVX1 _2235_ (
    .A(_1342_),
    .Y(_1343_)
);

FILL FILL_3_CLKBUF1_insert30 (
);

FILL FILL_3_CLKBUF1_insert31 (
);

FILL FILL_3_CLKBUF1_insert32 (
);

FILL FILL_3_CLKBUF1_insert33 (
);

FILL FILL_3_CLKBUF1_insert34 (
);

FILL FILL_3_CLKBUF1_insert35 (
);

FILL FILL_3_CLKBUF1_insert36 (
);

FILL FILL_2__1928_ (
);

FILL FILL_0__1910_ (
);

FILL FILL_1__2397_ (
);

FILL FILL_3__3264_ (
);

FILL FILL_6__2894_ (
);

FILL FILL_6__2474_ (
);

OAI21X1 _3193_ (
    .A(_737_),
    .B(_789_),
    .C(_791_),
    .Y(_78_)
);

FILL FILL_6__2054_ (
);

FILL FILL_2__2886_ (
);

FILL FILL_2__2466_ (
);

FILL FILL_2__2046_ (
);

NOR2X1 _1926_ (
    .A(_1042_),
    .B(_1027__bF$buf0),
    .Y(_1043_)
);

FILL FILL_7__1850_ (
);

FILL FILL_6__3259_ (
);

FILL FILL_3__1750_ (
);

FILL FILL_0__3653_ (
);

FILL FILL_0__3233_ (
);

FILL FILL_7__2635_ (
);

FILL FILL_3__2955_ (
);

FILL FILL_3__2535_ (
);

FILL FILL_3__2115_ (
);

FILL FILL_6__1745_ (
);

NAND2X1 _2884_ (
    .A(_1348_),
    .B(_1330_),
    .Y(_537_)
);

INVX1 _2464_ (
    .A(D),
    .Y(_164_)
);

INVX1 _2044_ (
    .A(NMI_edge),
    .Y(_1153_)
);

FILL FILL_4__2604_ (
);

OAI21X1 _3669_ (
    .A(_1629_),
    .B(_1626_),
    .C(RDY_bF$buf7),
    .Y(_1693_)
);

AND2X2 _3249_ (
    .A(_1200_),
    .B(_824_),
    .Y(_825_)
);

FILL FILL_7__3593_ (
);

FILL FILL_0__2924_ (
);

FILL FILL_0__2504_ (
);

FILL FILL_3__3493_ (
);

FILL FILL_3__3073_ (
);

FILL FILL_7__1906_ (
);

FILL FILL_0__3709_ (
);

FILL FILL_3__1806_ (
);

FILL FILL_6__2283_ (
);

FILL FILL_2__2695_ (
);

FILL FILL_2__2275_ (
);

FILL FILL_4__3562_ (
);

FILL FILL_4__3142_ (
);

FILL FILL_6__3488_ (
);

FILL FILL_6__3068_ (
);

FILL FILL_0__3462_ (
);

FILL FILL_0__3042_ (
);

FILL FILL_1__1897_ (
);

FILL FILL_7__2864_ (
);

FILL FILL_7__2024_ (
);

FILL FILL_3__2764_ (
);

FILL FILL_3__2344_ (
);

FILL FILL_5__3631_ (
);

FILL FILL_5__3211_ (
);

FILL FILL_1__3623_ (
);

FILL FILL_1__3203_ (
);

FILL FILL_3__3549_ (
);

FILL FILL_3__3129_ (
);

FILL FILL_6__1974_ (
);

NAND3X1 _2693_ (
    .A(_1027__bF$buf4),
    .B(_148_),
    .C(_197_),
    .Y(_364_)
);

OR2X2 _2273_ (
    .A(_1380_),
    .B(_1373_),
    .Y(_1381_)
);

FILL FILL_2__1966_ (
);

FILL FILL_4__2833_ (
);

FILL FILL_4__2413_ (
);

FILL FILL_6__2759_ (
);

OAI21X1 _3478_ (
    .A(_1723_),
    .B(_1721_),
    .C(_1715_),
    .Y(_1724_)
);

FILL FILL_6__2339_ (
);

OAI21X1 _3058_ (
    .A(_1027__bF$buf2),
    .B(_671_),
    .C(_657_),
    .Y(_672_)
);

FILL FILL_0__2733_ (
);

FILL FILL_0__2313_ (
);

FILL FILL_6__3700_ (
);

FILL FILL_4__3618_ (
);

FILL FILL_0__3518_ (
);

FILL FILL_6__2092_ (
);

FILL FILL_5__2902_ (
);

FILL FILL_2__2084_ (
);

NOR2X1 _1964_ (
    .A(_1080_),
    .B(_959_),
    .Y(_1081_)
);

FILL FILL_6__3297_ (
);

FILL FILL_0__3691_ (
);

FILL FILL_2__3289_ (
);

FILL FILL_0__3271_ (
);

AOI21X1 _2749_ (
    .A(_413_),
    .B(_414_),
    .C(_374_),
    .Y(_415_)
);

OAI21X1 _2329_ (
    .A(RDY_bF$buf8),
    .B(_1233_),
    .C(_1435_),
    .Y(_1436_)
);

FILL FILL_7__2253_ (
);

FILL FILL_3__2993_ (
);

FILL FILL_3__2573_ (
);

FILL FILL_3__2153_ (
);

FILL FILL_5__2499_ (
);

FILL FILL_5__2079_ (
);

FILL FILL_7__3458_ (
);

FILL FILL_5__3020_ (
);

FILL FILL_7__3038_ (
);

FILL FILL_1__3012_ (
);

FILL FILL_6__1783_ (
);

NOR2X1 _2082_ (
    .A(_1175_),
    .B(_1190_),
    .Y(_1191_)
);

FILL FILL_5_BUFX2_insert60 (
);

FILL FILL_5_BUFX2_insert61 (
);

FILL FILL_5_BUFX2_insert62 (
);

FILL FILL_5_BUFX2_insert63 (
);

FILL FILL_5_BUFX2_insert64 (
);

FILL FILL_2__1775_ (
);

FILL FILL_5_BUFX2_insert65 (
);

FILL FILL_5_BUFX2_insert66 (
);

FILL FILL_5_BUFX2_insert67 (
);

FILL FILL_5_BUFX2_insert68 (
);

FILL FILL_5_BUFX2_insert69 (
);

FILL FILL_4__2642_ (
);

FILL FILL_4__2222_ (
);

FILL FILL_6__2988_ (
);

FILL FILL_6__2568_ (
);

NAND2X1 _3287_ (
    .A(ABL[1]),
    .B(_860_),
    .Y(_862_)
);

FILL FILL_6__2148_ (
);

FILL FILL_0__2962_ (
);

FILL FILL_0__2542_ (
);

FILL FILL_0__2122_ (
);

FILL FILL_2__3501_ (
);

FILL FILL_4__3007_ (
);

FILL FILL_3__1844_ (
);

FILL FILL_5__2711_ (
);

FILL FILL_7__2729_ (
);

FILL FILL_7__2309_ (
);

FILL FILL_1__2703_ (
);

FILL FILL_3__2629_ (
);

FILL FILL_3__2209_ (
);

NAND2X1 _1773_ (
    .A(state[1]),
    .B(state[0]),
    .Y(_899_)
);

FILL FILL_4__3180_ (
);

FILL FILL_0__3080_ (
);

FILL FILL_2__3098_ (
);

FILL FILL_4__1913_ (
);

FILL FILL_6__1839_ (
);

OAI21X1 _2978_ (
    .A(_1149__bF$buf1),
    .B(_607_),
    .C(_608_),
    .Y(_46_)
);

AOI21X1 _2558_ (
    .A(_1116_),
    .B(_195_),
    .C(_248_),
    .Y(_249_)
);

AOI21X1 _2138_ (
    .A(_1231_),
    .B(_1230_),
    .C(_1246_),
    .Y(_1247_)
);

FILL FILL_7__2482_ (
);

FILL FILL_0__1813_ (
);

FILL FILL_3__2382_ (
);

FILL FILL_7__3267_ (
);

FILL FILL_1__3661_ (
);

FILL FILL_1__3241_ (
);

FILL FILL_3__3587_ (
);

FILL FILL_3__3167_ (
);

FILL FILL_4__2871_ (
);

FILL FILL_4__2451_ (
);

FILL FILL_4__2031_ (
);

FILL FILL_6__2797_ (
);

FILL FILL_6__2377_ (
);

NOR2X1 _3096_ (
    .A(plp),
    .B(clc),
    .Y(_706_)
);

FILL FILL_2__2789_ (
);

FILL FILL_0__2771_ (
);

FILL FILL_2__2369_ (
);

FILL FILL_0__2351_ (
);

FILL FILL_2__3310_ (
);

INVX1 _1829_ (
    .A(_954_),
    .Y(_955_)
);

FILL FILL_7__1753_ (
);

FILL FILL_4__3656_ (
);

FILL FILL_4__3236_ (
);

FILL FILL_0__3556_ (
);

FILL FILL_0__3136_ (
);

FILL FILL_5__1999_ (
);

FILL FILL_5__2940_ (
);

FILL FILL_5__2520_ (
);

FILL FILL_7__2538_ (
);

FILL FILL_5__2100_ (
);

FILL FILL_1__2932_ (
);

FILL FILL_1__2512_ (
);

FILL FILL_3__2858_ (
);

FILL FILL_3__2438_ (
);

FILL FILL_3__2018_ (
);

FILL FILL_5__3305_ (
);

OAI21X1 _2787_ (
    .A(_285_),
    .B(_352_),
    .C(_450_),
    .Y(_451_)
);

NAND2X1 _2367_ (
    .A(_1472_),
    .B(_1466_),
    .Y(_1473_)
);

FILL FILL_3__2191_ (
);

FILL FILL_4__2927_ (
);

FILL FILL_4__2507_ (
);

FILL FILL_7__3496_ (
);

FILL FILL_0__2827_ (
);

FILL FILL_0__2407_ (
);

FILL FILL_1__3470_ (
);

FILL FILL_1__3050_ (
);

FILL FILL_7__1809_ (
);

FILL FILL_4__2680_ (
);

FILL FILL_4__2260_ (
);

FILL FILL_6__2186_ (
);

FILL FILL_2__2598_ (
);

FILL FILL_0__2580_ (
);

FILL FILL_0__2160_ (
);

FILL FILL_2__2178_ (
);

FILL FILL_7__1982_ (
);

FILL FILL_4__3465_ (
);

FILL FILL_4__3045_ (
);

FILL FILL_3__1882_ (
);

FILL FILL_7__2767_ (
);

FILL FILL_1__2741_ (
);

FILL FILL_1__2321_ (
);

FILL FILL_3__2667_ (
);

FILL FILL_3__2247_ (
);

FILL FILL_5__3534_ (
);

FILL FILL_5__3114_ (
);

FILL FILL_1__3526_ (
);

FILL FILL_1__3106_ (
);

FILL FILL_4__1951_ (
);

FILL FILL_6__1877_ (
);

AOI22X1 _2596_ (
    .A(ADD[2]),
    .B(_198_),
    .C(_272_),
    .D(DIMUX[2]),
    .Y(_281_)
);

AOI22X1 _2176_ (
    .A(_886__bF$buf1),
    .B(_1201_),
    .C(_1284_),
    .D(_1283_),
    .Y(_1285_)
);

FILL FILL_2__1869_ (
);

FILL FILL_0__1851_ (
);

FILL FILL_2__2810_ (
);

FILL FILL_4__2736_ (
);

FILL FILL_4__2316_ (
);

FILL FILL_0__2636_ (
);

FILL FILL_6__3603_ (
);

FILL FILL_0__2216_ (
);

FILL FILL_3__1938_ (
);

FILL FILL_5__2805_ (
);

INVX1 _1867_ (
    .A(_989_),
    .Y(_992_)
);

FILL FILL_4__3694_ (
);

FILL FILL_4__3274_ (
);

FILL FILL_0__3594_ (
);

FILL FILL_0__3174_ (
);

FILL FILL_7__2996_ (
);

FILL FILL_7__2156_ (
);

FILL FILL_0__1907_ (
);

FILL FILL_1__2970_ (
);

FILL FILL_1__2550_ (
);

FILL FILL_1__2130_ (
);

FILL FILL_3__2896_ (
);

FILL FILL_3__2476_ (
);

FILL FILL_3__2056_ (
);

FILL FILL_4__1760_ (
);

FILL FILL_4__2965_ (
);

FILL FILL_4__2545_ (
);

FILL FILL_4__2125_ (
);

FILL FILL_0__2865_ (
);

FILL FILL_0__2445_ (
);

FILL FILL_0__2025_ (
);

FILL FILL_7__1847_ (
);

FILL FILL_1__1821_ (
);

FILL FILL_3__1747_ (
);

FILL FILL_5__2614_ (
);

FILL FILL_1__2606_ (
);

FILL FILL_4__3083_ (
);

FILL FILL_4__1816_ (
);

FILL FILL_7__2385_ (
);

DFFSR _3402_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_71_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[0] [2])
);

FILL FILL_3__2285_ (
);

FILL FILL_5__3572_ (
);

FILL FILL_5__3152_ (
);

FILL FILL_1__3564_ (
);

FILL FILL_1__3144_ (
);

FILL FILL_4__2774_ (
);

FILL FILL_4__2354_ (
);

FILL FILL_0__2674_ (
);

FILL FILL_6__3641_ (
);

FILL FILL_0__2254_ (
);

FILL FILL_6__3221_ (
);

FILL FILL_2__3633_ (
);

FILL FILL_2__3213_ (
);

FILL FILL_4__3559_ (
);

FILL FILL_4__3139_ (
);

FILL FILL_3__1976_ (
);

FILL FILL_0__3459_ (
);

FILL FILL_0__3039_ (
);

FILL FILL_5__2843_ (
);

FILL FILL_5__2423_ (
);

FILL FILL_5__2003_ (
);

FILL FILL_1__2835_ (
);

FILL FILL_1__2415_ (
);

FILL FILL_3__3702_ (
);

FILL FILL_5__3628_ (
);

FILL FILL_5__3208_ (
);

FILL FILL_0__1945_ (
);

FILL FILL_6__2912_ (
);

NAND2X1 _3631_ (
    .A(_1639_),
    .B(_1660_),
    .Y(_1661_)
);

NOR2X1 _3211_ (
    .A(\AXYS[2] [2]),
    .B(_798_),
    .Y(_801_)
);

FILL FILL_3__2094_ (
);

FILL FILL_2__2904_ (
);

FILL FILL_3__3299_ (
);

FILL FILL_4__2583_ (
);

FILL FILL_4__2163_ (
);

FILL FILL_6__2089_ (
);

FILL FILL_0__2483_ (
);

FILL FILL_6__3450_ (
);

FILL FILL_0__2063_ (
);

FILL FILL_6__3030_ (
);

FILL FILL_2__3022_ (
);

FILL FILL_7__1885_ (
);

OAI21X1 _2902_ (
    .A(_886__bF$buf5),
    .B(_1027__bF$buf0),
    .C(clv),
    .Y(_549_)
);

FILL FILL_3__1785_ (
);

FILL FILL_0__3268_ (
);

FILL FILL_5__2652_ (
);

FILL FILL_5__2232_ (
);

FILL FILL_1__2644_ (
);

FILL FILL_7__3611_ (
);

FILL FILL_1__2224_ (
);

FILL FILL_3__3511_ (
);

FILL FILL_5__3017_ (
);

FILL FILL_1__3009_ (
);

FILL FILL_4__1854_ (
);

NOR2X1 _2499_ (
    .A(_193_),
    .B(_135_),
    .Y(_194_)
);

NAND2X1 _2079_ (
    .A(_1185_),
    .B(_1187_),
    .Y(_1188_)
);

FILL FILL_0__1754_ (
);

FILL FILL_6__2721_ (
);

DFFSR _3440_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_108_),
    .CLK(clk_bF$buf1),
    .Q(ABL[7])
);

FILL FILL_6__2301_ (
);

AND2X2 _3020_ (
    .A(_1027__bF$buf4),
    .B(res),
    .Y(_52_)
);

FILL FILL_2__2713_ (
);

FILL FILL_4__2639_ (
);

FILL FILL_4__2219_ (
);

FILL FILL_5__3190_ (
);

FILL FILL_0__2959_ (
);

FILL FILL_0__2539_ (
);

FILL FILL_6__3506_ (
);

FILL FILL_0__2119_ (
);

FILL FILL_1__3182_ (
);

FILL FILL_5__1923_ (
);

FILL FILL_1__1915_ (
);

FILL FILL_4__2392_ (
);

FILL FILL_5__2708_ (
);

FILL FILL_0__2292_ (
);

FILL FILL_2__3671_ (
);

FILL FILL_2__3251_ (
);

FILL FILL_4__3597_ (
);

FILL FILL_4__3177_ (
);

OAI21X1 _2711_ (
    .A(_179_),
    .B(_326_),
    .C(_380_),
    .Y(_381_)
);

FILL FILL_0__3497_ (
);

FILL FILL_0__3077_ (
);

FILL FILL_5__2881_ (
);

FILL FILL_7__2899_ (
);

FILL FILL_7__2479_ (
);

FILL FILL_5__2461_ (
);

FILL FILL_7__2059_ (
);

FILL FILL_5__2041_ (
);

FILL FILL_1__2873_ (
);

FILL FILL_1__2453_ (
);

FILL FILL_1__2033_ (
);

FILL FILL_3__2799_ (
);

FILL FILL_3__2379_ (
);

FILL FILL_5__3666_ (
);

FILL FILL_5__3246_ (
);

FILL FILL_1__3658_ (
);

FILL FILL_1__3238_ (
);

FILL FILL_0__1983_ (
);

FILL FILL_6__2950_ (
);

FILL FILL_6__2530_ (
);

FILL FILL_6__2110_ (
);

FILL FILL_2__2942_ (
);

FILL FILL_2__2522_ (
);

FILL FILL_2__2102_ (
);

FILL FILL_4__2868_ (
);

FILL FILL_4__2448_ (
);

FILL FILL_4__2028_ (
);

FILL FILL_0__2768_ (
);

FILL FILL_0__2348_ (
);

FILL FILL_6__3315_ (
);

FILL FILL_2__3307_ (
);

FILL FILL_5__2937_ (
);

FILL FILL_5__2517_ (
);

FILL FILL_1__2929_ (
);

FILL FILL_1__2509_ (
);

FILL FILL_0_BUFX2_insert10 (
);

FILL FILL_0_BUFX2_insert11 (
);

FILL FILL_2__3480_ (
);

FILL FILL_0_BUFX2_insert12 (
);

OAI21X1 _1999_ (
    .A(_1074_),
    .B(_1109_),
    .C(_1112_),
    .Y(AI[3])
);

FILL FILL_0_BUFX2_insert13 (
);

FILL FILL_2__3060_ (
);

FILL FILL_0_BUFX2_insert14 (
);

FILL FILL_0_BUFX2_insert15 (
);

FILL FILL_0_BUFX2_insert16 (
);

FILL FILL_0_BUFX2_insert17 (
);

FILL FILL_0_BUFX2_insert18 (
);

FILL FILL_0_BUFX2_insert19 (
);

FILL FILL_6__1801_ (
);

AOI21X1 _2940_ (
    .A(_543_),
    .B(_577_),
    .C(_582_),
    .Y(_583_)
);

NOR2X1 _2520_ (
    .A(_212_),
    .B(_214_),
    .Y(_215_)
);

NOR2X1 _2100_ (
    .A(_1208_),
    .B(_1206_),
    .Y(_1209_)
);

FILL FILL169950x50550 (
);

FILL FILL_5__2690_ (
);

FILL FILL_5__2270_ (
);

FILL FILL_7__2288_ (
);

OAI21X1 _3305_ (
    .A(_1091_),
    .B(_869_),
    .C(_871_),
    .Y(_110_)
);

FILL FILL_1__2682_ (
);

FILL FILL_1__2262_ (
);

FILL FILL_3__2188_ (
);

FILL FILL_5__3475_ (
);

FILL FILL_5__3055_ (
);

FILL FILL_1__3467_ (
);

FILL FILL_1__3047_ (
);

FILL FILL_4__1892_ (
);

FILL FILL_0__1792_ (
);

FILL FILL_2__2751_ (
);

FILL FILL_2__2331_ (
);

FILL FILL_4__2677_ (
);

FILL FILL_4__2257_ (
);

FILL FILL_0__2997_ (
);

FILL FILL_0__2577_ (
);

FILL FILL_6__3544_ (
);

FILL FILL_0__2157_ (
);

FILL FILL_6__3124_ (
);

FILL FILL_2__3536_ (
);

FILL FILL_2__3116_ (
);

FILL FILL_7__1979_ (
);

FILL FILL_5__1961_ (
);

FILL FILL168750x32550 (
);

FILL FILL_1__1953_ (
);

FILL FILL_7__2920_ (
);

FILL FILL_7__2500_ (
);

FILL FILL_3__1879_ (
);

FILL FILL_3__2820_ (
);

FILL FILL_3__2400_ (
);

FILL FILL_5__2746_ (
);

FILL FILL_5__2326_ (
);

FILL FILL_1__2738_ (
);

FILL FILL_7__3705_ (
);

FILL FILL_1__2318_ (
);

FILL FILL_3__3605_ (
);

FILL FILL_4__1948_ (
);

FILL FILL_0__1848_ (
);

FILL FILL_6__2815_ (
);

AOI22X1 _3534_ (
    .A(_1716_),
    .B(BI[1]),
    .C(_1563_),
    .D(_1717_),
    .Y(_1564_)
);

NAND3X1 _3114_ (
    .A(_1051_),
    .B(_721_),
    .C(_1053_),
    .Y(_722_)
);

FILL FILL_1__2491_ (
);

FILL FILL_1__2071_ (
);

FILL FILL_2__2807_ (
);

FILL FILL_5__3284_ (
);

FILL FILL_1__3696_ (
);

FILL FILL_1__3276_ (
);

FILL FILL_2__2980_ (
);

FILL FILL_2__2560_ (
);

FILL FILL_2__2140_ (
);

FILL FILL_4__2486_ (
);

FILL FILL_4__2066_ (
);

FILL FILL_0__2386_ (
);

FILL FILL_7__1788_ (
);

FILL FILL_5__1770_ (
);

NOR2X1 _2805_ (
    .A(_362_),
    .B(_340_),
    .Y(_468_)
);

FILL FILL_1__1762_ (
);

FILL FILL_5__2975_ (
);

FILL FILL_5__2555_ (
);

FILL FILL_5__2135_ (
);

FILL FILL_1__2967_ (
);

FILL FILL_1__2547_ (
);

FILL FILL_7__3514_ (
);

FILL FILL_1__2127_ (
);

FILL FILL_2__1831_ (
);

FILL FILL_4__1757_ (
);

FILL FILL_6__2624_ (
);

DFFSR _3343_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_20_),
    .CLK(clk_bF$buf8),
    .Q(cond_code[1])
);

FILL FILL_6__2204_ (
);

FILL FILL_2__2616_ (
);

FILL FILL_5__3093_ (
);

FILL FILL_1__3085_ (
);

FILL FILL_3__1900_ (
);

FILL FILL_5__1826_ (
);

FILL FILL_1__1818_ (
);

FILL FILL_4__2295_ (
);

FILL FILL_6__3582_ (
);

FILL FILL_0__2195_ (
);

FILL FILL_6__3162_ (
);

FILL FILL_2__3574_ (
);

FILL FILL_2__3154_ (
);

INVX1 _2614_ (
    .A(ABH[5]),
    .Y(_296_)
);

FILL FILL_1__1991_ (
);

FILL FILL_5__2784_ (
);

FILL FILL_5__2364_ (
);

FILL FILL_1__2776_ (
);

FILL FILL_1__2356_ (
);

BUFX2 BUFX2_insert20 (
    .A(_1_),
    .Y(_1__bF$buf0)
);

BUFX2 BUFX2_insert21 (
    .A(_914_),
    .Y(_914__bF$buf4)
);

BUFX2 BUFX2_insert22 (
    .A(_914_),
    .Y(_914__bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .A(_914_),
    .Y(_914__bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .A(_914_),
    .Y(_914__bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .A(_914_),
    .Y(_914__bF$buf0)
);

FILL FILL_3__3643_ (
);

FILL FILL_3__3223_ (
);

FILL FILL_5__3569_ (
);

FILL FILL_5__3149_ (
);

FILL FILL_4__1986_ (
);

FILL FILL_0__1886_ (
);

FILL FILL_6__2853_ (
);

OAI21X1 _3572_ (
    .A(_1545_),
    .B(_1549_),
    .C(_1601_),
    .Y(_1602_)
);

FILL FILL_6__2433_ (
);

FILL FILL_6__2013_ (
);

OAI21X1 _3152_ (
    .A(_931__bF$buf2),
    .B(_1075_),
    .C(_173_),
    .Y(_756_)
);

FILL FILL_2__2845_ (
);

FILL FILL_2__2425_ (
);

FILL FILL_2__2005_ (
);

FILL FILL_4__3712_ (
);

FILL FILL_6__3638_ (
);

FILL FILL_6__3218_ (
);

FILL FILL_0__3612_ (
);

FILL FILL_3__2914_ (
);

AND2X2 _2843_ (
    .A(_502_),
    .B(_503_),
    .Y(_504_)
);

NAND3X1 _2423_ (
    .A(_1027__bF$buf3),
    .B(_130_),
    .C(_129_),
    .Y(_131_)
);

NAND3X1 _2003_ (
    .A(_1115_),
    .B(_1113_),
    .C(_1114_),
    .Y(_1116_)
);

FILL FILL_5__2593_ (
);

FILL FILL_5__2173_ (
);

FILL FILL_6__2909_ (
);

OR2X2 _3628_ (
    .A(_1656_),
    .B(_1657_),
    .Y(_1658_)
);

AOI21X1 _3208_ (
    .A(_724_),
    .B(_798_),
    .C(_799_),
    .Y(_85_)
);

FILL FILL_1__2585_ (
);

FILL FILL_1__2165_ (
);

FILL FILL_7__3132_ (
);

FILL FILL_3__3452_ (
);

FILL FILL_3__3032_ (
);

FILL FILL_4__1795_ (
);

FILL FILL_6__2662_ (
);

DFFSR _3381_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(DIMUX[6]),
    .CLK(clk_bF$buf3),
    .Q(DIHOLD[6])
);

FILL FILL_6__2242_ (
);

FILL FILL_2__2654_ (
);

FILL FILL_2__2234_ (
);

FILL FILL_4__3521_ (
);

FILL FILL_4__3101_ (
);

FILL FILL_6__3027_ (
);

FILL FILL_2__3019_ (
);

FILL FILL_0__3001_ (
);

FILL FILL_5__1864_ (
);

FILL FILL_1__1856_ (
);

FILL FILL_7__2403_ (
);

FILL FILL_3__2723_ (
);

FILL FILL_3__2303_ (
);

FILL FILL_5__2649_ (
);

FILL FILL_5__2229_ (
);

FILL FILL_7__3608_ (
);

FILL FILL_2__3192_ (
);

FILL FILL_3__3508_ (
);

FILL FILL_6__1933_ (
);

OAI21X1 _2652_ (
    .A(_914__bF$buf4),
    .B(_954_),
    .C(_1027__bF$buf3),
    .Y(_327_)
);

AOI21X1 _2232_ (
    .A(_886__bF$buf4),
    .B(_1304_),
    .C(_1339_),
    .Y(_1340_)
);

FILL FILL_2__1925_ (
);

FILL FILL_6__2718_ (
);

DFFSR _3437_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(_105_),
    .CLK(clk_bF$buf3),
    .Q(ABL[4])
);

NAND3X1 _3017_ (
    .A(_642_),
    .B(_641_),
    .C(_639_),
    .Y(_643_)
);

FILL FILL_1__2394_ (
);

FILL FILL_3__3261_ (
);

FILL FILL_1_BUFX2_insert80 (
);

FILL FILL_1_BUFX2_insert81 (
);

FILL FILL_1_BUFX2_insert82 (
);

FILL FILL_1_BUFX2_insert83 (
);

FILL FILL_5__3187_ (
);

FILL FILL_1__3599_ (
);

FILL FILL_1__3179_ (
);

FILL FILL_6__2891_ (
);

FILL FILL_6__2471_ (
);

OAI21X1 _3190_ (
    .A(_720__bF$buf3),
    .B(_687_),
    .C(\AXYS[1] [0]),
    .Y(_790_)
);

FILL FILL_6__2051_ (
);

FILL FILL_2__2883_ (
);

FILL FILL_2__2463_ (
);

FILL FILL_2__2043_ (
);

FILL FILL_4__2389_ (
);

OAI21X1 _1923_ (
    .A(_1017_),
    .B(_1036_),
    .C(_1039_),
    .Y(_1040_)
);

FILL FILL_6__3676_ (
);

FILL FILL_0__2289_ (
);

FILL FILL_6__3256_ (
);

FILL FILL_2__3668_ (
);

FILL FILL_0__3650_ (
);

FILL FILL_0__3230_ (
);

FILL FILL_2__3248_ (
);

INVX2 _2708_ (
    .A(_323_),
    .Y(_378_)
);

FILL FILL_7__2632_ (
);

FILL FILL_3__2952_ (
);

FILL FILL_3__2532_ (
);

FILL FILL_3__2112_ (
);

FILL FILL_5__2878_ (
);

FILL FILL_5__2458_ (
);

FILL FILL_5__2038_ (
);

FILL FILL_3__3317_ (
);

NAND2X1 _2881_ (
    .A(_1393_),
    .B(_534_),
    .Y(_535_)
);

NAND3X1 _2461_ (
    .A(_159_),
    .B(_160_),
    .C(_161_),
    .Y(_162_)
);

INVX8 _2041_ (
    .A(_1149__bF$buf0),
    .Y(_1150_)
);

FILL FILL_4__2601_ (
);

FILL FILL_6__2947_ (
);

OAI21X1 _3666_ (
    .A(_1714__bF$buf3),
    .B(_1664_),
    .C(_1690_),
    .Y(_1520_)
);

FILL FILL_6__2527_ (
);

AND2X2 _3246_ (
    .A(_819_),
    .B(_821_),
    .Y(_822_)
);

FILL FILL_6__2107_ (
);

FILL FILL_7__3590_ (
);

FILL FILL_7__3170_ (
);

FILL FILL_0__2921_ (
);

FILL FILL_2__2939_ (
);

FILL FILL_2__2519_ (
);

FILL FILL_0__2501_ (
);

FILL FILL_3__3490_ (
);

FILL FILL_3__3070_ (
);

FILL FILL_7__1903_ (
);

FILL FILL_0__3706_ (
);

FILL FILL_3__1803_ (
);

FILL FILL_6__2280_ (
);

FILL FILL_2__2692_ (
);

FILL FILL_2__2272_ (
);

FILL FILL_4__2198_ (
);

FILL FILL_6__3485_ (
);

FILL FILL_0__2098_ (
);

FILL FILL_6__3065_ (
);

FILL FILL_2__3477_ (
);

FILL FILL_2__3057_ (
);

OR2X2 _2937_ (
    .A(_578_),
    .B(_579_),
    .Y(_580_)
);

NAND3X1 _2517_ (
    .A(_210_),
    .B(_211_),
    .C(_1226_),
    .Y(_212_)
);

FILL FILL_1__1894_ (
);

FILL FILL_7__2861_ (
);

FILL FILL_7__2021_ (
);

FILL FILL_3__2761_ (
);

FILL FILL_3__2341_ (
);

FILL FILL_5__2687_ (
);

FILL FILL_5__2267_ (
);

FILL FILL_1__2679_ (
);

FILL FILL_7__3646_ (
);

FILL FILL_1__2259_ (
);

FILL FILL_1__3620_ (
);

FILL FILL_1__3200_ (
);

FILL FILL_3__3546_ (
);

FILL FILL_3__3126_ (
);

FILL FILL_6__1971_ (
);

OAI22X1 _2690_ (
    .A(_345_),
    .B(_361_),
    .C(_354_),
    .D(_357_),
    .Y(_362_)
);

NAND2X1 _2270_ (
    .A(C),
    .B(cond_code[2]),
    .Y(_1378_)
);

FILL FILL_2__1963_ (
);

FILL FILL_4__1889_ (
);

FILL FILL_4__2830_ (
);

FILL FILL_4__2410_ (
);

FILL FILL_0__1789_ (
);

FILL FILL_6__2756_ (
);

AOI22X1 _3475_ (
    .A(BI[7]),
    .B(_1716_),
    .C(_1720_),
    .D(_1717_),
    .Y(_1721_)
);

FILL FILL_6__2336_ (
);

OAI21X1 _3055_ (
    .A(_1374_),
    .B(_664_),
    .C(_669_),
    .Y(_62_)
);

FILL FILL_2__2748_ (
);

FILL FILL_0__2730_ (
);

FILL FILL_2__2328_ (
);

FILL FILL_0__2310_ (
);

FILL FILL_4__3615_ (
);

FILL FILL_0__3515_ (
);

FILL FILL_5__1958_ (
);

FILL FILL_7__2917_ (
);

FILL FILL_2__2081_ (
);

FILL FILL_3__2817_ (
);

NOR2X1 _1961_ (
    .A(_899_),
    .B(_934_),
    .Y(_1078_)
);

FILL FILL_6__3294_ (
);

FILL FILL_2__3286_ (
);

OAI22X1 _2746_ (
    .A(RDY_bF$buf0),
    .B(_268_),
    .C(_412_),
    .D(_411_),
    .Y(_10_)
);

NAND2X1 _2326_ (
    .A(_886__bF$buf0),
    .B(_990_),
    .Y(_1433_)
);

FILL FILL_7__2670_ (
);

FILL FILL_7__2250_ (
);

FILL FILL_3__2990_ (
);

FILL FILL_3__2570_ (
);

FILL FILL_3__2150_ (
);

FILL FILL_5__2496_ (
);

FILL FILL_5__2076_ (
);

FILL FILL_1__2488_ (
);

FILL FILL_1__2068_ (
);

FILL FILL_7__3035_ (
);

FILL FILL_6__1780_ (
);

FILL FILL169050x32550 (
);

FILL FILL_2__1772_ (
);

FILL FILL_5_BUFX2_insert37 (
);

FILL FILL_5_BUFX2_insert38 (
);

FILL FILL_5_BUFX2_insert39 (
);

FILL FILL_6__2985_ (
);

FILL FILL_6__2565_ (
);

NAND2X1 _3284_ (
    .A(RDY_bF$buf2),
    .B(_859_),
    .Y(_860_)
);

FILL FILL_6__2145_ (
);

FILL FILL_2__2977_ (
);

FILL FILL_2__2557_ (
);

FILL FILL_2__2137_ (
);

FILL FILL_4__3004_ (
);

FILL FILL_3__1841_ (
);

FILL FILL_5__1767_ (
);

FILL FILL_1__1759_ (
);

FILL FILL_7__2306_ (
);

FILL FILL_1__2700_ (
);

FILL FILL_3__2626_ (
);

FILL FILL_3__2206_ (
);

INVX1 _1770_ (
    .A(state[2]),
    .Y(_896_)
);

FILL FILL_2__3095_ (
);

FILL FILL_4__1910_ (
);

FILL FILL_6__1836_ (
);

NOR2X1 _2975_ (
    .A(_1178_),
    .B(_605_),
    .Y(_606_)
);

AOI21X1 _2555_ (
    .A(_216_),
    .B(ADD[4]),
    .C(_245_),
    .Y(_246_)
);

NOR2X1 _2135_ (
    .A(_886__bF$buf6),
    .B(_1241_),
    .Y(_1244_)
);

FILL FILL_0__1810_ (
);

FILL FILL_2__1828_ (
);

FILL FILL_1__2297_ (
);

FILL FILL_7__3264_ (
);

FILL FILL_3__3584_ (
);

FILL FILL_3__3164_ (
);

FILL FILL_6__2794_ (
);

FILL FILL_6__2374_ (
);

NOR2X1 _3093_ (
    .A(adc_sbc),
    .B(compare),
    .Y(_703_)
);

FILL FILL_2__2786_ (
);

FILL FILL_2__2366_ (
);

NOR2X1 _1826_ (
    .A(_904_),
    .B(_924_),
    .Y(_952_)
);

FILL FILL_7__1750_ (
);

FILL FILL_4__3653_ (
);

FILL FILL_4__3233_ (
);

FILL FILL_6__3579_ (
);

FILL FILL_6__3159_ (
);

FILL FILL_0__3553_ (
);

FILL FILL_0__3133_ (
);

FILL FILL_5__1996_ (
);

FILL FILL_1__1988_ (
);

FILL FILL_7__2535_ (
);

FILL FILL_3__2855_ (
);

FILL FILL_3__2435_ (
);

FILL FILL_3__2015_ (
);

FILL FILL_5__3302_ (
);

FILL FILL_1__3714_ (
);

INVX1 _2784_ (
    .A(ABH[3]),
    .Y(_448_)
);

NAND2X1 _2364_ (
    .A(_929_),
    .B(_1031_),
    .Y(_1470_)
);

FILL FILL_4__2924_ (
);

FILL FILL_4__2504_ (
);

INVX1 _3569_ (
    .A(_1598_),
    .Y(_1599_)
);

MUX2X1 _3149_ (
    .A(_753_),
    .B(DIMUX[3]),
    .S(_1018_),
    .Y(_754_)
);

FILL FILL_7__3493_ (
);

FILL FILL_0__2824_ (
);

FILL FILL_0__2404_ (
);

FILL FILL_4__3709_ (
);

FILL FILL_7__1806_ (
);

FILL FILL_0__3609_ (
);

FILL FILL_6__2183_ (
);

FILL FILL_2__2595_ (
);

FILL FILL_2__2175_ (
);

FILL FILL_4__3462_ (
);

FILL FILL_4__3042_ (
);

FILL FILL_6_BUFX2_insert80 (
);

FILL FILL_6_BUFX2_insert81 (
);

FILL FILL_6_BUFX2_insert82 (
);

FILL FILL_6_BUFX2_insert83 (
);

FILL FILL_1__1797_ (
);

FILL FILL_7__2764_ (
);

FILL FILL_3__2664_ (
);

FILL FILL_3__2244_ (
);

FILL FILL_5__3531_ (
);

FILL FILL_5__3111_ (
);

FILL FILL_1__3523_ (
);

FILL FILL_1__3103_ (
);

FILL FILL_3__3449_ (
);

FILL FILL_3__3029_ (
);

FILL FILL_6__1874_ (
);

AOI21X1 _2593_ (
    .A(_272_),
    .B(DIMUX[1]),
    .C(_278_),
    .Y(_279_)
);

OAI21X1 _2173_ (
    .A(RDY_bF$buf8),
    .B(_982_),
    .C(_1281_),
    .Y(_1282_)
);

FILL FILL_2__1866_ (
);

FILL FILL169350x75750 (
);

FILL FILL_4__2733_ (
);

FILL FILL_4__2313_ (
);

FILL FILL_6__2659_ (
);

DFFSR _3378_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(DIMUX[3]),
    .CLK(clk_bF$buf5),
    .Q(DIHOLD[3])
);

FILL FILL_6__2239_ (
);

FILL FILL_0__2633_ (
);

FILL FILL_6__3600_ (
);

FILL FILL_0__2213_ (
);

FILL FILL_4__3518_ (
);

FILL FILL_3__1935_ (
);

FILL FILL_5__2802_ (
);

NAND2X1 _1864_ (
    .A(_927_),
    .B(_910_),
    .Y(_989_)
);

FILL FILL_4__3691_ (
);

FILL FILL_4__3271_ (
);

FILL FILL_6__3197_ (
);

FILL FILL_0__3591_ (
);

FILL FILL_0__3171_ (
);

FILL FILL_2__3189_ (
);

AOI22X1 _2649_ (
    .A(ABL[0]),
    .B(_323_),
    .C(_322_),
    .D(ADD[0]),
    .Y(_324_)
);

NAND2X1 _2229_ (
    .A(_903__bF$buf2),
    .B(_941_),
    .Y(_1337_)
);

FILL FILL_7__2993_ (
);

FILL FILL_7__2153_ (
);

FILL FILL_0__1904_ (
);

FILL FILL_3__2893_ (
);

FILL FILL_3__2473_ (
);

FILL FILL_3__2053_ (
);

FILL FILL_5__2399_ (
);

FILL FILL_3__3678_ (
);

FILL FILL_3__3258_ (
);

FILL FILL_4__2962_ (
);

FILL FILL_4__2542_ (
);

FILL FILL_4__2122_ (
);

FILL FILL_6__2888_ (
);

FILL FILL_6__2468_ (
);

NAND2X1 _3187_ (
    .A(\AXYS[0] [7]),
    .B(_722_),
    .Y(_788_)
);

FILL FILL_6__2048_ (
);

FILL FILL_0__2862_ (
);

FILL FILL_0__2442_ (
);

FILL FILL_0__2022_ (
);

FILL FILL_3__1744_ (
);

FILL FILL_0__3647_ (
);

FILL FILL_0__3227_ (
);

FILL FILL_5__2611_ (
);

FILL FILL_7__2629_ (
);

FILL FILL_7__2209_ (
);

FILL FILL_1__2603_ (
);

FILL FILL_3__2949_ (
);

FILL FILL_3__2529_ (
);

FILL FILL_3__2109_ (
);

FILL FILL_4__3080_ (
);

FILL FILL_4__1813_ (
);

OAI21X1 _2878_ (
    .A(_529_),
    .B(_1150__bF$buf2),
    .C(_532_),
    .Y(_22_)
);

NAND2X1 _2458_ (
    .A(ADD[2]),
    .B(_144_),
    .Y(_159_)
);

AOI21X1 _2038_ (
    .A(_1082_),
    .B(AN),
    .C(_1147_),
    .Y(_1148_)
);

FILL FILL_7__2382_ (
);

FILL FILL_3__2282_ (
);

FILL FILL_7__3587_ (
);

FILL FILL_7__3167_ (
);

FILL FILL_0__2918_ (
);

FILL FILL_1__3561_ (
);

FILL FILL_1__3141_ (
);

FILL FILL_3__3487_ (
);

FILL FILL_3__3067_ (
);

FILL FILL_4__2771_ (
);

FILL FILL_4__2351_ (
);

FILL FILL_6__2697_ (
);

FILL FILL_6__2277_ (
);

FILL FILL_2__2689_ (
);

FILL FILL_0__2671_ (
);

FILL FILL_2__2269_ (
);

FILL FILL_0__2251_ (
);

FILL FILL_2__3630_ (
);

FILL FILL_2__3210_ (
);

FILL FILL169650x100950 (
);

FILL FILL_4__3556_ (
);

FILL FILL_4__3136_ (
);

FILL FILL_3__1973_ (
);

FILL FILL_0__3456_ (
);

FILL FILL_0__3036_ (
);

FILL FILL_5__1899_ (
);

FILL FILL_5__2840_ (
);

FILL FILL_7__2438_ (
);

FILL FILL_5__2420_ (
);

FILL FILL_5__2000_ (
);

FILL FILL_1__2832_ (
);

FILL FILL_1__2412_ (
);

FILL FILL_3__2758_ (
);

FILL FILL_3__2338_ (
);

FILL FILL_5__3625_ (
);

FILL FILL_5__3205_ (
);

FILL FILL_1__3617_ (
);

FILL FILL_6__1968_ (
);

INVX1 _2687_ (
    .A(_358_),
    .Y(_359_)
);

NAND2X1 _2267_ (
    .A(cond_code[2]),
    .B(Z),
    .Y(_1375_)
);

FILL FILL_0__1942_ (
);

FILL FILL_3__2091_ (
);

FILL FILL_2__2901_ (
);

FILL FILL_4__2827_ (
);

FILL FILL_4__2407_ (
);

FILL FILL_0__2727_ (
);

FILL FILL_0__2307_ (
);

FILL FILL_3__3296_ (
);

FILL FILL_4__2580_ (
);

FILL FILL_4__2160_ (
);

FILL FILL_6__2086_ (
);

FILL FILL_0__2480_ (
);

FILL FILL_2__2498_ (
);

FILL FILL_0__2060_ (
);

FILL FILL_2__2078_ (
);

NAND2X1 _1958_ (
    .A(_948_),
    .B(_957_),
    .Y(_1075_)
);

FILL FILL_7__1882_ (
);

FILL FILL_3__1782_ (
);

FILL FILL_0__3265_ (
);

FILL FILL_7__2667_ (
);

FILL FILL_1__2641_ (
);

FILL FILL_1__2221_ (
);

FILL FILL_3__2987_ (
);

FILL FILL_3__2567_ (
);

FILL FILL_3__2147_ (
);

FILL FILL_5__3014_ (
);

FILL FILL_1__3006_ (
);

FILL FILL_4__1851_ (
);

FILL FILL_6__1777_ (
);

INVX1 _2496_ (
    .A(_191_),
    .Y(_192_)
);

NAND2X1 _2076_ (
    .A(_1167_),
    .B(_1184_),
    .Y(_1185_)
);

FILL FILL_0__1751_ (
);

FILL FILL_2__1769_ (
);

FILL FILL_2__2710_ (
);

FILL FILL_4__2636_ (
);

FILL FILL_4__2216_ (
);

FILL FILL_0__2956_ (
);

FILL FILL_0__2536_ (
);

FILL FILL_6__3503_ (
);

FILL FILL_0__2116_ (
);

FILL FILL_5__1920_ (
);

FILL FILL_7__1938_ (
);

FILL FILL_1__1912_ (
);

FILL FILL_3__1838_ (
);

FILL FILL_5__2705_ (
);

INVX1 _1767_ (
    .A(_893_),
    .Y(DIMUX[7])
);

FILL FILL_4__3594_ (
);

FILL FILL_4__3174_ (
);

FILL FILL_0__3494_ (
);

FILL FILL_0__3074_ (
);

FILL FILL_4__1907_ (
);

FILL FILL_7__2896_ (
);

FILL FILL_7__2056_ (
);

FILL FILL_0__1807_ (
);

FILL FILL_1__2870_ (
);

FILL FILL_1__2450_ (
);

FILL FILL_1__2030_ (
);

FILL FILL_3__2796_ (
);

FILL FILL_3__2376_ (
);

FILL FILL_5__3663_ (
);

FILL FILL_5__3243_ (
);

FILL FILL_1__3655_ (
);

FILL FILL_1__3235_ (
);

FILL FILL_0__1980_ (
);

FILL FILL_2__1998_ (
);

FILL FILL_4__2865_ (
);

FILL FILL_4__2445_ (
);

FILL FILL_4__2025_ (
);

FILL FILL_0__2765_ (
);

FILL FILL_0__2345_ (
);

FILL FILL_6__3312_ (
);

FILL FILL_2__3304_ (
);

FILL FILL_7__1747_ (
);

FILL FILL_1_CLKBUF1_insert26 (
);

FILL FILL_1_CLKBUF1_insert27 (
);

FILL FILL_1_CLKBUF1_insert28 (
);

FILL FILL_1_CLKBUF1_insert29 (
);

FILL FILL_5__2934_ (
);

FILL FILL_5__2514_ (
);

FILL FILL_1__2926_ (
);

FILL FILL_1__2506_ (
);

NAND2X1 _1996_ (
    .A(ABH[3]),
    .B(_925_),
    .Y(_1110_)
);

FILL FILL_7__2285_ (
);

NAND2X1 _3302_ (
    .A(_1741_[8]),
    .B(_869_),
    .Y(_870_)
);

FILL FILL_3__2185_ (
);

FILL FILL_5__3472_ (
);

FILL FILL_5__3052_ (
);

FILL FILL_1__3464_ (
);

FILL FILL_1__3044_ (
);

FILL FILL_4__2674_ (
);

FILL FILL_4__2254_ (
);

FILL FILL_0__2994_ (
);

FILL FILL_0__2574_ (
);

FILL FILL_6__3541_ (
);

FILL FILL_0__2154_ (
);

FILL FILL_6__3121_ (
);

FILL FILL_2__3533_ (
);

FILL FILL_2__3113_ (
);

FILL FILL_7__1976_ (
);

FILL FILL_4__3459_ (
);

FILL FILL_4__3039_ (
);

FILL FILL_1__1950_ (
);

FILL FILL_3__1876_ (
);

FILL FILL_5__2743_ (
);

FILL FILL_5__2323_ (
);

FILL FILL_1__2735_ (
);

FILL FILL_7__3702_ (
);

FILL FILL_1__2315_ (
);

FILL FILL_3__3602_ (
);

FILL FILL_5__3528_ (
);

FILL FILL_5__3108_ (
);

FILL FILL_4__1945_ (
);

FILL FILL_0__1845_ (
);

FILL FILL_6__2812_ (
);

NAND2X1 _3531_ (
    .A(_1560_),
    .B(_1557_),
    .Y(_1561_)
);

NOR2X1 _3111_ (
    .A(_633_),
    .B(_662_),
    .Y(_719_)
);

FILL FILL_2__2804_ (
);

FILL FILL_7__3299_ (
);

FILL FILL_5__3281_ (
);

FILL FILL_1__3693_ (
);

FILL FILL_1__3273_ (
);

FILL FILL_3__3199_ (
);

FILL FILL_4__2483_ (
);

FILL FILL_4__2063_ (
);

FILL FILL_0__2383_ (
);

FILL FILL_7__1785_ (
);

FILL FILL_4__3268_ (
);

NOR2X1 _2802_ (
    .A(_464_),
    .B(_463_),
    .Y(_465_)
);

FILL FILL_0__3588_ (
);

FILL FILL_0__3168_ (
);

FILL FILL_5__2972_ (
);

FILL FILL_5__2552_ (
);

FILL FILL_5__2132_ (
);

FILL FILL_1__2964_ (
);

FILL FILL_1__2544_ (
);

FILL FILL_7__3511_ (
);

FILL FILL_1__2124_ (
);

FILL FILL_4__1754_ (
);

INVX1 _2399_ (
    .A(_1466_),
    .Y(_1504_)
);

FILL FILL_6__2621_ (
);

DFFSR _3340_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(NMI),
    .CLK(clk_bF$buf4),
    .Q(NMI_1)
);

FILL FILL_6__2201_ (
);

FILL FILL_2__2613_ (
);

FILL FILL_4__2959_ (
);

FILL FILL_4__2539_ (
);

FILL FILL_4__2119_ (
);

FILL FILL_5__3090_ (
);

FILL FILL_0__2859_ (
);

FILL FILL_0__2439_ (
);

FILL FILL_0__2019_ (
);

FILL FILL_1__3082_ (
);

FILL FILL_5__1823_ (
);

FILL FILL_1__1815_ (
);

FILL FILL_4__2292_ (
);

FILL FILL_5__2608_ (
);

FILL FILL_0__2192_ (
);

FILL FILL_2__3571_ (
);

FILL FILL_2__3151_ (
);

FILL FILL_4__3497_ (
);

FILL FILL_4__3077_ (
);

AOI21X1 _2611_ (
    .A(_272_),
    .B(DIMUX[4]),
    .C(_293_),
    .Y(_294_)
);

FILL FILL_7__2799_ (
);

FILL FILL_5__2781_ (
);

FILL FILL_5__2361_ (
);

FILL FILL_7__2379_ (
);

FILL FILL_1__2773_ (
);

FILL FILL_1__2353_ (
);

FILL FILL_3__2699_ (
);

FILL FILL_3__2279_ (
);

FILL FILL_3__3640_ (
);

FILL FILL_3__3220_ (
);

FILL FILL_5__3566_ (
);

FILL FILL_5__3146_ (
);

FILL FILL_1__3558_ (
);

FILL FILL_1__3138_ (
);

FILL FILL_4__1983_ (
);

FILL FILL_0__1883_ (
);

FILL FILL_6__2850_ (
);

FILL FILL_6__2430_ (
);

FILL FILL_6__2010_ (
);

FILL FILL168150x150 (
);

FILL FILL_2__2842_ (
);

FILL FILL_2__2422_ (
);

FILL FILL_2__2002_ (
);

FILL FILL_4__2768_ (
);

FILL FILL_4__2348_ (
);

FILL FILL_0__2668_ (
);

FILL FILL_6__3635_ (
);

FILL FILL_0__2248_ (
);

FILL FILL_6__3215_ (
);

FILL FILL_2__3627_ (
);

FILL FILL_2__3207_ (
);

FILL FILL_3__2911_ (
);

FILL FILL_5__2837_ (
);

FILL FILL_5__2417_ (
);

FILL FILL_1__2829_ (
);

FILL FILL_1__2409_ (
);

OAI22X1 _1899_ (
    .A(_1016_),
    .B(_968_),
    .C(_893_),
    .D(_1004_),
    .Y(BI[7])
);

NOR2X1 _2840_ (
    .A(_300_),
    .B(_418_),
    .Y(_501_)
);

INVX1 _2420_ (
    .A(op[0]),
    .Y(_128_)
);

NAND2X1 _2000_ (
    .A(\AXYS[1] [4]),
    .B(_1047_),
    .Y(_1113_)
);

FILL FILL_5__2590_ (
);

FILL FILL_7__2188_ (
);

FILL FILL_5__2170_ (
);

FILL FILL_0__1939_ (
);

FILL FILL_6__2906_ (
);

NAND2X1 _3625_ (
    .A(_1654_),
    .B(_1639_),
    .Y(_1655_)
);

OAI21X1 _3205_ (
    .A(_787_),
    .B(_789_),
    .C(_797_),
    .Y(_84_)
);

FILL FILL_1__2582_ (
);

FILL FILL_1__2162_ (
);

FILL FILL_3__2088_ (
);

FILL FILL_4__1792_ (
);

FILL FILL_2__2651_ (
);

FILL FILL_2__2231_ (
);

FILL FILL_4__2997_ (
);

FILL FILL_4__2577_ (
);

FILL FILL_4__2157_ (
);

FILL FILL_0__2897_ (
);

FILL FILL_0__2477_ (
);

FILL FILL_0__2057_ (
);

FILL FILL_6__3024_ (
);

FILL FILL_2__3016_ (
);

FILL FILL_7__1879_ (
);

FILL FILL_5__1861_ (
);

FILL FILL_1__1853_ (
);

FILL FILL_7__2820_ (
);

FILL FILL_7__2400_ (
);

FILL FILL_3__1779_ (
);

FILL FILL_3__2720_ (
);

FILL FILL_3__2300_ (
);

FILL FILL_5__2646_ (
);

FILL FILL_5__2226_ (
);

FILL FILL_1__2638_ (
);

FILL FILL_1__2218_ (
);

FILL FILL_3__3505_ (
);

FILL FILL_6__1930_ (
);

FILL FILL_2__1922_ (
);

FILL FILL_4__1848_ (
);

FILL FILL_0__1748_ (
);

FILL FILL_6__2715_ (
);

DFFSR _3434_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_102_),
    .CLK(clk_bF$buf1),
    .Q(ABL[1])
);

INVX1 _3014_ (
    .A(_551_),
    .Y(_640_)
);

FILL FILL_1__2391_ (
);

FILL FILL_2__2707_ (
);

FILL FILL_1_BUFX2_insert50 (
);

FILL FILL_1_BUFX2_insert51 (
);

FILL FILL_1_BUFX2_insert52 (
);

FILL FILL_1_BUFX2_insert53 (
);

FILL FILL_5__3184_ (
);

FILL FILL_1_BUFX2_insert54 (
);

FILL FILL_1_BUFX2_insert55 (
);

FILL FILL_1_BUFX2_insert56 (
);

FILL FILL_1_BUFX2_insert57 (
);

FILL FILL_1_BUFX2_insert58 (
);

FILL FILL_1_BUFX2_insert59 (
);

FILL FILL_1__3596_ (
);

FILL FILL_1__3176_ (
);

FILL FILL_0_CLKBUF1_insert30 (
);

FILL FILL_0_CLKBUF1_insert31 (
);

FILL FILL_5__1917_ (
);

FILL FILL_0_CLKBUF1_insert32 (
);

FILL FILL_0_CLKBUF1_insert33 (
);

FILL FILL_0_CLKBUF1_insert34 (
);

FILL FILL_0_CLKBUF1_insert35 (
);

FILL FILL_0_CLKBUF1_insert36 (
);

FILL FILL_1__1909_ (
);

FILL FILL_2__2880_ (
);

FILL FILL_2__2460_ (
);

FILL FILL_2__2040_ (
);

FILL FILL_4__2386_ (
);

INVX1 _1920_ (
    .A(_1027__bF$buf0),
    .Y(_1037_)
);

FILL FILL_6__3673_ (
);

FILL FILL_0__2286_ (
);

FILL FILL_6__3253_ (
);

FILL FILL_2__3665_ (
);

FILL FILL_2__3245_ (
);

OAI21X1 _2705_ (
    .A(_374_),
    .B(_370_),
    .C(RDY_bF$buf3),
    .Y(_376_)
);

FILL FILL_5__2875_ (
);

FILL FILL_5__2455_ (
);

FILL FILL_5__2035_ (
);

FILL FILL_1__2867_ (
);

FILL FILL_1__2447_ (
);

FILL FILL_1__2027_ (
);

FILL FILL_3__3314_ (
);

FILL FILL_0__1977_ (
);

FILL FILL_6__2944_ (
);

NAND2X1 _3663_ (
    .A(ADD[2]),
    .B(_1714__bF$buf1),
    .Y(_1689_)
);

FILL FILL_6__2524_ (
);

NOR2X1 _3243_ (
    .A(_818_),
    .B(_817_),
    .Y(_819_)
);

FILL FILL_6__2104_ (
);

FILL FILL_2__2936_ (
);

FILL FILL_2__2516_ (
);

FILL FILL_7__1900_ (
);

FILL FILL_6__3309_ (
);

FILL FILL_3__1800_ (
);

FILL FILL_0__3703_ (
);

FILL FILL_4__2195_ (
);

FILL FILL_6__3482_ (
);

FILL FILL_0__2095_ (
);

FILL FILL_6__3062_ (
);

FILL FILL_2__3474_ (
);

FILL FILL_2__3054_ (
);

OAI21X1 _2934_ (
    .A(_1181_),
    .B(_576_),
    .C(_1215_),
    .Y(_577_)
);

NAND2X1 _2514_ (
    .A(_208_),
    .B(_206_),
    .Y(_209_)
);

FILL FILL_1__1891_ (
);

FILL FILL_5__2684_ (
);

FILL FILL_5__2264_ (
);

FILL FILL_1__2676_ (
);

FILL FILL_7__3643_ (
);

FILL FILL_1__2256_ (
);

FILL FILL_3__3543_ (
);

FILL FILL_3__3123_ (
);

FILL FILL_5__3469_ (
);

FILL FILL_5__3049_ (
);

FILL FILL_2__1960_ (
);

FILL FILL_4__1886_ (
);

FILL FILL_0__1786_ (
);

FILL FILL_6__2753_ (
);

INVX2 _3472_ (
    .A(alu_op[0]),
    .Y(_1718_)
);

FILL FILL_6__2333_ (
);

OAI21X1 _3052_ (
    .A(_1027__bF$buf3),
    .B(_666_),
    .C(_665_),
    .Y(_667_)
);

FILL FILL_2__2745_ (
);

FILL FILL_2__2325_ (
);

FILL FILL_4__3612_ (
);

FILL FILL_6__3538_ (
);

FILL FILL_6__3118_ (
);

FILL FILL_0__3512_ (
);

FILL FILL_5__1955_ (
);

FILL FILL_1__1947_ (
);

FILL FILL_7__2914_ (
);

FILL FILL_3__2814_ (
);

FILL FILL_6__3291_ (
);

FILL FILL_2__3283_ (
);

INVX1 _2743_ (
    .A(_409_),
    .Y(_410_)
);

INVX1 _2323_ (
    .A(_1384_),
    .Y(_1430_)
);

FILL FILL_5__2493_ (
);

FILL FILL_5__2073_ (
);

FILL FILL_6__2809_ (
);

NOR2X1 _3528_ (
    .A(alu_op[3]),
    .B(alu_op[2]),
    .Y(_1558_)
);

OAI21X1 _3108_ (
    .A(RDY_bF$buf9),
    .B(_715_),
    .C(_716_),
    .Y(_68_)
);

FILL FILL_1__2485_ (
);

FILL FILL_1__2065_ (
);

FILL FILL_7__3032_ (
);

FILL FILL_5__3698_ (
);

FILL FILL_5__3278_ (
);

FILL FILL_6__2982_ (
);

FILL FILL_6__2562_ (
);

OAI21X1 _3281_ (
    .A(state[4]),
    .B(_981_),
    .C(_856_),
    .Y(_857_)
);

FILL FILL_6__2142_ (
);

FILL FILL_2__2974_ (
);

FILL FILL_2__2554_ (
);

FILL FILL_2__2134_ (
);

FILL FILL_4__3001_ (
);

FILL FILL_5__1764_ (
);

FILL FILL_1__1756_ (
);

FILL FILL_7__2303_ (
);

FILL FILL_3__2623_ (
);

FILL FILL_3__2203_ (
);

FILL FILL_5__2969_ (
);

FILL FILL_5__2549_ (
);

FILL FILL_5__2129_ (
);

FILL FILL_7__3508_ (
);

FILL FILL_2__3092_ (
);

FILL FILL_6__1833_ (
);

OAI21X1 _2972_ (
    .A(_1405_),
    .B(_603_),
    .C(_534_),
    .Y(_604_)
);

NAND2X1 _2552_ (
    .A(ADD[4]),
    .B(_209_),
    .Y(_243_)
);

OR2X2 _2132_ (
    .A(CO),
    .B(store),
    .Y(_1241_)
);

FILL FILL_2__1825_ (
);

FILL FILL_6__2618_ (
);

DFFSR _3337_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_15_),
    .CLK(clk_bF$buf2),
    .Q(PC[13])
);

FILL FILL_1__2294_ (
);

FILL FILL_7__3261_ (
);

FILL FILL_3__3581_ (
);

FILL FILL_3__3161_ (
);

FILL FILL_5__3087_ (
);

FILL FILL_1__3499_ (
);

FILL FILL_1__3079_ (
);

FILL FILL_6__2791_ (
);

FILL FILL_6__2371_ (
);

MUX2X1 _3090_ (
    .A(_700_),
    .B(AZ),
    .S(_1227_),
    .Y(_701_)
);

FILL FILL_2__2783_ (
);

FILL FILL_2__2363_ (
);

FILL FILL_4__2289_ (
);

NAND2X1 _1823_ (
    .A(_910_),
    .B(_948_),
    .Y(_949_)
);

FILL FILL_4__3650_ (
);

FILL FILL_4__3230_ (
);

FILL FILL_0__2189_ (
);

FILL FILL_6__3576_ (
);

FILL FILL_6__3156_ (
);

FILL FILL_2__3568_ (
);

FILL FILL_0__3550_ (
);

FILL FILL_2__3148_ (
);

FILL FILL_0__3130_ (
);

FILL FILL_5__1993_ (
);

INVX1 _2608_ (
    .A(ABH[4]),
    .Y(_291_)
);

FILL FILL_1__1985_ (
);

FILL FILL_7__2532_ (
);

FILL FILL_3__2852_ (
);

FILL FILL_3__2432_ (
);

FILL FILL_3__2012_ (
);

FILL FILL_5__2778_ (
);

FILL FILL_5__2358_ (
);

FILL FILL_7__3317_ (
);

FILL FILL_1__3711_ (
);

FILL FILL_3__3637_ (
);

FILL FILL_3__3217_ (
);

OAI21X1 _2781_ (
    .A(_1291_),
    .B(_325_),
    .C(DIMUX[3]),
    .Y(_445_)
);

NAND2X1 _2361_ (
    .A(_903__bF$buf3),
    .B(_1031_),
    .Y(_1467_)
);

FILL FILL_4__2921_ (
);

FILL FILL_4__2501_ (
);

FILL FILL_6__2847_ (
);

NAND2X1 _3566_ (
    .A(_1725_),
    .B(_1560_),
    .Y(_1596_)
);

FILL FILL_6__2427_ (
);

FILL FILL_6__2007_ (
);

AND2X2 _3146_ (
    .A(_747_),
    .B(_750_),
    .Y(_751_)
);

FILL FILL_7__3490_ (
);

FILL FILL_7__3070_ (
);

FILL FILL_2__2839_ (
);

FILL FILL_0__2821_ (
);

FILL FILL_2__2419_ (
);

FILL FILL_0__2401_ (
);

FILL FILL_4__3706_ (
);

FILL FILL_7__1803_ (
);

FILL FILL_0__3606_ (
);

FILL FILL_6__2180_ (
);

FILL FILL_2__2592_ (
);

FILL FILL_2__2172_ (
);

FILL FILL_4__2098_ (
);

FILL FILL_3__2908_ (
);

FILL FILL_6_BUFX2_insert50 (
);

FILL FILL_6_BUFX2_insert51 (
);

FILL FILL_6_BUFX2_insert52 (
);

FILL FILL_6_BUFX2_insert53 (
);

FILL FILL_6_BUFX2_insert54 (
);

FILL FILL_6_BUFX2_insert55 (
);

FILL FILL_6_BUFX2_insert56 (
);

FILL FILL_6_BUFX2_insert57 (
);

FILL FILL_6_BUFX2_insert58 (
);

FILL FILL_6_BUFX2_insert59 (
);

OAI21X1 _2837_ (
    .A(_498_),
    .B(_496_),
    .C(RDY_bF$buf4),
    .Y(_499_)
);

NAND2X1 _2417_ (
    .A(_1282_),
    .B(_125_),
    .Y(_126_)
);

FILL FILL_1__1794_ (
);

FILL FILL_7__2761_ (
);

FILL FILL_3__2661_ (
);

FILL FILL_3__2241_ (
);

FILL FILL_5__2587_ (
);

FILL FILL_5__2167_ (
);

FILL FILL_1__2999_ (
);

FILL FILL_1__2579_ (
);

FILL FILL_7__3546_ (
);

FILL FILL_1__2159_ (
);

FILL FILL_1__3520_ (
);

FILL FILL_1__3100_ (
);

FILL FILL_3__3026_ (
);

FILL FILL_6__1871_ (
);

INVX1 _2590_ (
    .A(PC[9]),
    .Y(_276_)
);

NOR2X1 _2170_ (
    .A(_1266_),
    .B(_1278_),
    .Y(_1279_)
);

FILL FILL_2__1863_ (
);

FILL FILL_4__1789_ (
);

FILL FILL_4__2730_ (
);

FILL FILL_4__2310_ (
);

FILL FILL_6__2656_ (
);

DFFSR _3375_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(DIMUX[0]),
    .CLK(clk_bF$buf5),
    .Q(DIHOLD[0])
);

FILL FILL_6__2236_ (
);

FILL FILL_2__2648_ (
);

FILL FILL_0__2630_ (
);

FILL FILL_0__2210_ (
);

FILL FILL_2__2228_ (
);

FILL FILL_4__3515_ (
);

FILL FILL_3__1932_ (
);

FILL FILL_5__1858_ (
);

FILL FILL_7__2817_ (
);

FILL FILL_3__2717_ (
);

INVX1 _1861_ (
    .A(_985_),
    .Y(_986_)
);

FILL FILL_6__3194_ (
);

FILL FILL_2__3186_ (
);

FILL FILL_6__1927_ (
);

OAI22X1 _2646_ (
    .A(_903__bF$buf1),
    .B(_969_),
    .C(_1221_),
    .D(_1427_),
    .Y(_321_)
);

NOR2X1 _2226_ (
    .A(_914__bF$buf0),
    .B(_1075_),
    .Y(_1334_)
);

FILL FILL_7__2990_ (
);

FILL FILL_7__2570_ (
);

FILL FILL_7__2150_ (
);

FILL FILL_0__1901_ (
);

FILL FILL_2__1919_ (
);

FILL FILL_3__2890_ (
);

FILL FILL_3__2470_ (
);

FILL FILL_3__2050_ (
);

FILL FILL_5__2396_ (
);

FILL FILL_1__2388_ (
);

FILL FILL_3__3675_ (
);

FILL FILL_3__3255_ (
);

FILL FILL_6__2885_ (
);

FILL FILL_6__2465_ (
);

FILL FILL_6__2045_ (
);

OAI21X1 _3184_ (
    .A(_784_),
    .B(_780_),
    .C(_1018_),
    .Y(_785_)
);

FILL FILL_2__2877_ (
);

FILL FILL_2__2457_ (
);

FILL FILL_2__2037_ (
);

NOR2X1 _1917_ (
    .A(_1029_),
    .B(_1033_),
    .Y(_1034_)
);

FILL FILL_0__3644_ (
);

FILL FILL_0__3224_ (
);

FILL FILL169650x3750 (
);

FILL FILL_7__2206_ (
);

FILL FILL_1__2600_ (
);

FILL FILL_3__2946_ (
);

FILL FILL_3__2526_ (
);

FILL FILL_3__2106_ (
);

FILL FILL_4__1810_ (
);

INVX2 _2875_ (
    .A(_1251_),
    .Y(_530_)
);

NAND3X1 _2455_ (
    .A(_153_),
    .B(_156_),
    .C(_155_),
    .Y(_157_)
);

NOR2X1 _2035_ (
    .A(_1144_),
    .B(_1092_),
    .Y(_1145_)
);

FILL FILL_1__2197_ (
);

FILL FILL_7__3164_ (
);

FILL FILL_0__2915_ (
);

FILL FILL_3__3484_ (
);

FILL FILL_3__3064_ (
);

FILL FILL_6__2694_ (
);

FILL FILL_6__2274_ (
);

FILL FILL_2__2686_ (
);

FILL FILL_2__2266_ (
);

FILL FILL_4__3553_ (
);

FILL FILL_4__3133_ (
);

FILL FILL_6__3479_ (
);

FILL FILL_6__3059_ (
);

FILL FILL_3__1970_ (
);

FILL FILL_0__3453_ (
);

FILL FILL_0__3033_ (
);

FILL FILL_5__1896_ (
);

FILL FILL_1__1888_ (
);

FILL FILL_7__2435_ (
);

FILL FILL_3__2755_ (
);

FILL FILL_3__2335_ (
);

FILL FILL_5__3622_ (
);

FILL FILL_5__3202_ (
);

FILL FILL_1__3614_ (
);

FILL FILL_6__1965_ (
);

AOI21X1 _2684_ (
    .A(ABL[3]),
    .B(_323_),
    .C(_1334_),
    .Y(_356_)
);

OAI21X1 _2264_ (
    .A(RDY_bF$buf5),
    .B(_936_),
    .C(_1371_),
    .Y(_1372_)
);

FILL FILL_2__1957_ (
);

FILL FILL_4__2824_ (
);

FILL FILL_4__2404_ (
);

NAND2X1 _3469_ (
    .A(CI),
    .B(alu_shift_right),
    .Y(_1715_)
);

AOI21X1 _3049_ (
    .A(_308_),
    .B(_663_),
    .C(_660_),
    .Y(_664_)
);

FILL FILL_0__2724_ (
);

FILL FILL_0__2304_ (
);

FILL FILL_3__3293_ (
);

FILL FILL_4__3609_ (
);

FILL FILL_0__3509_ (
);

FILL FILL_6__2083_ (
);

FILL FILL_2__2495_ (
);

FILL FILL_2__2075_ (
);

NOR2X1 _1955_ (
    .A(_1029_),
    .B(_918_),
    .Y(_1072_)
);

FILL FILL_6__3288_ (
);

FILL FILL_0__3262_ (
);

FILL FILL_7__2664_ (
);

FILL FILL_3__2984_ (
);

FILL FILL_3__2564_ (
);

FILL FILL_3__2144_ (
);

FILL FILL_5__3011_ (
);

FILL FILL_1__3003_ (
);

FILL FILL_6__1774_ (
);

OAI21X1 _2493_ (
    .A(_1016_),
    .B(_136_),
    .C(_188_),
    .Y(_189_)
);

NOR2X1 _2073_ (
    .A(_1181_),
    .B(_1179_),
    .Y(_1182_)
);

FILL FILL_2__1766_ (
);

FILL FILL_4__2633_ (
);

FILL FILL_4__2213_ (
);

FILL FILL_6__2979_ (
);

BUFX2 _3698_ (
    .A(_1741_[15]),
    .Y(AB[15])
);

FILL FILL_6__2559_ (
);

NAND3X1 _3278_ (
    .A(_852_),
    .B(_853_),
    .C(_822_),
    .Y(_854_)
);

FILL FILL_6__2139_ (
);

FILL FILL_0__2953_ (
);

FILL FILL_0__2533_ (
);

FILL FILL_6__3500_ (
);

FILL FILL_0__2113_ (
);

FILL FILL_7__1935_ (
);

FILL FILL_3__1835_ (
);

FILL FILL_5__2702_ (
);

NAND2X1 _1764_ (
    .A(RDY_bF$buf9),
    .B(DI[6]),
    .Y(_892_)
);

FILL FILL_4__3591_ (
);

FILL FILL_4__3171_ (
);

FILL FILL_6__3097_ (
);

FILL FILL_0__3491_ (
);

FILL FILL_2__3089_ (
);

FILL FILL_0__3071_ (
);

FILL FILL_4__1904_ (
);

INVX1 _2969_ (
    .A(_589_),
    .Y(_601_)
);

OAI21X1 _2549_ (
    .A(_1009_),
    .B(_218_),
    .C(_240_),
    .Y(_241_)
);

NAND2X1 _2129_ (
    .A(RDY_bF$buf8),
    .B(_990_),
    .Y(_1238_)
);

FILL FILL_7__2893_ (
);

FILL FILL_7__2053_ (
);

FILL FILL_0__1804_ (
);

FILL FILL_3__2793_ (
);

FILL FILL_3__2373_ (
);

FILL FILL_5__2299_ (
);

FILL FILL_5__3660_ (
);

FILL FILL_5__3240_ (
);

FILL FILL_1__3652_ (
);

FILL FILL_1__3232_ (
);

FILL FILL_3__3578_ (
);

FILL FILL_3__3158_ (
);

FILL FILL_2__1995_ (
);

FILL FILL_4__2862_ (
);

FILL FILL_4__2442_ (
);

FILL FILL_4__2022_ (
);

FILL FILL_6__2788_ (
);

FILL FILL_6__2368_ (
);

AOI22X1 _3087_ (
    .A(_1227_),
    .B(_658_),
    .C(_689_),
    .D(_656_),
    .Y(_698_)
);

FILL FILL_0__2762_ (
);

FILL FILL_0__2342_ (
);

FILL FILL_2__3301_ (
);

FILL FILL_4__3647_ (
);

FILL FILL_4__3227_ (
);

FILL FILL_0__3547_ (
);

FILL FILL_0__3127_ (
);

FILL FILL_7__2949_ (
);

FILL FILL_5__2931_ (
);

FILL FILL_7__2529_ (
);

FILL FILL_5__2511_ (
);

FILL FILL_7__2109_ (
);

FILL FILL_1__2923_ (
);

FILL FILL_1__2503_ (
);

FILL FILL_3__2849_ (
);

FILL FILL_3__2429_ (
);

FILL FILL_3__2009_ (
);

NAND3X1 _1993_ (
    .A(\AXYS[0] [3]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1107_)
);

FILL FILL169350x61350 (
);

FILL FILL169950x100950 (
);

FILL FILL_1__3708_ (
);

OAI21X1 _2778_ (
    .A(_365_),
    .B(_442_),
    .C(_441_),
    .Y(_443_)
);

NOR2X1 _2358_ (
    .A(_931__bF$buf0),
    .B(_1272_),
    .Y(_1464_)
);

FILL FILL_7__2282_ (
);

FILL FILL_3__2182_ (
);

FILL FILL_4__2918_ (
);

FILL FILL_7__3487_ (
);

FILL FILL_7__3067_ (
);

FILL FILL_0__2818_ (
);

FILL FILL_1__3461_ (
);

FILL FILL_1__3041_ (
);

FILL FILL_4__2671_ (
);

FILL FILL_4__2251_ (
);

FILL FILL_6__2597_ (
);

FILL FILL_6__2177_ (
);

FILL FILL_0__2991_ (
);

FILL FILL_2__2589_ (
);

FILL FILL_0__2571_ (
);

FILL FILL_0__2151_ (
);

FILL FILL_2__2169_ (
);

FILL FILL_2__3530_ (
);

FILL FILL_2__3110_ (
);

FILL FILL_4__3456_ (
);

FILL FILL_4__3036_ (
);

FILL FILL_3__1873_ (
);

FILL FILL_5__1799_ (
);

FILL FILL_7__2758_ (
);

FILL FILL_5__2740_ (
);

FILL FILL_7__2338_ (
);

FILL FILL_5__2320_ (
);

FILL FILL_1__2732_ (
);

FILL FILL_1__2312_ (
);

FILL FILL_3__2658_ (
);

FILL FILL_3__2238_ (
);

FILL FILL_5__3525_ (
);

FILL FILL_5__3105_ (
);

FILL FILL_1__3517_ (
);

FILL FILL_4__1942_ (
);

FILL FILL_6__1868_ (
);

NAND3X1 _2587_ (
    .A(_1083_),
    .B(_194_),
    .C(_273_),
    .Y(_274_)
);

OAI21X1 _2167_ (
    .A(_914__bF$buf1),
    .B(_1272_),
    .C(RDY_bF$buf1),
    .Y(_1276_)
);

FILL FILL_0__1842_ (
);

FILL FILL_2__2801_ (
);

FILL FILL_4__2727_ (
);

FILL FILL_4__2307_ (
);

FILL FILL_7__3296_ (
);

FILL FILL_0__2627_ (
);

FILL FILL_0__2207_ (
);

FILL FILL_1__3270_ (
);

FILL FILL_3__3196_ (
);

FILL FILL_3__1929_ (
);

FILL FILL_4__2480_ (
);

FILL FILL_4__2060_ (
);

FILL FILL_2__2398_ (
);

FILL FILL_0__2380_ (
);

NOR2X1 _1858_ (
    .A(_967_),
    .B(_982_),
    .Y(_983_)
);

FILL FILL_7__1782_ (
);

FILL FILL_4__3265_ (
);

FILL FILL_0__3585_ (
);

FILL FILL_0__3165_ (
);

FILL FILL_7__2567_ (
);

FILL FILL_1__2961_ (
);

FILL FILL_1__2541_ (
);

FILL FILL_1__2121_ (
);

FILL FILL_3__2887_ (
);

FILL FILL_3__2467_ (
);

FILL FILL_3__2047_ (
);

FILL FILL_4__1751_ (
);

NOR2X1 _2396_ (
    .A(_1499_),
    .B(_1500_),
    .Y(_1501_)
);

FILL FILL_2__2610_ (
);

FILL FILL_4__2956_ (
);

FILL FILL_4__2536_ (
);

FILL FILL_4__2116_ (
);

FILL FILL_0__2856_ (
);

FILL FILL_0__2436_ (
);

FILL FILL_0__2016_ (
);

FILL FILL_7__1838_ (
);

FILL FILL_5__1820_ (
);

FILL FILL_1__1812_ (
);

FILL FILL_5__2605_ (
);

FILL FILL_4__3494_ (
);

FILL FILL_4__3074_ (
);

FILL FILL_4__1807_ (
);

FILL FILL_7__2796_ (
);

FILL FILL_1__2770_ (
);

FILL FILL_1__2350_ (
);

FILL FILL_3__2696_ (
);

FILL FILL_3__2276_ (
);

FILL FILL_5__3563_ (
);

FILL FILL_5__3143_ (
);

FILL FILL_1__3555_ (
);

FILL FILL_1__3135_ (
);

FILL FILL_4__1980_ (
);

FILL FILL_2__1898_ (
);

FILL FILL_0__1880_ (
);

FILL FILL_4__2765_ (
);

FILL FILL_4__2345_ (
);

FILL FILL_0__2665_ (
);

FILL FILL_6__3632_ (
);

FILL FILL_0__2245_ (
);

FILL FILL_6__3212_ (
);

FILL FILL_2__3624_ (
);

FILL FILL_2__3204_ (
);

FILL FILL_3__1967_ (
);

FILL FILL_5__2834_ (
);

FILL FILL_5__2414_ (
);

FILL FILL_1__2826_ (
);

FILL FILL_1__2406_ (
);

INVX2 _1896_ (
    .A(DIMUX[6]),
    .Y(_1015_)
);

FILL FILL_5__3619_ (
);

FILL FILL_7__2185_ (
);

FILL FILL_0__1936_ (
);

FILL FILL_6__2903_ (
);

INVX1 _3622_ (
    .A(_1651_),
    .Y(_1652_)
);

OAI21X1 _3202_ (
    .A(_720__bF$buf1),
    .B(_687_),
    .C(\AXYS[1] [6]),
    .Y(_796_)
);

FILL FILL_3__2085_ (
);

FILL FILL_4__2994_ (
);

FILL FILL_4__2574_ (
);

FILL FILL_4__2154_ (
);

FILL FILL_0__2894_ (
);

FILL FILL_0__2474_ (
);

FILL FILL_0__2054_ (
);

FILL FILL_6__3021_ (
);

FILL FILL_2__3013_ (
);

FILL FILL_7__1876_ (
);

FILL FILL_1__1850_ (
);

FILL FILL_3__1776_ (
);

FILL FILL_0__3259_ (
);

FILL FILL_5__2643_ (
);

FILL FILL_5__2223_ (
);

FILL FILL_1__2635_ (
);

FILL FILL_1__2215_ (
);

FILL FILL_3__3502_ (
);

FILL FILL_5__3008_ (
);

FILL FILL_4__1845_ (
);

FILL FILL_0__1745_ (
);

FILL FILL_6__2712_ (
);

DFFSR _3431_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_99_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[3] [6])
);

NOR2X1 _3011_ (
    .A(_636_),
    .B(_634_),
    .Y(_637_)
);

FILL FILL_2__2704_ (
);

FILL FILL_1_BUFX2_insert20 (
);

FILL FILL_1_BUFX2_insert21 (
);

FILL FILL_1_BUFX2_insert22 (
);

FILL FILL_1_BUFX2_insert23 (
);

FILL FILL_5__3181_ (
);

FILL FILL_7__3199_ (
);

FILL FILL_1_BUFX2_insert24 (
);

FILL FILL_1_BUFX2_insert25 (
);

FILL FILL_1__3593_ (
);

FILL FILL_1__3173_ (
);

FILL FILL_3__3099_ (
);

FILL FILL_5__1914_ (
);

FILL FILL_1__1906_ (
);

FILL FILL_4__2383_ (
);

FILL FILL_6__3670_ (
);

FILL FILL_0__2283_ (
);

FILL FILL_6__3250_ (
);

FILL FILL_2__3662_ (
);

FILL FILL_2__3242_ (
);

FILL FILL_4__3588_ (
);

FILL FILL_4__3168_ (
);

OAI21X1 _2702_ (
    .A(_173_),
    .B(_326_),
    .C(_372_),
    .Y(_373_)
);

FILL FILL_0__3488_ (
);

FILL FILL_0__3068_ (
);

FILL FILL_5__2872_ (
);

FILL FILL_5__2452_ (
);

FILL FILL_5__2032_ (
);

FILL FILL_1__2864_ (
);

FILL FILL_1__2444_ (
);

FILL FILL_1__2024_ (
);

FILL FILL_3__3311_ (
);

FILL FILL_5__3657_ (
);

FILL FILL_5__3237_ (
);

FILL FILL_1__3649_ (
);

FILL FILL_1__3229_ (
);

NOR2X1 _2299_ (
    .A(_1179_),
    .B(_1328_),
    .Y(_1406_)
);

FILL FILL_0__1974_ (
);

FILL FILL_6__2941_ (
);

OAI21X1 _3660_ (
    .A(_1685_),
    .B(_1687_),
    .C(_1684_),
    .Y(_1517_)
);

FILL FILL_6__2521_ (
);

OAI21X1 _3240_ (
    .A(_787_),
    .B(_807_),
    .C(_816_),
    .Y(_100_)
);

FILL FILL_6__2101_ (
);

FILL FILL_2__2933_ (
);

FILL FILL_2__2513_ (
);

FILL FILL_4__2859_ (
);

FILL FILL_4__2439_ (
);

FILL FILL_4__2019_ (
);

FILL FILL_0__2759_ (
);

FILL FILL_0__2339_ (
);

FILL FILL_6__3306_ (
);

FILL FILL_0__3700_ (
);

FILL FILL_4__2192_ (
);

FILL FILL_5__2928_ (
);

FILL FILL_5__2508_ (
);

FILL FILL_0__2092_ (
);

FILL FILL_2__3471_ (
);

FILL FILL_2__3051_ (
);

NOR2X1 _2931_ (
    .A(_1160_),
    .B(_573_),
    .Y(_574_)
);

NOR2X1 _2511_ (
    .A(_1020_),
    .B(_205_),
    .Y(_206_)
);

FILL FILL_0__3297_ (
);

FILL FILL_7__2699_ (
);

FILL FILL_5__2681_ (
);

FILL FILL_7__2279_ (
);

FILL FILL_5__2261_ (
);

FILL FILL_1__2673_ (
);

FILL FILL_7__3640_ (
);

FILL FILL_1__2253_ (
);

FILL FILL_7__3220_ (
);

FILL FILL_3__2599_ (
);

FILL FILL_3__2179_ (
);

FILL FILL_3__3540_ (
);

FILL FILL_3__3120_ (
);

FILL FILL_5__3466_ (
);

FILL FILL_5__3046_ (
);

FILL FILL_1__3458_ (
);

FILL FILL_1__3038_ (
);

FILL FILL_4__1883_ (
);

FILL FILL_0__1783_ (
);

FILL FILL_6__2750_ (
);

FILL FILL_6__2330_ (
);

FILL FILL_2__2742_ (
);

FILL FILL_2__2322_ (
);

FILL FILL_4__2668_ (
);

FILL FILL_4__2248_ (
);

FILL FILL_0__2988_ (
);

FILL FILL_0__2568_ (
);

FILL FILL_6__3535_ (
);

FILL FILL_0__2148_ (
);

FILL FILL_6__3115_ (
);

FILL FILL_2__3527_ (
);

FILL FILL_2__3107_ (
);

FILL FILL_5__1952_ (
);

FILL FILL_1__1944_ (
);

FILL FILL_7__2911_ (
);

FILL FILL_3__2811_ (
);

FILL FILL_5__2737_ (
);

FILL FILL_5__2317_ (
);

FILL FILL_2_BUFX2_insert70 (
);

FILL FILL_2_BUFX2_insert71 (
);

FILL FILL_2_BUFX2_insert72 (
);

FILL FILL_2_BUFX2_insert73 (
);

FILL FILL_2_BUFX2_insert74 (
);

FILL FILL_2_BUFX2_insert75 (
);

FILL FILL_2_BUFX2_insert76 (
);

FILL FILL_1__2729_ (
);

FILL FILL_2_BUFX2_insert77 (
);

FILL FILL_2_BUFX2_insert78 (
);

FILL FILL_1__2309_ (
);

FILL FILL_2_BUFX2_insert79 (
);

FILL FILL_2__3280_ (
);

NOR3X1 _1799_ (
    .A(_904_),
    .B(_914__bF$buf3),
    .C(_924_),
    .Y(_925_)
);

NAND3X1 _2740_ (
    .A(_148_),
    .B(_405_),
    .C(_406_),
    .Y(_407_)
);

NOR2X1 _2320_ (
    .A(_976_),
    .B(_934_),
    .Y(_1427_)
);

FILL FILL_4__1939_ (
);

FILL FILL_5__2490_ (
);

FILL FILL_7__2088_ (
);

FILL FILL_5__2070_ (
);

FILL FILL_0__1839_ (
);

FILL FILL_6__2806_ (
);

OAI21X1 _3525_ (
    .A(alu_op[0]),
    .B(_1553_),
    .C(_1554_),
    .Y(_1555_)
);

OAI21X1 _3105_ (
    .A(_709_),
    .B(_714_),
    .C(_710_),
    .Y(_67_)
);

FILL FILL_1__2482_ (
);

FILL FILL_1__2062_ (
);

FILL FILL_5__3695_ (
);

FILL FILL_5__3275_ (
);

FILL FILL_1__3267_ (
);

FILL FILL_2__2971_ (
);

FILL FILL_2__2551_ (
);

FILL FILL_2__2131_ (
);

FILL FILL_4__2897_ (
);

FILL FILL_4__2477_ (
);

FILL FILL_4__2057_ (
);

FILL FILL_0__2797_ (
);

FILL FILL_0__2377_ (
);

FILL FILL_5__1761_ (
);

FILL FILL_7__1779_ (
);

FILL FILL_1__1753_ (
);

FILL FILL_7__2720_ (
);

FILL FILL_7__2300_ (
);

FILL FILL_3__2620_ (
);

FILL FILL_3__2200_ (
);

FILL FILL_5__2966_ (
);

FILL FILL_5__2546_ (
);

FILL FILL_5__2126_ (
);

FILL FILL168450x18150 (
);

FILL FILL_1__2958_ (
);

FILL FILL_1__2538_ (
);

FILL FILL_1__2118_ (
);

FILL FILL_6__1830_ (
);

FILL FILL_2__1822_ (
);

FILL FILL_4__1748_ (
);

FILL FILL_6__2615_ (
);

DFFSR _3334_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_12_),
    .CLK(clk_bF$buf2),
    .Q(PC[10])
);

FILL FILL_1__2291_ (
);

FILL FILL_2__2607_ (
);

FILL FILL_5__3084_ (
);

FILL FILL_1__3496_ (
);

FILL FILL_1__3076_ (
);

FILL FILL_5__1817_ (
);

FILL FILL_1__1809_ (
);

FILL FILL_2__2780_ (
);

FILL FILL_2__2360_ (
);

FILL FILL_4__2286_ (
);

NAND2X1 _1820_ (
    .A(_926_),
    .B(_911_),
    .Y(_946_)
);

FILL FILL_6__3573_ (
);

FILL FILL_0__2186_ (
);

FILL FILL_6__3153_ (
);

FILL FILL_2__3565_ (
);

FILL FILL_2__3145_ (
);

FILL FILL_5__1990_ (
);

INVX1 _2605_ (
    .A(_288_),
    .Y(_289_)
);

FILL FILL_1__1982_ (
);

FILL FILL_5__2775_ (
);

FILL FILL_5__2355_ (
);

FILL FILL_1__2767_ (
);

FILL FILL_1__2347_ (
);

FILL FILL_7__3314_ (
);

FILL FILL_3__3634_ (
);

FILL FILL_3__3214_ (
);

FILL FILL_4__1977_ (
);

FILL FILL_0__1877_ (
);

FILL FILL_6__2844_ (
);

AOI22X1 _3563_ (
    .A(_1580_),
    .B(_1584_),
    .C(_1592_),
    .D(_1586_),
    .Y(_1593_)
);

FILL FILL_6__2424_ (
);

FILL FILL_6__2004_ (
);

OAI21X1 _3143_ (
    .A(HC),
    .B(_728_),
    .C(_355_),
    .Y(_748_)
);

FILL FILL_2__2836_ (
);

FILL FILL_2__2416_ (
);

FILL FILL_7__1800_ (
);

FILL FILL_4__3703_ (
);

FILL FILL_6__3629_ (
);

FILL FILL_6__3209_ (
);

FILL FILL_0__3603_ (
);

FILL FILL_4__2095_ (
);

FILL FILL_3__2905_ (
);

FILL FILL_6_BUFX2_insert20 (
);

FILL FILL_6_BUFX2_insert21 (
);

FILL FILL_6_BUFX2_insert22 (
);

FILL FILL_6_BUFX2_insert23 (
);

FILL FILL_6_BUFX2_insert24 (
);

FILL FILL_6_BUFX2_insert25 (
);

AOI21X1 _2834_ (
    .A(_466_),
    .B(_488_),
    .C(_495_),
    .Y(_496_)
);

NOR2X1 _2414_ (
    .A(_122_),
    .B(_1387_),
    .Y(_123_)
);

FILL FILL_1__1791_ (
);

FILL FILL_5__2584_ (
);

FILL FILL_5__2164_ (
);

INVX1 _3619_ (
    .A(_1648_),
    .Y(_1649_)
);

FILL FILL_1__2996_ (
);

FILL FILL_1__2576_ (
);

FILL FILL_7__3543_ (
);

FILL FILL_1__2156_ (
);

FILL FILL_3__3023_ (
);

FILL FILL169950x79350 (
);

FILL FILL_2__1860_ (
);

FILL FILL_4__1786_ (
);

FILL FILL_6__2653_ (
);

DFFSR _3372_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_49_),
    .CLK(clk_bF$buf10),
    .Q(dst_reg[0])
);

FILL FILL_6__2233_ (
);

FILL FILL_2__2645_ (
);

FILL FILL_2__2225_ (
);

FILL FILL_4__3512_ (
);

FILL FILL_6__3018_ (
);

FILL FILL_5__1855_ (
);

FILL FILL_1__1847_ (
);

FILL FILL_7__2814_ (
);

FILL FILL_3__2714_ (
);

FILL FILL_6__3191_ (
);

FILL FILL_2__3183_ (
);

FILL FILL_6__1924_ (
);

NOR2X1 _2643_ (
    .A(_1424_),
    .B(_1021_),
    .Y(_318_)
);

OAI21X1 _2223_ (
    .A(_1329_),
    .B(_1326_),
    .C(_1330_),
    .Y(_1331_)
);

FILL FILL_2__1916_ (
);

FILL FILL_5__2393_ (
);

FILL FILL_6__2709_ (
);

DFFSR _3428_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_96_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[3] [3])
);

OAI22X1 _3008_ (
    .A(_1179_),
    .B(_530_),
    .C(_578_),
    .D(_553_),
    .Y(_634_)
);

FILL FILL_1__2385_ (
);

FILL FILL_3__3672_ (
);

FILL FILL_3__3252_ (
);

FILL FILL_5__3598_ (
);

FILL FILL_5__3178_ (
);

FILL FILL_6__2882_ (
);

FILL FILL_6__2462_ (
);

NAND2X1 _3181_ (
    .A(AN),
    .B(_763_),
    .Y(_782_)
);

FILL FILL_6__2042_ (
);

FILL FILL_2__2874_ (
);

FILL FILL_2__2454_ (
);

FILL FILL_2__2034_ (
);

NOR2X1 _1914_ (
    .A(_898_),
    .B(_907_),
    .Y(_1031_)
);

FILL FILL_6__3667_ (
);

FILL FILL_6__3247_ (
);

FILL FILL_2__3659_ (
);

FILL FILL_0__3641_ (
);

FILL FILL_0__3221_ (
);

FILL FILL_2__3239_ (
);

FILL FILL_7__2203_ (
);

FILL FILL_3__2943_ (
);

FILL FILL_3__2523_ (
);

FILL FILL_3__2103_ (
);

FILL FILL_5__2869_ (
);

FILL FILL_5__2449_ (
);

FILL FILL_5__2029_ (
);

FILL FILL_3__3308_ (
);

NAND2X1 _2872_ (
    .A(cond_code[2]),
    .B(_886__bF$buf5),
    .Y(_528_)
);

NOR2X1 _2452_ (
    .A(_147_),
    .B(_1337_),
    .Y(_154_)
);

NAND3X1 _2032_ (
    .A(_1141_),
    .B(_1139_),
    .C(_1140_),
    .Y(_1142_)
);

FILL FILL_6__2938_ (
);

AOI21X1 _3657_ (
    .A(_1611_),
    .B(_1592_),
    .C(_1586_),
    .Y(_1685_)
);

FILL FILL_6__2518_ (
);

OAI21X1 _3237_ (
    .A(_720__bF$buf0),
    .B(_808_),
    .C(\AXYS[3] [6]),
    .Y(_815_)
);

FILL FILL_1__2194_ (
);

FILL FILL_7__3161_ (
);

FILL FILL_0__2912_ (
);

FILL FILL_3__3481_ (
);

FILL FILL_3__3061_ (
);

FILL FILL_6__2691_ (
);

FILL FILL_6__2271_ (
);

FILL FILL_2__2683_ (
);

FILL FILL_2__2263_ (
);

FILL FILL_4__2189_ (
);

FILL FILL_4__3550_ (
);

FILL FILL_4__3130_ (
);

FILL FILL_6__3476_ (
);

FILL FILL_0__2089_ (
);

FILL FILL_6__3056_ (
);

FILL FILL_2__3468_ (
);

FILL FILL_0__3450_ (
);

FILL FILL_2__3048_ (
);

FILL FILL_0__3030_ (
);

FILL FILL_5__1893_ (
);

INVX1 _2928_ (
    .A(op[2]),
    .Y(_571_)
);

NOR2X1 _2508_ (
    .A(_200_),
    .B(_202_),
    .Y(_203_)
);

FILL FILL_1__1885_ (
);

FILL FILL_7__2432_ (
);

FILL FILL_3__2752_ (
);

FILL FILL_3__2332_ (
);

FILL FILL_5__2678_ (
);

FILL FILL_5__2258_ (
);

FILL FILL_7__3637_ (
);

FILL FILL_7__3217_ (
);

FILL FILL_1__3611_ (
);

FILL FILL_3__3537_ (
);

FILL FILL_3__3117_ (
);

FILL FILL_6__1962_ (
);

INVX2 _2681_ (
    .A(_329_),
    .Y(_353_)
);

OAI21X1 _2261_ (
    .A(RDY_bF$buf5),
    .B(_1018_),
    .C(_1368_),
    .Y(_1369_)
);

FILL FILL_2__1954_ (
);

FILL FILL_4__2821_ (
);

FILL FILL_4__2401_ (
);

FILL FILL_6__2747_ (
);

NAND2X1 _3466_ (
    .A(_1711_),
    .B(_1713_),
    .Y(AV)
);

FILL FILL_6__2327_ (
);

NOR2X1 _3046_ (
    .A(plp),
    .B(_1027__bF$buf3),
    .Y(_661_)
);

FILL FILL_0__2721_ (
);

FILL FILL_2__2739_ (
);

FILL FILL_2__2319_ (
);

FILL FILL_0__2301_ (
);

FILL FILL_3__3290_ (
);

FILL FILL_4__3606_ (
);

FILL FILL_0__3506_ (
);

FILL FILL_5__1949_ (
);

FILL FILL_6__2080_ (
);

FILL FILL_2__2492_ (
);

FILL FILL_2__2072_ (
);

FILL FILL_3__2808_ (
);

INVX2 _1952_ (
    .A(_993_),
    .Y(_1069_)
);

FILL FILL_6__3285_ (
);

FILL FILL_2__3697_ (
);

FILL FILL_2__3277_ (
);

OAI21X1 _2737_ (
    .A(_268_),
    .B(_313_),
    .C(_1083_),
    .Y(_404_)
);

NOR2X1 _2317_ (
    .A(state[5]),
    .B(_954_),
    .Y(_1424_)
);

FILL FILL_7__2661_ (
);

FILL FILL_3__2981_ (
);

FILL FILL_3__2561_ (
);

FILL FILL_3__2141_ (
);

FILL FILL_5__2487_ (
);

FILL FILL_5__2067_ (
);

FILL FILL_1__2899_ (
);

FILL FILL_1__2479_ (
);

FILL FILL_1__2059_ (
);

FILL FILL_1__3000_ (
);

FILL FILL_6__1771_ (
);

INVX1 _2490_ (
    .A(_186_),
    .Y(_187_)
);

INVX2 _2070_ (
    .A(_1178_),
    .Y(_1179_)
);

FILL FILL_2__1763_ (
);

FILL FILL_4__2630_ (
);

FILL FILL_4__2210_ (
);

FILL FILL_6__2976_ (
);

BUFX2 _3695_ (
    .A(_1741_[12]),
    .Y(AB[12])
);

FILL FILL_6__2556_ (
);

OAI21X1 _3275_ (
    .A(_931__bF$buf2),
    .B(_984_),
    .C(_210_),
    .Y(_851_)
);

FILL FILL_6__2136_ (
);

FILL FILL_0__2950_ (
);

FILL FILL_2__2968_ (
);

FILL FILL_2__2548_ (
);

FILL FILL_0__2530_ (
);

FILL FILL_2__2128_ (
);

FILL FILL_0__2110_ (
);

FILL FILL_7__1932_ (
);

FILL FILL_3__1832_ (
);

FILL FILL_0__3315_ (
);

FILL FILL_5__1758_ (
);

FILL FILL_7__2717_ (
);

FILL FILL_3__2617_ (
);

NAND2X1 _1761_ (
    .A(RDY_bF$buf9),
    .B(DI[5]),
    .Y(_890_)
);

FILL FILL_6__3094_ (
);

FILL FILL_2__3086_ (
);

FILL FILL_4__1901_ (
);

FILL FILL_6__1827_ (
);

OAI21X1 _2966_ (
    .A(_1149__bF$buf1),
    .B(_551_),
    .C(_599_),
    .Y(_43_)
);

INVX1 _2546_ (
    .A(ABL[3]),
    .Y(_238_)
);

NOR2X1 _2126_ (
    .A(_902__bF$buf3),
    .B(_912_),
    .Y(_1235_)
);

FILL FILL_7__2890_ (
);

FILL FILL_7__2050_ (
);

FILL FILL_2__1819_ (
);

FILL FILL_0__1801_ (
);

FILL FILL_3__2790_ (
);

FILL FILL_3__2370_ (
);

FILL FILL_5__2296_ (
);

FILL FILL_7__3675_ (
);

FILL FILL_1__2288_ (
);

FILL FILL_3__3575_ (
);

FILL FILL_3__3155_ (
);

FILL FILL_2__1992_ (
);

FILL FILL_6__2785_ (
);

FILL FILL_6__2365_ (
);

NAND2X1 _3084_ (
    .A(_695_),
    .B(_690_),
    .Y(_696_)
);

FILL FILL_2__2777_ (
);

FILL FILL_2__2357_ (
);

NOR2X1 _1817_ (
    .A(_931__bF$buf0),
    .B(_942_),
    .Y(_943_)
);

FILL FILL_4__3644_ (
);

FILL FILL_4__3224_ (
);

FILL FILL_0__3544_ (
);

FILL FILL_0__3124_ (
);

FILL FILL_5__1987_ (
);

FILL FILL_1__1979_ (
);

FILL FILL_7__2946_ (
);

FILL FILL_7__2106_ (
);

FILL FILL_1__2920_ (
);

FILL FILL_1__2500_ (
);

FILL FILL_3__2846_ (
);

FILL FILL_3__2426_ (
);

FILL FILL_3__2006_ (
);

OAI21X1 _1990_ (
    .A(_1074_),
    .B(_1101_),
    .C(_1104_),
    .Y(AI[2])
);

FILL FILL_5__3713_ (
);

FILL FILL_1__3705_ (
);

NAND3X1 _2775_ (
    .A(_409_),
    .B(_423_),
    .C(_417_),
    .Y(_440_)
);

NAND3X1 _2355_ (
    .A(_1457_),
    .B(_1408_),
    .C(_1460_),
    .Y(_1461_)
);

FILL FILL_4__2915_ (
);

FILL FILL_7__3484_ (
);

FILL FILL_1__2097_ (
);

FILL FILL_7__3064_ (
);

FILL FILL_0__2815_ (
);

FILL FILL_6__2594_ (
);

FILL FILL_6__2174_ (
);

FILL FILL_2__2586_ (
);

FILL FILL_2__2166_ (
);

FILL FILL169350x82950 (
);

FILL FILL_4__3453_ (
);

FILL FILL_4__3033_ (
);

FILL FILL_3__1870_ (
);

FILL FILL_5__1796_ (
);

FILL FILL_1__1788_ (
);

FILL FILL_7__2335_ (
);

FILL FILL_3__2655_ (
);

FILL FILL_3__2235_ (
);

FILL FILL_5__3522_ (
);

FILL FILL_5__3102_ (
);

FILL FILL_1__3514_ (
);

FILL FILL_6__1865_ (
);

OAI21X1 _2584_ (
    .A(_269_),
    .B(_270_),
    .C(_206_),
    .Y(_271_)
);

OAI21X1 _2164_ (
    .A(_931__bF$buf4),
    .B(_1272_),
    .C(RDY_bF$buf6),
    .Y(_1273_)
);

FILL FILL_2__1857_ (
);

FILL FILL_4__2724_ (
);

FILL FILL_4__2304_ (
);

DFFSR _3369_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_46_),
    .CLK(clk_bF$buf9),
    .Q(index_y)
);

FILL FILL168150x64950 (
);

FILL FILL_7__3293_ (
);

FILL FILL_0__2624_ (
);

FILL FILL_0__2204_ (
);

FILL FILL_3__3193_ (
);

FILL FILL_4__3509_ (
);

FILL FILL_3__1926_ (
);

FILL FILL_2__2395_ (
);

NOR2X1 _1855_ (
    .A(_975_),
    .B(_979_),
    .Y(_980_)
);

FILL FILL_4__3262_ (
);

FILL FILL_6__3188_ (
);

FILL FILL_0__3582_ (
);

FILL FILL_0__3162_ (
);

FILL FILL_7__2564_ (
);

FILL FILL_3__2884_ (
);

FILL FILL_3__2464_ (
);

FILL FILL_3__2044_ (
);

FILL FILL_3__3669_ (
);

FILL FILL_3__3249_ (
);

AND2X2 _2393_ (
    .A(_1311_),
    .B(_1321_),
    .Y(_1498_)
);

FILL FILL_4__2953_ (
);

FILL FILL_4__2533_ (
);

FILL FILL_4__2113_ (
);

FILL FILL_6__2879_ (
);

INVX1 _3598_ (
    .A(_1627_),
    .Y(_1628_)
);

FILL FILL_6__2459_ (
);

FILL FILL_6__2039_ (
);

OAI21X1 _3178_ (
    .A(_722_),
    .B(_778_),
    .C(_779_),
    .Y(_75_)
);

FILL FILL_0__2853_ (
);

FILL FILL_0__2433_ (
);

FILL FILL_0__2013_ (
);

FILL FILL_7__1835_ (
);

FILL FILL_0__3638_ (
);

FILL FILL_0__3218_ (
);

FILL FILL_5__2602_ (
);

FILL FILL_4__3491_ (
);

FILL FILL_4__3071_ (
);

FILL FILL_4__1804_ (
);

OAI21X1 _2869_ (
    .A(RDY_bF$buf2),
    .B(_1373_),
    .C(_526_),
    .Y(_19_)
);

INVX1 _2449_ (
    .A(_151_),
    .Y(_152_)
);

NAND2X1 _2029_ (
    .A(\AXYS[1] [7]),
    .B(_1047_),
    .Y(_1139_)
);

FILL FILL_7__2793_ (
);

FILL FILL_3__2693_ (
);

FILL FILL_3__2273_ (
);

FILL FILL_5__2199_ (
);

FILL FILL_5__3560_ (
);

FILL FILL_5__3140_ (
);

FILL FILL_0__2909_ (
);

FILL FILL_1__3552_ (
);

FILL FILL_1__3132_ (
);

FILL FILL_3__3478_ (
);

FILL FILL_3__3058_ (
);

FILL FILL_2__1895_ (
);

FILL FILL_4__2762_ (
);

FILL FILL_4__2342_ (
);

FILL FILL_6__2688_ (
);

FILL FILL_6__2268_ (
);

FILL FILL_0__2662_ (
);

FILL FILL_0__2242_ (
);

FILL FILL_2__3621_ (
);

FILL FILL_2__3201_ (
);

FILL FILL_4__3547_ (
);

FILL FILL_4__3127_ (
);

FILL FILL_3__1964_ (
);

FILL FILL_0__3027_ (
);

FILL FILL_7__2849_ (
);

FILL FILL_5__2831_ (
);

FILL FILL_7__2429_ (
);

FILL FILL_5__2411_ (
);

FILL FILL_7__2009_ (
);

FILL FILL_1__2823_ (
);

FILL FILL_1__2403_ (
);

FILL FILL_3__2749_ (
);

FILL FILL_3__2329_ (
);

INVX2 _1893_ (
    .A(DIMUX[5]),
    .Y(_1013_)
);

FILL FILL_5__3616_ (
);

FILL FILL_1__3608_ (
);

FILL FILL_6__1959_ (
);

OAI22X1 _2678_ (
    .A(RDY_bF$buf3),
    .B(_1007_),
    .C(_350_),
    .D(_348_),
    .Y(_4_)
);

OAI21X1 _2258_ (
    .A(_1154_),
    .B(_1186_),
    .C(_1185_),
    .Y(_1366_)
);

FILL FILL_7__2182_ (
);

FILL FILL_0__1933_ (
);

FILL FILL_6__2900_ (
);

FILL FILL_3__2082_ (
);

FILL FILL_4__2818_ (
);

FILL FILL_0__2718_ (
);

FILL FILL_3__3287_ (
);

FILL FILL_4__2991_ (
);

FILL FILL_4__2571_ (
);

FILL FILL_4__2151_ (
);

FILL FILL_6__2497_ (
);

FILL FILL_6__2077_ (
);

FILL FILL_0__2891_ (
);

FILL FILL_2__2489_ (
);

FILL FILL_0__2471_ (
);

FILL FILL_2__2069_ (
);

FILL FILL_0__2051_ (
);

NOR2X1 _1949_ (
    .A(_1062_),
    .B(_1065_),
    .Y(_1066_)
);

FILL FILL_2__3010_ (
);

FILL FILL_0__3676_ (
);

FILL FILL_3__1773_ (
);

FILL FILL_0__3256_ (
);

FILL FILL_7__2658_ (
);

FILL FILL_5__2640_ (
);

FILL FILL_7__2238_ (
);

FILL FILL_5__2220_ (
);

FILL FILL_1__2632_ (
);

FILL FILL_1__2212_ (
);

FILL FILL_3__2978_ (
);

FILL FILL_3__2558_ (
);

FILL FILL_3__2138_ (
);

FILL FILL_5__3005_ (
);

FILL FILL_4__1842_ (
);

FILL FILL_6__1768_ (
);

OAI21X1 _2487_ (
    .A(_1014_),
    .B(_136_),
    .C(_183_),
    .Y(_184_)
);

NAND2X1 _2067_ (
    .A(IRHOLD_valid),
    .B(IRHOLD[4]),
    .Y(_1176_)
);

FILL FILL_2__2701_ (
);

FILL FILL_4__2627_ (
);

FILL FILL_4__2207_ (
);

FILL FILL_7__3196_ (
);

FILL FILL_0__2947_ (
);

FILL FILL_0__2527_ (
);

FILL FILL_0__2107_ (
);

FILL FILL_1__3590_ (
);

FILL FILL_1__3170_ (
);

FILL FILL_3__3096_ (
);

FILL FILL_5__1911_ (
);

FILL FILL_7__1929_ (
);

FILL FILL_1__1903_ (
);

FILL FILL_3__1829_ (
);

FILL FILL_4__2380_ (
);

FILL FILL_0__2280_ (
);

FILL FILL_2__2298_ (
);

OAI21X1 _1758_ (
    .A(_886__bF$buf3),
    .B(DI[4]),
    .C(_887_),
    .Y(_888_)
);

FILL FILL_4__3585_ (
);

FILL FILL_4__3165_ (
);

FILL FILL169350x14550 (
);

FILL FILL_0__3485_ (
);

FILL FILL_0__3065_ (
);

FILL FILL_7__2887_ (
);

FILL FILL_7__2467_ (
);

FILL FILL_1__2861_ (
);

FILL FILL_1__2441_ (
);

FILL FILL_1__2021_ (
);

FILL FILL_3__2787_ (
);

FILL FILL_3__2367_ (
);

FILL FILL_5__3654_ (
);

FILL FILL_5__3234_ (
);

FILL FILL_1__3646_ (
);

FILL FILL_1__3226_ (
);

FILL FILL_6__1997_ (
);

OAI21X1 _2296_ (
    .A(_1367_),
    .B(_1402_),
    .C(_1351_),
    .Y(_1403_)
);

FILL FILL_2__1989_ (
);

FILL FILL_0__1971_ (
);

FILL FILL_2__2930_ (
);

FILL FILL_2__2510_ (
);

FILL FILL_4__2856_ (
);

FILL FILL_4__2436_ (
);

FILL FILL_4__2016_ (
);

FILL FILL_0__2756_ (
);

FILL FILL_0__2336_ (
);

FILL FILL_6__3303_ (
);

FILL FILL_2__3715_ (
);

FILL FILL_5__2925_ (
);

FILL FILL_5__2505_ (
);

FILL FILL_1__2917_ (
);

INVX1 _1987_ (
    .A(ABH[2]),
    .Y(_1102_)
);

FILL FILL_0__3294_ (
);

FILL FILL_7__2696_ (
);

BUFX2 _3713_ (
    .A(_1742_[6]),
    .Y(DO[6])
);

FILL FILL_1__2670_ (
);

FILL FILL_1__2250_ (
);

FILL FILL_3__2596_ (
);

FILL FILL_3__2176_ (
);

FILL FILL_5__3463_ (
);

FILL FILL_5__3043_ (
);

FILL FILL_1__3455_ (
);

FILL FILL_1__3035_ (
);

FILL FILL_4__1880_ (
);

FILL FILL_2__1798_ (
);

FILL FILL_0__1780_ (
);

FILL FILL_4__2665_ (
);

FILL FILL_4__2245_ (
);

FILL FILL_0__2985_ (
);

FILL FILL_0__2565_ (
);

FILL FILL_6__3532_ (
);

FILL FILL_0__2145_ (
);

FILL FILL169050x136950 (
);

FILL FILL_6__3112_ (
);

FILL FILL_2__3524_ (
);

FILL FILL_2__3104_ (
);

FILL FILL_7__1967_ (
);

FILL FILL_1__1941_ (
);

FILL FILL_3__1867_ (
);

FILL FILL_5__2734_ (
);

FILL FILL_5__2314_ (
);

FILL FILL_2_BUFX2_insert40 (
);

FILL FILL_2_BUFX2_insert41 (
);

FILL FILL_2_BUFX2_insert42 (
);

FILL FILL_2_BUFX2_insert43 (
);

FILL FILL_2_BUFX2_insert44 (
);

FILL FILL_2_BUFX2_insert45 (
);

FILL FILL_2_BUFX2_insert46 (
);

FILL FILL_1__2726_ (
);

FILL FILL_2_BUFX2_insert47 (
);

FILL FILL_2_BUFX2_insert48 (
);

FILL FILL_1__2306_ (
);

FILL FILL_2_BUFX2_insert49 (
);

NAND2X1 _1796_ (
    .A(inc),
    .B(_895_),
    .Y(_922_)
);

FILL FILL_5__3519_ (
);

FILL FILL_4__1936_ (
);

FILL FILL_7__2085_ (
);

FILL FILL_0__1836_ (
);

FILL FILL_6__2803_ (
);

AOI22X1 _3522_ (
    .A(_1716_),
    .B(BI[2]),
    .C(_1551_),
    .D(_1717_),
    .Y(_1552_)
);

NAND2X1 _3102_ (
    .A(CO),
    .B(_704_),
    .Y(_712_)
);

FILL FILL_5__3692_ (
);

FILL FILL_5__3272_ (
);

FILL FILL_1__3264_ (
);

FILL FILL_4__2894_ (
);

FILL FILL_4__2474_ (
);

FILL FILL_4__2054_ (
);

FILL FILL_0__2794_ (
);

FILL FILL_0__2374_ (
);

FILL FILL_7__1776_ (
);

FILL FILL_4__3259_ (
);

FILL FILL_1__1750_ (
);

FILL FILL_0__3579_ (
);

FILL FILL_0__3159_ (
);

FILL FILL169650x57750 (
);

FILL FILL_5__2963_ (
);

FILL FILL_5__2543_ (
);

FILL FILL_5__2123_ (
);

FILL FILL_1__2955_ (
);

FILL FILL_1__2535_ (
);

FILL FILL_1__2115_ (
);

FILL FILL_4__1745_ (
);

FILL FILL_6__2612_ (
);

DFFSR _3331_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(_9_),
    .CLK(clk_bF$buf5),
    .Q(PC[7])
);

FILL FILL_2__2604_ (
);

FILL FILL_5__3081_ (
);

FILL FILL_7__3099_ (
);

FILL FILL_1__3493_ (
);

FILL FILL_1__3073_ (
);

FILL FILL_5__1814_ (
);

FILL FILL_1__1806_ (
);

FILL FILL168450x39750 (
);

FILL FILL_4__2283_ (
);

FILL FILL_6__3570_ (
);

FILL FILL_0__2183_ (
);

FILL FILL_6__3150_ (
);

FILL FILL_2__3562_ (
);

FILL FILL_2__3142_ (
);

FILL FILL_4__3488_ (
);

FILL FILL_4__3068_ (
);

AOI22X1 _2602_ (
    .A(ADD[3]),
    .B(_198_),
    .C(_272_),
    .D(DIMUX[3]),
    .Y(_286_)
);

FILL FILL_5__2772_ (
);

FILL FILL_5__2352_ (
);

FILL FILL_1__2764_ (
);

FILL FILL_1__2344_ (
);

FILL FILL_7__3311_ (
);

FILL FILL_3__3631_ (
);

FILL FILL_3__3211_ (
);

FILL FILL_5__3557_ (
);

FILL FILL_5__3137_ (
);

FILL FILL_1__3549_ (
);

FILL FILL_1__3129_ (
);

FILL FILL_4__1974_ (
);

OAI21X1 _2199_ (
    .A(RDY_bF$buf6),
    .B(_1020_),
    .C(_1307_),
    .Y(_1308_)
);

FILL FILL_0__1874_ (
);

FILL FILL_6__2841_ (
);

AOI21X1 _3560_ (
    .A(_1572_),
    .B(_1576_),
    .C(alu_shift_right),
    .Y(_1590_)
);

FILL FILL_6__2421_ (
);

FILL FILL_6__2001_ (
);

OAI21X1 _3140_ (
    .A(_722_),
    .B(_744_),
    .C(_745_),
    .Y(_71_)
);

FILL FILL_2__2833_ (
);

FILL FILL_2__2413_ (
);

FILL FILL_4__2759_ (
);

FILL FILL_4__2339_ (
);

FILL FILL_4__3700_ (
);

FILL FILL_0__2659_ (
);

FILL FILL_6__3626_ (
);

FILL FILL_0__2239_ (
);

FILL FILL_6__3206_ (
);

FILL FILL169950x108150 (
);

FILL FILL_0__3600_ (
);

FILL FILL_2__3618_ (
);

FILL FILL_4__2092_ (
);

FILL FILL_3__2902_ (
);

FILL FILL_5__2828_ (
);

FILL FILL_5__2408_ (
);

FILL FILL_4__3297_ (
);

OAI21X1 _2831_ (
    .A(_1013_),
    .B(_351_),
    .C(_492_),
    .Y(_493_)
);

NOR2X1 _2411_ (
    .A(_1289_),
    .B(_1270_),
    .Y(_120_)
);

FILL FILL_0__3197_ (
);

FILL FILL_5__2581_ (
);

FILL FILL_5__2161_ (
);

FILL FILL_7__2179_ (
);

OAI21X1 _3616_ (
    .A(alu_op[3]),
    .B(BI[6]),
    .C(_1740_),
    .Y(_1646_)
);

FILL FILL_1__2993_ (
);

FILL FILL_1__2573_ (
);

FILL FILL_7__3540_ (
);

FILL FILL_1__2153_ (
);

FILL FILL_7__3120_ (
);

FILL FILL_3__2499_ (
);

FILL FILL_3__2079_ (
);

FILL FILL_3__3020_ (
);

FILL FILL_4__1783_ (
);

FILL FILL_6__2650_ (
);

FILL FILL_6__2230_ (
);

FILL FILL_2__2642_ (
);

FILL FILL_2__2222_ (
);

FILL FILL_4__2988_ (
);

FILL FILL_4__2568_ (
);

FILL FILL_4__2148_ (
);

FILL FILL_0__2888_ (
);

FILL FILL_0__2468_ (
);

FILL FILL_0__2048_ (
);

FILL FILL_6__3015_ (
);

FILL FILL_2__3007_ (
);

FILL FILL_5__1852_ (
);

FILL FILL_1__1844_ (
);

FILL FILL_7__2811_ (
);

FILL FILL_3__2711_ (
);

FILL FILL_5__2637_ (
);

FILL FILL_5__2217_ (
);

FILL FILL_1__2629_ (
);

FILL FILL_1__2209_ (
);

FILL FILL_2__3180_ (
);

FILL FILL_6__1921_ (
);

OAI21X1 _2640_ (
    .A(_929_),
    .B(_314_),
    .C(_313_),
    .Y(_315_)
);

NAND2X1 _2220_ (
    .A(_1212_),
    .B(_1327_),
    .Y(_1328_)
);

FILL FILL_2__1913_ (
);

FILL FILL_4__1839_ (
);

FILL FILL_5__2390_ (
);

FILL FILL_6__2706_ (
);

DFFSR _3425_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_93_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[3] [0])
);

AOI22X1 _3005_ (
    .A(dst_reg[1]),
    .B(_1149__bF$buf0),
    .C(_531_),
    .D(_631_),
    .Y(_632_)
);

FILL FILL_1__2382_ (
);

FILL FILL169950x10950 (
);

FILL FILL_5__3595_ (
);

FILL FILL_5__3175_ (
);

FILL FILL_1__3587_ (
);

FILL FILL_1__3167_ (
);

FILL FILL_5__1908_ (
);

FILL FILL_2__2871_ (
);

FILL FILL_2__2451_ (
);

FILL FILL_2__2031_ (
);

FILL FILL_4__2797_ (
);

FILL FILL_4__2377_ (
);

NAND2X1 _1911_ (
    .A(_969_),
    .B(_900_),
    .Y(_1028_)
);

FILL FILL_0__2697_ (
);

FILL FILL_6__3664_ (
);

FILL FILL_0__2277_ (
);

FILL FILL_6__3244_ (
);

FILL FILL_2__3656_ (
);

FILL FILL_2__3236_ (
);

FILL FILL_7__2620_ (
);

FILL FILL_7__2200_ (
);

FILL FILL_3__1999_ (
);

FILL FILL_3__2940_ (
);

FILL FILL_3__2520_ (
);

FILL FILL_3__2100_ (
);

FILL FILL_5__2866_ (
);

FILL FILL_5__2446_ (
);

FILL FILL_5__2026_ (
);

FILL FILL_1__2858_ (
);

FILL FILL_1__2438_ (
);

FILL FILL_1__2018_ (
);

FILL FILL_3__3305_ (
);

FILL FILL_0__1968_ (
);

FILL FILL_6__2935_ (
);

NAND2X1 _3654_ (
    .A(HC),
    .B(_1714__bF$buf3),
    .Y(_1683_)
);

FILL FILL_6__2515_ (
);

OAI21X1 _3234_ (
    .A(_757_),
    .B(_807_),
    .C(_813_),
    .Y(_97_)
);

FILL FILL_1__2191_ (
);

FILL FILL_2__2927_ (
);

FILL FILL_2__2507_ (
);

FILL FILL_2__2680_ (
);

FILL FILL_2__2260_ (
);

FILL FILL_4__2186_ (
);

FILL FILL_6__3473_ (
);

FILL FILL_0__2086_ (
);

FILL FILL_6__3053_ (
);

FILL FILL_2__3465_ (
);

FILL FILL_2__3045_ (
);

FILL FILL_5__1890_ (
);

NOR2X1 _2925_ (
    .A(_1215_),
    .B(_568_),
    .Y(_569_)
);

INVX2 _2505_ (
    .A(_199_),
    .Y(_200_)
);

FILL FILL_1__1882_ (
);

FILL FILL_5__2675_ (
);

FILL FILL_5__2255_ (
);

FILL FILL_1__2667_ (
);

FILL FILL_1__2247_ (
);

FILL FILL_7__3214_ (
);

FILL FILL_3__3534_ (
);

FILL FILL_3__3114_ (
);

FILL FILL_2__1951_ (
);

FILL FILL_4__1877_ (
);

FILL FILL_0__1777_ (
);

FILL FILL_6__2744_ (
);

OAI21X1 _3463_ (
    .A(_1708_),
    .B(_1710_),
    .C(_1706_),
    .Y(_1711_)
);

FILL FILL_6__2324_ (
);

INVX1 _3043_ (
    .A(_657_),
    .Y(_658_)
);

FILL FILL_2__2736_ (
);

FILL FILL_2__2316_ (
);

FILL FILL_4__3603_ (
);

FILL FILL_6__3529_ (
);

FILL FILL_6__3109_ (
);

FILL FILL_0__3503_ (
);

FILL FILL_5__1946_ (
);

FILL FILL_1__1938_ (
);

FILL FILL_3__2805_ (
);

FILL FILL_6__3282_ (
);

FILL FILL_2__3694_ (
);

FILL FILL_2__3274_ (
);

NAND2X1 _2734_ (
    .A(RDY_bF$buf0),
    .B(_401_),
    .Y(_402_)
);

AND2X2 _2314_ (
    .A(_1419_),
    .B(_1420_),
    .Y(_1421_)
);

FILL FILL_5__2484_ (
);

FILL FILL_5__2064_ (
);

AND2X2 _3519_ (
    .A(_1548_),
    .B(_1546_),
    .Y(_1549_)
);

FILL FILL_1__2896_ (
);

FILL FILL_1__2476_ (
);

FILL FILL_1__2056_ (
);

FILL FILL_5__3269_ (
);

FILL FILL_2__1760_ (
);

FILL FILL_6__2973_ (
);

FILL FILL_6__2553_ (
);

BUFX2 _3692_ (
    .A(_1741_[1]),
    .Y(AB[1])
);

OAI21X1 _3272_ (
    .A(state[5]),
    .B(state[4]),
    .C(_1225_),
    .Y(_848_)
);

FILL FILL_6__2133_ (
);

FILL FILL_2__2965_ (
);

FILL FILL_2__2545_ (
);

FILL FILL_2__2125_ (
);

FILL FILL_0__3312_ (
);

FILL FILL_5__1755_ (
);

FILL FILL_1__1747_ (
);

FILL FILL_7__2714_ (
);

FILL FILL_3__2614_ (
);

FILL FILL_6__3091_ (
);

FILL FILL_2__3083_ (
);

FILL FILL_6__1824_ (
);

AOI22X1 _2963_ (
    .A(inc),
    .B(_1149__bF$buf4),
    .C(_531_),
    .D(_572_),
    .Y(_598_)
);

AOI21X1 _2543_ (
    .A(_1100_),
    .B(_195_),
    .C(_235_),
    .Y(_236_)
);

NAND2X1 _2123_ (
    .A(_886__bF$buf6),
    .B(_916_),
    .Y(_1232_)
);

FILL FILL_2__1816_ (
);

FILL FILL_5__2293_ (
);

FILL FILL_6__2609_ (
);

DFFSR _3328_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(_6_),
    .CLK(clk_bF$buf5),
    .Q(PC[4])
);

FILL FILL_7__3672_ (
);

FILL FILL_1__2285_ (
);

FILL FILL_7_BUFX2_insert61 (
);

FILL FILL_3__3572_ (
);

FILL FILL_7_BUFX2_insert63 (
);

FILL FILL_3__3152_ (
);

FILL FILL_7_BUFX2_insert64 (
);

FILL FILL_7_BUFX2_insert66 (
);

FILL FILL_7_BUFX2_insert67 (
);

FILL FILL_5__3498_ (
);

FILL FILL_5__3078_ (
);

FILL FILL_7_BUFX2_insert69 (
);

FILL FILL_6__2782_ (
);

FILL FILL_6__2362_ (
);

AOI21X1 _3081_ (
    .A(plp),
    .B(_692_),
    .C(_1027__bF$buf4),
    .Y(_693_)
);

FILL FILL_2__2774_ (
);

FILL FILL_2__2354_ (
);

NAND2X1 _1814_ (
    .A(_929_),
    .B(_939_),
    .Y(_940_)
);

FILL FILL_4__3641_ (
);

FILL FILL_4__3221_ (
);

FILL FILL_6__3567_ (
);

FILL FILL_6__3147_ (
);

FILL FILL_0__3541_ (
);

FILL FILL_2__3559_ (
);

FILL FILL_0__3121_ (
);

FILL FILL_2__3139_ (
);

FILL FILL_5__1984_ (
);

FILL FILL_1__1976_ (
);

FILL FILL_7__2943_ (
);

FILL FILL_7__2103_ (
);

FILL FILL_3__2843_ (
);

FILL FILL_3__2423_ (
);

FILL FILL_3__2003_ (
);

FILL FILL_5__2769_ (
);

FILL FILL_5__2349_ (
);

FILL FILL_5__3710_ (
);

FILL FILL_1__3702_ (
);

FILL FILL_3__3628_ (
);

FILL FILL_3__3208_ (
);

AND2X2 _2772_ (
    .A(_436_),
    .B(_433_),
    .Y(_437_)
);

OR2X2 _2352_ (
    .A(_1410_),
    .B(_1414_),
    .Y(_1458_)
);

FILL FILL_4__2912_ (
);

FILL FILL_6__2838_ (
);

MUX2X1 _3557_ (
    .A(alu_op[1]),
    .B(_1575_),
    .S(alu_op[0]),
    .Y(_1587_)
);

FILL FILL_6__2418_ (
);

AOI21X1 _3137_ (
    .A(_732_),
    .B(_741_),
    .C(_742_),
    .Y(_743_)
);

FILL FILL_1__2094_ (
);

FILL FILL_7__3061_ (
);

FILL FILL_0__2812_ (
);

FILL FILL_1__3299_ (
);

FILL FILL_6__2591_ (
);

FILL FILL_6__2171_ (
);

FILL FILL_2__2583_ (
);

FILL FILL_2__2163_ (
);

FILL FILL_4__2089_ (
);

FILL FILL_4__3450_ (
);

FILL FILL_4__3030_ (
);

FILL FILL_5__1793_ (
);

AOI21X1 _2828_ (
    .A(ADD[5]),
    .B(_1299_),
    .C(_1334_),
    .Y(_490_)
);

AND2X2 _2408_ (
    .A(_1511_),
    .B(_1285_),
    .Y(_117_)
);

FILL FILL_1__1785_ (
);

FILL FILL_7__2332_ (
);

FILL FILL_3__2652_ (
);

FILL FILL_3__2232_ (
);

FILL FILL_5__2998_ (
);

FILL FILL_5__2578_ (
);

FILL FILL_5__2158_ (
);

FILL FILL_7__3537_ (
);

FILL FILL_7__3117_ (
);

FILL FILL_1__3511_ (
);

FILL FILL_3__3017_ (
);

FILL FILL_6__1862_ (
);

INVX2 _2581_ (
    .A(PC[8]),
    .Y(_268_)
);

OAI21X1 _2161_ (
    .A(RDY_bF$buf6),
    .B(_1267_),
    .C(_1269_),
    .Y(_1270_)
);

FILL FILL_2__1854_ (
);

FILL FILL_4__2721_ (
);

FILL FILL_4__2301_ (
);

FILL FILL_6__2647_ (
);

FILL FILL_6__2227_ (
);

DFFSR _3366_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_43_),
    .CLK(clk_bF$buf9),
    .Q(load_only)
);

FILL FILL_7__3290_ (
);

FILL FILL_0__2621_ (
);

FILL FILL_2__2639_ (
);

FILL FILL_2__2219_ (
);

FILL FILL_0__2201_ (
);

FILL FILL_3__3190_ (
);

FILL FILL_4__3506_ (
);

FILL FILL_3__1923_ (
);

FILL FILL_5__1849_ (
);

FILL FILL_7__2808_ (
);

FILL FILL_2__2392_ (
);

FILL FILL_3__2708_ (
);

NOR2X1 _1852_ (
    .A(_904_),
    .B(_976_),
    .Y(_977_)
);

FILL FILL_6__3185_ (
);

FILL FILL_2__3597_ (
);

FILL FILL_2__3177_ (
);

FILL FILL_6__1918_ (
);

NOR2X1 _2637_ (
    .A(_1154_),
    .B(_1027__bF$buf4),
    .Y(_312_)
);

NAND2X1 _2217_ (
    .A(_1325_),
    .B(_1250_),
    .Y(_1512_[0])
);

FILL FILL_7__2561_ (
);

FILL FILL_3__2881_ (
);

FILL FILL_3__2461_ (
);

FILL FILL_3__2041_ (
);

FILL FILL_5__2387_ (
);

FILL FILL_1__2799_ (
);

FILL FILL_1__2379_ (
);

FILL FILL_3__3666_ (
);

FILL FILL_3__3246_ (
);

NOR2X1 _2390_ (
    .A(_1494_),
    .B(_1353_),
    .Y(_1495_)
);

FILL FILL_4__2950_ (
);

FILL FILL_4__2530_ (
);

FILL FILL_4__2110_ (
);

FILL FILL_6__2876_ (
);

NAND2X1 _3595_ (
    .A(_1601_),
    .B(_1604_),
    .Y(_1625_)
);

FILL FILL_6__2456_ (
);

FILL FILL_6__2036_ (
);

OAI21X1 _3175_ (
    .A(_1015_),
    .B(_1018_),
    .C(_776_),
    .Y(_777_)
);

FILL FILL_0__2850_ (
);

FILL FILL_2__2868_ (
);

FILL FILL_2__2448_ (
);

FILL FILL_0__2430_ (
);

FILL FILL_2__2028_ (
);

FILL FILL_0__2010_ (
);

NAND3X1 _1908_ (
    .A(_997_),
    .B(_1024_),
    .C(_951_),
    .Y(_1025_)
);

FILL FILL_7__1832_ (
);

FILL FILL_4__3315_ (
);

FILL FILL_0__3635_ (
);

FILL FILL_0__3215_ (
);

FILL FILL_7__2617_ (
);

FILL FILL_3__2937_ (
);

FILL FILL_3__2517_ (
);

FILL FILL_4__1801_ (
);

NAND3X1 _2866_ (
    .A(NMI),
    .B(_524_),
    .C(_1153_),
    .Y(_525_)
);

OAI21X1 _2446_ (
    .A(_147_),
    .B(_1337_),
    .C(_148_),
    .Y(_149_)
);

OAI21X1 _2026_ (
    .A(_1015_),
    .B(_983_),
    .C(_1136_),
    .Y(_1137_)
);

FILL FILL_7__2790_ (
);

FILL FILL_3__2690_ (
);

FILL FILL_3__2270_ (
);

FILL FILL_5__2196_ (
);

FILL FILL_7__3575_ (
);

FILL FILL_1__2188_ (
);

FILL FILL_0__2906_ (
);

FILL FILL_3__3475_ (
);

FILL FILL_3__3055_ (
);

FILL FILL_2__1892_ (
);

FILL FILL_6__2685_ (
);

FILL FILL_6__2265_ (
);

FILL FILL_2__2677_ (
);

FILL FILL_2__2257_ (
);

FILL FILL_4__3544_ (
);

FILL FILL_4__3124_ (
);

FILL FILL_3__1961_ (
);

FILL FILL_0__3024_ (
);

FILL FILL_5__1887_ (
);

FILL FILL_1__1879_ (
);

FILL FILL_7__2846_ (
);

FILL FILL_7__2006_ (
);

FILL FILL_1__2820_ (
);

FILL FILL_1__2400_ (
);

FILL FILL_3__2746_ (
);

FILL FILL_3__2326_ (
);

INVX1 _1890_ (
    .A(PC[4]),
    .Y(_1011_)
);

FILL FILL_5__3613_ (
);

FILL FILL_1__3605_ (
);

FILL FILL_6__1956_ (
);

NOR2X1 _2675_ (
    .A(_347_),
    .B(_342_),
    .Y(_348_)
);

NAND3X1 _2255_ (
    .A(_1359_),
    .B(_1361_),
    .C(_1362_),
    .Y(_1363_)
);

FILL FILL_2__1948_ (
);

FILL FILL_0__1930_ (
);

FILL FILL_4__2815_ (
);

FILL FILL_0__2715_ (
);

FILL FILL_3__3284_ (
);

FILL FILL_6__2494_ (
);

FILL FILL_6__2074_ (
);

FILL FILL_2__2486_ (
);

FILL FILL_2__2066_ (
);

NOR2X1 _1946_ (
    .A(_902__bF$buf1),
    .B(_974_),
    .Y(_1063_)
);

FILL FILL_6__3699_ (
);

FILL FILL_6__3279_ (
);

FILL FILL_0__3673_ (
);

FILL FILL_3__1770_ (
);

FILL FILL_0__3253_ (
);

FILL FILL_7__2235_ (
);

FILL FILL_3__2975_ (
);

FILL FILL_3__2555_ (
);

FILL FILL_3__2135_ (
);

FILL FILL_5__3002_ (
);

FILL FILL_6__1765_ (
);

NOR2X1 _2484_ (
    .A(_178_),
    .B(_181_),
    .Y(_182_)
);

NAND2X1 _2064_ (
    .A(_1164_),
    .B(_1172_),
    .Y(_1173_)
);

FILL FILL_2__1757_ (
);

FILL FILL168450x150 (
);

FILL FILL_4__2624_ (
);

FILL FILL_4__2204_ (
);

DFFSR _3689_ (
    .R(_1513_),
    .S(vdd),
    .D(_1524_),
    .CLK(clk_bF$buf6),
    .Q(AN)
);

AND2X2 _3269_ (
    .A(_917_),
    .B(_1019_),
    .Y(_845_)
);

FILL FILL_7__3193_ (
);

FILL FILL_0__2944_ (
);

FILL FILL_0__2524_ (
);

FILL FILL_0__2104_ (
);

FILL FILL_3__3093_ (
);

FILL FILL_7__1926_ (
);

FILL FILL_1__1900_ (
);

FILL FILL_3__1826_ (
);

FILL FILL_0__3309_ (
);

FILL FILL_2__2295_ (
);

OAI21X1 _1755_ (
    .A(RDY_bF$buf9),
    .B(_884_),
    .C(_885_),
    .Y(DIMUX[3])
);

FILL FILL_4__3582_ (
);

FILL FILL_4__3162_ (
);

FILL FILL_6__3088_ (
);

FILL FILL_0__3482_ (
);

FILL FILL_0__3062_ (
);

FILL FILL_7__2464_ (
);

FILL FILL_3__2784_ (
);

FILL FILL_3__2364_ (
);

FILL FILL_7__3669_ (
);

FILL FILL_5__3651_ (
);

FILL FILL_5__3231_ (
);

FILL FILL_7__3249_ (
);

FILL FILL_1__3643_ (
);

FILL FILL_1__3223_ (
);

FILL FILL_3__3569_ (
);

FILL FILL_3__3149_ (
);

FILL FILL_6__1994_ (
);

MUX2X1 _2293_ (
    .A(_1219_),
    .B(_1399_),
    .S(_1178_),
    .Y(_1400_)
);

FILL FILL_2__1986_ (
);

FILL FILL_4__2853_ (
);

FILL FILL_4__2433_ (
);

FILL FILL_4__2013_ (
);

FILL FILL_6__2779_ (
);

NAND2X1 _3498_ (
    .A(alu_shift_right),
    .B(AI[5]),
    .Y(_1528_)
);

FILL FILL_6__2359_ (
);

AOI21X1 _3078_ (
    .A(_1227_),
    .B(_660_),
    .C(_689_),
    .Y(_690_)
);

FILL FILL_0__2753_ (
);

FILL FILL_0__2333_ (
);

FILL FILL_6__3300_ (
);

FILL FILL_2__3712_ (
);

FILL FILL_4__3638_ (
);

FILL FILL_4__3218_ (
);

FILL FILL_0__3538_ (
);

FILL FILL_0__3118_ (
);

FILL FILL_5__2922_ (
);

FILL FILL_5__2502_ (
);

FILL FILL_1__2914_ (
);

NAND3X1 _1984_ (
    .A(\AXYS[0] [2]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1099_)
);

FILL FILL_5__3707_ (
);

FILL FILL_0__3291_ (
);

OAI21X1 _2769_ (
    .A(_1291_),
    .B(_325_),
    .C(DIMUX[2]),
    .Y(_434_)
);

NOR3X1 _2349_ (
    .A(_1455_),
    .B(_1249_),
    .C(_1454_),
    .Y(_1456_)
);

FILL FILL_7__2693_ (
);

BUFX2 _3710_ (
    .A(_1742_[3]),
    .Y(DO[3])
);

FILL FILL_3__2593_ (
);

FILL FILL_3__2173_ (
);

FILL FILL_5__2099_ (
);

FILL FILL_4__2909_ (
);

FILL FILL_5__3460_ (
);

FILL FILL_5__3040_ (
);

FILL FILL_0__2809_ (
);

FILL FILL_1__3452_ (
);

FILL FILL_1__3032_ (
);

FILL FILL_2__1795_ (
);

FILL FILL_4__2662_ (
);

FILL FILL_4__2242_ (
);

FILL FILL_6__2588_ (
);

FILL FILL_6__2168_ (
);

FILL FILL_0__2982_ (
);

FILL FILL_0__2562_ (
);

FILL FILL_0__2142_ (
);

FILL FILL_2__3521_ (
);

FILL FILL_2__3101_ (
);

FILL FILL_7__1964_ (
);

FILL FILL_4__3027_ (
);

FILL FILL_3__1864_ (
);

FILL FILL_7__2749_ (
);

FILL FILL_5__2731_ (
);

FILL FILL_7__2329_ (
);

FILL FILL_5__2311_ (
);

FILL FILL_2_BUFX2_insert10 (
);

FILL FILL_2_BUFX2_insert11 (
);

FILL FILL_2_BUFX2_insert12 (
);

FILL FILL_2_BUFX2_insert13 (
);

FILL FILL_2_BUFX2_insert14 (
);

FILL FILL_2_BUFX2_insert15 (
);

FILL FILL_2_BUFX2_insert16 (
);

FILL FILL_1__2723_ (
);

FILL FILL_2_BUFX2_insert17 (
);

FILL FILL_2_BUFX2_insert18 (
);

FILL FILL_1__2303_ (
);

FILL FILL_2_BUFX2_insert19 (
);

FILL FILL_3__2649_ (
);

FILL FILL_3__2229_ (
);

AOI22X1 _1793_ (
    .A(rotate),
    .B(_915_),
    .C(_918_),
    .D(_895_),
    .Y(_919_)
);

FILL FILL_5__3516_ (
);

FILL FILL_1__3508_ (
);

FILL FILL_4__1933_ (
);

FILL FILL_6__1859_ (
);

OAI21X1 _2998_ (
    .A(_551_),
    .B(_625_),
    .C(_615_),
    .Y(_626_)
);

OAI21X1 _2578_ (
    .A(_1016_),
    .B(_218_),
    .C(_265_),
    .Y(_266_)
);

NAND2X1 _2158_ (
    .A(_1030_),
    .B(_1225_),
    .Y(_1267_)
);

FILL FILL_7__2082_ (
);

FILL FILL_0__1833_ (
);

FILL FILL_6__2800_ (
);

FILL FILL_4__2718_ (
);

FILL FILL_0__2618_ (
);

FILL FILL_1__3261_ (
);

FILL FILL_3__3187_ (
);

FILL FILL_4__2891_ (
);

FILL FILL_4__2471_ (
);

FILL FILL_4__2051_ (
);

FILL FILL_6__2397_ (
);

FILL FILL_0__2791_ (
);

FILL FILL_0__2371_ (
);

FILL FILL_2__2389_ (
);

NAND2X1 _1849_ (
    .A(_973_),
    .B(_911_),
    .Y(_974_)
);

FILL FILL_4__3676_ (
);

FILL FILL_4__3256_ (
);

FILL FILL_0__3576_ (
);

FILL FILL_0__3156_ (
);

FILL FILL_5__2960_ (
);

FILL FILL_7__2978_ (
);

FILL FILL_7__2558_ (
);

FILL FILL_5__2540_ (
);

FILL FILL_5__2120_ (
);

FILL FILL_7__2138_ (
);

FILL FILL_1__2952_ (
);

FILL FILL_1__2532_ (
);

FILL FILL_1__2112_ (
);

FILL FILL_3__2878_ (
);

FILL FILL_3__2458_ (
);

FILL FILL_3__2038_ (
);

FILL FILL_1__3317_ (
);

NOR2X1 _2387_ (
    .A(_1492_),
    .B(_1442_),
    .Y(_1493_)
);

FILL FILL_2__2601_ (
);

FILL FILL_4__2947_ (
);

FILL FILL_4__2527_ (
);

FILL FILL_4__2107_ (
);

FILL FILL_7__3096_ (
);

FILL FILL_0__2847_ (
);

FILL FILL_0__2427_ (
);

FILL FILL_0__2007_ (
);

FILL FILL_1__3490_ (
);

FILL FILL_1__3070_ (
);

FILL FILL_7__1829_ (
);

FILL FILL_5__1811_ (
);

FILL FILL_1__1803_ (
);

FILL FILL_4__2280_ (
);

FILL FILL_0__2180_ (
);

FILL FILL_2__2198_ (
);

FILL FILL_4__3485_ (
);

FILL FILL_4__3065_ (
);

FILL FILL_7__2787_ (
);

FILL FILL_7__2367_ (
);

FILL FILL_1__2761_ (
);

FILL FILL_1__2341_ (
);

FILL FILL_3__2687_ (
);

FILL FILL_3__2267_ (
);

FILL FILL_5__3554_ (
);

FILL FILL_5__3134_ (
);

FILL FILL_1__3546_ (
);

FILL FILL_1__3126_ (
);

FILL FILL_4__1971_ (
);

FILL FILL_6__1897_ (
);

OAI21X1 _2196_ (
    .A(_914__bF$buf1),
    .B(_981_),
    .C(_886__bF$buf2),
    .Y(_1305_)
);

FILL FILL_2__1889_ (
);

FILL FILL_0__1871_ (
);

FILL FILL_2__2830_ (
);

FILL FILL_2__2410_ (
);

FILL FILL_4__2756_ (
);

FILL FILL_4__2336_ (
);

FILL FILL_0__2656_ (
);

FILL FILL_6__3623_ (
);

FILL FILL_0__2236_ (
);

FILL FILL_6__3203_ (
);

FILL FILL_2__3615_ (
);

FILL FILL_3__1958_ (
);

FILL FILL_5__2825_ (
);

FILL FILL_5__2405_ (
);

FILL FILL_1__2817_ (
);

INVX2 _1887_ (
    .A(PC[3]),
    .Y(_1009_)
);

FILL FILL_4__3294_ (
);

FILL FILL169350x136950 (
);

FILL FILL_0__3194_ (
);

FILL FILL169950x162150 (
);

FILL FILL_7__2596_ (
);

FILL FILL_0__1927_ (
);

AOI22X1 _3613_ (
    .A(_1716_),
    .B(BI[6]),
    .C(_1642_),
    .D(_1717_),
    .Y(_1643_)
);

FILL FILL_1__2990_ (
);

FILL FILL_1__2570_ (
);

FILL FILL_1__2150_ (
);

FILL FILL_3__2496_ (
);

FILL FILL_3__2076_ (
);

FILL FILL169950x129750 (
);

FILL FILL_4__1780_ (
);

FILL FILL_4__2985_ (
);

FILL FILL_4__2565_ (
);

FILL FILL_4__2145_ (
);

FILL FILL_0__2885_ (
);

FILL FILL_0__2465_ (
);

FILL FILL_0__2045_ (
);

FILL FILL_6__3012_ (
);

FILL FILL_2__3004_ (
);

FILL FILL_7__1867_ (
);

FILL FILL_1__1841_ (
);

FILL FILL_3__1767_ (
);

FILL FILL_5__2634_ (
);

FILL FILL_5__2214_ (
);

FILL FILL_1__2626_ (
);

FILL FILL169050x3750 (
);

FILL FILL_1__2206_ (
);

FILL FILL_2__1910_ (
);

FILL FILL_4__1836_ (
);

FILL FILL_6__2703_ (
);

DFFSR _3422_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_91_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[2] [6])
);

OAI21X1 _3002_ (
    .A(_1396_),
    .B(_551_),
    .C(_580_),
    .Y(_629_)
);

FILL FILL_5__3592_ (
);

FILL FILL_5__3172_ (
);

FILL FILL_1__3584_ (
);

FILL FILL_1__3164_ (
);

FILL FILL_5__1905_ (
);

FILL FILL_4__2794_ (
);

FILL FILL_4__2374_ (
);

FILL FILL_0__2694_ (
);

FILL FILL_6__3661_ (
);

FILL FILL_0__2274_ (
);

FILL FILL_6__3241_ (
);

FILL FILL_2__3653_ (
);

FILL FILL_2__3233_ (
);

FILL FILL_4__3579_ (
);

FILL FILL_4__3159_ (
);

FILL FILL_3__1996_ (
);

FILL FILL_0__3479_ (
);

FILL FILL_0__3059_ (
);

FILL FILL_5__2863_ (
);

FILL FILL_5__2443_ (
);

FILL FILL_5__2023_ (
);

FILL FILL_1__2855_ (
);

FILL FILL_1__2435_ (
);

FILL FILL_1__2015_ (
);

FILL FILL_3__3302_ (
);

FILL FILL_5__3648_ (
);

FILL FILL_5__3228_ (
);

FILL FILL_0__1965_ (
);

FILL FILL_6__2932_ (
);

AOI21X1 _3651_ (
    .A(_1680_),
    .B(_1678_),
    .C(_1608_),
    .Y(_1681_)
);

FILL FILL_6__2512_ (
);

OAI21X1 _3231_ (
    .A(_720__bF$buf2),
    .B(_808_),
    .C(\AXYS[3] [3]),
    .Y(_812_)
);

FILL FILL_3_BUFX2_insert80 (
);

FILL FILL_3_BUFX2_insert81 (
);

FILL FILL_3_BUFX2_insert82 (
);

FILL FILL_3_BUFX2_insert83 (
);

FILL FILL_2__2924_ (
);

FILL FILL_2__2504_ (
);

FILL FILL_2__3709_ (
);

FILL FILL169650x115350 (
);

FILL FILL_4__2183_ (
);

FILL FILL_5__2919_ (
);

FILL FILL_6__3470_ (
);

FILL FILL_0__2083_ (
);

FILL FILL_6__3050_ (
);

FILL FILL_2__3462_ (
);

FILL FILL_2__3042_ (
);

AOI21X1 _2922_ (
    .A(_566_),
    .B(_565_),
    .C(_1149__bF$buf2),
    .Y(_567_)
);

NAND2X1 _2502_ (
    .A(_929_),
    .B(_955_),
    .Y(_197_)
);

FILL FILL_0__3288_ (
);

FILL FILL_5__2672_ (
);

FILL FILL_5__2252_ (
);

BUFX2 _3707_ (
    .A(_1742_[0]),
    .Y(DO[0])
);

FILL FILL_1__2664_ (
);

FILL FILL_1__2244_ (
);

FILL FILL_7__3211_ (
);

FILL FILL_3__3531_ (
);

FILL FILL_3__3111_ (
);

FILL FILL_5__3457_ (
);

FILL FILL_5__3037_ (
);

FILL FILL_1__3449_ (
);

FILL FILL_1__3029_ (
);

FILL FILL_4__1874_ (
);

NAND2X1 _2099_ (
    .A(RDY_bF$buf8),
    .B(_1207_),
    .Y(_1208_)
);

FILL FILL_0__1774_ (
);

FILL FILL_6__2741_ (
);

NOR2X1 _3460_ (
    .A(\u_ALU8.BI7 ),
    .B(_1707_),
    .Y(_1708_)
);

FILL FILL_6__2321_ (
);

OAI21X1 _3040_ (
    .A(_1168_),
    .B(_1150__bF$buf1),
    .C(_645_),
    .Y(_61_)
);

FILL FILL_2__2733_ (
);

FILL FILL_2__2313_ (
);

FILL FILL_4__2659_ (
);

FILL FILL_4__2239_ (
);

FILL FILL_4__3600_ (
);

FILL FILL_0__2979_ (
);

FILL FILL_0__2559_ (
);

FILL FILL_6__3526_ (
);

FILL FILL_0__2139_ (
);

FILL FILL_6__3106_ (
);

FILL FILL_2__3518_ (
);

FILL FILL_0__3500_ (
);

FILL FILL_5__1943_ (
);

FILL FILL_1__1935_ (
);

FILL FILL_3__2802_ (
);

FILL FILL_5__2728_ (
);

FILL FILL_5__2308_ (
);

FILL FILL_2__3691_ (
);

FILL FILL_2__3271_ (
);

FILL FILL_4__3197_ (
);

OAI21X1 _2731_ (
    .A(_1016_),
    .B(_330_),
    .C(_398_),
    .Y(_399_)
);

NOR2X1 _2311_ (
    .A(_1417_),
    .B(_1332_),
    .Y(_1418_)
);

FILL FILL_0__3097_ (
);

FILL FILL_5__2481_ (
);

FILL FILL_5__2061_ (
);

FILL FILL_7__2079_ (
);

INVX1 _3516_ (
    .A(_1728_),
    .Y(_1546_)
);

FILL FILL_1__2893_ (
);

FILL FILL_1__2473_ (
);

FILL FILL_1__2053_ (
);

FILL FILL_7__3020_ (
);

FILL FILL_3__2399_ (
);

FILL FILL_5__3266_ (
);

FILL FILL_1__3678_ (
);

FILL FILL_1__3258_ (
);

FILL FILL_6__2970_ (
);

FILL FILL_6__2550_ (
);

FILL FILL_6__2130_ (
);

FILL FILL_2__2962_ (
);

FILL FILL_2__2542_ (
);

FILL FILL_2__2122_ (
);

FILL FILL_4__2888_ (
);

FILL FILL_4__2468_ (
);

FILL FILL_4__2048_ (
);

FILL FILL_0__2788_ (
);

FILL FILL_0__2368_ (
);

FILL FILL_5__1752_ (
);

FILL FILL_1__1744_ (
);

FILL FILL_7__2711_ (
);

FILL FILL_3__2611_ (
);

FILL FILL_5__2957_ (
);

FILL FILL_5__2537_ (
);

FILL FILL_5__2117_ (
);

FILL FILL_1__2949_ (
);

FILL FILL_1__2529_ (
);

FILL FILL_1__2109_ (
);

FILL FILL_2__3080_ (
);

OAI21X1 _2960_ (
    .A(_308_),
    .B(_593_),
    .C(_595_),
    .Y(_41_)
);

FILL FILL_6__1821_ (
);

AOI22X1 _2540_ (
    .A(DIMUX[2]),
    .B(_227_),
    .C(_200_),
    .D(ABL[2]),
    .Y(_233_)
);

NOR2X1 _2120_ (
    .A(_1223_),
    .B(_1228_),
    .Y(_1229_)
);

FILL FILL_2__1813_ (
);

FILL FILL_5__2290_ (
);

FILL FILL_6__2606_ (
);

DFFSR _3325_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(_3_),
    .CLK(clk_bF$buf3),
    .Q(PC[1])
);

FILL FILL_1__2282_ (
);

FILL FILL_7_BUFX2_insert37 (
);

FILL FILL_5__3495_ (
);

FILL FILL_7_BUFX2_insert38 (
);

FILL FILL_5__3075_ (
);

FILL FILL_1__3487_ (
);

FILL FILL_1__3067_ (
);

FILL FILL_5__1808_ (
);

FILL FILL_2__2771_ (
);

FILL FILL_2__2351_ (
);

FILL FILL_4__2697_ (
);

FILL FILL_4__2277_ (
);

AND2X2 _1811_ (
    .A(state[1]),
    .B(state[0]),
    .Y(_937_)
);

FILL FILL_0__2597_ (
);

FILL FILL_6__3564_ (
);

FILL FILL_0__2177_ (
);

FILL FILL_6__3144_ (
);

FILL FILL_2__3556_ (
);

FILL FILL_2__3136_ (
);

FILL FILL_5__1981_ (
);

FILL FILL_1__1973_ (
);

FILL FILL_7__2940_ (
);

FILL FILL_7__2100_ (
);

FILL FILL_3__1899_ (
);

FILL FILL_3__2840_ (
);

FILL FILL_3__2420_ (
);

FILL FILL_3__2000_ (
);

FILL FILL_5__2766_ (
);

FILL FILL_5__2346_ (
);

FILL FILL_1__2758_ (
);

FILL FILL_1__2338_ (
);

FILL FILL_3__3625_ (
);

FILL FILL_3__3205_ (
);

FILL FILL_4__1968_ (
);

FILL FILL_0__1868_ (
);

FILL FILL_6__2835_ (
);

OAI21X1 _3554_ (
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1583_),
    .Y(_1584_)
);

FILL FILL_6__2415_ (
);

NOR2X1 _3134_ (
    .A(ADD[2]),
    .B(_730_),
    .Y(_740_)
);

FILL FILL_1__2091_ (
);

FILL FILL_2__2827_ (
);

FILL FILL_2__2407_ (
);

FILL FILL_1__3296_ (
);

FILL FILL169950x86550 (
);

FILL FILL_2__2580_ (
);

FILL FILL_2__2160_ (
);

FILL FILL_4__2086_ (
);

FILL FILL_5__1790_ (
);

OAI21X1 _2825_ (
    .A(_886__bF$buf3),
    .B(_487_),
    .C(_458_),
    .Y(_14_)
);

NOR2X1 _2405_ (
    .A(_1469_),
    .B(_1508_),
    .Y(_1509_)
);

FILL FILL_1__1782_ (
);

FILL FILL_5__2995_ (
);

FILL FILL_5__2575_ (
);

FILL FILL_5__2155_ (
);

FILL FILL_1__2987_ (
);

FILL FILL_1__2567_ (
);

FILL FILL_1__2147_ (
);

FILL FILL_7__3114_ (
);

FILL FILL_3__3014_ (
);

FILL FILL_2__1851_ (
);

FILL FILL_4__1777_ (
);

FILL FILL_6__2644_ (
);

DFFSR _3363_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_40_),
    .CLK(clk_bF$buf10),
    .Q(adc_bcd)
);

FILL FILL_6__2224_ (
);

FILL FILL_2__2636_ (
);

FILL FILL_2__2216_ (
);

FILL FILL_4__3503_ (
);

FILL FILL_6__3009_ (
);

FILL FILL_3__1920_ (
);

FILL FILL_5__1846_ (
);

FILL FILL_1__1838_ (
);

FILL FILL_3__2705_ (
);

FILL FILL_6__3182_ (
);

FILL FILL_2__3594_ (
);

FILL FILL_2__3174_ (
);

FILL FILL_6__1915_ (
);

NOR2X1 _2634_ (
    .A(_310_),
    .B(_129_),
    .Y(alu_shift_right)
);

NOR2X1 _2214_ (
    .A(_1312_),
    .B(_1322_),
    .Y(_1323_)
);

FILL FILL_2__1907_ (
);

FILL FILL_5__2384_ (
);

DFFSR _3419_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_88_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[2] [3])
);

FILL FILL_1__2796_ (
);

FILL FILL_1__2376_ (
);

FILL FILL_3__3663_ (
);

FILL FILL_3__3243_ (
);

FILL FILL_5__3589_ (
);

FILL FILL_5__3169_ (
);

FILL FILL_6__2873_ (
);

NAND2X1 _3592_ (
    .A(_1593_),
    .B(_1621_),
    .Y(_1622_)
);

FILL FILL_6__2453_ (
);

INVX1 _3172_ (
    .A(_773_),
    .Y(_774_)
);

FILL FILL_6__2033_ (
);

FILL FILL_2__2865_ (
);

FILL FILL_2__2445_ (
);

FILL FILL_2__2025_ (
);

NOR2X1 _1905_ (
    .A(_1020_),
    .B(_1021_),
    .Y(_1022_)
);

FILL FILL_4__3312_ (
);

FILL FILL_6__3658_ (
);

FILL FILL_6__3238_ (
);

FILL FILL_0__3632_ (
);

FILL FILL_0__3212_ (
);

FILL FILL_7__2614_ (
);

FILL FILL_3__2934_ (
);

FILL FILL_3__2514_ (
);

AOI21X1 _2863_ (
    .A(_522_),
    .B(_521_),
    .C(_886__bF$buf3),
    .Y(_523_)
);

OAI21X1 _2443_ (
    .A(_1319__bF$buf2),
    .B(_1263_),
    .C(PC[8]),
    .Y(_146_)
);

INVX1 _2023_ (
    .A(ABH[6]),
    .Y(_1134_)
);

FILL FILL_5__2193_ (
);

FILL FILL_6__2929_ (
);

NAND2X1 _3648_ (
    .A(_1676_),
    .B(_1677_),
    .Y(_1678_)
);

FILL FILL_6__2509_ (
);

OAI21X1 _3228_ (
    .A(_737_),
    .B(_807_),
    .C(_810_),
    .Y(_94_)
);

FILL FILL_7__3572_ (
);

FILL FILL_1__2185_ (
);

FILL FILL_0__2903_ (
);

FILL FILL_3__3472_ (
);

FILL FILL_3__3052_ (
);

FILL FILL_6__2682_ (
);

FILL FILL_6__2262_ (
);

FILL FILL_2__2674_ (
);

FILL FILL_2__2254_ (
);

FILL FILL_4__3541_ (
);

FILL FILL_4__3121_ (
);

FILL FILL_6__3467_ (
);

FILL FILL_6__3047_ (
);

FILL FILL_2__3459_ (
);

FILL FILL_2__3039_ (
);

FILL FILL_0__3021_ (
);

FILL FILL_5__1884_ (
);

NOR2X1 _2919_ (
    .A(_1217_),
    .B(_1396_),
    .Y(_564_)
);

FILL FILL_1__1876_ (
);

FILL FILL_7__2843_ (
);

FILL FILL_7__2003_ (
);

FILL FILL_3__2743_ (
);

FILL FILL_3__2323_ (
);

FILL FILL_5__2669_ (
);

FILL FILL_5__2249_ (
);

FILL FILL_5__3610_ (
);

FILL FILL_1__3602_ (
);

FILL FILL_3__3528_ (
);

FILL FILL_3__3108_ (
);

FILL FILL_6__1953_ (
);

NAND2X1 _2672_ (
    .A(_343_),
    .B(_344_),
    .Y(_345_)
);

NOR2X1 _2252_ (
    .A(state[4]),
    .B(_949_),
    .Y(_1360_)
);

FILL FILL_2__1945_ (
);

FILL FILL_4__2812_ (
);

FILL FILL_6__2738_ (
);

NOR2X1 _3457_ (
    .A(CO),
    .B(_1703_),
    .Y(_1705_)
);

FILL FILL_6__2318_ (
);

OAI21X1 _3037_ (
    .A(_1015_),
    .B(_647_),
    .C(_654_),
    .Y(_59_)
);

FILL FILL_0__2712_ (
);

FILL FILL_3__3281_ (
);

FILL FILL_1__3199_ (
);

FILL FILL_6__2491_ (
);

FILL FILL_6__2071_ (
);

FILL FILL_2__2483_ (
);

FILL FILL_2__2063_ (
);

INVX1 _1943_ (
    .A(_1059_),
    .Y(_1060_)
);

FILL FILL_6__3696_ (
);

FILL FILL_6__3276_ (
);

FILL FILL_0__3670_ (
);

FILL FILL_0__3250_ (
);

FILL FILL_2__3268_ (
);

INVX1 _2728_ (
    .A(ABL[7]),
    .Y(_396_)
);

NOR2X1 _2308_ (
    .A(_1414_),
    .B(_1410_),
    .Y(_1415_)
);

FILL FILL_7__2232_ (
);

FILL FILL_3__2972_ (
);

FILL FILL_3__2552_ (
);

FILL FILL_3__2132_ (
);

FILL FILL_5__2898_ (
);

FILL FILL_5__2478_ (
);

FILL FILL_5__2058_ (
);

FILL FILL_7__3017_ (
);

FILL FILL_6__1762_ (
);

INVX1 _2481_ (
    .A(ADD[5]),
    .Y(_179_)
);

NAND2X1 _2061_ (
    .A(_1168_),
    .B(DIMUX[2]),
    .Y(_1170_)
);

FILL FILL_2__1754_ (
);

FILL FILL_4__2621_ (
);

FILL FILL_4__2201_ (
);

FILL FILL_6__2967_ (
);

DFFSR _3686_ (
    .R(_1513_),
    .S(vdd),
    .D(_1521_),
    .CLK(clk_bF$buf3),
    .Q(ADD[4])
);

FILL FILL_6__2547_ (
);

NOR2X1 _3266_ (
    .A(_841_),
    .B(_838_),
    .Y(_842_)
);

FILL FILL_6__2127_ (
);

FILL FILL_7__3190_ (
);

FILL FILL_2__2959_ (
);

FILL FILL_0__2941_ (
);

FILL FILL_2__2539_ (
);

FILL FILL_0__2521_ (
);

FILL FILL_2__2119_ (
);

FILL FILL_0__2101_ (
);

FILL FILL_3__3090_ (
);

FILL FILL_3__1823_ (
);

FILL FILL_0__3306_ (
);

FILL FILL_5__1749_ (
);

FILL FILL_7__2708_ (
);

FILL FILL_2__2292_ (
);

FILL FILL_3__2608_ (
);

OAI21X1 _1752_ (
    .A(RDY_bF$buf0),
    .B(_882_),
    .C(_883_),
    .Y(DIMUX[2])
);

FILL FILL169950x18150 (
);

FILL FILL_6__3085_ (
);

FILL FILL_2__3497_ (
);

FILL FILL_2__3077_ (
);

NAND2X1 _2957_ (
    .A(D),
    .B(_1185_),
    .Y(_594_)
);

FILL FILL_6__1818_ (
);

AOI21X1 _2537_ (
    .A(_1089_),
    .B(_195_),
    .C(_230_),
    .Y(_231_)
);

NAND2X1 _2117_ (
    .A(_969_),
    .B(_1225_),
    .Y(_1226_)
);

FILL FILL_7__2461_ (
);

FILL FILL_3__2781_ (
);

FILL FILL_3__2361_ (
);

FILL FILL_5__2287_ (
);

FILL FILL_1__2699_ (
);

FILL FILL_7__3666_ (
);

FILL FILL_1__2279_ (
);

FILL FILL_7__3246_ (
);

FILL FILL_1__3640_ (
);

FILL FILL_1__3220_ (
);

FILL FILL_3__3566_ (
);

FILL FILL_3__3146_ (
);

FILL FILL_6__1991_ (
);

NOR2X1 _2290_ (
    .A(_1213_),
    .B(_1396_),
    .Y(_1397_)
);

FILL FILL_2__1983_ (
);

FILL FILL_4__2850_ (
);

FILL FILL_4__2430_ (
);

FILL FILL_4__2010_ (
);

FILL FILL_6__2776_ (
);

INVX2 _3495_ (
    .A(alu_op[2]),
    .Y(_1740_)
);

FILL FILL_6__2356_ (
);

NAND2X1 _3075_ (
    .A(_1051_),
    .B(_686_),
    .Y(_687_)
);

FILL FILL_0__2750_ (
);

FILL FILL_2__2768_ (
);

FILL FILL_0__2330_ (
);

FILL FILL_2__2348_ (
);

NAND2X1 _1808_ (
    .A(state[3]),
    .B(_896_),
    .Y(_934_)
);

FILL FILL_4__3635_ (
);

FILL FILL_4__3215_ (
);

FILL FILL_0__3535_ (
);

FILL FILL_0__3115_ (
);

FILL FILL_5__1978_ (
);

FILL FILL_7__2937_ (
);

FILL FILL_7__2517_ (
);

FILL FILL_1__2911_ (
);

FILL FILL_3__2837_ (
);

FILL FILL_3__2417_ (
);

OAI21X1 _1981_ (
    .A(_1074_),
    .B(_1090_),
    .C(_1096_),
    .Y(AI[1])
);

FILL FILL_5__3704_ (
);

INVX1 _2766_ (
    .A(ADD[2]),
    .Y(_431_)
);

NOR2X1 _2346_ (
    .A(_1389_),
    .B(_1452_),
    .Y(_1453_)
);

FILL FILL_7__2690_ (
);

FILL FILL_3__2590_ (
);

FILL FILL_3__2170_ (
);

FILL FILL_5__2096_ (
);

FILL FILL_4__2906_ (
);

FILL FILL_7__3475_ (
);

FILL FILL_1__2088_ (
);

FILL FILL_0__2806_ (
);

FILL FILL168150x136950 (
);

FILL FILL_2__1792_ (
);

FILL FILL_6__2585_ (
);

FILL FILL_6__2165_ (
);

FILL FILL_2__2997_ (
);

FILL FILL_2__2577_ (
);

FILL FILL_2__2157_ (
);

FILL FILL_7__1961_ (
);

FILL FILL_4__3024_ (
);

FILL FILL_3__1861_ (
);

FILL FILL_5__1787_ (
);

FILL FILL_1__1779_ (
);

FILL FILL_7__2746_ (
);

FILL FILL_1__2720_ (
);

FILL FILL_1__2300_ (
);

FILL FILL_3__2646_ (
);

FILL FILL_3__2226_ (
);

NOR2X1 _1790_ (
    .A(_914__bF$buf3),
    .B(_912_),
    .Y(_916_)
);

FILL FILL_5__3513_ (
);

FILL FILL_1__3505_ (
);

FILL FILL_4__1930_ (
);

FILL FILL_6__1856_ (
);

NOR2X1 _2995_ (
    .A(_620_),
    .B(_623_),
    .Y(_624_)
);

OAI21X1 _2575_ (
    .A(_216_),
    .B(_209_),
    .C(AN),
    .Y(_263_)
);

OAI21X1 _2155_ (
    .A(_914__bF$buf1),
    .B(_984_),
    .C(_886__bF$buf2),
    .Y(_1264_)
);

FILL FILL_0__1830_ (
);

FILL FILL_2__1848_ (
);

FILL FILL_4__2715_ (
);

FILL FILL_0__2615_ (
);

FILL FILL_3__3184_ (
);

FILL FILL_3__1917_ (
);

FILL FILL_6__2394_ (
);

FILL FILL_2__2386_ (
);

NOR2X1 _1846_ (
    .A(_970_),
    .B(_924_),
    .Y(_971_)
);

FILL FILL_4__3673_ (
);

FILL FILL_4__3253_ (
);

FILL FILL_6__3599_ (
);

FILL FILL_6__3179_ (
);

FILL FILL_0__3573_ (
);

FILL FILL_0__3153_ (
);

FILL FILL_7__2975_ (
);

FILL FILL_7__2135_ (
);

FILL FILL_3__2875_ (
);

FILL FILL_3__2455_ (
);

FILL FILL_3__2035_ (
);

FILL FILL_1__3314_ (
);

NOR3X1 _2384_ (
    .A(_1288_),
    .B(_1322_),
    .C(_1489_),
    .Y(_1490_)
);

FILL FILL_4__2944_ (
);

FILL FILL_4__2524_ (
);

FILL FILL_4__2104_ (
);

NAND3X1 _3589_ (
    .A(_1571_),
    .B(_1598_),
    .C(_1618_),
    .Y(_1619_)
);

NOR2X1 _3169_ (
    .A(ADD[6]),
    .B(_762_),
    .Y(_771_)
);

FILL FILL_7__3093_ (
);

FILL FILL_0__2844_ (
);

FILL FILL_0__2424_ (
);

FILL FILL_0__2004_ (
);

FILL FILL_7__1826_ (
);

FILL FILL_4__3309_ (
);

FILL FILL_1__1800_ (
);

FILL FILL_0__3629_ (
);

FILL FILL_0__3209_ (
);

FILL FILL_2__2195_ (
);

FILL FILL_4__3482_ (
);

FILL FILL_4__3062_ (
);

FILL FILL_7__2364_ (
);

FILL FILL_3__2684_ (
);

FILL FILL_3__2264_ (
);

FILL FILL_7__3569_ (
);

FILL FILL_5__3551_ (
);

FILL FILL_7__3149_ (
);

FILL FILL_5__3131_ (
);

FILL FILL_1__3543_ (
);

FILL FILL_1__3123_ (
);

FILL FILL_3__3469_ (
);

FILL FILL_3__3049_ (
);

FILL FILL_6__1894_ (
);

NOR2X1 _2193_ (
    .A(_1301_),
    .B(_1288_),
    .Y(_1302_)
);

FILL FILL_2__1886_ (
);

FILL FILL_4__2753_ (
);

FILL FILL_4__2333_ (
);

FILL FILL_6__2679_ (
);

DFFSR _3398_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_67_),
    .CLK(clk_bF$buf6),
    .Q(C)
);

FILL FILL_6__2259_ (
);

FILL FILL_0__2653_ (
);

FILL FILL_6__3620_ (
);

FILL FILL_0__2233_ (
);

FILL FILL_6__3200_ (
);

FILL FILL_2__3612_ (
);

FILL FILL_4__3538_ (
);

FILL FILL_4__3118_ (
);

FILL FILL_3__1955_ (
);

FILL FILL_0__3018_ (
);

FILL FILL_5__2822_ (
);

FILL FILL_5__2402_ (
);

FILL FILL_1__2814_ (
);

INVX2 _1884_ (
    .A(PC[2]),
    .Y(_1007_)
);

FILL FILL_4__3291_ (
);

FILL FILL_5__3607_ (
);

FILL FILL_0__3191_ (
);

INVX1 _2669_ (
    .A(_340_),
    .Y(_342_)
);

NAND2X1 _2249_ (
    .A(_1356_),
    .B(_1251_),
    .Y(_1357_)
);

FILL FILL_7__2593_ (
);

FILL FILL_0__1924_ (
);

NAND2X1 _3610_ (
    .A(AI[7]),
    .B(alu_shift_right),
    .Y(_1640_)
);

FILL FILL_3__2493_ (
);

FILL FILL_3__2073_ (
);

FILL FILL_4__2809_ (
);

FILL FILL_0__2709_ (
);

FILL FILL_3__3698_ (
);

FILL FILL_3__3278_ (
);

FILL FILL_4__2982_ (
);

FILL FILL_4__2562_ (
);

FILL FILL_4__2142_ (
);

FILL FILL_6__2488_ (
);

FILL FILL_6__2068_ (
);

FILL FILL_0__2882_ (
);

FILL FILL_0__2462_ (
);

FILL FILL_0__2042_ (
);

FILL FILL_2__3001_ (
);

FILL FILL_7__1864_ (
);

FILL FILL_3__1764_ (
);

FILL FILL_0__3667_ (
);

FILL FILL_0__3247_ (
);

FILL FILL_5__2631_ (
);

FILL FILL_7__2229_ (
);

FILL FILL_5__2211_ (
);

FILL FILL_1__2623_ (
);

FILL FILL_1__2203_ (
);

FILL FILL_3__2969_ (
);

FILL FILL_3__2549_ (
);

FILL FILL_3__2129_ (
);

FILL FILL_4__1833_ (
);

FILL FILL_6__1759_ (
);

NAND2X1 _2898_ (
    .A(_1189_),
    .B(_1251_),
    .Y(_547_)
);

NOR2X1 _2478_ (
    .A(_176_),
    .B(_172_),
    .Y(_177_)
);

OAI21X1 _2058_ (
    .A(_1165_),
    .B(NMI_edge),
    .C(_1166_),
    .Y(_1167_)
);

FILL FILL_6__2700_ (
);

FILL FILL_4__2618_ (
);

FILL FILL_0__2938_ (
);

FILL FILL_0__2518_ (
);

FILL FILL_1__3581_ (
);

FILL FILL_1__3161_ (
);

FILL FILL_3__3087_ (
);

FILL FILL_5__1902_ (
);

FILL FILL_4__2791_ (
);

FILL FILL_4__2371_ (
);

FILL FILL_6__2297_ (
);

FILL FILL_0__2691_ (
);

FILL FILL_0__2271_ (
);

FILL FILL_2__2289_ (
);

FILL FILL_2__3650_ (
);

FILL FILL_2__3230_ (
);

OAI21X1 _1749_ (
    .A(RDY_bF$buf9),
    .B(_880_),
    .C(_881_),
    .Y(DIMUX[1])
);

FILL FILL_4__3576_ (
);

FILL FILL_4__3156_ (
);

FILL FILL_3__1993_ (
);

FILL FILL_0__3476_ (
);

FILL FILL_0__3056_ (
);

FILL FILL_5__2860_ (
);

FILL FILL_7__2878_ (
);

FILL FILL_7__2458_ (
);

FILL FILL_5__2440_ (
);

FILL FILL_7__2038_ (
);

FILL FILL_5__2020_ (
);

FILL FILL_1__2852_ (
);

FILL FILL_1__2432_ (
);

FILL FILL_1__2012_ (
);

FILL FILL_3__2778_ (
);

FILL FILL_3__2358_ (
);

FILL FILL_5__3645_ (
);

FILL FILL_5__3225_ (
);

FILL FILL_1__3637_ (
);

FILL FILL_1__3217_ (
);

FILL FILL_6__1988_ (
);

INVX1 _2287_ (
    .A(_1393_),
    .Y(_1394_)
);

FILL FILL_0__1962_ (
);

FILL FILL_3_BUFX2_insert50 (
);

FILL FILL_3_BUFX2_insert51 (
);

FILL FILL_3_BUFX2_insert52 (
);

FILL FILL_3_BUFX2_insert53 (
);

FILL FILL_2__2921_ (
);

FILL FILL_2__2501_ (
);

FILL FILL_3_BUFX2_insert54 (
);

FILL FILL_3_BUFX2_insert55 (
);

FILL FILL_3_BUFX2_insert56 (
);

FILL FILL_3_BUFX2_insert57 (
);

FILL FILL_4__2847_ (
);

FILL FILL_3_BUFX2_insert58 (
);

FILL FILL_4__2427_ (
);

FILL FILL_3_BUFX2_insert59 (
);

FILL FILL_4__2007_ (
);

FILL FILL_0__2747_ (
);

FILL FILL_6__3714_ (
);

FILL FILL_0__2327_ (
);

FILL FILL_2__3706_ (
);

FILL FILL_4__2180_ (
);

FILL FILL_5__2916_ (
);

FILL FILL_0__2080_ (
);

FILL FILL_2__2098_ (
);

FILL FILL_1__2908_ (
);

INVX1 _1978_ (
    .A(_1093_),
    .Y(_1094_)
);

FILL FILL_0__3285_ (
);

FILL FILL_7__2687_ (
);

FILL FILL_7__2267_ (
);

BUFX2 _3704_ (
    .A(_1741_[7]),
    .Y(AB[7])
);

FILL FILL_1__2661_ (
);

FILL FILL_1__2241_ (
);

FILL FILL_3__2587_ (
);

FILL FILL_3__2167_ (
);

FILL FILL_5__3454_ (
);

FILL FILL_5__3034_ (
);

FILL FILL169650x136950 (
);

FILL FILL_1__3026_ (
);

FILL FILL_4__1871_ (
);

FILL FILL_6__1797_ (
);

OAI21X1 _2096_ (
    .A(_913_),
    .B(_1200_),
    .C(_1204_),
    .Y(_1205_)
);

FILL FILL_2__1789_ (
);

FILL FILL_0__1771_ (
);

FILL FILL_2__2730_ (
);

FILL FILL_2__2310_ (
);

FILL FILL_4__2656_ (
);

FILL FILL_4__2236_ (
);

FILL FILL_0__2976_ (
);

FILL FILL_0__2556_ (
);

FILL FILL_6__3523_ (
);

FILL FILL_0__2136_ (
);

FILL FILL_6__3103_ (
);

FILL FILL_2__3515_ (
);

FILL FILL_5__1940_ (
);

FILL FILL_7__1958_ (
);

FILL FILL_1__1932_ (
);

FILL FILL_3__1858_ (
);

FILL FILL_5__2725_ (
);

FILL FILL_5__2305_ (
);

FILL FILL_1__2717_ (
);

INVX2 _1787_ (
    .A(state[5]),
    .Y(_913_)
);

FILL FILL_4__3194_ (
);

FILL FILL_0__3094_ (
);

FILL FILL169950x7350 (
);

FILL FILL_4__1927_ (
);

FILL FILL_7__2496_ (
);

FILL FILL_0__1827_ (
);

AOI21X1 _3513_ (
    .A(_1540_),
    .B(_1539_),
    .C(alu_shift_right),
    .Y(_1543_)
);

FILL FILL_1__2890_ (
);

FILL FILL_1__2470_ (
);

FILL FILL_1__2050_ (
);

FILL FILL_3__2396_ (
);

FILL FILL169650x64950 (
);

FILL FILL_5__3263_ (
);

FILL FILL_1__3675_ (
);

FILL FILL_1__3255_ (
);

FILL FILL_4__2885_ (
);

FILL FILL_4__2465_ (
);

FILL FILL_4__2045_ (
);

FILL FILL_0__2785_ (
);

FILL FILL_0__2365_ (
);

FILL FILL_5__2954_ (
);

FILL FILL_5__2534_ (
);

FILL FILL_5__2114_ (
);

FILL FILL_1__2946_ (
);

FILL FILL_1__2526_ (
);

FILL FILL_1__2106_ (
);

FILL FILL_2__1810_ (
);

FILL FILL_6__2603_ (
);

DFFSR _3322_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_1512_[4]),
    .CLK(clk_bF$buf6),
    .Q(state[4])
);

FILL FILL_5__3492_ (
);

FILL FILL_5__3072_ (
);

FILL FILL_1__3484_ (
);

FILL FILL_1__3064_ (
);

FILL FILL_5__1805_ (
);

FILL FILL_4__2694_ (
);

FILL FILL_4__2274_ (
);

FILL FILL_0__2594_ (
);

FILL FILL_6__3561_ (
);

FILL FILL_0__2174_ (
);

FILL FILL_6__3141_ (
);

FILL FILL_2__3553_ (
);

FILL FILL_2__3133_ (
);

FILL FILL_7__1996_ (
);

FILL FILL_4__3479_ (
);

FILL FILL_4__3059_ (
);

FILL FILL_1__1970_ (
);

FILL FILL_3__1896_ (
);

FILL FILL169950x115350 (
);

FILL FILL_5__2763_ (
);

FILL FILL_5__2343_ (
);

FILL FILL_1__2755_ (
);

FILL FILL_1__2335_ (
);

FILL FILL_3__3622_ (
);

FILL FILL_3__3202_ (
);

FILL FILL_5__3548_ (
);

FILL FILL_5__3128_ (
);

FILL FILL_4__1965_ (
);

FILL FILL_0__1865_ (
);

FILL FILL_6__2832_ (
);

OAI21X1 _3551_ (
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1725_),
    .Y(_1581_)
);

FILL FILL_6__2412_ (
);

NAND2X1 _3131_ (
    .A(\AXYS[0] [1]),
    .B(_722_),
    .Y(_738_)
);

FILL FILL_2__2824_ (
);

FILL FILL_2__2404_ (
);

FILL FILL_6__3617_ (
);

FILL FILL_1__3293_ (
);

FILL FILL_2__3609_ (
);

FILL FILL_4__2083_ (
);

FILL FILL_5__2819_ (
);

FILL FILL_4__3288_ (
);

NAND3X1 _2822_ (
    .A(_468_),
    .B(_470_),
    .C(_484_),
    .Y(_485_)
);

INVX1 _2402_ (
    .A(_1192_),
    .Y(_1506_)
);

FILL FILL_0__3188_ (
);

FILL FILL_5__2992_ (
);

FILL FILL_5__2572_ (
);

FILL FILL_5__2152_ (
);

OAI21X1 _3607_ (
    .A(_1727_),
    .B(_1728_),
    .C(_1724_),
    .Y(_1637_)
);

FILL FILL_1__2984_ (
);

FILL FILL_1__2564_ (
);

FILL FILL_1__2144_ (
);

FILL FILL_7__3111_ (
);

FILL FILL_3__3011_ (
);

FILL FILL_4__1774_ (
);

FILL FILL_6__2641_ (
);

DFFSR _3360_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_37_),
    .CLK(clk_bF$buf9),
    .Q(shift_right)
);

FILL FILL_6__2221_ (
);

FILL FILL_2__2633_ (
);

FILL FILL_2__2213_ (
);

FILL FILL_4__2979_ (
);

FILL FILL_4__2559_ (
);

FILL FILL_4__2139_ (
);

FILL FILL_4__3500_ (
);

FILL FILL_0__2879_ (
);

FILL FILL_0__2459_ (
);

FILL FILL_0__2039_ (
);

FILL FILL_6__3006_ (
);

FILL FILL_5__1843_ (
);

FILL FILL_1__1835_ (
);

FILL FILL_3__2702_ (
);

FILL FILL_5__2628_ (
);

FILL FILL_5__2208_ (
);

FILL FILL_2__3591_ (
);

FILL FILL_2__3171_ (
);

FILL FILL_4__3097_ (
);

FILL FILL_6__1912_ (
);

INVX1 _2631_ (
    .A(adc_bcd),
    .Y(_309_)
);

OAI21X1 _2211_ (
    .A(_931__bF$buf0),
    .B(_958_),
    .C(_886__bF$buf4),
    .Y(_1320_)
);

FILL FILL_2__1904_ (
);

FILL FILL_5__2381_ (
);

DFFSR _3416_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_85_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[2] [0])
);

FILL FILL_1__2793_ (
);

FILL FILL_1__2373_ (
);

FILL FILL_3__2299_ (
);

FILL FILL_3__3660_ (
);

FILL FILL_3__3240_ (
);

FILL FILL_5__3586_ (
);

FILL FILL_5__3166_ (
);

FILL FILL_1__3578_ (
);

FILL FILL_1__3158_ (
);

FILL FILL_6__2870_ (
);

FILL FILL_6__2450_ (
);

FILL FILL_6__2030_ (
);

FILL FILL_2__2862_ (
);

FILL FILL_2__2442_ (
);

FILL FILL_2__2022_ (
);

FILL FILL_4__2788_ (
);

FILL FILL_4__2368_ (
);

OAI21X1 _1902_ (
    .A(_903__bF$buf2),
    .B(_969_),
    .C(_992_),
    .Y(_1019_)
);

FILL FILL_0__2688_ (
);

FILL FILL_6__3655_ (
);

FILL FILL_0__2268_ (
);

FILL FILL_6__3235_ (
);

FILL FILL_2__3647_ (
);

FILL FILL_2__3227_ (
);

FILL FILL_7__2611_ (
);

FILL FILL_3__2931_ (
);

FILL FILL_3__2511_ (
);

FILL FILL_5__2857_ (
);

FILL FILL_5__2437_ (
);

FILL FILL_5__2017_ (
);

FILL FILL_1__2849_ (
);

FILL FILL_1__2429_ (
);

FILL FILL_1__2009_ (
);

NAND3X1 _2860_ (
    .A(_509_),
    .B(_519_),
    .C(_513_),
    .Y(_520_)
);

OAI21X1 _2440_ (
    .A(_902__bF$buf0),
    .B(_949_),
    .C(_138_),
    .Y(_143_)
);

NAND3X1 _2020_ (
    .A(\AXYS[0] [6]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1131_)
);

FILL FILL_5__2190_ (
);

FILL FILL_0__1959_ (
);

FILL FILL_6__2926_ (
);

AND2X2 _3645_ (
    .A(_1661_),
    .B(_1674_),
    .Y(_1675_)
);

FILL FILL_6__2506_ (
);

OAI21X1 _3225_ (
    .A(_720__bF$buf3),
    .B(_808_),
    .C(\AXYS[3] [0]),
    .Y(_809_)
);

FILL FILL_1__2182_ (
);

FILL FILL_2__2918_ (
);

FILL FILL_0__2900_ (
);

FILL FILL_2__2671_ (
);

FILL FILL_2__2251_ (
);

FILL FILL_4__2597_ (
);

FILL FILL_4__2177_ (
);

FILL FILL_0__2497_ (
);

FILL FILL_6__3464_ (
);

FILL FILL_0__2077_ (
);

FILL FILL_6__3044_ (
);

FILL FILL_2__3456_ (
);

FILL FILL_2__3036_ (
);

FILL FILL_5__1881_ (
);

AND2X2 _2916_ (
    .A(_560_),
    .B(_1405_),
    .Y(_561_)
);

FILL FILL_1__1873_ (
);

FILL FILL_7__2840_ (
);

FILL FILL_7__2000_ (
);

FILL FILL_3__1799_ (
);

FILL FILL_3__2740_ (
);

FILL FILL_3__2320_ (
);

FILL FILL_5__2666_ (
);

FILL FILL_5__2246_ (
);

FILL FILL_1__2658_ (
);

FILL FILL_7__3625_ (
);

FILL FILL_1__2238_ (
);

FILL FILL_3__3525_ (
);

FILL FILL_3__3105_ (
);

FILL FILL_6__1950_ (
);

FILL FILL_2__1942_ (
);

FILL FILL_4__1868_ (
);

FILL FILL_0__1768_ (
);

FILL FILL_6__2735_ (
);

NOR2X1 _3454_ (
    .A(_1698_),
    .B(_1702_),
    .Y(AZ)
);

FILL FILL_6__2315_ (
);

OAI21X1 _3034_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[5]),
    .Y(_653_)
);

FILL FILL_2__2727_ (
);

FILL FILL_2__2307_ (
);

FILL FILL_1__3196_ (
);

FILL FILL_5__1937_ (
);

FILL FILL_1__1929_ (
);

FILL FILL_2__2480_ (
);

FILL FILL_2__2060_ (
);

AOI22X1 _1940_ (
    .A(_1048_),
    .B(_1039_),
    .C(_1052_),
    .D(_1056_),
    .Y(_1057_)
);

FILL FILL_6__3693_ (
);

FILL FILL_6__3273_ (
);

FILL FILL_2__3265_ (
);

INVX1 _2725_ (
    .A(_392_),
    .Y(_394_)
);

INVX2 _2305_ (
    .A(_1187_),
    .Y(_1412_)
);

FILL FILL_5__2895_ (
);

FILL FILL_5__2475_ (
);

FILL FILL_5__2055_ (
);

FILL FILL_1__2887_ (
);

FILL FILL_1__2467_ (
);

FILL FILL_1__2047_ (
);

FILL FILL_7__3014_ (
);

FILL FILL_2__1751_ (
);

FILL FILL_0__1997_ (
);

FILL FILL_6__2964_ (
);

DFFSR _3683_ (
    .R(_1513_),
    .S(vdd),
    .D(_1518_),
    .CLK(clk_bF$buf5),
    .Q(ADD[1])
);

FILL FILL_6__2544_ (
);

OAI21X1 _3263_ (
    .A(_952_),
    .B(_1360_),
    .C(_823_),
    .Y(_839_)
);

FILL FILL_6__2124_ (
);

FILL FILL_2__2956_ (
);

FILL FILL_2__2536_ (
);

FILL FILL_2__2116_ (
);

FILL FILL_3__1820_ (
);

FILL FILL_0__3303_ (
);

FILL FILL_5__1746_ (
);

FILL FILL_3__2605_ (
);

FILL FILL_6__3082_ (
);

FILL FILL_2__3494_ (
);

FILL FILL_2__3074_ (
);

FILL FILL_6__1815_ (
);

OAI22X1 _2954_ (
    .A(_895_),
    .B(_1150__bF$buf1),
    .C(_1174_),
    .D(_591_),
    .Y(_39_)
);

AOI22X1 _2534_ (
    .A(DIMUX[1]),
    .B(_227_),
    .C(_200_),
    .D(ABL[1]),
    .Y(_228_)
);

OAI21X1 _2114_ (
    .A(_902__bF$buf3),
    .B(_912_),
    .C(_1222_),
    .Y(_1223_)
);

FILL FILL_2__1807_ (
);

FILL FILL_5__2284_ (
);

DFFSR _3319_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_1512_[1]),
    .CLK(clk_bF$buf6),
    .Q(state[1])
);

FILL FILL_1__2696_ (
);

FILL FILL_1__2276_ (
);

FILL FILL_7__3243_ (
);

FILL FILL_3__3563_ (
);

FILL FILL_3__3143_ (
);

FILL FILL169950x72150 (
);

FILL FILL_5__3489_ (
);

FILL FILL_5__3069_ (
);

FILL FILL_2__1980_ (
);

FILL FILL_6__2773_ (
);

OAI21X1 _3492_ (
    .A(AI[5]),
    .B(_1734_),
    .C(_1722_),
    .Y(_1737_)
);

FILL FILL_6__2353_ (
);

FILL FILL169950x39750 (
);

NAND2X1 _3072_ (
    .A(I),
    .B(_680_),
    .Y(_685_)
);

FILL FILL_2__2765_ (
);

FILL FILL_2__2345_ (
);

NAND2X1 _1805_ (
    .A(state[4]),
    .B(_913_),
    .Y(_931_)
);

FILL FILL_4__3632_ (
);

FILL FILL_4__3212_ (
);

FILL FILL_6__3558_ (
);

FILL FILL_6__3138_ (
);

FILL FILL_0__3532_ (
);

FILL FILL_0__3112_ (
);

FILL FILL_5__1975_ (
);

FILL FILL_1__1967_ (
);

FILL FILL_7__2514_ (
);

FILL FILL_3__2834_ (
);

FILL FILL_3__2414_ (
);

FILL FILL_5__3701_ (
);

FILL FILL_3__3619_ (
);

OAI21X1 _2763_ (
    .A(_428_),
    .B(_401_),
    .C(RDY_bF$buf4),
    .Y(_429_)
);

NAND3X1 _2343_ (
    .A(_1448_),
    .B(_1449_),
    .C(_1446_),
    .Y(_1450_)
);

FILL FILL_5__2093_ (
);

FILL FILL_4__2903_ (
);

FILL FILL_6__2829_ (
);

NAND2X1 _3548_ (
    .A(_1722_),
    .B(_1577_),
    .Y(_1578_)
);

FILL FILL_6__2409_ (
);

OAI21X1 _3128_ (
    .A(ADD[1]),
    .B(_729_),
    .C(_734_),
    .Y(_735_)
);

FILL FILL_7__3472_ (
);

FILL FILL_1__2085_ (
);

FILL FILL_0__2803_ (
);

FILL FILL_5__3298_ (
);

FILL FILL_6__2582_ (
);

FILL FILL_6__2162_ (
);

FILL FILL_2__2994_ (
);

FILL FILL_2__2574_ (
);

FILL FILL_2__2154_ (
);

FILL FILL_4__3021_ (
);

FILL FILL_5__1784_ (
);

NOR2X1 _2819_ (
    .A(_285_),
    .B(_352_),
    .Y(_482_)
);

FILL FILL_1__1776_ (
);

FILL FILL_7__2743_ (
);

FILL FILL_3__2643_ (
);

FILL FILL_3__2223_ (
);

FILL FILL_5__2989_ (
);

FILL FILL_5__2569_ (
);

FILL FILL_5__2149_ (
);

FILL FILL_5__3510_ (
);

FILL FILL_1__3502_ (
);

FILL FILL_3__3008_ (
);

FILL FILL_6__1853_ (
);

NAND2X1 _2992_ (
    .A(_1402_),
    .B(_559_),
    .Y(_621_)
);

OAI21X1 _2572_ (
    .A(_1014_),
    .B(_218_),
    .C(_260_),
    .Y(_261_)
);

OAI21X1 _2152_ (
    .A(_931__bF$buf1),
    .B(_984_),
    .C(_886__bF$buf0),
    .Y(_1261_)
);

FILL FILL_2__1845_ (
);

FILL FILL_4__2712_ (
);

FILL FILL_6__2638_ (
);

DFFSR _3357_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_34_),
    .CLK(clk_bF$buf9),
    .Q(op[2])
);

FILL FILL_6__2218_ (
);

FILL FILL_0__2612_ (
);

FILL FILL_3__3181_ (
);

FILL FILL_1__3099_ (
);

FILL FILL_3__1914_ (
);

FILL FILL_6__2391_ (
);

FILL FILL_2__2383_ (
);

INVX2 _1843_ (
    .A(_967_),
    .Y(_968_)
);

FILL FILL_4__3670_ (
);

FILL FILL_4__3250_ (
);

FILL FILL_6__3596_ (
);

FILL FILL_6__3176_ (
);

FILL FILL_2__3588_ (
);

FILL FILL_0__3570_ (
);

FILL FILL_2__3168_ (
);

FILL FILL_0__3150_ (
);

FILL FILL_7_CLKBUF1_insert27 (
);

FILL FILL_7_CLKBUF1_insert29 (
);

FILL FILL_6__1909_ (
);

OAI21X1 _2628_ (
    .A(_304_),
    .B(_218_),
    .C(_307_),
    .Y(_1741_[15])
);

AND2X2 _2208_ (
    .A(_1315_),
    .B(_1316_),
    .Y(_1317_)
);

FILL FILL_7__2972_ (
);

FILL FILL_7__2132_ (
);

FILL FILL_3__2872_ (
);

FILL FILL_3__2452_ (
);

FILL FILL_3__2032_ (
);

FILL FILL_5__2798_ (
);

FILL FILL_5__2378_ (
);

FILL FILL_1__3311_ (
);

FILL FILL_3__3657_ (
);

FILL FILL_3__3237_ (
);

NOR2X1 _2381_ (
    .A(_1369_),
    .B(_1372_),
    .Y(_1487_)
);

FILL FILL_4__2941_ (
);

FILL FILL_4__2521_ (
);

FILL FILL_4__2101_ (
);

FILL FILL_6__2867_ (
);

OAI21X1 _3586_ (
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1615_),
    .Y(_1616_)
);

FILL FILL_6__2447_ (
);

FILL FILL_6__2027_ (
);

OAI21X1 _3166_ (
    .A(_722_),
    .B(_767_),
    .C(_768_),
    .Y(_74_)
);

FILL FILL_7__3090_ (
);

FILL FILL_2__2859_ (
);

FILL FILL_0__2841_ (
);

FILL FILL_0__2421_ (
);

FILL FILL_2__2439_ (
);

FILL FILL_2__2019_ (
);

FILL FILL_0__2001_ (
);

FILL FILL_4__3306_ (
);

FILL FILL_0__3626_ (
);

FILL FILL_0__3206_ (
);

FILL FILL_7__2608_ (
);

FILL FILL_2__2192_ (
);

FILL FILL_3__2928_ (
);

FILL FILL_3__2508_ (
);

AND2X2 _2857_ (
    .A(_515_),
    .B(_516_),
    .Y(_517_)
);

OAI21X1 _2437_ (
    .A(_931__bF$buf3),
    .B(_946_),
    .C(_1204_),
    .Y(_141_)
);

OAI21X1 _2017_ (
    .A(_1074_),
    .B(_1125_),
    .C(_1128_),
    .Y(AI[5])
);

FILL FILL_7__2361_ (
);

FILL FILL_3__2681_ (
);

FILL FILL_3__2261_ (
);

FILL FILL_5__2187_ (
);

FILL FILL_1__2599_ (
);

FILL FILL_7__3566_ (
);

FILL FILL_1__2179_ (
);

FILL FILL_7__3146_ (
);

FILL FILL_1__3540_ (
);

FILL FILL_1__3120_ (
);

FILL FILL_3__3466_ (
);

FILL FILL_3__3046_ (
);

FILL FILL_6__1891_ (
);

NOR2X1 _2190_ (
    .A(_914__bF$buf4),
    .B(_954_),
    .Y(_1299_)
);

FILL FILL_2__1883_ (
);

FILL FILL_4__2750_ (
);

FILL FILL_4__2330_ (
);

FILL FILL_6__2676_ (
);

DFFSR _3395_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_64_),
    .CLK(clk_bF$buf1),
    .Q(I)
);

FILL FILL_6__2256_ (
);

FILL FILL_2__2668_ (
);

FILL FILL_0__2650_ (
);

FILL FILL_0__2230_ (
);

FILL FILL_2__2248_ (
);

FILL FILL_4__3535_ (
);

FILL FILL_4__3115_ (
);

FILL FILL168450x136950 (
);

FILL FILL_3__1952_ (
);

FILL FILL_0__3015_ (
);

FILL FILL_5__1878_ (
);

FILL FILL_7__2837_ (
);

FILL FILL_7__2417_ (
);

FILL FILL_1__2811_ (
);

FILL FILL_3__2737_ (
);

FILL FILL_3__2317_ (
);

INVX1 _1881_ (
    .A(PC[1]),
    .Y(_1005_)
);

FILL FILL_5__3604_ (
);

FILL FILL_6__1947_ (
);

NAND3X1 _2666_ (
    .A(_320_),
    .B(_331_),
    .C(_338_),
    .Y(_340_)
);

INVX1 _2246_ (
    .A(_1353_),
    .Y(_1354_)
);

FILL FILL_7__2590_ (
);

FILL FILL_0__1921_ (
);

FILL FILL_2__1939_ (
);

FILL FILL_3__2490_ (
);

FILL FILL_3__2070_ (
);

FILL FILL_4__2806_ (
);

FILL FILL_0__2706_ (
);

FILL FILL_3__3695_ (
);

FILL FILL_3__3275_ (
);

FILL FILL_6__2485_ (
);

FILL FILL_6__2065_ (
);

FILL FILL_2__2897_ (
);

FILL FILL_2__2477_ (
);

FILL FILL_2__2057_ (
);

NAND3X1 _1937_ (
    .A(\AXYS[0] [0]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1054_)
);

FILL FILL_7__1861_ (
);

FILL FILL_3__1761_ (
);

FILL FILL_0__3664_ (
);

FILL FILL_0__3244_ (
);

FILL FILL_7__2646_ (
);

FILL FILL_1__2620_ (
);

FILL FILL_1__2200_ (
);

FILL FILL_3__2966_ (
);

FILL FILL_3__2546_ (
);

FILL FILL_3__2126_ (
);

FILL FILL_4__1830_ (
);

INVX1 _2895_ (
    .A(sed),
    .Y(_545_)
);

FILL FILL_6__1756_ (
);

OAI21X1 _2475_ (
    .A(_971_),
    .B(_941_),
    .C(_903__bF$buf2),
    .Y(_174_)
);

OAI21X1 _2055_ (
    .A(IRHOLD_valid),
    .B(DIMUX[3]),
    .C(_1163_),
    .Y(_1164_)
);

FILL FILL_2__1748_ (
);

FILL FILL_4__2615_ (
);

FILL FILL_0__2935_ (
);

FILL FILL_0__2515_ (
);

FILL FILL_3__3084_ (
);

FILL FILL_7__1917_ (
);

FILL FILL_3__1817_ (
);

FILL FILL_6__2294_ (
);

FILL FILL_2__2286_ (
);

OAI21X1 _1746_ (
    .A(RDY_bF$buf0),
    .B(_878_),
    .C(_879_),
    .Y(DIMUX[0])
);

FILL FILL_4__3573_ (
);

FILL FILL_4__3153_ (
);

FILL FILL_6__3499_ (
);

FILL FILL_6__3079_ (
);

FILL FILL_3__1990_ (
);

FILL FILL_0__3473_ (
);

FILL FILL_0__3053_ (
);

FILL FILL_7__2875_ (
);

FILL FILL_7__2035_ (
);

FILL FILL_3__2775_ (
);

FILL FILL_3__2355_ (
);

FILL FILL_5__3642_ (
);

FILL FILL_5__3222_ (
);

FILL FILL_1__3634_ (
);

FILL FILL_1__3214_ (
);

FILL FILL_6__1985_ (
);

NOR2X1 _2284_ (
    .A(_1324_),
    .B(_1391_),
    .Y(_1392_)
);

FILL FILL_2__1977_ (
);

FILL FILL_3_BUFX2_insert20 (
);

FILL FILL_3_BUFX2_insert21 (
);

FILL FILL_3_BUFX2_insert22 (
);

FILL FILL_3_BUFX2_insert23 (
);

FILL FILL_3_BUFX2_insert24 (
);

FILL FILL_3_BUFX2_insert25 (
);

FILL FILL_4__2844_ (
);

FILL FILL_4__2424_ (
);

FILL FILL_4__2004_ (
);

AND2X2 _3489_ (
    .A(_1718_),
    .B(BI[5]),
    .Y(_1734_)
);

OAI21X1 _3069_ (
    .A(_681_),
    .B(_677_),
    .C(_956_),
    .Y(_682_)
);

FILL FILL_0__2744_ (
);

FILL FILL_6__3711_ (
);

FILL FILL_0__2324_ (
);

FILL FILL_2__3703_ (
);

FILL FILL_4__3629_ (
);

FILL FILL_4__3209_ (
);

FILL FILL_0__3529_ (
);

FILL FILL_0__3109_ (
);

FILL FILL_5__2913_ (
);

FILL FILL_2__2095_ (
);

FILL FILL_1__2905_ (
);

INVX1 _1975_ (
    .A(ABH[1]),
    .Y(_1091_)
);

FILL FILL_0__3282_ (
);

FILL FILL_7__2264_ (
);

BUFX2 _3701_ (
    .A(_1741_[4]),
    .Y(AB[4])
);

FILL FILL_3__2584_ (
);

FILL FILL_3__2164_ (
);

FILL FILL_5__3451_ (
);

FILL FILL_7__3469_ (
);

FILL FILL_7__3049_ (
);

FILL FILL_5__3031_ (
);

FILL FILL_1__3023_ (
);

FILL FILL_6__1794_ (
);

NAND2X1 _2093_ (
    .A(_929_),
    .B(_908_),
    .Y(_1202_)
);

FILL FILL_2__1786_ (
);

FILL FILL_4__2653_ (
);

FILL FILL_4__2233_ (
);

FILL FILL_6__2999_ (
);

FILL FILL_6__2579_ (
);

OAI21X1 _3298_ (
    .A(_262_),
    .B(_860_),
    .C(_867_),
    .Y(_107_)
);

FILL FILL_6__2159_ (
);

FILL FILL_0__2973_ (
);

FILL FILL_0__2553_ (
);

FILL FILL_6__3520_ (
);

FILL FILL_0__2133_ (
);

FILL FILL_6__3100_ (
);

FILL FILL_2__3512_ (
);

FILL FILL_7__1955_ (
);

FILL FILL_4__3018_ (
);

FILL FILL_3__1855_ (
);

FILL FILL_5__2722_ (
);

FILL FILL_5__2302_ (
);

FILL FILL_1__2714_ (
);

AND2X2 _1784_ (
    .A(state[2]),
    .B(state[3]),
    .Y(_910_)
);

FILL FILL_4__3191_ (
);

FILL FILL_5__3507_ (
);

FILL FILL_0__3091_ (
);

FILL FILL_4__1924_ (
);

NAND2X1 _2989_ (
    .A(_1150__bF$buf4),
    .B(_618_),
    .Y(_619_)
);

OAI21X1 _2569_ (
    .A(_216_),
    .B(_209_),
    .C(ADD[6]),
    .Y(_258_)
);

OAI21X1 _2149_ (
    .A(_902__bF$buf2),
    .B(_984_),
    .C(_886__bF$buf6),
    .Y(_1258_)
);

FILL FILL_7__2493_ (
);

FILL FILL_0__1824_ (
);

NAND2X1 _3510_ (
    .A(BI[3]),
    .B(_1718_),
    .Y(_1540_)
);

FILL FILL_3__2393_ (
);

FILL FILL_4__2709_ (
);

FILL FILL_5__3260_ (
);

FILL FILL_7__3278_ (
);

FILL FILL_0__2609_ (
);

FILL FILL_1__3672_ (
);

FILL FILL_1__3252_ (
);

FILL FILL_3__3598_ (
);

FILL FILL_3__3178_ (
);

FILL FILL_4__2882_ (
);

FILL FILL_4__2462_ (
);

FILL FILL_4__2042_ (
);

FILL FILL_6__2388_ (
);

FILL FILL_0__2782_ (
);

FILL FILL_0__2362_ (
);

FILL FILL_7__1764_ (
);

FILL FILL_4__3667_ (
);

FILL FILL_4__3247_ (
);

FILL FILL_0__3567_ (
);

FILL FILL_0__3147_ (
);

FILL FILL_4_BUFX2_insert70 (
);

FILL FILL_4_BUFX2_insert71 (
);

FILL FILL_4_BUFX2_insert72 (
);

FILL FILL_4_BUFX2_insert73 (
);

FILL FILL_4_BUFX2_insert74 (
);

FILL FILL_4_BUFX2_insert75 (
);

FILL FILL_4_BUFX2_insert76 (
);

FILL FILL_4_BUFX2_insert77 (
);

FILL FILL_4_BUFX2_insert78 (
);

FILL FILL_4_BUFX2_insert79 (
);

FILL FILL_5__2951_ (
);

FILL FILL_7__2969_ (
);

FILL FILL_5__2531_ (
);

FILL FILL_7__2129_ (
);

FILL FILL_5__2111_ (
);

FILL FILL_1__2943_ (
);

FILL FILL_1__2523_ (
);

FILL FILL_1__2103_ (
);

FILL FILL_3__2869_ (
);

FILL FILL_3__2449_ (
);

FILL FILL_3__2029_ (
);

FILL FILL_5__3316_ (
);

FILL FILL_1__3308_ (
);

OAI21X1 _2798_ (
    .A(_291_),
    .B(_378_),
    .C(_460_),
    .Y(_461_)
);

NAND3X1 _2378_ (
    .A(_1325_),
    .B(_1250_),
    .C(_1483_),
    .Y(_1484_)
);

FILL FILL_6__2600_ (
);

FILL FILL_4__2938_ (
);

FILL FILL_4__2518_ (
);

FILL FILL_0__2838_ (
);

FILL FILL_0__2418_ (
);

FILL FILL_1__3481_ (
);

FILL FILL_1__3061_ (
);

FILL FILL_5__1802_ (
);

FILL FILL_4__2691_ (
);

FILL FILL_4__2271_ (
);

FILL FILL_6__2197_ (
);

FILL FILL_0__2591_ (
);

FILL FILL_2__2189_ (
);

FILL FILL_0__2171_ (
);

FILL FILL_2__3550_ (
);

FILL FILL_2__3130_ (
);

FILL FILL_7__1993_ (
);

FILL FILL_4__3476_ (
);

FILL FILL_4__3056_ (
);

FILL FILL_3__1893_ (
);

FILL FILL_7__2778_ (
);

FILL FILL_5__2760_ (
);

FILL FILL_7__2358_ (
);

FILL FILL_5__2340_ (
);

FILL FILL_1__2752_ (
);

FILL FILL_1__2332_ (
);

FILL FILL_3__2678_ (
);

FILL FILL_3__2258_ (
);

FILL FILL_5__3545_ (
);

FILL FILL_5__3125_ (
);

FILL FILL_1__3537_ (
);

FILL FILL_1__3117_ (
);

FILL FILL_4__1962_ (
);

FILL FILL_6__1888_ (
);

OR2X2 _2187_ (
    .A(CO),
    .B(backwards),
    .Y(_1296_)
);

FILL FILL_0__1862_ (
);

FILL FILL_2__2821_ (
);

FILL FILL_2__2401_ (
);

FILL FILL_4__2747_ (
);

FILL FILL_4__2327_ (
);

FILL FILL_0__2647_ (
);

FILL FILL_6__3614_ (
);

FILL FILL_0__2227_ (
);

FILL FILL_1__3290_ (
);

FILL FILL_2__3606_ (
);

FILL FILL169950x136950 (
);

FILL FILL_3__1949_ (
);

FILL FILL_4__2080_ (
);

FILL FILL_5__2816_ (
);

FILL FILL_1__2808_ (
);

NOR2X1 _1878_ (
    .A(_995_),
    .B(_1002_),
    .Y(_1003_)
);

FILL FILL_4__3285_ (
);

FILL FILL_0__3185_ (
);

FILL FILL_7__2587_ (
);

FILL FILL_7__2167_ (
);

FILL FILL_0__1918_ (
);

OAI21X1 _3604_ (
    .A(_1738_),
    .B(_1633_),
    .C(_1631_),
    .Y(_1634_)
);

FILL FILL_1__2981_ (
);

FILL FILL_1__2561_ (
);

FILL FILL_1__2141_ (
);

FILL FILL_3__2487_ (
);

FILL FILL_3__2067_ (
);

FILL FILL_4__1771_ (
);

FILL FILL167550x133350 (
);

FILL FILL_2__2630_ (
);

FILL FILL_2__2210_ (
);

FILL FILL_4__2976_ (
);

FILL FILL_4__2556_ (
);

FILL FILL_4__2136_ (
);

FILL FILL_0__2876_ (
);

FILL FILL_0__2456_ (
);

FILL FILL_0__2036_ (
);

FILL FILL_6__3003_ (
);

FILL FILL_5__1840_ (
);

FILL FILL_7__1858_ (
);

FILL FILL_1__1832_ (
);

FILL FILL_3__1758_ (
);

FILL FILL_5__2625_ (
);

FILL FILL_5__2205_ (
);

FILL FILL_1__2617_ (
);

FILL FILL_4__3094_ (
);

FILL FILL_2__1901_ (
);

FILL FILL_4__1827_ (
);

FILL FILL_7__2396_ (
);

DFFSR _3413_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_82_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[1] [5])
);

FILL FILL_1__2790_ (
);

FILL FILL_1__2370_ (
);

FILL FILL_3__2296_ (
);

FILL FILL_5__3583_ (
);

FILL FILL_5__3163_ (
);

FILL FILL_1__3575_ (
);

FILL FILL_1__3155_ (
);

FILL FILL_4__2785_ (
);

FILL FILL_4__2365_ (
);

FILL FILL_0__2685_ (
);

FILL FILL_6__3652_ (
);

FILL FILL_0__2265_ (
);

FILL FILL_6__3232_ (
);

FILL FILL_2__3644_ (
);

FILL FILL_2__3224_ (
);

FILL FILL_3__1987_ (
);

FILL FILL_5__2854_ (
);

FILL FILL_5__2434_ (
);

FILL FILL_5__2014_ (
);

FILL FILL_1__2846_ (
);

FILL FILL_1__2426_ (
);

FILL FILL_1__2006_ (
);

FILL FILL_3__3713_ (
);

FILL FILL_5__3639_ (
);

FILL FILL_5__3219_ (
);

FILL FILL_0__1956_ (
);

FILL FILL_6__2923_ (
);

OAI21X1 _3642_ (
    .A(_1634_),
    .B(_1671_),
    .C(_1631_),
    .Y(_1672_)
);

FILL FILL_6__2503_ (
);

AOI21X1 _3222_ (
    .A(_787_),
    .B(_798_),
    .C(_806_),
    .Y(_92_)
);

FILL FILL_2__2915_ (
);

FILL FILL_6__3708_ (
);

FILL FILL_4__2594_ (
);

FILL FILL_4__2174_ (
);

FILL FILL_0__2494_ (
);

FILL FILL_6__3461_ (
);

FILL FILL_0__2074_ (
);

FILL FILL_6__3041_ (
);

FILL FILL_2__3453_ (
);

FILL FILL_2__3033_ (
);

OAI21X1 _2913_ (
    .A(_1149__bF$buf2),
    .B(_557_),
    .C(_558_),
    .Y(_31_)
);

FILL FILL_1__1870_ (
);

FILL FILL_3__1796_ (
);

FILL FILL_0__3699_ (
);

FILL FILL_0__3279_ (
);

FILL FILL_5__2663_ (
);

FILL FILL_5__2243_ (
);

FILL FILL_1__2655_ (
);

FILL FILL_7__3622_ (
);

FILL FILL_1__2235_ (
);

FILL FILL_3__3522_ (
);

FILL FILL_3__3102_ (
);

FILL FILL_5__3028_ (
);

FILL FILL_4__1865_ (
);

FILL FILL_0__1765_ (
);

FILL FILL_6__2732_ (
);

NOR2X1 _3451_ (
    .A(AN),
    .B(ADD[6]),
    .Y(_1700_)
);

FILL FILL_6__2312_ (
);

OAI21X1 _3031_ (
    .A(_1010_),
    .B(_647_),
    .C(_651_),
    .Y(_56_)
);

FILL FILL_2__2724_ (
);

FILL FILL_2__2304_ (
);

FILL FILL_6__3517_ (
);

FILL FILL_1__3193_ (
);

FILL FILL_2__3509_ (
);

FILL FILL_5__1934_ (
);

FILL FILL_1__1926_ (
);

FILL FILL168450x32550 (
);

FILL FILL_5__2719_ (
);

FILL FILL_6__3270_ (
);

FILL FILL_2__3262_ (
);

FILL FILL_4__3188_ (
);

AOI21X1 _2722_ (
    .A(_322_),
    .B(ADD[6]),
    .C(_390_),
    .Y(_391_)
);

INVX1 _2302_ (
    .A(_1351_),
    .Y(_1409_)
);

FILL FILL_0__3088_ (
);

FILL FILL_5__2892_ (
);

FILL FILL_5__2472_ (
);

FILL FILL_5__2052_ (
);

INVX1 _3507_ (
    .A(AI[4]),
    .Y(_1537_)
);

FILL FILL_1__2884_ (
);

FILL FILL_1__2464_ (
);

FILL FILL_1__2044_ (
);

FILL FILL_7__3011_ (
);

FILL FILL_5__3677_ (
);

FILL FILL_5__3257_ (
);

FILL FILL_1__3669_ (
);

FILL FILL_1__3249_ (
);

FILL FILL_0__1994_ (
);

FILL FILL_6__2961_ (
);

FILL FILL_6__2541_ (
);

DFFSR _3680_ (
    .R(_1513_),
    .S(vdd),
    .D(_1515_),
    .CLK(clk_bF$buf6),
    .Q(CO)
);

AOI21X1 _3260_ (
    .A(_1221_),
    .B(_969_),
    .C(_1424_),
    .Y(_836_)
);

FILL FILL_6__2121_ (
);

FILL FILL_2__2953_ (
);

FILL FILL_2__2533_ (
);

FILL FILL_2__2113_ (
);

FILL FILL_4__2879_ (
);

FILL FILL_4__2459_ (
);

FILL FILL_4__2039_ (
);

FILL FILL_0__2779_ (
);

FILL FILL_0__2359_ (
);

FILL FILL_0__3300_ (
);

FILL FILL_3__2602_ (
);

FILL FILL_5__2948_ (
);

FILL FILL_5__2528_ (
);

FILL FILL_5__2108_ (
);

FILL FILL_2__3491_ (
);

FILL FILL_2__3071_ (
);

FILL FILL_6__1812_ (
);

AOI22X1 _2951_ (
    .A(compare),
    .B(_1149__bF$buf4),
    .C(_569_),
    .D(_589_),
    .Y(_590_)
);

INVX1 _2531_ (
    .A(_225_),
    .Y(_1741_[0])
);

NAND3X1 _2111_ (
    .A(_1150__bF$buf0),
    .B(_1178_),
    .C(_1219_),
    .Y(_1220_)
);

FILL FILL_2__1804_ (
);

FILL FILL_5__2281_ (
);

NAND2X1 _3316_ (
    .A(_1741_[15]),
    .B(_869_),
    .Y(_877_)
);

FILL FILL_1__2693_ (
);

FILL FILL_1__2273_ (
);

FILL FILL_7__3240_ (
);

FILL FILL_3__2199_ (
);

FILL FILL_3__3560_ (
);

FILL FILL_3__3140_ (
);

FILL FILL_5__3486_ (
);

FILL FILL_5__3066_ (
);

FILL FILL_1__3478_ (
);

FILL FILL_1__3058_ (
);

FILL FILL_6__2770_ (
);

FILL FILL_6__2350_ (
);

FILL FILL_2__2762_ (
);

FILL FILL_2__2342_ (
);

FILL FILL_4__2688_ (
);

FILL FILL_4__2268_ (
);

NAND2X1 _1802_ (
    .A(_927_),
    .B(_926_),
    .Y(_928_)
);

FILL FILL_0__2588_ (
);

FILL FILL_6__3555_ (
);

FILL FILL_0__2168_ (
);

FILL FILL_6__3135_ (
);

FILL FILL_2__3547_ (
);

FILL FILL_2__3127_ (
);

FILL FILL_5__1972_ (
);

FILL FILL_1__1964_ (
);

FILL FILL_7__2511_ (
);

FILL FILL_3__2831_ (
);

FILL FILL_3__2411_ (
);

FILL FILL_5__2757_ (
);

FILL FILL_5__2337_ (
);

FILL FILL169950x93750 (
);

FILL FILL_1__2749_ (
);

FILL FILL_1__2329_ (
);

FILL FILL_3__3616_ (
);

OAI21X1 _2760_ (
    .A(_966_),
    .B(_351_),
    .C(_425_),
    .Y(_426_)
);

OAI21X1 _2340_ (
    .A(_931__bF$buf1),
    .B(_928_),
    .C(_886__bF$buf0),
    .Y(_1447_)
);

FILL FILL_4__1959_ (
);

FILL FILL_5__2090_ (
);

FILL FILL_4__2900_ (
);

FILL FILL168750x150 (
);

FILL FILL_0__1859_ (
);

FILL FILL_6__2826_ (
);

INVX1 _3545_ (
    .A(BI[0]),
    .Y(_1575_)
);

FILL FILL_6__2406_ (
);

OAI21X1 _3125_ (
    .A(_731_),
    .B(_730_),
    .C(ADD[1]),
    .Y(_732_)
);

FILL FILL_1__2082_ (
);

FILL FILL_0__2800_ (
);

FILL FILL_2__2818_ (
);

FILL FILL_5__3295_ (
);

FILL FILL_1__3287_ (
);

FILL FILL_2__2991_ (
);

FILL FILL_2__2571_ (
);

FILL FILL_2__2151_ (
);

FILL FILL_4__2497_ (
);

FILL FILL_4__2077_ (
);

FILL FILL168750x75750 (
);

FILL FILL_0__2397_ (
);

FILL FILL_5__1781_ (
);

AND2X2 _2816_ (
    .A(_445_),
    .B(_1110_),
    .Y(_479_)
);

FILL FILL_1__1773_ (
);

FILL FILL_7__2740_ (
);

FILL FILL_3__2640_ (
);

FILL FILL_3__2220_ (
);

FILL FILL_5__2986_ (
);

FILL FILL_5__2566_ (
);

FILL FILL_5__2146_ (
);

FILL FILL_1__2978_ (
);

FILL FILL_1__2558_ (
);

FILL FILL_7__3525_ (
);

FILL FILL_1__2138_ (
);

FILL FILL_3__3005_ (
);

FILL FILL_6__1850_ (
);

FILL FILL_2__1842_ (
);

FILL FILL_4__1768_ (
);

FILL FILL_6__2635_ (
);

DFFSR _3354_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_31_),
    .CLK(clk_bF$buf10),
    .Q(bit_ins)
);

FILL FILL_6__2215_ (
);

FILL FILL_2__2627_ (
);

FILL FILL_2__2207_ (
);

FILL FILL_1__3096_ (
);

FILL FILL_3__1911_ (
);

FILL FILL_5__1837_ (
);

FILL FILL_1__1829_ (
);

FILL FILL_2__2380_ (
);

INVX1 _1840_ (
    .A(PC[0]),
    .Y(_965_)
);

FILL FILL_6__3593_ (
);

FILL FILL_6__3173_ (
);

FILL FILL_2__3585_ (
);

FILL FILL_2__3165_ (
);

FILL FILL_6__1906_ (
);

AOI21X1 _2625_ (
    .A(_198_),
    .B(AN),
    .C(_1145_),
    .Y(_305_)
);

OAI21X1 _2205_ (
    .A(RDY_bF$buf1),
    .B(_1021_),
    .C(_1313_),
    .Y(_1314_)
);

FILL FILL_5__2795_ (
);

FILL FILL_5__2375_ (
);

FILL FILL_1__2787_ (
);

FILL FILL_1__2367_ (
);

FILL FILL_3__3654_ (
);

FILL FILL_3__3234_ (
);

FILL FILL_4__1997_ (
);

FILL FILL_0__1897_ (
);

FILL FILL_6__2864_ (
);

NOR2X1 _3583_ (
    .A(_1610_),
    .B(_1580_),
    .Y(_1613_)
);

FILL FILL_6__2444_ (
);

FILL FILL_6__2024_ (
);

NOR2X1 _3163_ (
    .A(_1319__bF$buf1),
    .B(_765_),
    .Y(_766_)
);

FILL FILL_2__2856_ (
);

FILL FILL_2__2436_ (
);

FILL FILL_2__2016_ (
);

FILL FILL_4__3303_ (
);

FILL FILL_6__3649_ (
);

FILL FILL_6__3229_ (
);

FILL FILL_0__3623_ (
);

FILL FILL_0__3203_ (
);

FILL FILL_3__2925_ (
);

FILL FILL_3__2505_ (
);

NOR2X1 _2854_ (
    .A(_304_),
    .B(_418_),
    .Y(_514_)
);

NAND2X1 _2434_ (
    .A(_139_),
    .B(_138_),
    .Y(alu_op[2])
);

NAND2X1 _2014_ (
    .A(ABH[5]),
    .B(_925_),
    .Y(_1126_)
);

FILL FILL_5__2184_ (
);

OAI21X1 _3639_ (
    .A(_1667_),
    .B(_1664_),
    .C(_1668_),
    .Y(_1669_)
);

NOR2X1 _3219_ (
    .A(\AXYS[2] [6]),
    .B(_798_),
    .Y(_805_)
);

FILL FILL_1__2596_ (
);

FILL FILL_7__3563_ (
);

FILL FILL_1__2176_ (
);

FILL FILL_7__3143_ (
);

FILL FILL_3__3463_ (
);

FILL FILL_3__3043_ (
);

FILL FILL_2__1880_ (
);

FILL FILL_6__2673_ (
);

DFFSR _3392_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_61_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD_valid)
);

FILL FILL_6__2253_ (
);

FILL FILL_2__2665_ (
);

FILL FILL_2__2245_ (
);

FILL FILL_4__3532_ (
);

FILL FILL_4__3112_ (
);

FILL FILL_6__3458_ (
);

FILL FILL_6__3038_ (
);

FILL FILL_0__3012_ (
);

FILL FILL_5__1875_ (
);

FILL FILL_1__1867_ (
);

FILL FILL_7__2414_ (
);

FILL FILL_3__2734_ (
);

FILL FILL_3__2314_ (
);

FILL FILL_5__3601_ (
);

FILL FILL_7__3619_ (
);

FILL FILL_3__3519_ (
);

FILL FILL_6__1944_ (
);

AOI21X1 _2663_ (
    .A(_322_),
    .B(ADD[1]),
    .C(_336_),
    .Y(_337_)
);

NOR2X1 _2243_ (
    .A(_1160_),
    .B(_1328_),
    .Y(_1351_)
);

FILL FILL_2__1936_ (
);

FILL FILL_4__2803_ (
);

FILL FILL_6__2729_ (
);

DFFSR _3448_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_116_),
    .CLK(clk_bF$buf0),
    .Q(ABH[7])
);

FILL FILL_6__2309_ (
);

OAI21X1 _3028_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[2]),
    .Y(_650_)
);

FILL FILL_0__2703_ (
);

FILL FILL_3__3692_ (
);

FILL FILL_3__3272_ (
);

FILL FILL_5__3198_ (
);

FILL FILL_6__2482_ (
);

FILL FILL_6__2062_ (
);

FILL FILL_2__2894_ (
);

FILL FILL_2__2474_ (
);

FILL FILL_2__2054_ (
);

AND2X2 _1934_ (
    .A(_1048_),
    .B(_1039_),
    .Y(_1051_)
);

FILL FILL_6__3267_ (
);

FILL FILL_0__3661_ (
);

FILL FILL_2__3259_ (
);

FILL FILL_0__3241_ (
);

OAI21X1 _2719_ (
    .A(RDY_bF$buf3),
    .B(_1012_),
    .C(_388_),
    .Y(_7_)
);

FILL FILL_7__2643_ (
);

FILL FILL_3__2963_ (
);

FILL FILL_3__2543_ (
);

FILL FILL_3__2123_ (
);

FILL FILL_5__2889_ (
);

FILL FILL_5__2469_ (
);

FILL FILL_5__2049_ (
);

FILL FILL_6__1753_ (
);

NOR2X1 _2892_ (
    .A(_1185_),
    .B(_1412_),
    .Y(_543_)
);

AOI21X1 _2472_ (
    .A(PC[4]),
    .B(_1080_),
    .C(_154_),
    .Y(_171_)
);

INVX1 _2052_ (
    .A(_1160_),
    .Y(_1161_)
);

FILL FILL169950x25350 (
);

FILL FILL_2__1745_ (
);

FILL FILL_4__2612_ (
);

FILL FILL_6__2958_ (
);

NAND2X1 _3677_ (
    .A(AI[7]),
    .B(RDY_bF$buf7),
    .Y(_1697_)
);

FILL FILL_6__2538_ (
);

FILL FILL_6__2118_ (
);

NOR2X1 _3257_ (
    .A(_950_),
    .B(_832_),
    .Y(_833_)
);

FILL FILL_0__2932_ (
);

FILL FILL_0__2512_ (
);

FILL FILL_3__3081_ (
);

FILL FILL_7__1914_ (
);

FILL FILL_3__1814_ (
);

FILL FILL_6__2291_ (
);

FILL FILL_2__2283_ (
);

FILL FILL_4__3570_ (
);

FILL FILL_4__3150_ (
);

FILL FILL_6__3496_ (
);

FILL FILL_6__3076_ (
);

FILL FILL_2__3488_ (
);

FILL FILL_0__3470_ (
);

FILL FILL_0__3050_ (
);

FILL FILL_2__3068_ (
);

FILL FILL_6__1809_ (
);

OAI22X1 _2948_ (
    .A(_920_),
    .B(_1150__bF$buf2),
    .C(_588_),
    .D(_565_),
    .Y(_36_)
);

AND2X2 _2528_ (
    .A(_219_),
    .B(_222_),
    .Y(_223_)
);

INVX2 _2108_ (
    .A(_1185_),
    .Y(_1217_)
);

FILL FILL_7__2872_ (
);

FILL FILL_7__2032_ (
);

FILL FILL_3__2772_ (
);

FILL FILL_3__2352_ (
);

FILL FILL_5__2698_ (
);

FILL FILL_5__2278_ (
);

FILL FILL_1__3631_ (
);

FILL FILL_1__3211_ (
);

FILL FILL_3__3557_ (
);

FILL FILL_3__3137_ (
);

FILL FILL_6__1982_ (
);

OAI21X1 _2281_ (
    .A(RDY_bF$buf6),
    .B(_1092_),
    .C(_1388_),
    .Y(_1389_)
);

FILL FILL_2__1974_ (
);

FILL FILL_4__2841_ (
);

FILL FILL_4__2421_ (
);

FILL FILL_4__2001_ (
);

FILL FILL_6__2767_ (
);

OAI21X1 _3486_ (
    .A(_1714__bF$buf2),
    .B(_1730_),
    .C(_1731_),
    .Y(_1514_)
);

FILL FILL_6__2347_ (
);

AOI21X1 _3066_ (
    .A(_658_),
    .B(_1344_),
    .C(_661_),
    .Y(_679_)
);

FILL FILL_0__2741_ (
);

FILL FILL_2__2759_ (
);

FILL FILL_0__2321_ (
);

FILL FILL_2__2339_ (
);

FILL FILL_2__3700_ (
);

FILL FILL_4__3626_ (
);

FILL FILL_4__3206_ (
);

FILL FILL_0__3526_ (
);

FILL FILL_0__3106_ (
);

FILL FILL_5__1969_ (
);

FILL FILL_7__2928_ (
);

FILL FILL_5__2910_ (
);

FILL FILL_7__2508_ (
);

FILL FILL_2__2092_ (
);

FILL FILL_1__2902_ (
);

FILL FILL_3__2828_ (
);

FILL FILL_3__2408_ (
);

NAND3X1 _1972_ (
    .A(\AXYS[0] [1]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1088_)
);

FILL FILL_2__3297_ (
);

FILL FILL168750x136950 (
);

OAI21X1 _2757_ (
    .A(_276_),
    .B(_418_),
    .C(_422_),
    .Y(_423_)
);

INVX1 _2337_ (
    .A(_988_),
    .Y(_1444_)
);

FILL FILL_7__2261_ (
);

FILL FILL_3__2581_ (
);

FILL FILL_3__2161_ (
);

FILL FILL_5__2087_ (
);

FILL FILL_1__2499_ (
);

FILL FILL_7__3466_ (
);

FILL FILL_1__2079_ (
);

FILL FILL_7__3046_ (
);

FILL FILL_1__3020_ (
);

FILL FILL_6__1791_ (
);

NOR2X1 _2090_ (
    .A(_901_),
    .B(_974_),
    .Y(_1199_)
);

FILL FILL_2__1783_ (
);

FILL FILL_4__2650_ (
);

FILL FILL_4__2230_ (
);

FILL FILL_6__2996_ (
);

FILL FILL_6__2576_ (
);

NAND2X1 _3295_ (
    .A(ABL[5]),
    .B(_860_),
    .Y(_866_)
);

FILL FILL_6__2156_ (
);

FILL FILL_0__2970_ (
);

FILL FILL_2__2988_ (
);

FILL FILL_0__2550_ (
);

FILL FILL_2__2568_ (
);

FILL FILL_2__2148_ (
);

FILL FILL_0__2130_ (
);

FILL FILL_4__3015_ (
);

FILL FILL_3__1852_ (
);

FILL FILL_5__1778_ (
);

FILL FILL_7__2737_ (
);

FILL FILL_7__2317_ (
);

FILL FILL_1__2711_ (
);

FILL FILL_3__2637_ (
);

FILL FILL_3__2217_ (
);

NAND2X1 _1781_ (
    .A(_905_),
    .B(_906_),
    .Y(_907_)
);

FILL FILL_5__3504_ (
);

FILL FILL_4__1921_ (
);

FILL FILL_6__1847_ (
);

OAI21X1 _2986_ (
    .A(_530_),
    .B(_612_),
    .C(_615_),
    .Y(_616_)
);

OAI21X1 _2566_ (
    .A(_1012_),
    .B(_218_),
    .C(_255_),
    .Y(_256_)
);

NOR2X1 _2146_ (
    .A(_1178_),
    .B(_1175_),
    .Y(_1255_)
);

FILL FILL_7__2490_ (
);

FILL FILL_2__1839_ (
);

FILL FILL_0__1821_ (
);

FILL FILL_3__2390_ (
);

FILL FILL169050x75750 (
);

FILL FILL_4__2706_ (
);

FILL FILL_7__3695_ (
);

FILL FILL_7__3275_ (
);

FILL FILL_0__2606_ (
);

FILL FILL_3__3595_ (
);

FILL FILL_3__3175_ (
);

FILL FILL_3__1908_ (
);

FILL FILL_6__2385_ (
);

FILL FILL_2__2797_ (
);

FILL FILL_2__2377_ (
);

NAND2X1 _1837_ (
    .A(_933_),
    .B(_962_),
    .Y(_963_)
);

FILL FILL_7__1761_ (
);

FILL FILL_4__3664_ (
);

FILL FILL_4__3244_ (
);

FILL FILL_0__3564_ (
);

FILL FILL_0__3144_ (
);

FILL FILL_4_BUFX2_insert40 (
);

FILL FILL_4_BUFX2_insert41 (
);

FILL FILL_4_BUFX2_insert42 (
);

FILL FILL_4_BUFX2_insert43 (
);

FILL FILL_4_BUFX2_insert44 (
);

FILL FILL_4_BUFX2_insert45 (
);

FILL FILL_4_BUFX2_insert46 (
);

FILL FILL_4_BUFX2_insert47 (
);

FILL FILL_1__1999_ (
);

FILL FILL_4_BUFX2_insert48 (
);

FILL FILL_4_BUFX2_insert49 (
);

FILL FILL_7__2966_ (
);

FILL FILL_7__2546_ (
);

FILL FILL_1__2940_ (
);

FILL FILL_1__2520_ (
);

FILL FILL_1__2100_ (
);

FILL FILL_3__2866_ (
);

FILL FILL_3__2446_ (
);

FILL FILL_3__2026_ (
);

FILL FILL_5__3313_ (
);

FILL FILL_1__3305_ (
);

NAND2X1 _2795_ (
    .A(PC[12]),
    .B(_886__bF$buf3),
    .Y(_458_)
);

OR2X2 _2375_ (
    .A(_1408_),
    .B(_1149__bF$buf3),
    .Y(_1481_)
);

FILL FILL_4__2935_ (
);

FILL FILL_4__2515_ (
);

FILL FILL_0__2835_ (
);

FILL FILL_0__2415_ (
);

FILL FILL_6__2194_ (
);

FILL FILL_2__2186_ (
);

FILL FILL_7__1990_ (
);

FILL FILL_4__3473_ (
);

FILL FILL_4__3053_ (
);

FILL FILL_3__1890_ (
);

FILL FILL_7__2775_ (
);

FILL FILL_3__2675_ (
);

FILL FILL_3__2255_ (
);

FILL FILL_5__3542_ (
);

FILL FILL_5__3122_ (
);

FILL FILL_1__3534_ (
);

FILL FILL_1__3114_ (
);

FILL FILL_6__1885_ (
);

OAI21X1 _2184_ (
    .A(_886__bF$buf4),
    .B(_1290_),
    .C(_1292_),
    .Y(_1293_)
);

FILL FILL_2__1877_ (
);

FILL FILL_4__2744_ (
);

FILL FILL_4__2324_ (
);

DFFPOSX1 _3389_ (
    .D(_58_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD[5])
);

FILL FILL_0__2644_ (
);

FILL FILL_6__3611_ (
);

FILL FILL_0__2224_ (
);

FILL FILL_2__3603_ (
);

FILL FILL_4__3529_ (
);

FILL FILL_4__3109_ (
);

FILL FILL_3__1946_ (
);

FILL FILL_0__3009_ (
);

FILL FILL_6_CLKBUF1_insert26 (
);

FILL FILL_6_CLKBUF1_insert27 (
);

FILL FILL_6_CLKBUF1_insert28 (
);

FILL FILL_6_CLKBUF1_insert29 (
);

FILL FILL_5__2813_ (
);

FILL FILL_1__2805_ (
);

OR2X2 _1875_ (
    .A(_999_),
    .B(_998_),
    .Y(_1000_)
);

FILL FILL_4__3282_ (
);

FILL FILL_0__3182_ (
);

FILL FILL_7__2164_ (
);

FILL FILL_0__1915_ (
);

NAND2X1 _3601_ (
    .A(_1527_),
    .B(_1738_),
    .Y(_1631_)
);

FILL FILL_3__2484_ (
);

FILL FILL_3__2064_ (
);

FILL FILL_3__3269_ (
);

FILL FILL_4__2973_ (
);

FILL FILL_4__2553_ (
);

FILL FILL_4__2133_ (
);

FILL FILL_6__2899_ (
);

FILL FILL_6__2479_ (
);

OAI21X1 _3198_ (
    .A(_720__bF$buf0),
    .B(_687_),
    .C(\AXYS[1] [4]),
    .Y(_794_)
);

FILL FILL_6__2059_ (
);

FILL FILL_0__2873_ (
);

FILL FILL_0__2453_ (
);

FILL FILL_0__2033_ (
);

FILL FILL_6__3000_ (
);

FILL FILL_7__1855_ (
);

FILL FILL_0__3658_ (
);

FILL FILL_3__1755_ (
);

FILL FILL_0__3238_ (
);

FILL FILL_5__2622_ (
);

FILL FILL_5__2202_ (
);

FILL FILL_1__2614_ (
);

FILL FILL_4__3091_ (
);

FILL FILL_4__1824_ (
);

NAND2X1 _2889_ (
    .A(_1179_),
    .B(_540_),
    .Y(_541_)
);

OAI21X1 _2469_ (
    .A(_164_),
    .B(_165_),
    .C(_168_),
    .Y(_169_)
);

AOI21X1 _2049_ (
    .A(_1157_),
    .B(IRHOLD_valid),
    .C(_1154_),
    .Y(_1158_)
);

FILL FILL_7__2393_ (
);

DFFSR _3410_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_79_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[1] [2])
);

FILL FILL_3__2293_ (
);

FILL FILL_4__2609_ (
);

FILL FILL_7__3598_ (
);

FILL FILL_5__3580_ (
);

FILL FILL_5__3160_ (
);

FILL FILL_7__3178_ (
);

FILL FILL_0__2929_ (
);

FILL FILL_0__2509_ (
);

FILL FILL_1__3572_ (
);

FILL FILL_1__3152_ (
);

FILL FILL_3__3498_ (
);

FILL FILL_3__3078_ (
);

FILL FILL_4__2782_ (
);

FILL FILL_4__2362_ (
);

FILL FILL_6__2288_ (
);

FILL FILL_0__2682_ (
);

FILL FILL_0__2262_ (
);

FILL FILL_2__3641_ (
);

FILL FILL_2__3221_ (
);

FILL FILL_4__3567_ (
);

FILL FILL_4__3147_ (
);

FILL FILL_3__1984_ (
);

FILL FILL_0__3467_ (
);

FILL FILL_0__3047_ (
);

FILL FILL_5__2851_ (
);

FILL FILL_7__2869_ (
);

FILL FILL_5__2431_ (
);

FILL FILL_5__2011_ (
);

FILL FILL_7__2029_ (
);

FILL FILL_1__2843_ (
);

FILL FILL_1__2423_ (
);

FILL FILL_1__2003_ (
);

FILL FILL_3__2769_ (
);

FILL FILL_3__2349_ (
);

FILL FILL_3__3710_ (
);

FILL FILL_5__3636_ (
);

FILL FILL_5__3216_ (
);

FILL FILL_1__3628_ (
);

FILL FILL_1__3208_ (
);

FILL FILL_6__1979_ (
);

AOI22X1 _2698_ (
    .A(_367_),
    .B(_368_),
    .C(_346_),
    .D(_366_),
    .Y(_369_)
);

INVX1 _2278_ (
    .A(_1385_),
    .Y(_1386_)
);

FILL FILL_0__1953_ (
);

FILL FILL_6__2920_ (
);

FILL FILL_6__2500_ (
);

FILL FILL_2__2912_ (
);

FILL FILL_4__2838_ (
);

FILL FILL_4__2418_ (
);

FILL FILL_0__2738_ (
);

FILL FILL_6__3705_ (
);

FILL FILL_0__2318_ (
);

FILL FILL_4__2591_ (
);

FILL FILL_4__2171_ (
);

FILL FILL_6__2097_ (
);

FILL FILL_5__2907_ (
);

FILL FILL_0__2491_ (
);

FILL FILL_0__2071_ (
);

FILL FILL_2__2089_ (
);

FILL FILL_2__3450_ (
);

OAI21X1 _1969_ (
    .A(_1074_),
    .B(_1060_),
    .C(_1085_),
    .Y(AI[0])
);

FILL FILL_2__3030_ (
);

FILL FILL_7__1893_ (
);

NOR2X1 _2910_ (
    .A(_555_),
    .B(_554_),
    .Y(_556_)
);

FILL FILL_0__3696_ (
);

FILL FILL_3__1793_ (
);

FILL FILL_0__3276_ (
);

FILL FILL_5__2660_ (
);

FILL FILL_7__2258_ (
);

FILL FILL_5__2240_ (
);

FILL FILL_1__2652_ (
);

FILL FILL_1__2232_ (
);

FILL FILL_3__2998_ (
);

FILL FILL_3__2578_ (
);

FILL FILL_3__2158_ (
);

FILL FILL_5__3025_ (
);

FILL FILL_1__3017_ (
);

FILL FILL_4__1862_ (
);

FILL FILL_6__1788_ (
);

NOR2X1 _2087_ (
    .A(_931__bF$buf3),
    .B(_946_),
    .Y(_1196_)
);

FILL FILL_0__1762_ (
);

FILL FILL_2__2721_ (
);

FILL FILL_2__2301_ (
);

FILL FILL_4__2647_ (
);

FILL FILL_4__2227_ (
);

FILL FILL_0__2967_ (
);

FILL FILL_0__2547_ (
);

FILL FILL_6__3514_ (
);

FILL FILL_0__2127_ (
);

FILL FILL_1__3190_ (
);

FILL FILL_2__3506_ (
);

FILL FILL_5__1931_ (
);

FILL FILL167850x133350 (
);

FILL FILL_1__1923_ (
);

FILL FILL_3__1849_ (
);

FILL FILL_5__2716_ (
);

FILL FILL_1__2708_ (
);

NAND2X1 _1778_ (
    .A(state[2]),
    .B(_897_),
    .Y(_904_)
);

FILL FILL_4__3185_ (
);

FILL FILL_0__3085_ (
);

FILL FILL_4__1918_ (
);

FILL FILL_7__2487_ (
);

FILL FILL_7__2067_ (
);

FILL FILL_0__1818_ (
);

OAI21X1 _3504_ (
    .A(alu_op[3]),
    .B(BI[4]),
    .C(_1740_),
    .Y(_1534_)
);

FILL FILL_1__2881_ (
);

FILL FILL_1__2461_ (
);

FILL FILL_1__2041_ (
);

FILL FILL_3__2387_ (
);

FILL FILL_5__3674_ (
);

FILL FILL_5__3254_ (
);

FILL FILL_1__3666_ (
);

FILL FILL_1__3246_ (
);

FILL FILL_0__1991_ (
);

FILL FILL_2__2950_ (
);

FILL FILL_2__2530_ (
);

FILL FILL_2__2110_ (
);

FILL FILL_4__2876_ (
);

FILL FILL_4__2456_ (
);

FILL FILL_4__2036_ (
);

FILL FILL_0__2776_ (
);

FILL FILL_0__2356_ (
);

FILL FILL_2__3315_ (
);

FILL FILL_7__1758_ (
);

FILL FILL_5__2945_ (
);

FILL FILL_5__2525_ (
);

FILL FILL_5__2105_ (
);

FILL FILL_1__2937_ (
);

FILL FILL_1__2517_ (
);

FILL FILL_2__1801_ (
);

FILL FILL_7__2296_ (
);

OAI21X1 _3313_ (
    .A(_296_),
    .B(_869_),
    .C(_875_),
    .Y(_114_)
);

FILL FILL_1__2690_ (
);

FILL FILL_1__2270_ (
);

FILL FILL_3__2196_ (
);

FILL FILL169950x122550 (
);

FILL FILL_5__3483_ (
);

FILL FILL_5__3063_ (
);

FILL FILL_1__3475_ (
);

FILL FILL_1__3055_ (
);

FILL FILL_5_CLKBUF1_insert30 (
);

FILL FILL_5_CLKBUF1_insert31 (
);

FILL FILL_5_CLKBUF1_insert32 (
);

FILL FILL_5_CLKBUF1_insert33 (
);

FILL FILL_5_CLKBUF1_insert34 (
);

FILL FILL_5_CLKBUF1_insert35 (
);

FILL FILL_5_CLKBUF1_insert36 (
);

FILL FILL_4__2685_ (
);

FILL FILL_4__2265_ (
);

FILL FILL_0__2585_ (
);

FILL FILL_6__3552_ (
);

FILL FILL_0__2165_ (
);

FILL FILL_6__3132_ (
);

FILL FILL_2__3544_ (
);

FILL FILL_2__3124_ (
);

FILL FILL_7__1987_ (
);

FILL FILL_1__1961_ (
);

FILL FILL_3__1887_ (
);

FILL FILL_5__2754_ (
);

FILL FILL_5__2334_ (
);

FILL FILL_1__2746_ (
);

FILL FILL_7__3713_ (
);

FILL FILL_1__2326_ (
);

FILL FILL_3__3613_ (
);

FILL FILL_5__3539_ (
);

FILL FILL_5__3119_ (
);

FILL FILL_4__1956_ (
);

FILL FILL_0__1856_ (
);

FILL FILL_6__2823_ (
);

NAND2X1 _3542_ (
    .A(BI[0]),
    .B(_1718_),
    .Y(_1572_)
);

FILL FILL_6__2403_ (
);

OAI21X1 _3122_ (
    .A(HC),
    .B(_728_),
    .C(_727_),
    .Y(_729_)
);

FILL FILL_2__2815_ (
);

FILL FILL_5__3292_ (
);

FILL FILL_6__3608_ (
);

FILL FILL_1__3284_ (
);

FILL FILL_4__2494_ (
);

FILL FILL_4__2074_ (
);

FILL FILL_0__2394_ (
);

FILL FILL_4__3699_ (
);

FILL FILL_4__3279_ (
);

AOI21X1 _2813_ (
    .A(PC[9]),
    .B(_312_),
    .C(_1093_),
    .Y(_476_)
);

FILL FILL_1__1770_ (
);

FILL FILL_0__3599_ (
);

FILL FILL_0__3179_ (
);

FILL FILL_5__2983_ (
);

FILL FILL_5__2563_ (
);

FILL FILL_5__2143_ (
);

FILL FILL_1__2975_ (
);

FILL FILL_1__2555_ (
);

FILL FILL_7__3522_ (
);

FILL FILL_1__2135_ (
);

FILL FILL_3__3002_ (
);

FILL FILL_4__1765_ (
);

FILL FILL_6__2632_ (
);

FILL FILL_6__2212_ (
);

DFFSR _3351_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_28_),
    .CLK(clk_bF$buf6),
    .Q(cli)
);

FILL FILL_2__2624_ (
);

FILL FILL_2__2204_ (
);

FILL FILL_1__3093_ (
);

FILL FILL_5__1834_ (
);

FILL FILL_1__1826_ (
);

FILL FILL_5__2619_ (
);

FILL FILL_6__3590_ (
);

FILL FILL_6__3170_ (
);

FILL FILL_2__3582_ (
);

FILL FILL_2__3162_ (
);

FILL FILL_4__3088_ (
);

FILL FILL_6__1903_ (
);

AOI21X1 _2622_ (
    .A(_272_),
    .B(DIMUX[6]),
    .C(_302_),
    .Y(_303_)
);

OAI21X1 _2202_ (
    .A(RDY_bF$buf1),
    .B(_1309_),
    .C(_1310_),
    .Y(_1311_)
);

FILL FILL_5__2792_ (
);

FILL FILL_5__2372_ (
);

DFFSR _3407_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_76_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[0] [7])
);

FILL FILL_1__2784_ (
);

FILL FILL_1__2364_ (
);

FILL FILL_3__3651_ (
);

FILL FILL_3__3231_ (
);

FILL FILL_5__3577_ (
);

FILL FILL_5__3157_ (
);

FILL FILL_1__3569_ (
);

FILL FILL_1__3149_ (
);

FILL FILL_4__1994_ (
);

FILL FILL_0__1894_ (
);

FILL FILL_6__2861_ (
);

AOI21X1 _3580_ (
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1581_),
    .Y(_1610_)
);

FILL FILL_6__2441_ (
);

NOR2X1 _3160_ (
    .A(CO),
    .B(_728_),
    .Y(_763_)
);

FILL FILL_6__2021_ (
);

FILL FILL_2__2853_ (
);

FILL FILL_2__2433_ (
);

FILL FILL_2__2013_ (
);

FILL FILL_4__2779_ (
);

FILL FILL_4__2359_ (
);

FILL FILL_4__3300_ (
);

FILL FILL_0__2679_ (
);

FILL FILL_6__3646_ (
);

FILL FILL_0__2259_ (
);

FILL FILL_6__3226_ (
);

FILL FILL_2__3638_ (
);

FILL FILL_0__3620_ (
);

FILL FILL_0__3200_ (
);

FILL FILL_2__3218_ (
);

FILL FILL_3__2922_ (
);

FILL FILL_3__2502_ (
);

FILL FILL_5__2848_ (
);

FILL FILL_5__2428_ (
);

FILL FILL_5__2008_ (
);

FILL FILL_3__3707_ (
);

NAND2X1 _2851_ (
    .A(_886__bF$buf3),
    .B(_300_),
    .Y(_512_)
);

OAI21X1 _2431_ (
    .A(state[5]),
    .B(_1075_),
    .C(_136_),
    .Y(_137_)
);

NAND3X1 _2011_ (
    .A(\AXYS[0] [5]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1123_)
);

FILL FILL_5__2181_ (
);

FILL FILL_6__2917_ (
);

OAI21X1 _3636_ (
    .A(_1665_),
    .B(_1600_),
    .C(_1623_),
    .Y(_1666_)
);

AOI21X1 _3216_ (
    .A(_757_),
    .B(_798_),
    .C(_803_),
    .Y(_89_)
);

FILL FILL_1__2593_ (
);

FILL FILL_1__2173_ (
);

FILL FILL_7__3140_ (
);

FILL FILL_3__2099_ (
);

FILL FILL_2__2909_ (
);

FILL FILL_3__3460_ (
);

FILL FILL_3__3040_ (
);

FILL FILL_6__2670_ (
);

FILL FILL_6__2250_ (
);

FILL FILL_2__2662_ (
);

FILL FILL_2__2242_ (
);

FILL FILL_4__2588_ (
);

FILL FILL_4__2168_ (
);

FILL FILL_0__2488_ (
);

FILL FILL_6__3455_ (
);

FILL FILL_0__2068_ (
);

FILL FILL_6__3035_ (
);

FILL FILL_2__3027_ (
);

FILL FILL_5__1872_ (
);

OAI21X1 _2907_ (
    .A(_553_),
    .B(_533_),
    .C(_549_),
    .Y(_30_)
);

FILL FILL_1__1864_ (
);

FILL FILL_7__2411_ (
);

FILL FILL_3__2731_ (
);

FILL FILL_3__2311_ (
);

FILL FILL_5__2657_ (
);

FILL FILL_5__2237_ (
);

FILL FILL_1__2649_ (
);

FILL FILL_7__3616_ (
);

FILL FILL_1__2229_ (
);

FILL FILL_3__3516_ (
);

FILL FILL_6__1941_ (
);

OAI22X1 _2660_ (
    .A(RDY_bF$buf7),
    .B(_965_),
    .C(_332_),
    .D(_334_),
    .Y(_2_)
);

INVX1 _2240_ (
    .A(_1181_),
    .Y(_1348_)
);

FILL FILL_2__1933_ (
);

FILL FILL_4__1859_ (
);

FILL FILL_4__2800_ (
);

FILL FILL_0__1759_ (
);

FILL FILL_6__2726_ (
);

DFFSR _3445_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_113_),
    .CLK(clk_bF$buf0),
    .Q(ABH[4])
);

FILL FILL_6__2306_ (
);

OAI21X1 _3025_ (
    .A(_966_),
    .B(_647_),
    .C(_648_),
    .Y(_53_)
);

FILL FILL_2__2718_ (
);

FILL FILL_0__2700_ (
);

FILL FILL_5__3195_ (
);

FILL FILL_1__3187_ (
);

FILL FILL_5__1928_ (
);

FILL FILL_2__2891_ (
);

FILL FILL_2__2471_ (
);

FILL FILL_2__2051_ (
);

FILL FILL_4__2397_ (
);

NAND3X1 _1931_ (
    .A(src_reg[1]),
    .B(_1035_),
    .C(_1026_),
    .Y(_1048_)
);

FILL FILL_0__2297_ (
);

FILL FILL_6__3264_ (
);

FILL FILL_2__3676_ (
);

FILL FILL_2__3256_ (
);

NOR3X1 _2716_ (
    .A(_362_),
    .B(_385_),
    .C(_340_),
    .Y(_386_)
);

FILL FILL_7__2640_ (
);

FILL FILL_3__2960_ (
);

FILL FILL_3__2540_ (
);

FILL FILL_3__2120_ (
);

FILL FILL_5__2886_ (
);

FILL FILL_5__2466_ (
);

FILL FILL_5__2046_ (
);

FILL FILL_1__2878_ (
);

FILL FILL_1__2458_ (
);

FILL FILL_1__2038_ (
);

FILL FILL_6__1750_ (
);

FILL FILL_0__1988_ (
);

FILL FILL_6__2955_ (
);

OAI21X1 _3674_ (
    .A(_1714__bF$buf2),
    .B(_1680_),
    .C(_1695_),
    .Y(_1523_)
);

FILL FILL_6__2535_ (
);

NOR2X1 _3254_ (
    .A(_1070_),
    .B(_829_),
    .Y(_830_)
);

FILL FILL_6__2115_ (
);

FILL FILL_2__2947_ (
);

FILL FILL_2__2527_ (
);

FILL FILL_2__2107_ (
);

FILL FILL_7__1911_ (
);

FILL FILL_0__3714_ (
);

FILL FILL_3__1811_ (
);

FILL FILL_2__2280_ (
);

FILL FILL_6__3493_ (
);

FILL FILL_6__3073_ (
);

FILL FILL_0_BUFX2_insert60 (
);

FILL FILL_0_BUFX2_insert61 (
);

FILL FILL_0_BUFX2_insert62 (
);

FILL FILL_2__3485_ (
);

FILL FILL_0_BUFX2_insert63 (
);

FILL FILL_2__3065_ (
);

FILL FILL_0_BUFX2_insert64 (
);

FILL FILL_0_BUFX2_insert65 (
);

FILL FILL_0_BUFX2_insert66 (
);

FILL FILL_0_BUFX2_insert67 (
);

FILL FILL_0_BUFX2_insert68 (
);

FILL FILL_0_BUFX2_insert69 (
);

INVX1 _2945_ (
    .A(_567_),
    .Y(_587_)
);

FILL FILL_6__1806_ (
);

OAI21X1 _2525_ (
    .A(_196_),
    .B(_198_),
    .C(ABL[0]),
    .Y(_220_)
);

INVX1 _2105_ (
    .A(_1159_),
    .Y(_1214_)
);

FILL FILL_5__2695_ (
);

FILL FILL_5__2275_ (
);

FILL FILL_1__2687_ (
);

FILL FILL_7__3654_ (
);

FILL FILL_1__2267_ (
);

FILL FILL_3__3554_ (
);

FILL FILL_3__3134_ (
);

FILL FILL_2__1971_ (
);

FILL FILL_4__1897_ (
);

FILL FILL168750x61350 (
);

FILL FILL_0__1797_ (
);

FILL FILL_6__2764_ (
);

OR2X2 _3483_ (
    .A(_1727_),
    .B(_1728_),
    .Y(_1729_)
);

FILL FILL_6__2344_ (
);

OAI21X1 _3063_ (
    .A(_672_),
    .B(_676_),
    .C(_673_),
    .Y(_63_)
);

FILL FILL_2__2756_ (
);

FILL FILL_2__2336_ (
);

FILL FILL_4__3623_ (
);

FILL FILL_4__3203_ (
);

FILL FILL_6__3549_ (
);

FILL FILL_6__3129_ (
);

FILL FILL_0__3523_ (
);

FILL FILL_0__3103_ (
);

FILL FILL_5__1966_ (
);

FILL FILL_1__1958_ (
);

FILL FILL_7__2925_ (
);

FILL FILL_3__2825_ (
);

FILL FILL_3__2405_ (
);

FILL FILL_2__3294_ (
);

AOI22X1 _2754_ (
    .A(ADD[1]),
    .B(_1299_),
    .C(_323_),
    .D(ABH[1]),
    .Y(_420_)
);

AOI21X1 _2334_ (
    .A(_1423_),
    .B(_1429_),
    .C(_1440_),
    .Y(_1441_)
);

FILL FILL169350x7350 (
);

FILL FILL_5__2084_ (
);

OAI21X1 _3539_ (
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1725_),
    .Y(_1569_)
);

AND2X2 _3119_ (
    .A(adj_bcd),
    .B(adc_bcd),
    .Y(_726_)
);

FILL FILL_1__2496_ (
);

FILL FILL_7__3463_ (
);

FILL FILL_1__2076_ (
);

FILL FILL_7__3043_ (
);

FILL FILL_5__3289_ (
);

FILL FILL_2__1780_ (
);

FILL FILL_6__2993_ (
);

FILL FILL_6__2573_ (
);

OAI21X1 _3292_ (
    .A(_860_),
    .B(_242_),
    .C(_864_),
    .Y(_104_)
);

FILL FILL_6__2153_ (
);

FILL FILL_2__2985_ (
);

FILL FILL_2__2565_ (
);

FILL FILL_2__2145_ (
);

FILL FILL_4__3012_ (
);

FILL FILL_5__1775_ (
);

FILL FILL_1__1767_ (
);

FILL FILL_7__2314_ (
);

FILL FILL_3__2634_ (
);

FILL FILL_3__2214_ (
);

FILL FILL_7__3519_ (
);

FILL FILL_5__3501_ (
);

FILL FILL_6__1844_ (
);

NAND2X1 _2983_ (
    .A(_1217_),
    .B(_1182_),
    .Y(_613_)
);

AOI21X1 _2563_ (
    .A(_216_),
    .B(ADD[5]),
    .C(_252_),
    .Y(_253_)
);

NAND3X1 _2143_ (
    .A(_1182_),
    .B(_1185_),
    .C(_1251_),
    .Y(_1252_)
);

FILL FILL_2__1836_ (
);

FILL FILL_4__2703_ (
);

FILL FILL_6__2629_ (
);

FILL FILL_6__2209_ (
);

DFFSR _3348_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_25_),
    .CLK(clk_bF$buf9),
    .Q(sec)
);

FILL FILL_7__3692_ (
);

FILL FILL_7__3272_ (
);

FILL FILL_0__2603_ (
);

FILL FILL_3__3592_ (
);

FILL FILL_3__3172_ (
);

FILL FILL_5__3098_ (
);

FILL FILL_3__1905_ (
);

FILL FILL_6__2382_ (
);

FILL FILL_2__2794_ (
);

FILL FILL_2__2374_ (
);

INVX1 _1834_ (
    .A(_959_),
    .Y(_960_)
);

FILL FILL_4__3661_ (
);

FILL FILL_4__3241_ (
);

FILL FILL_6__3587_ (
);

FILL FILL_6__3167_ (
);

FILL FILL_2__3579_ (
);

FILL FILL_0__3561_ (
);

FILL FILL_2__3159_ (
);

FILL FILL_0__3141_ (
);

FILL FILL_4_BUFX2_insert10 (
);

FILL FILL_4_BUFX2_insert11 (
);

FILL FILL_4_BUFX2_insert12 (
);

FILL FILL_4_BUFX2_insert13 (
);

FILL FILL_4_BUFX2_insert14 (
);

FILL FILL_4_BUFX2_insert15 (
);

FILL FILL_4_BUFX2_insert16 (
);

INVX1 _2619_ (
    .A(PC[14]),
    .Y(_300_)
);

FILL FILL_4_BUFX2_insert17 (
);

FILL FILL_1__1996_ (
);

FILL FILL_4_BUFX2_insert18 (
);

FILL FILL_4_BUFX2_insert19 (
);

FILL FILL_7__2543_ (
);

FILL FILL_3__2863_ (
);

FILL FILL_3__2443_ (
);

FILL FILL_3__2023_ (
);

FILL FILL_5__2789_ (
);

FILL FILL_5__2369_ (
);

FILL FILL_5__3310_ (
);

BUFX2 BUFX2_insert70 (
    .A(_886_),
    .Y(_886__bF$buf0)
);

BUFX2 BUFX2_insert71 (
    .A(_1149_),
    .Y(_1149__bF$buf4)
);

BUFX2 BUFX2_insert72 (
    .A(_1149_),
    .Y(_1149__bF$buf3)
);

BUFX2 BUFX2_insert73 (
    .A(_1149_),
    .Y(_1149__bF$buf2)
);

BUFX2 BUFX2_insert74 (
    .A(_1149_),
    .Y(_1149__bF$buf1)
);

FILL FILL_1__3302_ (
);

BUFX2 BUFX2_insert75 (
    .A(_1149_),
    .Y(_1149__bF$buf0)
);

BUFX2 BUFX2_insert76 (
    .A(_903_),
    .Y(_903__bF$buf3)
);

BUFX2 BUFX2_insert77 (
    .A(_903_),
    .Y(_903__bF$buf2)
);

BUFX2 BUFX2_insert78 (
    .A(_903_),
    .Y(_903__bF$buf1)
);

FILL FILL_3__3648_ (
);

BUFX2 BUFX2_insert79 (
    .A(_903_),
    .Y(_903__bF$buf0)
);

FILL FILL_3__3228_ (
);

NAND3X1 _2792_ (
    .A(_455_),
    .B(_423_),
    .C(_438_),
    .Y(_456_)
);

OAI21X1 _2372_ (
    .A(RDY_bF$buf1),
    .B(_1257_),
    .C(_1477_),
    .Y(_1478_)
);

FILL FILL_4__2932_ (
);

FILL FILL_4__2512_ (
);

FILL FILL_6__2858_ (
);

NAND2X1 _3577_ (
    .A(_1606_),
    .B(_1603_),
    .Y(_1607_)
);

FILL FILL_6__2438_ (
);

OAI21X1 _3157_ (
    .A(CO),
    .B(_728_),
    .C(_759_),
    .Y(_760_)
);

FILL FILL_6__2018_ (
);

FILL FILL_0__2832_ (
);

FILL FILL_0__2412_ (
);

FILL FILL_7__1814_ (
);

FILL FILL_0__3617_ (
);

FILL FILL_6__2191_ (
);

FILL FILL_2__2183_ (
);

FILL FILL_3__2919_ (
);

FILL FILL_4__3470_ (
);

FILL FILL_4__3050_ (
);

INVX1 _2848_ (
    .A(_506_),
    .Y(_509_)
);

NOR2X1 _2428_ (
    .A(_133_),
    .B(_1263_),
    .Y(_134_)
);

OAI21X1 _2008_ (
    .A(_1074_),
    .B(_1117_),
    .C(_1120_),
    .Y(AI[4])
);

FILL FILL_7__2772_ (
);

FILL FILL_3__2672_ (
);

FILL FILL_3__2252_ (
);

FILL FILL_5__2598_ (
);

FILL FILL_5__2178_ (
);

FILL FILL_1__3531_ (
);

FILL FILL_1__3111_ (
);

FILL FILL_3__3457_ (
);

FILL FILL_3__3037_ (
);

FILL FILL_6__1882_ (
);

NAND2X1 _2181_ (
    .A(_969_),
    .B(_952_),
    .Y(_1290_)
);

FILL FILL_2__1874_ (
);

FILL FILL_4__2741_ (
);

FILL FILL_4__2321_ (
);

FILL FILL_6__2667_ (
);

DFFPOSX1 _3386_ (
    .D(_55_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD[2])
);

FILL FILL_6__2247_ (
);

FILL FILL_2__2659_ (
);

FILL FILL_0__2641_ (
);

FILL FILL_2__2239_ (
);

FILL FILL_0__2221_ (
);

FILL FILL_2__3600_ (
);

FILL FILL_4__3526_ (
);

FILL FILL_4__3106_ (
);

FILL FILL_3__1943_ (
);

FILL FILL_0__3006_ (
);

FILL FILL_5__1869_ (
);

FILL FILL_5__2810_ (
);

FILL FILL_7__2828_ (
);

FILL FILL_7__2408_ (
);

FILL FILL_1__2802_ (
);

FILL FILL_3__2728_ (
);

FILL FILL_3__2308_ (
);

OAI21X1 _1872_ (
    .A(_935_),
    .B(_941_),
    .C(_903__bF$buf3),
    .Y(_997_)
);

FILL FILL_2__3197_ (
);

FILL FILL_6__1938_ (
);

NOR2X1 _2657_ (
    .A(_320_),
    .B(_331_),
    .Y(_332_)
);

OAI21X1 _2237_ (
    .A(_931__bF$buf1),
    .B(_984_),
    .C(_1344_),
    .Y(_1345_)
);

FILL FILL_7__2161_ (
);

FILL FILL_0__1912_ (
);

FILL FILL_3__2481_ (
);

FILL FILL_3__2061_ (
);

FILL FILL_1__2399_ (
);

FILL FILL_3__3266_ (
);

FILL FILL_4__2970_ (
);

FILL FILL_4__2550_ (
);

FILL FILL_4__2130_ (
);

FILL FILL_6__2896_ (
);

FILL FILL_6__2476_ (
);

FILL FILL_6__2056_ (
);

OAI21X1 _3195_ (
    .A(_744_),
    .B(_789_),
    .C(_792_),
    .Y(_79_)
);

FILL FILL_0__2870_ (
);

FILL FILL_2__2888_ (
);

FILL FILL_2__2468_ (
);

FILL FILL_0__2450_ (
);

FILL FILL_0__2030_ (
);

FILL FILL_2__2048_ (
);

AND2X2 _1928_ (
    .A(_1044_),
    .B(_1041_),
    .Y(_1045_)
);

FILL FILL_3__1752_ (
);

FILL FILL_0__3655_ (
);

FILL FILL_0__3235_ (
);

FILL FILL_7__2637_ (
);

FILL FILL_7__2217_ (
);

FILL FILL_1__2611_ (
);

FILL FILL_3__2957_ (
);

FILL FILL_3__2537_ (
);

FILL FILL_3__2117_ (
);

FILL FILL_4__1821_ (
);

FILL FILL_6__1747_ (
);

OAI21X1 _2886_ (
    .A(_537_),
    .B(_538_),
    .C(_536_),
    .Y(_24_)
);

OAI21X1 _2466_ (
    .A(_1319__bF$buf2),
    .B(_1263_),
    .C(PC[11]),
    .Y(_166_)
);

AOI21X1 _2046_ (
    .A(IRHOLD_valid),
    .B(_1151_),
    .C(_1154_),
    .Y(_1155_)
);

FILL FILL_7__2390_ (
);

FILL FILL_3__2290_ (
);

FILL FILL_4__2606_ (
);

FILL FILL_7__3595_ (
);

FILL FILL_7__3175_ (
);

FILL FILL_0__2926_ (
);

FILL FILL_0__2506_ (
);

FILL FILL_3__3495_ (
);

FILL FILL_3__3075_ (
);

FILL FILL_7__1908_ (
);

FILL FILL_3__1808_ (
);

FILL FILL_6__2285_ (
);

FILL FILL_2__2697_ (
);

FILL FILL_2__2277_ (
);

FILL FILL_4__3564_ (
);

FILL FILL_4__3144_ (
);

FILL FILL_3__1981_ (
);

FILL FILL_0__3464_ (
);

FILL FILL_0__3044_ (
);

FILL FILL_1__1899_ (
);

FILL FILL_7__2866_ (
);

FILL FILL_7__2446_ (
);

FILL FILL_7__2026_ (
);

FILL FILL_1__2840_ (
);

FILL FILL_1__2420_ (
);

FILL FILL_1__2000_ (
);

FILL FILL_3__2766_ (
);

FILL FILL_3__2346_ (
);

FILL FILL_5__3633_ (
);

FILL FILL_5__3213_ (
);

FILL FILL_1__3625_ (
);

FILL FILL_1__3205_ (
);

FILL FILL_6__1976_ (
);

OAI21X1 _2695_ (
    .A(_329_),
    .B(_365_),
    .C(PC[2]),
    .Y(_366_)
);

NAND2X1 _2275_ (
    .A(_1382_),
    .B(_1381_),
    .Y(_1383_)
);

FILL FILL_2__1968_ (
);

FILL FILL_0__1950_ (
);

FILL FILL_4__2835_ (
);

FILL FILL_4__2415_ (
);

FILL FILL_0__2735_ (
);

FILL FILL_6__3702_ (
);

FILL FILL_0__2315_ (
);

FILL FILL_6__2094_ (
);

FILL FILL_5__2904_ (
);

FILL FILL_2__2086_ (
);

NAND2X1 _1966_ (
    .A(ABH[0]),
    .B(_925_),
    .Y(_1083_)
);

FILL FILL_7__1890_ (
);

FILL FILL_6__3299_ (
);

FILL FILL_0__3693_ (
);

FILL FILL_3__1790_ (
);

FILL FILL_0__3273_ (
);

FILL FILL169050x61350 (
);

FILL FILL_7__2675_ (
);

FILL FILL_3__2995_ (
);

FILL FILL_3__2575_ (
);

FILL FILL_3__2155_ (
);

FILL FILL_5__3022_ (
);

FILL FILL_1__3014_ (
);

FILL FILL_6__1785_ (
);

NOR2X1 _2084_ (
    .A(_931__bF$buf1),
    .B(_928_),
    .Y(_1193_)
);

FILL FILL_5_BUFX2_insert80 (
);

FILL FILL_5_BUFX2_insert81 (
);

FILL FILL_5_BUFX2_insert82 (
);

FILL FILL_5_BUFX2_insert83 (
);

FILL FILL_2__1777_ (
);

FILL FILL_4__2644_ (
);

FILL FILL_4__2224_ (
);

NAND2X1 _3289_ (
    .A(ABL[2]),
    .B(_860_),
    .Y(_863_)
);

FILL FILL_0__2964_ (
);

FILL FILL_0__2544_ (
);

FILL FILL_6__3511_ (
);

FILL FILL_0__2124_ (
);

FILL FILL_2__3503_ (
);

FILL FILL_4__3009_ (
);

FILL FILL_1__1920_ (
);

FILL FILL_3__1846_ (
);

FILL FILL_5__2713_ (
);

FILL FILL_1__2705_ (
);

INVX2 _1775_ (
    .A(state[4]),
    .Y(_901_)
);

FILL FILL_4__3182_ (
);

FILL FILL_0__3082_ (
);

FILL FILL_4__1915_ (
);

FILL FILL_7__2064_ (
);

FILL FILL_0__1815_ (
);

AOI22X1 _3501_ (
    .A(_1716_),
    .B(BI[4]),
    .C(_1530_),
    .D(_1717_),
    .Y(_1531_)
);

FILL FILL_3__2384_ (
);

FILL FILL_5__3671_ (
);

FILL FILL_7__3269_ (
);

FILL FILL_5__3251_ (
);

FILL FILL_1__3663_ (
);

FILL FILL_1__3243_ (
);

FILL FILL_3__3589_ (
);

FILL FILL_3__3169_ (
);

FILL FILL_4__2873_ (
);

FILL FILL_4__2453_ (
);

FILL FILL_4__2033_ (
);

FILL FILL_6__2799_ (
);

FILL FILL_6__2379_ (
);

OAI21X1 _3098_ (
    .A(_895_),
    .B(_1227_),
    .C(_956_),
    .Y(_708_)
);

FILL FILL_0__2773_ (
);

FILL FILL_0__2353_ (
);

FILL FILL_2__3312_ (
);

FILL FILL_4__3658_ (
);

FILL FILL_7__1755_ (
);

FILL FILL_4__3238_ (
);

FILL FILL_0__3558_ (
);

FILL FILL_0__3138_ (
);

FILL FILL_5__2942_ (
);

FILL FILL_5__2522_ (
);

FILL FILL_5__2102_ (
);

FILL FILL_1__2934_ (
);

FILL FILL_1__2514_ (
);

FILL FILL_5__3307_ (
);

NAND2X1 _2789_ (
    .A(PC[8]),
    .B(_365_),
    .Y(_453_)
);

NAND2X1 _2369_ (
    .A(_886__bF$buf6),
    .B(_1260_),
    .Y(_1475_)
);

FILL FILL_7__2293_ (
);

NAND2X1 _3310_ (
    .A(_1741_[12]),
    .B(_869_),
    .Y(_874_)
);

FILL FILL_3__2193_ (
);

FILL FILL_4__2929_ (
);

FILL FILL_4__2509_ (
);

FILL FILL_7__3498_ (
);

FILL FILL_5__3480_ (
);

FILL FILL_7__3078_ (
);

FILL FILL_5__3060_ (
);

FILL FILL_0__2829_ (
);

FILL FILL_0__2409_ (
);

FILL FILL_1__3472_ (
);

FILL FILL_1__3052_ (
);

FILL FILL_4__2682_ (
);

FILL FILL_4__2262_ (
);

FILL FILL_6__2188_ (
);

FILL FILL_0__2582_ (
);

FILL FILL_0__2162_ (
);

FILL FILL_2__3541_ (
);

FILL FILL_2__3121_ (
);

FILL FILL_7__1984_ (
);

FILL FILL_4__3467_ (
);

FILL FILL_4__3047_ (
);

FILL FILL_3__1884_ (
);

FILL FILL_5__2751_ (
);

FILL FILL_7__2769_ (
);

FILL FILL_5__2331_ (
);

FILL FILL_1__2743_ (
);

FILL FILL_7__3710_ (
);

FILL FILL_1__2323_ (
);

FILL FILL_3__2669_ (
);

FILL FILL_3__2249_ (
);

FILL FILL_3__3610_ (
);

FILL FILL_5__3536_ (
);

FILL FILL_5__3116_ (
);

FILL FILL_1__3528_ (
);

FILL FILL_1__3108_ (
);

FILL FILL_4__1953_ (
);

FILL FILL_6__1879_ (
);

NAND2X1 _2598_ (
    .A(_282_),
    .B(_281_),
    .Y(_283_)
);

OAI21X1 _2178_ (
    .A(RDY_bF$buf5),
    .B(_998_),
    .C(_1286_),
    .Y(_1287_)
);

FILL FILL_0__1853_ (
);

FILL FILL_6__2820_ (
);

FILL FILL_6__2400_ (
);

FILL FILL_2__2812_ (
);

FILL FILL_4__2738_ (
);

FILL FILL_4__2318_ (
);

FILL FILL_0__2638_ (
);

FILL FILL_6__3605_ (
);

FILL FILL_0__2218_ (
);

FILL FILL_1__3281_ (
);

FILL FILL_4__2491_ (
);

FILL FILL_4__2071_ (
);

FILL FILL_5__2807_ (
);

FILL FILL_0__2391_ (
);

OAI21X1 _1869_ (
    .A(_993_),
    .B(_992_),
    .C(_929_),
    .Y(_994_)
);

FILL FILL_4__3696_ (
);

FILL FILL_7__1793_ (
);

FILL FILL_4__3276_ (
);

INVX1 _2810_ (
    .A(ADD[1]),
    .Y(_473_)
);

FILL FILL_0__3596_ (
);

FILL FILL_0__3176_ (
);

FILL FILL_7__2998_ (
);

FILL FILL_5__2980_ (
);

FILL FILL_5__2560_ (
);

FILL FILL_7__2158_ (
);

FILL FILL_5__2140_ (
);

FILL FILL_0__1909_ (
);

FILL FILL_1__2972_ (
);

FILL FILL_1__2552_ (
);

FILL FILL_1__2132_ (
);

FILL FILL_3__2898_ (
);

FILL FILL_3__2478_ (
);

FILL FILL_3__2058_ (
);

FILL FILL_4__1762_ (
);

FILL FILL_2__2621_ (
);

FILL FILL_2__2201_ (
);

FILL FILL_4__2967_ (
);

FILL FILL_4__2547_ (
);

FILL FILL_4__2127_ (
);

FILL FILL_0__2867_ (
);

FILL FILL_0__2447_ (
);

FILL FILL_0__2027_ (
);

FILL FILL_1__3090_ (
);

FILL FILL_5__1831_ (
);

FILL FILL_1__1823_ (
);

FILL FILL_3__1749_ (
);

FILL FILL_5__2616_ (
);

FILL FILL_1__2608_ (
);

FILL FILL_4__3085_ (
);

FILL FILL_6__1900_ (
);

FILL FILL_4__1818_ (
);

FILL FILL_7__2387_ (
);

DFFSR _3404_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_73_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[0] [4])
);

FILL FILL_1__2781_ (
);

FILL FILL_1__2361_ (
);

FILL FILL_3__2287_ (
);

FILL FILL_5__3574_ (
);

FILL FILL_5__3154_ (
);

FILL FILL_1__3566_ (
);

FILL FILL_1__3146_ (
);

FILL FILL_4__1991_ (
);

FILL FILL_0__1891_ (
);

FILL FILL_2__2850_ (
);

FILL FILL_2__2430_ (
);

FILL FILL_2__2010_ (
);

FILL FILL_4__2776_ (
);

FILL FILL_4__2356_ (
);

FILL FILL_0__2676_ (
);

FILL FILL_6__3643_ (
);

FILL FILL_0__2256_ (
);

FILL FILL_6__3223_ (
);

FILL FILL_2__3635_ (
);

FILL FILL_2__3215_ (
);

FILL FILL_3__1978_ (
);

FILL FILL_5__2845_ (
);

FILL FILL_5__2425_ (
);

FILL FILL_5__2005_ (
);

FILL FILL_1__2837_ (
);

FILL FILL_1__2417_ (
);

FILL FILL_3__3704_ (
);

FILL FILL_7__2196_ (
);

FILL FILL_0__1947_ (
);

FILL FILL_6__2914_ (
);

OAI21X1 _3633_ (
    .A(_1562_),
    .B(_1600_),
    .C(_1605_),
    .Y(_1663_)
);

NOR2X1 _3213_ (
    .A(\AXYS[2] [3]),
    .B(_798_),
    .Y(_802_)
);

FILL FILL_1__2590_ (
);

FILL FILL_1__2170_ (
);

FILL FILL_3__2096_ (
);

FILL FILL_2__2906_ (
);

FILL FILL_4__2585_ (
);

FILL FILL_4__2165_ (
);

FILL FILL_0__2485_ (
);

FILL FILL_6__3452_ (
);

FILL FILL_0__2065_ (
);

FILL FILL_6__3032_ (
);

FILL FILL_2__3024_ (
);

FILL FILL_7__1887_ (
);

NAND2X1 _2904_ (
    .A(_1181_),
    .B(_550_),
    .Y(_551_)
);

FILL FILL_1__1861_ (
);

FILL FILL_3__1787_ (
);

FILL FILL_5__2654_ (
);

FILL FILL_5__2234_ (
);

FILL FILL_1__2646_ (
);

FILL FILL_1__2226_ (
);

FILL FILL_3__3513_ (
);

FILL FILL_5__3019_ (
);

FILL FILL_2__1930_ (
);

FILL FILL_4__1856_ (
);

FILL FILL_0__1756_ (
);

FILL FILL_6__2723_ (
);

DFFSR _3442_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_110_),
    .CLK(clk_bF$buf2),
    .Q(ABH[1])
);

FILL FILL_6__2303_ (
);

NOR2X1 _3022_ (
    .A(reset),
    .B(_645_),
    .Y(_646_)
);

FILL FILL_2__2715_ (
);

FILL FILL_5__3192_ (
);

FILL FILL_6__3508_ (
);

FILL FILL_1__3184_ (
);

FILL FILL_5__1925_ (
);

FILL FILL_1__1917_ (
);

FILL FILL169050x150 (
);

FILL FILL_4__2394_ (
);

FILL FILL_0__2294_ (
);

FILL FILL_6__3261_ (
);

FILL FILL_2__3673_ (
);

FILL FILL_2__3253_ (
);

FILL FILL_4__3599_ (
);

FILL FILL_4__3179_ (
);

OAI21X1 _2713_ (
    .A(_374_),
    .B(_370_),
    .C(_382_),
    .Y(_383_)
);

FILL FILL_0__3499_ (
);

FILL FILL_0__3079_ (
);

FILL FILL_5__2883_ (
);

FILL FILL_5__2463_ (
);

FILL FILL_5__2043_ (
);

FILL FILL_1__2875_ (
);

FILL FILL_1__2455_ (
);

FILL FILL_1__2035_ (
);

FILL FILL_5__3668_ (
);

FILL FILL_5__3248_ (
);

FILL FILL_0__1985_ (
);

FILL FILL_6__2952_ (
);

NAND2X1 _3671_ (
    .A(ADD[5]),
    .B(_1714__bF$buf0),
    .Y(_1694_)
);

FILL FILL_6__2532_ (
);

FILL FILL_6__2112_ (
);

OR2X2 _3251_ (
    .A(_1257_),
    .B(_818_),
    .Y(_827_)
);

FILL FILL_2__2944_ (
);

FILL FILL_2__2524_ (
);

FILL FILL_2__2104_ (
);

FILL FILL_6__3317_ (
);

FILL FILL_0__3711_ (
);

FILL FILL_2__3309_ (
);

FILL FILL_5__2939_ (
);

FILL FILL_5__2519_ (
);

FILL FILL_6__3490_ (
);

FILL FILL_6__3070_ (
);

FILL FILL_2__3482_ (
);

FILL FILL_2__3062_ (
);

FILL FILL_0_BUFX2_insert37 (
);

FILL FILL_0_BUFX2_insert38 (
);

FILL FILL_0_BUFX2_insert39 (
);

FILL FILL_6__1803_ (
);

AOI21X1 _2942_ (
    .A(_1395_),
    .B(_1189_),
    .C(_1149__bF$buf1),
    .Y(_585_)
);

NOR2X1 _2522_ (
    .A(_216_),
    .B(_209_),
    .Y(_217_)
);

OAI21X1 _2102_ (
    .A(_1168_),
    .B(IRHOLD[3]),
    .C(_1167_),
    .Y(_1211_)
);

FILL FILL_5__2692_ (
);

FILL FILL_5__2272_ (
);

OAI21X1 _3307_ (
    .A(_1102_),
    .B(_869_),
    .C(_872_),
    .Y(_111_)
);

FILL FILL_1__2684_ (
);

FILL FILL_7__3651_ (
);

FILL FILL_1__2264_ (
);

FILL FILL_3__3551_ (
);

FILL FILL_3__3131_ (
);

FILL FILL_5__3477_ (
);

FILL FILL_5__3057_ (
);

FILL FILL_1__3469_ (
);

FILL FILL_1__3049_ (
);

FILL FILL_4__1894_ (
);

FILL FILL_0__1794_ (
);

FILL FILL_6__2761_ (
);

OAI21X1 _3480_ (
    .A(BI[7]),
    .B(alu_op[2]),
    .C(_1725_),
    .Y(_1726_)
);

FILL FILL_6__2341_ (
);

INVX1 _3060_ (
    .A(_670_),
    .Y(_674_)
);

FILL FILL_2__2753_ (
);

FILL FILL_2__2333_ (
);

FILL FILL_4__2679_ (
);

FILL FILL_4__2259_ (
);

FILL FILL_4__3620_ (
);

FILL FILL_4__3200_ (
);

FILL FILL_0__2999_ (
);

FILL FILL_0__2579_ (
);

FILL FILL_6__3546_ (
);

FILL FILL_0__2159_ (
);

FILL FILL_6__3126_ (
);

FILL FILL_0__3520_ (
);

FILL FILL_2__3538_ (
);

FILL FILL_2__3118_ (
);

FILL FILL_0__3100_ (
);

FILL FILL_5__1963_ (
);

FILL FILL_1__1955_ (
);

FILL FILL_7__2922_ (
);

FILL FILL_3__2822_ (
);

FILL FILL_3__2402_ (
);

FILL FILL169050x158550 (
);

FILL FILL_5__2748_ (
);

FILL FILL_5__2328_ (
);

FILL FILL_7__3707_ (
);

FILL FILL_2__3291_ (
);

FILL FILL_3__3607_ (
);

NOR2X1 _2751_ (
    .A(_416_),
    .B(_370_),
    .Y(_417_)
);

NOR2X1 _2331_ (
    .A(_1434_),
    .B(_1437_),
    .Y(_1438_)
);

FILL FILL_5__2081_ (
);

FILL FILL_6__2817_ (
);

NOR2X1 _3536_ (
    .A(alu_op[0]),
    .B(_1565_),
    .Y(_1566_)
);

OAI21X1 _3116_ (
    .A(ADD[0]),
    .B(_1319__bF$buf3),
    .C(_723_),
    .Y(_724_)
);

FILL FILL_1__2493_ (
);

FILL FILL_1__2073_ (
);

FILL FILL_7__3040_ (
);

FILL FILL_2__2809_ (
);

FILL FILL_5__3286_ (
);

FILL FILL_1__3698_ (
);

FILL FILL_1__3278_ (
);

FILL FILL_6__2990_ (
);

FILL FILL_6__2570_ (
);

FILL FILL_6__2150_ (
);

FILL FILL_2__2982_ (
);

FILL FILL_2__2562_ (
);

FILL FILL_2__2142_ (
);

FILL FILL_4__2488_ (
);

FILL FILL_4__2068_ (
);

FILL FILL_0__2388_ (
);

FILL FILL_5__1772_ (
);

NOR2X1 _2807_ (
    .A(_385_),
    .B(_469_),
    .Y(_470_)
);

FILL FILL_1__1764_ (
);

FILL FILL_7__2311_ (
);

FILL FILL_3__2631_ (
);

FILL FILL_3__2211_ (
);

FILL FILL_5__2977_ (
);

FILL FILL_5__2557_ (
);

FILL FILL_5__2137_ (
);

FILL FILL_1__2969_ (
);

FILL FILL_1__2549_ (
);

FILL FILL_7__3516_ (
);

FILL FILL_1__2129_ (
);

FILL FILL_6__1841_ (
);

INVX1 _2980_ (
    .A(_609_),
    .Y(_610_)
);

NAND2X1 _2560_ (
    .A(ADD[5]),
    .B(_209_),
    .Y(_250_)
);

OR2X2 _2140_ (
    .A(_1198_),
    .B(_1248_),
    .Y(_1249_)
);

FILL FILL_2__1833_ (
);

FILL FILL_4__1759_ (
);

FILL FILL_4__2700_ (
);

FILL FILL_6__2626_ (
);

DFFSR _3345_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_22_),
    .CLK(clk_bF$buf9),
    .Q(plp)
);

FILL FILL_6__2206_ (
);

FILL FILL_0__2600_ (
);

FILL FILL_2__2618_ (
);

FILL FILL_5__3095_ (
);

FILL FILL_1__3087_ (
);

FILL FILL_3__1902_ (
);

FILL FILL_5__1828_ (
);

FILL FILL_2__2791_ (
);

FILL FILL_2__2371_ (
);

FILL FILL_4__2297_ (
);

NOR2X1 _1831_ (
    .A(state[2]),
    .B(_897_),
    .Y(_957_)
);

FILL FILL_6__3584_ (
);

FILL FILL_0__2197_ (
);

FILL FILL_6__3164_ (
);

FILL FILL_2__3576_ (
);

FILL FILL_2__3156_ (
);

OAI21X1 _2616_ (
    .A(_296_),
    .B(_270_),
    .C(_297_),
    .Y(_298_)
);

FILL FILL_1__1993_ (
);

FILL FILL_7__2540_ (
);

FILL FILL_3__2860_ (
);

FILL FILL_3__2440_ (
);

FILL FILL_3__2020_ (
);

FILL FILL_5__2786_ (
);

FILL FILL_5__2366_ (
);

FILL FILL_1__2778_ (
);

FILL FILL_1__2358_ (
);

BUFX2 BUFX2_insert40 (
    .A(_720_),
    .Y(_720__bF$buf0)
);

BUFX2 BUFX2_insert41 (
    .A(_902_),
    .Y(_902__bF$buf3)
);

BUFX2 BUFX2_insert42 (
    .A(_902_),
    .Y(_902__bF$buf2)
);

BUFX2 BUFX2_insert43 (
    .A(_902_),
    .Y(_902__bF$buf1)
);

BUFX2 BUFX2_insert44 (
    .A(_902_),
    .Y(_902__bF$buf0)
);

BUFX2 BUFX2_insert45 (
    .A(_1027_),
    .Y(_1027__bF$buf4)
);

BUFX2 BUFX2_insert46 (
    .A(_1027_),
    .Y(_1027__bF$buf3)
);

BUFX2 BUFX2_insert47 (
    .A(_1027_),
    .Y(_1027__bF$buf2)
);

BUFX2 BUFX2_insert48 (
    .A(_1027_),
    .Y(_1027__bF$buf1)
);

FILL FILL_3__3645_ (
);

BUFX2 BUFX2_insert49 (
    .A(_1027_),
    .Y(_1027__bF$buf0)
);

FILL FILL_3__3225_ (
);

FILL FILL_4__1988_ (
);

FILL FILL_0__1888_ (
);

FILL FILL_6__2855_ (
);

AOI21X1 _3574_ (
    .A(_1595_),
    .B(_1599_),
    .C(_1562_),
    .Y(_1604_)
);

FILL FILL_6__2435_ (
);

FILL FILL_6__2015_ (
);

NAND2X1 _3154_ (
    .A(\AXYS[0] [4]),
    .B(_722_),
    .Y(_758_)
);

FILL FILL_2__2847_ (
);

FILL FILL_2__2427_ (
);

FILL FILL_2__2007_ (
);

FILL FILL_4__3714_ (
);

FILL FILL_7__1811_ (
);

FILL FILL_0__3614_ (
);

FILL FILL_2__2180_ (
);

FILL FILL_3__2916_ (
);

NOR2X1 _2845_ (
    .A(_505_),
    .B(_501_),
    .Y(_506_)
);

INVX1 _2425_ (
    .A(op[1]),
    .Y(_132_)
);

NAND2X1 _2005_ (
    .A(ABH[4]),
    .B(_925_),
    .Y(_1118_)
);

FILL FILL_5__2595_ (
);

FILL FILL_5__2175_ (
);

FILL FILL_1__2587_ (
);

FILL FILL_7__3554_ (
);

FILL FILL_1__2167_ (
);

FILL FILL_3__3454_ (
);

FILL FILL_3__3034_ (
);

FILL FILL_2__1871_ (
);

FILL FILL_4__1797_ (
);

FILL FILL_6__2664_ (
);

DFFSR _3383_ (
    .R(vdd),
    .S(_1__bF$buf4),
    .D(_52_),
    .CLK(clk_bF$buf2),
    .Q(res)
);

FILL FILL_6__2244_ (
);

FILL FILL_2__2656_ (
);

FILL FILL_2__2236_ (
);

FILL FILL_4__3523_ (
);

FILL FILL_4__3103_ (
);

FILL FILL_6__3449_ (
);

FILL FILL_6__3029_ (
);

FILL FILL_3__1940_ (
);

FILL FILL_0__3003_ (
);

FILL FILL_5__1866_ (
);

FILL FILL_1__1858_ (
);

FILL FILL_7__2825_ (
);

FILL FILL_3__2725_ (
);

FILL FILL_3__2305_ (
);

FILL FILL_2__3194_ (
);

FILL FILL_6__1935_ (
);

OAI21X1 _2654_ (
    .A(_1027__bF$buf4),
    .B(_1154_),
    .C(_197_),
    .Y(_329_)
);

NAND3X1 _2234_ (
    .A(_1331_),
    .B(_1333_),
    .C(_1341_),
    .Y(_1342_)
);

FILL FILL_3_CLKBUF1_insert26 (
);

FILL FILL_2__1927_ (
);

FILL FILL_3_CLKBUF1_insert27 (
);

FILL FILL_3_CLKBUF1_insert28 (
);

FILL FILL_3_CLKBUF1_insert29 (
);

DFFSR _3439_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_107_),
    .CLK(clk_bF$buf1),
    .Q(ABL[6])
);

AOI22X1 _3019_ (
    .A(_633_),
    .B(_1149__bF$buf0),
    .C(_637_),
    .D(_644_),
    .Y(_51_)
);

FILL FILL_1__2396_ (
);

FILL FILL_3__3263_ (
);

FILL FILL_5__3189_ (
);

FILL FILL_6__2893_ (
);

FILL FILL_6__2473_ (
);

OAI21X1 _3192_ (
    .A(_720__bF$buf2),
    .B(_687_),
    .C(\AXYS[1] [1]),
    .Y(_791_)
);

FILL FILL_6__2053_ (
);

FILL FILL169950x32550 (
);

FILL FILL_2__2885_ (
);

FILL FILL_2__2465_ (
);

FILL FILL_2__2045_ (
);

INVX1 _1925_ (
    .A(dst_reg[0]),
    .Y(_1042_)
);

FILL FILL_6__3678_ (
);

FILL FILL_6__3258_ (
);

FILL FILL_0__3652_ (
);

FILL FILL_0__3232_ (
);

FILL FILL_7__2214_ (
);

FILL FILL_3__2954_ (
);

FILL FILL_3__2534_ (
);

FILL FILL_3__2114_ (
);

FILL FILL_6__1744_ (
);

OAI21X1 _2883_ (
    .A(_886__bF$buf4),
    .B(_1027__bF$buf2),
    .C(clc),
    .Y(_536_)
);

OAI21X1 _2463_ (
    .A(_143_),
    .B(_1101_),
    .C(_163_),
    .Y(_1742_[2])
);

INVX1 _2043_ (
    .A(IRQ),
    .Y(_1152_)
);

FILL FILL168750x14550 (
);

FILL FILL_4__2603_ (
);

FILL FILL_6__2949_ (
);

NOR2X1 _3668_ (
    .A(_1670_),
    .B(_1669_),
    .Y(_1692_)
);

FILL FILL_6__2529_ (
);

OAI21X1 _3248_ (
    .A(_935_),
    .B(_941_),
    .C(_823_),
    .Y(_824_)
);

FILL FILL_6__2109_ (
);

FILL FILL_7__3592_ (
);

FILL FILL_7__3172_ (
);

FILL FILL_0__2923_ (
);

FILL FILL_0__2503_ (
);

FILL FILL_3__3492_ (
);

FILL FILL_3__3072_ (
);

FILL FILL_7__1905_ (
);

FILL FILL_0__3708_ (
);

FILL FILL_3__1805_ (
);

FILL FILL_6__2282_ (
);

FILL FILL_2__2694_ (
);

FILL FILL_2__2274_ (
);

FILL FILL_4__3561_ (
);

FILL FILL_4__3141_ (
);

FILL FILL_6__3487_ (
);

FILL FILL_6__3067_ (
);

FILL FILL_2__3479_ (
);

FILL FILL_0__3461_ (
);

FILL FILL_2__3059_ (
);

FILL FILL_0__3041_ (
);

OAI21X1 _2939_ (
    .A(_530_),
    .B(_581_),
    .C(_580_),
    .Y(_582_)
);

OR2X2 _2519_ (
    .A(_932_),
    .B(_213_),
    .Y(_214_)
);

FILL FILL_1__1896_ (
);

FILL FILL_7__2443_ (
);

FILL FILL_3__2763_ (
);

FILL FILL_3__2343_ (
);

FILL FILL_5__2689_ (
);

FILL FILL_5__2269_ (
);

FILL FILL_7__3648_ (
);

FILL FILL_5__3630_ (
);

FILL FILL_7__3228_ (
);

FILL FILL_5__3210_ (
);

FILL FILL_1__3622_ (
);

FILL FILL_1__3202_ (
);

FILL FILL_3__3548_ (
);

FILL FILL_3__3128_ (
);

FILL FILL_6__1973_ (
);

OAI22X1 _2692_ (
    .A(RDY_bF$buf3),
    .B(_1009_),
    .C(_363_),
    .D(_360_),
    .Y(_5_)
);

MUX2X1 _2272_ (
    .A(_1376_),
    .B(_1379_),
    .S(cond_code[1]),
    .Y(_1380_)
);

FILL FILL_2__1965_ (
);

FILL FILL_4__2832_ (
);

FILL FILL_4__2412_ (
);

FILL FILL_6__2758_ (
);

OAI21X1 _3477_ (
    .A(AI[7]),
    .B(_1719_),
    .C(_1722_),
    .Y(_1723_)
);

FILL FILL_6__2338_ (
);

NAND2X1 _3057_ (
    .A(_545_),
    .B(_670_),
    .Y(_671_)
);

FILL FILL_0__2732_ (
);

FILL FILL_0__2312_ (
);

FILL FILL_4__3617_ (
);

FILL FILL_0__3517_ (
);

FILL FILL_6__2091_ (
);

FILL FILL_7__2919_ (
);

FILL FILL_5__2901_ (
);

FILL FILL_2__2083_ (
);

FILL FILL_3__2819_ (
);

OAI21X1 _1963_ (
    .A(_914__bF$buf3),
    .B(_984_),
    .C(_1079_),
    .Y(_1080_)
);

FILL FILL_6__3296_ (
);

FILL FILL_2__3288_ (
);

FILL FILL_0__3270_ (
);

AOI21X1 _2748_ (
    .A(_322_),
    .B(ADD[5]),
    .C(_379_),
    .Y(_414_)
);

OAI21X1 _2328_ (
    .A(_902__bF$buf3),
    .B(_958_),
    .C(RDY_bF$buf8),
    .Y(_1435_)
);

FILL FILL_7__2672_ (
);

FILL FILL_3__2992_ (
);

FILL FILL_3__2572_ (
);

FILL FILL_3__2152_ (
);

FILL FILL_5__2498_ (
);

FILL FILL_5__2078_ (
);

FILL FILL_1__3011_ (
);

FILL FILL_6__1782_ (
);

NAND2X1 _2081_ (
    .A(_1189_),
    .B(_1182_),
    .Y(_1190_)
);

FILL FILL_5_BUFX2_insert50 (
);

FILL FILL_5_BUFX2_insert51 (
);

FILL FILL_5_BUFX2_insert52 (
);

FILL FILL_5_BUFX2_insert53 (
);

FILL FILL_5_BUFX2_insert54 (
);

FILL FILL_2__1774_ (
);

FILL FILL_5_BUFX2_insert55 (
);

FILL FILL_5_BUFX2_insert56 (
);

FILL FILL_5_BUFX2_insert57 (
);

FILL FILL_5_BUFX2_insert58 (
);

FILL FILL_5_BUFX2_insert59 (
);

FILL FILL_4__2641_ (
);

FILL FILL_4__2221_ (
);

FILL FILL_6__2987_ (
);

FILL FILL_6__2567_ (
);

OAI21X1 _3286_ (
    .A(_860_),
    .B(_225_),
    .C(_861_),
    .Y(_101_)
);

FILL FILL_6__2147_ (
);

FILL FILL_0__2961_ (
);

FILL FILL_2__2979_ (
);

FILL FILL_0__2541_ (
);

FILL FILL_2__2559_ (
);

FILL FILL_0__2121_ (
);

FILL FILL_2__2139_ (
);

FILL FILL_2__3500_ (
);

FILL FILL_7__1943_ (
);

FILL FILL_4__3006_ (
);

FILL FILL_3__1843_ (
);

FILL FILL_5__1769_ (
);

FILL FILL_5__2710_ (
);

FILL FILL_7__2308_ (
);

FILL FILL_1__2702_ (
);

FILL FILL_3__2628_ (
);

FILL FILL_3__2208_ (
);

NAND2X1 _1772_ (
    .A(_896_),
    .B(_897_),
    .Y(_898_)
);

FILL FILL_2__3097_ (
);

FILL FILL_4__1912_ (
);

FILL FILL_6__1838_ (
);

AOI22X1 _2977_ (
    .A(index_y),
    .B(_1149__bF$buf3),
    .C(_1332_),
    .D(_1330_),
    .Y(_608_)
);

OAI21X1 _2557_ (
    .A(_1011_),
    .B(_218_),
    .C(_247_),
    .Y(_248_)
);

NAND3X1 _2137_ (
    .A(_1232_),
    .B(_1245_),
    .C(_1240_),
    .Y(_1246_)
);

FILL FILL_7__2061_ (
);

FILL FILL_0__1812_ (
);

FILL FILL_3__2381_ (
);

FILL FILL_1__2299_ (
);

FILL FILL_1__3660_ (
);

FILL FILL_1__3240_ (
);

FILL FILL_3__3586_ (
);

FILL FILL_3__3166_ (
);

FILL FILL_4__2870_ (
);

FILL FILL_4__2450_ (
);

FILL FILL_4__2030_ (
);

FILL FILL_6__2796_ (
);

FILL FILL_6__2376_ (
);

INVX1 _3095_ (
    .A(_704_),
    .Y(_705_)
);

FILL FILL_2__2788_ (
);

FILL FILL_0__2770_ (
);

FILL FILL_2__2368_ (
);

FILL FILL_0__2350_ (
);

NAND3X1 _1828_ (
    .A(state[2]),
    .B(_897_),
    .C(_937_),
    .Y(_954_)
);

FILL FILL_4__3655_ (
);

FILL FILL_4__3235_ (
);

FILL FILL_0__3555_ (
);

FILL FILL_0__3135_ (
);

FILL FILL_5__1998_ (
);

FILL FILL_7__2957_ (
);

FILL FILL_7__2537_ (
);

FILL FILL_7__2117_ (
);

FILL FILL_1__2931_ (
);

FILL FILL_1__2511_ (
);

FILL FILL_3__2857_ (
);

FILL FILL_3__2437_ (
);

FILL FILL_3__2017_ (
);

FILL FILL_5__3304_ (
);

AOI21X1 _2786_ (
    .A(_1037_),
    .B(_449_),
    .C(_447_),
    .Y(_450_)
);

NOR2X1 _2366_ (
    .A(_1471_),
    .B(_1469_),
    .Y(_1472_)
);

FILL FILL_7__2290_ (
);

FILL FILL_3__2190_ (
);

FILL FILL_4__2926_ (
);

FILL FILL_4__2506_ (
);

FILL FILL_7__3495_ (
);

FILL FILL_7__3075_ (
);

FILL FILL_0__2826_ (
);

FILL FILL_0__2406_ (
);

FILL FILL_7__1808_ (
);

FILL FILL_6__2185_ (
);

FILL FILL_2__2597_ (
);

FILL FILL_2__2177_ (
);

FILL FILL_4__3464_ (
);

FILL FILL_4__3044_ (
);

FILL FILL_3__1881_ (
);

FILL FILL_2_CLKBUF1_insert30 (
);

FILL FILL_2_CLKBUF1_insert31 (
);

FILL FILL_2_CLKBUF1_insert32 (
);

FILL FILL_2_CLKBUF1_insert33 (
);

FILL FILL_2_CLKBUF1_insert34 (
);

FILL FILL_2_CLKBUF1_insert35 (
);

FILL FILL_2_CLKBUF1_insert36 (
);

FILL FILL_1__1799_ (
);

FILL FILL_7__2766_ (
);

FILL FILL_7__2346_ (
);

FILL FILL_1__2740_ (
);

FILL FILL_1__2320_ (
);

FILL FILL_3__2666_ (
);

FILL FILL_3__2246_ (
);

FILL FILL_5__3533_ (
);

FILL FILL_5__3113_ (
);

FILL FILL_1__3525_ (
);

FILL FILL_1__3105_ (
);

FILL FILL_4__1950_ (
);

FILL FILL_6__1876_ (
);

INVX1 _2595_ (
    .A(PC[10]),
    .Y(_280_)
);

NOR2X1 _2175_ (
    .A(_1149__bF$buf1),
    .B(_1179_),
    .Y(_1284_)
);

FILL FILL_0__1850_ (
);

FILL FILL_2__1868_ (
);

FILL FILL_4__2735_ (
);

FILL FILL_4__2315_ (
);

FILL FILL_0__2635_ (
);

FILL FILL_6__3602_ (
);

FILL FILL_0__2215_ (
);

FILL FILL_3__1937_ (
);

FILL FILL_5__2804_ (
);

NOR2X1 _1866_ (
    .A(_990_),
    .B(_988_),
    .Y(_991_)
);

FILL FILL_4__3693_ (
);

FILL FILL_7__1790_ (
);

FILL FILL_4__3273_ (
);

FILL FILL_6__3199_ (
);

FILL FILL_0__3593_ (
);

FILL FILL_0__3173_ (
);

FILL FILL_7__2995_ (
);

FILL FILL_7__2575_ (
);

FILL FILL_7__2155_ (
);

FILL FILL_0__1906_ (
);

FILL FILL_3__2895_ (
);

FILL FILL_3__2475_ (
);

FILL FILL_3__2055_ (
);

FILL FILL_4__2964_ (
);

FILL FILL_4__2544_ (
);

FILL FILL_4__2124_ (
);

NAND2X1 _3189_ (
    .A(_721_),
    .B(_1047_),
    .Y(_789_)
);

FILL FILL_0__2864_ (
);

FILL FILL_0__2444_ (
);

FILL FILL_0__2024_ (
);

FILL FILL_1__1820_ (
);

FILL FILL_3__1746_ (
);

FILL FILL_0__3649_ (
);

FILL FILL_0__3229_ (
);

FILL FILL_5__2613_ (
);

FILL FILL_1__2605_ (
);

FILL FILL_4__3082_ (
);

FILL FILL_4__1815_ (
);

DFFSR _3401_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_70_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[0] [1])
);

FILL FILL_3__2284_ (
);

FILL FILL_5__3571_ (
);

FILL FILL_7__3169_ (
);

FILL FILL_5__3151_ (
);

FILL FILL_1__3563_ (
);

FILL FILL_1__3143_ (
);

FILL FILL_3__3489_ (
);

FILL FILL_3__3069_ (
);

FILL FILL_4__2773_ (
);

FILL FILL_4__2353_ (
);

FILL FILL_6__2699_ (
);

FILL FILL_6__2279_ (
);

FILL FILL_0__2673_ (
);

FILL FILL_6__3640_ (
);

FILL FILL_0__2253_ (
);

FILL FILL_6__3220_ (
);

FILL FILL_2__3632_ (
);

FILL FILL_2__3212_ (
);

FILL FILL_4__3558_ (
);

FILL FILL_4__3138_ (
);

FILL FILL_3__1975_ (
);

FILL FILL_0__3458_ (
);

FILL FILL_0__3038_ (
);

FILL FILL169050x14550 (
);

FILL FILL_5__2842_ (
);

FILL FILL_5__2422_ (
);

FILL FILL_5__2002_ (
);

FILL FILL_1__2834_ (
);

FILL FILL_1__2414_ (
);

FILL FILL_3__3701_ (
);

FILL FILL_5__3627_ (
);

FILL FILL_5__3207_ (
);

FILL FILL_1__3619_ (
);

AOI21X1 _2689_ (
    .A(_352_),
    .B(_353_),
    .C(_1007_),
    .Y(_361_)
);

INVX1 _2269_ (
    .A(N),
    .Y(_1377_)
);

FILL FILL_7__2193_ (
);

FILL FILL_0__1944_ (
);

FILL FILL_6__2911_ (
);

OAI21X1 _3630_ (
    .A(_1653_),
    .B(_1636_),
    .C(_1648_),
    .Y(_1660_)
);

AOI21X1 _3210_ (
    .A(_737_),
    .B(_798_),
    .C(_800_),
    .Y(_86_)
);

FILL FILL_3__2093_ (
);

FILL FILL_2__2903_ (
);

FILL FILL_4__2829_ (
);

FILL FILL_4__2409_ (
);

FILL FILL_0__2729_ (
);

FILL FILL_0__2309_ (
);

FILL FILL_3__3298_ (
);

FILL FILL_4__2582_ (
);

FILL FILL_4__2162_ (
);

FILL FILL_6__2088_ (
);

FILL FILL_0__2482_ (
);

FILL FILL_0__2062_ (
);

FILL FILL_2__3021_ (
);

FILL FILL_7__1884_ (
);

OAI22X1 _2901_ (
    .A(_548_),
    .B(_1150__bF$buf2),
    .C(_541_),
    .D(_547_),
    .Y(_29_)
);

FILL FILL_3__1784_ (
);

FILL FILL_0__3267_ (
);

FILL FILL_7__2669_ (
);

FILL FILL_5__2651_ (
);

FILL FILL_5__2231_ (
);

FILL FILL_1__2643_ (
);

FILL FILL_1__2223_ (
);

FILL FILL_3__2989_ (
);

FILL FILL_3__2569_ (
);

FILL FILL_3__2149_ (
);

FILL FILL_3__3510_ (
);

FILL FILL_5__3016_ (
);

FILL FILL_1__3008_ (
);

FILL FILL_4__1853_ (
);

FILL FILL_6__1779_ (
);

OAI21X1 _2498_ (
    .A(_902__bF$buf0),
    .B(_946_),
    .C(_1067_),
    .Y(_193_)
);

NOR2X1 _2078_ (
    .A(_1154_),
    .B(_1186_),
    .Y(_1187_)
);

FILL FILL_0__1753_ (
);

FILL FILL_6__2720_ (
);

FILL FILL_6__2300_ (
);

FILL FILL_2__2712_ (
);

FILL FILL_4__2638_ (
);

FILL FILL_4__2218_ (
);

FILL FILL_0__2958_ (
);

FILL FILL_0__2538_ (
);

FILL FILL_6__3505_ (
);

FILL FILL_0__2118_ (
);

FILL FILL_1__3181_ (
);

FILL FILL_5__1922_ (
);

FILL FILL_1__1914_ (
);

FILL FILL_4__2391_ (
);

FILL FILL_5__2707_ (
);

FILL FILL_0__2291_ (
);

FILL FILL_2__3670_ (
);

FILL FILL_2__3250_ (
);

INVX1 _1769_ (
    .A(shift),
    .Y(_895_)
);

FILL FILL_4__3596_ (
);

FILL FILL_4__3176_ (
);

INVX1 _2710_ (
    .A(_379_),
    .Y(_380_)
);

FILL FILL_0__3496_ (
);

FILL FILL_0__3076_ (
);

FILL FILL_4__1909_ (
);

FILL FILL_5__2880_ (
);

FILL FILL_7__2898_ (
);

FILL FILL_5__2460_ (
);

FILL FILL_7__2058_ (
);

FILL FILL_5__2040_ (
);

FILL FILL_0__1809_ (
);

FILL FILL_1__2872_ (
);

FILL FILL_1__2452_ (
);

FILL FILL_1__2032_ (
);

FILL FILL_3__2798_ (
);

FILL FILL_3__2378_ (
);

FILL FILL_5__3665_ (
);

FILL FILL_5__3245_ (
);

FILL FILL_1__3657_ (
);

FILL FILL_1__3237_ (
);

FILL FILL_0__1982_ (
);

FILL FILL_2__2941_ (
);

FILL FILL_2__2521_ (
);

FILL FILL_2__2101_ (
);

FILL FILL_4__2867_ (
);

FILL FILL_4__2447_ (
);

FILL FILL_4__2027_ (
);

FILL FILL_0__2767_ (
);

FILL FILL_0__2347_ (
);

FILL FILL_6__3314_ (
);

FILL FILL_2__3306_ (
);

FILL FILL_5__2936_ (
);

FILL FILL_5__2516_ (
);

FILL FILL169350x57750 (
);

FILL FILL_1__2928_ (
);

FILL FILL_1__2508_ (
);

AOI21X1 _1998_ (
    .A(_1082_),
    .B(ADD[3]),
    .C(_1111_),
    .Y(_1112_)
);

FILL FILL_6__1800_ (
);

FILL FILL_7__2287_ (
);

NAND2X1 _3304_ (
    .A(_1741_[9]),
    .B(_869_),
    .Y(_871_)
);

FILL FILL_1__2681_ (
);

FILL FILL_1__2261_ (
);

FILL FILL_3__2187_ (
);

FILL FILL_5__3474_ (
);

FILL FILL_5__3054_ (
);

FILL FILL_1__3466_ (
);

FILL FILL_1__3046_ (
);

FILL FILL_4__1891_ (
);

FILL FILL_0__1791_ (
);

FILL FILL_2__2750_ (
);

FILL FILL_2__2330_ (
);

FILL FILL168150x39750 (
);

FILL FILL_4__2676_ (
);

FILL FILL_4__2256_ (
);

FILL FILL_0__2996_ (
);

FILL FILL_0__2576_ (
);

FILL FILL_6__3543_ (
);

FILL FILL_0__2156_ (
);

FILL FILL_6__3123_ (
);

FILL FILL_2__3535_ (
);

FILL FILL_2__3115_ (
);

FILL FILL_5__1960_ (
);

FILL FILL_1__1952_ (
);

FILL FILL_3__1878_ (
);

FILL FILL_5__2745_ (
);

FILL FILL_5__2325_ (
);

FILL FILL_1__2737_ (
);

FILL FILL_1__2317_ (
);

FILL FILL_3__3604_ (
);

FILL FILL_4__1947_ (
);

FILL FILL_7__2096_ (
);

FILL FILL_0__1847_ (
);

FILL FILL_6__2814_ (
);

NAND3X1 _3533_ (
    .A(BI[1]),
    .B(AI[1]),
    .C(_1718_),
    .Y(_1563_)
);

INVX1 _3113_ (
    .A(_720__bF$buf2),
    .Y(_721_)
);

FILL FILL_1__2490_ (
);

FILL FILL_1__2070_ (
);

FILL FILL_2__2806_ (
);

FILL FILL_5__3283_ (
);

FILL FILL_1__3695_ (
);

FILL FILL_1__3275_ (
);

FILL FILL_4__2485_ (
);

FILL FILL_4__2065_ (
);

FILL FILL_0__2385_ (
);

FILL FILL_7__1787_ (
);

NAND2X1 _2804_ (
    .A(_465_),
    .B(_466_),
    .Y(_467_)
);

FILL FILL_1__1761_ (
);

FILL FILL_5__2974_ (
);

FILL FILL_5__2554_ (
);

FILL FILL_5__2134_ (
);

FILL FILL_1__2966_ (
);

FILL FILL_1__2546_ (
);

FILL FILL_7__3513_ (
);

FILL FILL_1__2126_ (
);

FILL FILL_2__1830_ (
);

FILL FILL_4__1756_ (
);

FILL FILL_6__2623_ (
);

DFFSR _3342_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_19_),
    .CLK(clk_bF$buf10),
    .Q(cond_code[0])
);

FILL FILL_6__2203_ (
);

FILL FILL_2__2615_ (
);

FILL FILL_5__3092_ (
);

FILL FILL_1__3084_ (
);

FILL FILL_5__1825_ (
);

FILL FILL_1__1817_ (
);

FILL FILL_4__2294_ (
);

FILL FILL_6__3581_ (
);

FILL FILL_0__2194_ (
);

FILL FILL_6__3161_ (
);

FILL FILL_2__3573_ (
);

FILL FILL_2__3153_ (
);

FILL FILL_4__3499_ (
);

FILL FILL_4__3079_ (
);

INVX1 _2613_ (
    .A(PC[13]),
    .Y(_295_)
);

FILL FILL_1__1990_ (
);

FILL FILL_5__2783_ (
);

FILL FILL_5__2363_ (
);

FILL FILL_1__2775_ (
);

FILL FILL_1__2355_ (
);

BUFX2 BUFX2_insert10 (
    .A(_1_),
    .Y(_1__bF$buf10)
);

BUFX2 BUFX2_insert11 (
    .A(_1_),
    .Y(_1__bF$buf9)
);

BUFX2 BUFX2_insert12 (
    .A(_1_),
    .Y(_1__bF$buf8)
);

BUFX2 BUFX2_insert13 (
    .A(_1_),
    .Y(_1__bF$buf7)
);

BUFX2 BUFX2_insert14 (
    .A(_1_),
    .Y(_1__bF$buf6)
);

BUFX2 BUFX2_insert15 (
    .A(_1_),
    .Y(_1__bF$buf5)
);

BUFX2 BUFX2_insert16 (
    .A(_1_),
    .Y(_1__bF$buf4)
);

BUFX2 BUFX2_insert17 (
    .A(_1_),
    .Y(_1__bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .A(_1_),
    .Y(_1__bF$buf2)
);

FILL FILL_3__3642_ (
);

BUFX2 BUFX2_insert19 (
    .A(_1_),
    .Y(_1__bF$buf1)
);

FILL FILL_3__3222_ (
);

FILL FILL169650x10950 (
);

FILL FILL_5__3568_ (
);

FILL FILL_5__3148_ (
);

FILL FILL_4__1985_ (
);

FILL FILL_0__1885_ (
);

FILL FILL_6__2852_ (
);

NAND2X1 _3571_ (
    .A(_1548_),
    .B(_1545_),
    .Y(_1601_)
);

FILL FILL_6__2432_ (
);

FILL FILL_6__2012_ (
);

OAI21X1 _3151_ (
    .A(_722_),
    .B(_754_),
    .C(_755_),
    .Y(_72_)
);

FILL FILL_2__2844_ (
);

FILL FILL_2__2424_ (
);

FILL FILL_2__2004_ (
);

FILL FILL_4__3711_ (
);

FILL FILL_6__3637_ (
);

FILL FILL_6__3217_ (
);

FILL FILL_0__3611_ (
);

FILL FILL_2__3629_ (
);

FILL FILL_2__3209_ (
);

FILL FILL_3__2913_ (
);

FILL FILL_5__2839_ (
);

FILL FILL_5__2419_ (
);

AOI22X1 _2842_ (
    .A(ADD[6]),
    .B(_1299_),
    .C(_323_),
    .D(ABH[6]),
    .Y(_503_)
);

INVX1 _2422_ (
    .A(_1275_),
    .Y(_130_)
);

NAND3X1 _2002_ (
    .A(\AXYS[0] [4]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1115_)
);

FILL FILL_5__2592_ (
);

FILL FILL_5__2172_ (
);

FILL FILL_6__2908_ (
);

NOR2X1 _3627_ (
    .A(_1722_),
    .B(_1576_),
    .Y(_1657_)
);

NOR2X1 _3207_ (
    .A(\AXYS[2] [0]),
    .B(_798_),
    .Y(_799_)
);

FILL FILL_1__2584_ (
);

FILL FILL_7__3551_ (
);

FILL FILL_1__2164_ (
);

FILL FILL169350x158550 (
);

FILL FILL_3__3451_ (
);

FILL FILL_3__3031_ (
);

FILL FILL_4__1794_ (
);

FILL FILL_6__2661_ (
);

DFFSR _3380_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(DIMUX[5]),
    .CLK(clk_bF$buf2),
    .Q(DIHOLD[5])
);

FILL FILL_6__2241_ (
);

FILL FILL_2__2653_ (
);

FILL FILL_2__2233_ (
);

FILL FILL_4__2999_ (
);

FILL FILL_4__2579_ (
);

FILL FILL_4__2159_ (
);

FILL FILL_4__3520_ (
);

FILL FILL_4__3100_ (
);

FILL FILL_0__2899_ (
);

FILL FILL_0__2479_ (
);

FILL FILL_0__2059_ (
);

FILL FILL_6__3026_ (
);

FILL FILL_2__3018_ (
);

FILL FILL_0__3000_ (
);

FILL FILL_5__1863_ (
);

FILL FILL_1__1855_ (
);

FILL FILL_7__2822_ (
);

FILL FILL_3__2722_ (
);

FILL FILL_3__2302_ (
);

FILL FILL_5__2648_ (
);

FILL FILL_5__2228_ (
);

FILL FILL_2__3191_ (
);

FILL FILL_3__3507_ (
);

FILL FILL_6__1932_ (
);

NOR3X1 _2651_ (
    .A(_925_),
    .B(_1291_),
    .C(_325_),
    .Y(_326_)
);

OAI21X1 _2231_ (
    .A(RDY_bF$buf2),
    .B(_1337_),
    .C(_1338_),
    .Y(_1339_)
);

FILL FILL_2__1924_ (
);

FILL FILL_6__2717_ (
);

DFFSR _3436_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_104_),
    .CLK(clk_bF$buf1),
    .Q(ABL[3])
);

OAI21X1 _3016_ (
    .A(_1181_),
    .B(_1185_),
    .C(_1405_),
    .Y(_642_)
);

FILL FILL_1__2393_ (
);

FILL FILL_2__2709_ (
);

FILL FILL_3__3260_ (
);

FILL FILL_1_BUFX2_insert70 (
);

FILL FILL_1_BUFX2_insert71 (
);

FILL FILL_1_BUFX2_insert72 (
);

FILL FILL_1_BUFX2_insert73 (
);

FILL FILL_5__3186_ (
);

FILL FILL_1_BUFX2_insert74 (
);

FILL FILL_1_BUFX2_insert75 (
);

FILL FILL_1_BUFX2_insert76 (
);

FILL FILL_1_BUFX2_insert77 (
);

FILL FILL_1_BUFX2_insert78 (
);

FILL FILL_1_BUFX2_insert79 (
);

FILL FILL_1__3598_ (
);

FILL FILL_1__3178_ (
);

FILL FILL_5__1919_ (
);

FILL FILL_6__2890_ (
);

FILL FILL_6__2470_ (
);

FILL FILL_6__2050_ (
);

FILL FILL_2__2882_ (
);

FILL FILL_2__2462_ (
);

FILL FILL_2__2042_ (
);

FILL FILL_4__2388_ (
);

AOI21X1 _1922_ (
    .A(dst_reg[1]),
    .B(_1037_),
    .C(_1038_),
    .Y(_1039_)
);

FILL FILL_6__3675_ (
);

FILL FILL_0__2288_ (
);

FILL FILL_6__3255_ (
);

FILL FILL_2__3667_ (
);

FILL FILL_2__3247_ (
);

AOI21X1 _2707_ (
    .A(_352_),
    .B(_353_),
    .C(_1012_),
    .Y(_377_)
);

FILL FILL_7__2211_ (
);

FILL FILL_3__2951_ (
);

FILL FILL_3__2531_ (
);

FILL FILL_3__2111_ (
);

FILL FILL_5__2877_ (
);

FILL FILL_5__2457_ (
);

FILL FILL_5__2037_ (
);

FILL FILL_1__2869_ (
);

FILL FILL_1__2449_ (
);

FILL FILL_1__2029_ (
);

FILL FILL_3__3316_ (
);

NOR2X1 _2880_ (
    .A(_1187_),
    .B(_1181_),
    .Y(_534_)
);

AOI22X1 _2460_ (
    .A(PC[2]),
    .B(_1080_),
    .C(_149_),
    .D(I),
    .Y(_161_)
);

NAND2X1 _2040_ (
    .A(RDY_bF$buf2),
    .B(_1037_),
    .Y(_1149_)
);

FILL FILL_4__2600_ (
);

FILL FILL_0__1979_ (
);

FILL FILL_6__2946_ (
);

NAND2X1 _3665_ (
    .A(ADD[3]),
    .B(_1714__bF$buf3),
    .Y(_1690_)
);

FILL FILL_6__2526_ (
);

AOI21X1 _3245_ (
    .A(_901_),
    .B(_993_),
    .C(_820_),
    .Y(_821_)
);

FILL FILL_6__2106_ (
);

FILL FILL_0__2920_ (
);

FILL FILL_2__2938_ (
);

FILL FILL_0__2500_ (
);

FILL FILL_2__2518_ (
);

FILL FILL_0__3705_ (
);

FILL FILL_3__1802_ (
);

FILL FILL169050x144150 (
);

FILL FILL_2__2691_ (
);

FILL FILL_2__2271_ (
);

FILL FILL_4__2197_ (
);

FILL FILL_6__3484_ (
);

FILL FILL_0__2097_ (
);

FILL FILL_6__3064_ (
);

FILL FILL_2__3476_ (
);

FILL FILL_2__3056_ (
);

NAND2X1 _2936_ (
    .A(_543_),
    .B(_1182_),
    .Y(_579_)
);

INVX1 _2516_ (
    .A(_1291_),
    .Y(_211_)
);

FILL FILL_1__1893_ (
);

FILL FILL_7__2440_ (
);

FILL FILL_3__2760_ (
);

FILL FILL_3__2340_ (
);

FILL FILL_5__2686_ (
);

FILL FILL_5__2266_ (
);

FILL FILL_1__2678_ (
);

FILL FILL_7__3645_ (
);

FILL FILL_1__2258_ (
);

FILL FILL_7__3225_ (
);

FILL FILL_3__3545_ (
);

FILL FILL_3__3125_ (
);

FILL FILL_6__1970_ (
);

FILL FILL_2__1962_ (
);

FILL FILL_4__1888_ (
);

FILL FILL_0__1788_ (
);

FILL FILL_6__2755_ (
);

NAND2X1 _3474_ (
    .A(AI[7]),
    .B(_1719_),
    .Y(_1720_)
);

FILL FILL_6__2335_ (
);

OAI21X1 _3054_ (
    .A(_667_),
    .B(_668_),
    .C(_664_),
    .Y(_669_)
);

FILL FILL_2__2747_ (
);

FILL FILL_2__2327_ (
);

FILL FILL_4__3614_ (
);

FILL FILL_0__3514_ (
);

FILL FILL_5__1957_ (
);

FILL FILL_1__1949_ (
);

FILL FILL_7__2916_ (
);

FILL FILL_2__2080_ (
);

FILL FILL_3__2816_ (
);

INVX1 _1960_ (
    .A(_1076_),
    .Y(_1077_)
);

FILL FILL_6__3293_ (
);

FILL FILL_2__3285_ (
);

OAI21X1 _2745_ (
    .A(_410_),
    .B(_401_),
    .C(RDY_bF$buf0),
    .Y(_412_)
);

NAND2X1 _2325_ (
    .A(_1297_),
    .B(_925_),
    .Y(_1432_)
);

FILL FILL_5__2495_ (
);

FILL FILL_5__2075_ (
);

FILL FILL_1__2487_ (
);

FILL FILL_7__3454_ (
);

FILL FILL_1__2067_ (
);

FILL FILL_5_BUFX2_insert20 (
);

FILL FILL_5_BUFX2_insert21 (
);

FILL FILL_5_BUFX2_insert22 (
);

FILL FILL_5_BUFX2_insert23 (
);

FILL FILL_5_BUFX2_insert24 (
);

FILL FILL_5_BUFX2_insert25 (
);

FILL FILL_2__1771_ (
);

FILL FILL_6__2984_ (
);

FILL FILL_6__2564_ (
);

NAND2X1 _3283_ (
    .A(_858_),
    .B(_855_),
    .Y(_859_)
);

FILL FILL_6__2144_ (
);

FILL FILL_2__2976_ (
);

FILL FILL_2__2556_ (
);

FILL FILL_2__2136_ (
);

FILL FILL_7__1940_ (
);

FILL FILL_4__3003_ (
);

FILL FILL_3__1840_ (
);

FILL FILL_5__1766_ (
);

FILL FILL_1__1758_ (
);

FILL FILL_7__2725_ (
);

FILL FILL_3__2625_ (
);

FILL FILL_3__2205_ (
);

FILL FILL_2__3094_ (
);

FILL FILL_6__1835_ (
);

INVX1 _2974_ (
    .A(_550_),
    .Y(_605_)
);

OAI22X1 _2554_ (
    .A(_888_),
    .B(_201_),
    .C(_244_),
    .D(_199_),
    .Y(_245_)
);

NOR2X1 _2134_ (
    .A(_886__bF$buf6),
    .B(_930_),
    .Y(_1243_)
);

FILL FILL_2__1827_ (
);

DFFSR _3339_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_17_),
    .CLK(clk_bF$buf2),
    .Q(PC[15])
);

FILL FILL_1__2296_ (
);

FILL FILL_3__3583_ (
);

FILL FILL_3__3163_ (
);

FILL FILL_5__3089_ (
);

FILL FILL_6__2793_ (
);

FILL FILL_6__2373_ (
);

NOR2X1 _3092_ (
    .A(write_back),
    .B(_1027__bF$buf1),
    .Y(_702_)
);

FILL FILL_2__2785_ (
);

FILL FILL_2__2365_ (
);

NOR2X1 _1825_ (
    .A(_950_),
    .B(_947_),
    .Y(_951_)
);

FILL FILL_4__3652_ (
);

FILL FILL_4__3232_ (
);

FILL FILL_6__3578_ (
);

FILL FILL_6__3158_ (
);

FILL FILL_0__3552_ (
);

FILL FILL_0__3132_ (
);

FILL FILL_5__1995_ (
);

FILL FILL_1__1987_ (
);

FILL FILL_7__2954_ (
);

FILL FILL_7__2114_ (
);

FILL FILL_3__2854_ (
);

FILL FILL_3__2434_ (
);

FILL FILL_3__2014_ (
);

FILL FILL_5__3301_ (
);

FILL FILL_1__3713_ (
);

FILL FILL_3__3639_ (
);

FILL FILL_3__3219_ (
);

NAND3X1 _2783_ (
    .A(_1110_),
    .B(_445_),
    .C(_446_),
    .Y(_447_)
);

OAI21X1 _2363_ (
    .A(RDY_bF$buf6),
    .B(_1467_),
    .C(_1468_),
    .Y(_1469_)
);

FILL FILL_4__2923_ (
);

FILL FILL_4__2503_ (
);

FILL FILL_6__2849_ (
);

OAI21X1 _3568_ (
    .A(_1557_),
    .B(_1597_),
    .C(_1561_),
    .Y(_1598_)
);

FILL FILL_6__2429_ (
);

FILL FILL_6__2009_ (
);

NOR2X1 _3148_ (
    .A(_752_),
    .B(_751_),
    .Y(_753_)
);

FILL FILL_7__3492_ (
);

FILL FILL_7__3072_ (
);

FILL FILL_0__2823_ (
);

FILL FILL_0__2403_ (
);

FILL FILL_4__3708_ (
);

FILL FILL_7__1805_ (
);

FILL FILL_0__3608_ (
);

FILL FILL_6__2182_ (
);

FILL FILL_2__2594_ (
);

FILL FILL_2__2174_ (
);

FILL FILL_4__3461_ (
);

FILL FILL_4__3041_ (
);

FILL FILL_6_BUFX2_insert70 (
);

FILL FILL_6_BUFX2_insert71 (
);

FILL FILL_6_BUFX2_insert72 (
);

FILL FILL_6_BUFX2_insert73 (
);

FILL FILL_6_BUFX2_insert74 (
);

FILL FILL_6_BUFX2_insert75 (
);

FILL FILL_6_BUFX2_insert76 (
);

FILL FILL_6_BUFX2_insert77 (
);

FILL FILL_6_BUFX2_insert78 (
);

FILL FILL_6_BUFX2_insert79 (
);

NOR2X1 _2839_ (
    .A(_465_),
    .B(_495_),
    .Y(_500_)
);

NAND3X1 _2419_ (
    .A(_1507_),
    .B(_127_),
    .C(_118_),
    .Y(_1512_[5])
);

FILL FILL_1__1796_ (
);

FILL FILL_7__2343_ (
);

FILL FILL_3__2663_ (
);

FILL FILL_3__2243_ (
);

FILL FILL_5__2589_ (
);

FILL FILL_5__2169_ (
);

FILL FILL_5__3530_ (
);

FILL FILL_7__3548_ (
);

FILL FILL_7__3128_ (
);

FILL FILL_5__3110_ (
);

FILL FILL_1__3522_ (
);

FILL FILL_1__3102_ (
);

FILL FILL_3__3028_ (
);

FILL FILL_6__1873_ (
);

OAI21X1 _2592_ (
    .A(_1091_),
    .B(_270_),
    .C(_277_),
    .Y(_278_)
);

OAI21X1 _2172_ (
    .A(_1207_),
    .B(_1206_),
    .C(RDY_bF$buf8),
    .Y(_1281_)
);

FILL FILL_2__1865_ (
);

FILL FILL_4__2732_ (
);

FILL FILL_4__2312_ (
);

FILL FILL_6__2658_ (
);

DFFSR _3377_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(DIMUX[2]),
    .CLK(clk_bF$buf5),
    .Q(DIHOLD[2])
);

FILL FILL_6__2238_ (
);

FILL FILL_0__2632_ (
);

FILL FILL_0__2212_ (
);

FILL FILL_4__3517_ (
);

FILL FILL_3__1934_ (
);

FILL FILL_7__2819_ (
);

FILL FILL_5__2801_ (
);

FILL FILL_3__2719_ (
);

NOR2X1 _1863_ (
    .A(_902__bF$buf2),
    .B(_928_),
    .Y(_988_)
);

FILL FILL_4__3270_ (
);

FILL FILL_6__3196_ (
);

FILL FILL_0__3590_ (
);

FILL FILL_0__3170_ (
);

FILL FILL_2__3188_ (
);

FILL FILL_6__1929_ (
);

NOR2X1 _2648_ (
    .A(_1027__bF$buf4),
    .B(_1167_),
    .Y(_323_)
);

OAI21X1 _2228_ (
    .A(RDY_bF$buf6),
    .B(_1334_),
    .C(_1335_),
    .Y(_1336_)
);

FILL FILL_7__2572_ (
);

FILL FILL_0__1903_ (
);

FILL FILL_3__2892_ (
);

FILL FILL_3__2472_ (
);

FILL FILL_3__2052_ (
);

FILL FILL_5__2398_ (
);

FILL FILL_3__3677_ (
);

FILL FILL_3__3257_ (
);

FILL FILL_4__2961_ (
);

FILL FILL_4__2541_ (
);

FILL FILL_4__2121_ (
);

FILL FILL_6__2887_ (
);

FILL FILL_6__2467_ (
);

AOI21X1 _3186_ (
    .A(DIMUX[7]),
    .B(_1319__bF$buf1),
    .C(_786_),
    .Y(_787_)
);

FILL FILL_6__2047_ (
);

FILL FILL_0__2861_ (
);

FILL FILL_2__2879_ (
);

FILL FILL_2__2459_ (
);

FILL FILL_0__2441_ (
);

FILL FILL_2__2039_ (
);

FILL FILL_0__2021_ (
);

NAND2X1 _1919_ (
    .A(_1035_),
    .B(_1026_),
    .Y(_1036_)
);

FILL FILL_7__1843_ (
);

FILL FILL_0__3646_ (
);

FILL FILL_0__3226_ (
);

FILL FILL_5__2610_ (
);

FILL FILL_7__2208_ (
);

FILL FILL_1__2602_ (
);

FILL FILL_3__2948_ (
);

FILL FILL_3__2528_ (
);

FILL FILL_3__2108_ (
);

FILL FILL_4__1812_ (
);

NAND2X1 _2877_ (
    .A(_1367_),
    .B(_531_),
    .Y(_532_)
);

OAI21X1 _2457_ (
    .A(_143_),
    .B(_1090_),
    .C(_158_),
    .Y(_1742_[1])
);

OAI21X1 _2037_ (
    .A(_893_),
    .B(_983_),
    .C(_1146_),
    .Y(_1147_)
);

FILL FILL_3__2281_ (
);

FILL FILL_1__2199_ (
);

FILL FILL_0__2917_ (
);

FILL FILL_1__3560_ (
);

FILL FILL_1__3140_ (
);

FILL FILL_3__3486_ (
);

FILL FILL_3__3066_ (
);

FILL FILL_4__2770_ (
);

FILL FILL_4__2350_ (
);

FILL FILL_6__2696_ (
);

FILL FILL_6__2276_ (
);

FILL FILL_2__2688_ (
);

FILL FILL_0__2670_ (
);

FILL FILL_2__2268_ (
);

FILL FILL_0__2250_ (
);

FILL FILL_4__3555_ (
);

FILL FILL_4__3135_ (
);

FILL FILL_3__1972_ (
);

FILL FILL_0__3455_ (
);

FILL FILL_0__3035_ (
);

FILL FILL_5__1898_ (
);

FILL FILL_7__2857_ (
);

FILL FILL_7__2437_ (
);

FILL FILL_7__2017_ (
);

FILL FILL_1__2831_ (
);

FILL FILL_1__2411_ (
);

FILL FILL_3__2757_ (
);

FILL FILL_3__2337_ (
);

FILL FILL_5__3624_ (
);

FILL FILL_5__3204_ (
);

FILL FILL_1__3616_ (
);

FILL FILL_6__1967_ (
);

NOR2X1 _2686_ (
    .A(_357_),
    .B(_354_),
    .Y(_358_)
);

INVX1 _2266_ (
    .A(V),
    .Y(_1374_)
);

FILL FILL_7__2190_ (
);

FILL FILL_0__1941_ (
);

FILL FILL_2__1959_ (
);

FILL FILL_3__2090_ (
);

FILL FILL_2__2900_ (
);

FILL FILL_4__2826_ (
);

FILL FILL_4__2406_ (
);

FILL FILL_0__2726_ (
);

FILL FILL_0__2306_ (
);

FILL FILL_3__3295_ (
);

FILL FILL_6__2085_ (
);

FILL FILL_2__2497_ (
);

FILL FILL_2__2077_ (
);

INVX2 _1957_ (
    .A(_1073_),
    .Y(_1074_)
);

FILL FILL_3__1781_ (
);

FILL FILL_0__3264_ (
);

FILL FILL_7__2666_ (
);

FILL FILL_7__2246_ (
);

FILL FILL_1__2640_ (
);

FILL FILL_1__2220_ (
);

FILL FILL_3__2986_ (
);

FILL FILL_3__2566_ (
);

FILL FILL_3__2146_ (
);

FILL FILL_5__3013_ (
);

FILL FILL_1__3005_ (
);

FILL FILL_4__1850_ (
);

FILL FILL_6__1776_ (
);

OAI21X1 _2495_ (
    .A(_1377_),
    .B(_165_),
    .C(_190_),
    .Y(_191_)
);

OAI21X1 _2075_ (
    .A(IRHOLD_valid),
    .B(_893_),
    .C(_1183_),
    .Y(_1184_)
);

FILL FILL_0__1750_ (
);

FILL FILL_2__1768_ (
);

FILL FILL_4__2635_ (
);

FILL FILL_4__2215_ (
);

FILL FILL_0__2955_ (
);

FILL FILL_0__2535_ (
);

FILL FILL_6__3502_ (
);

FILL FILL_0__2115_ (
);

FILL FILL_7__1937_ (
);

FILL FILL_1__1911_ (
);

FILL FILL_3__1837_ (
);

FILL FILL_5__2704_ (
);

MUX2X1 _1766_ (
    .A(DI[7]),
    .B(DIHOLD[7]),
    .S(RDY_bF$buf7),
    .Y(_893_)
);

FILL FILL_4__3593_ (
);

FILL FILL_4__3173_ (
);

FILL FILL_6__3099_ (
);

FILL FILL_0__3493_ (
);

FILL FILL_0__3073_ (
);

FILL FILL_4__1906_ (
);

FILL FILL_7__2895_ (
);

FILL FILL_7__2475_ (
);

FILL FILL_7__2055_ (
);

FILL FILL_0__1806_ (
);

FILL FILL_3__2795_ (
);

FILL FILL_3__2375_ (
);

FILL FILL_5__3662_ (
);

FILL FILL_5__3242_ (
);

FILL FILL_1__3654_ (
);

FILL FILL_1__3234_ (
);

FILL FILL_2__1997_ (
);

FILL FILL_4__2864_ (
);

FILL FILL_4__2444_ (
);

FILL FILL_4__2024_ (
);

MUX2X1 _3089_ (
    .A(_699_),
    .B(_1006_),
    .S(_956_),
    .Y(_700_)
);

FILL FILL_0__2764_ (
);

FILL FILL_0__2344_ (
);

FILL FILL_6__3311_ (
);

FILL FILL_2__3303_ (
);

FILL FILL_4__3649_ (
);

FILL FILL_4__3229_ (
);

FILL FILL_0__3549_ (
);

FILL FILL_0__3129_ (
);

FILL FILL_5__2933_ (
);

FILL FILL_5__2513_ (
);

FILL FILL_1__2925_ (
);

FILL FILL_1__2505_ (
);

INVX1 _1995_ (
    .A(_1108_),
    .Y(_1109_)
);

AOI21X1 _3301_ (
    .A(_855_),
    .B(_858_),
    .C(_886__bF$buf3),
    .Y(_869_)
);

FILL FILL_3__2184_ (
);

FILL FILL_5__3471_ (
);

FILL FILL_5__3051_ (
);

FILL FILL_7__3069_ (
);

FILL FILL_1__3463_ (
);

FILL FILL_1__3043_ (
);

FILL FILL_4__2673_ (
);

FILL FILL_4__2253_ (
);

FILL FILL_6__2599_ (
);

FILL FILL_6__2179_ (
);

FILL FILL168150x158550 (
);

FILL FILL_0__2993_ (
);

FILL FILL_0__2573_ (
);

FILL FILL_6__3540_ (
);

FILL FILL_0__2153_ (
);

FILL FILL_6__3120_ (
);

FILL FILL_2__3532_ (
);

FILL FILL_2__3112_ (
);

FILL FILL_4__3458_ (
);

FILL FILL_4__3038_ (
);

FILL FILL_3__1875_ (
);

FILL FILL_5__2742_ (
);

FILL FILL_5__2322_ (
);

FILL FILL_1__2734_ (
);

FILL FILL_1__2314_ (
);

FILL FILL_3__3601_ (
);

FILL FILL_5__3527_ (
);

FILL FILL_5__3107_ (
);

FILL FILL_1__3519_ (
);

FILL FILL_4__1944_ (
);

OAI21X1 _2589_ (
    .A(_268_),
    .B(_218_),
    .C(_275_),
    .Y(_1741_[8])
);

NAND2X1 _2169_ (
    .A(_1277_),
    .B(_1274_),
    .Y(_1278_)
);

FILL FILL_7__2093_ (
);

FILL FILL_0__1844_ (
);

FILL FILL_6__2811_ (
);

AOI21X1 _3530_ (
    .A(_1553_),
    .B(_1558_),
    .C(_1559_),
    .Y(_1560_)
);

NAND3X1 _3110_ (
    .A(_204_),
    .B(_717_),
    .C(_1022_),
    .Y(_718_)
);

FILL FILL_2__2803_ (
);

FILL FILL_4__2729_ (
);

FILL FILL_4__2309_ (
);

FILL FILL_7__3298_ (
);

FILL FILL_5__3280_ (
);

FILL FILL_0__2629_ (
);

FILL FILL_0__2209_ (
);

FILL FILL_1__3692_ (
);

FILL FILL_1__3272_ (
);

FILL FILL_3__3198_ (
);

FILL FILL_4__2482_ (
);

FILL FILL_4__2062_ (
);

FILL FILL_0__2382_ (
);

FILL FILL_7__1784_ (
);

FILL FILL_4__3267_ (
);

NOR2X1 _2801_ (
    .A(_290_),
    .B(_352_),
    .Y(_464_)
);

FILL FILL_0__3587_ (
);

FILL FILL_0__3167_ (
);

FILL FILL167850x75750 (
);

FILL FILL_5__2971_ (
);

FILL FILL_7__2569_ (
);

FILL FILL_5__2551_ (
);

FILL FILL_5__2131_ (
);

FILL FILL_1__2963_ (
);

FILL FILL_1__2543_ (
);

FILL FILL_1__2123_ (
);

FILL FILL_3__2889_ (
);

FILL FILL_3__2469_ (
);

FILL FILL_3__2049_ (
);

FILL FILL_4__1753_ (
);

NOR2X1 _2398_ (
    .A(_1369_),
    .B(_1502_),
    .Y(_1503_)
);

FILL FILL_6__2620_ (
);

FILL FILL_6__2200_ (
);

FILL FILL_2__2612_ (
);

FILL FILL_4__2958_ (
);

FILL FILL_4__2538_ (
);

FILL FILL_4__2118_ (
);

FILL FILL_0__2858_ (
);

FILL FILL_0__2438_ (
);

FILL FILL_0__2018_ (
);

FILL FILL_1__3081_ (
);

FILL FILL_5__1822_ (
);

FILL FILL_1__1814_ (
);

FILL FILL_4__2291_ (
);

FILL FILL_5__2607_ (
);

FILL FILL_0__2191_ (
);

FILL FILL_2__3570_ (
);

FILL FILL_2__3150_ (
);

FILL FILL_4__3496_ (
);

FILL FILL_4__3076_ (
);

OAI21X1 _2610_ (
    .A(_291_),
    .B(_270_),
    .C(_292_),
    .Y(_293_)
);

FILL FILL_4__1809_ (
);

FILL FILL_5__2780_ (
);

FILL FILL_7__2798_ (
);

FILL FILL_5__2360_ (
);

FILL FILL_1__2772_ (
);

FILL FILL_1__2352_ (
);

FILL FILL_3__2698_ (
);

FILL FILL_3__2278_ (
);

FILL FILL_5__3565_ (
);

FILL FILL_5__3145_ (
);

FILL FILL_1__3557_ (
);

FILL FILL_1__3137_ (
);

FILL FILL_4__1982_ (
);

FILL FILL_0__1882_ (
);

FILL FILL_2__2841_ (
);

FILL FILL_2__2421_ (
);

FILL FILL_2__2001_ (
);

FILL FILL_4__2767_ (
);

FILL FILL_4__2347_ (
);

FILL FILL_0__2667_ (
);

FILL FILL_6__3634_ (
);

FILL FILL_0__2247_ (
);

FILL FILL_6__3214_ (
);

FILL FILL_2__3626_ (
);

FILL FILL_2__3206_ (
);

FILL FILL_3__1969_ (
);

FILL FILL_3__2910_ (
);

FILL FILL_5__2836_ (
);

FILL FILL_5__2416_ (
);

FILL FILL_1__2828_ (
);

FILL FILL_1__2408_ (
);

INVX2 _1898_ (
    .A(PC[7]),
    .Y(_1016_)
);

FILL FILL_7__2187_ (
);

FILL FILL_0__1938_ (
);

FILL FILL_6__2905_ (
);

INVX1 _3624_ (
    .A(_1653_),
    .Y(_1654_)
);

OAI21X1 _3204_ (
    .A(_720__bF$buf1),
    .B(_687_),
    .C(\AXYS[1] [7]),
    .Y(_797_)
);

FILL FILL_1__2581_ (
);

FILL FILL_1__2161_ (
);

FILL FILL_3__2087_ (
);

FILL FILL_4__1791_ (
);

FILL FILL_2__2650_ (
);

FILL FILL_2__2230_ (
);

FILL FILL_4__2996_ (
);

FILL FILL_4__2576_ (
);

FILL FILL_4__2156_ (
);

FILL FILL_0__2896_ (
);

FILL FILL_0__2476_ (
);

FILL FILL_0__2056_ (
);

FILL FILL_6__3023_ (
);

FILL FILL_2__3015_ (
);

FILL FILL_5__1860_ (
);

FILL FILL_1__1852_ (
);

FILL FILL_3__1778_ (
);

FILL FILL_5__2645_ (
);

FILL FILL_5__2225_ (
);

FILL FILL_1__2637_ (
);

FILL FILL_7__3604_ (
);

FILL FILL_1__2217_ (
);

FILL FILL_3__3504_ (
);

FILL FILL_2__1921_ (
);

FILL FILL_4__1847_ (
);

FILL FILL_0__1747_ (
);

FILL FILL_6__2714_ (
);

DFFSR _3433_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_101_),
    .CLK(clk_bF$buf1),
    .Q(ABL[0])
);

NAND2X1 _3013_ (
    .A(_638_),
    .B(_609_),
    .Y(_639_)
);

FILL FILL_1__2390_ (
);

FILL FILL_2__2706_ (
);

FILL FILL_1_BUFX2_insert40 (
);

FILL FILL_1_BUFX2_insert41 (
);

FILL FILL_1_BUFX2_insert42 (
);

FILL FILL_1_BUFX2_insert43 (
);

FILL FILL_5__3183_ (
);

FILL FILL_1_BUFX2_insert44 (
);

FILL FILL_1_BUFX2_insert45 (
);

FILL FILL_1_BUFX2_insert46 (
);

FILL FILL_1_BUFX2_insert47 (
);

FILL FILL_1_BUFX2_insert48 (
);

FILL FILL_1_BUFX2_insert49 (
);

FILL FILL_1__3595_ (
);

FILL FILL_1__3175_ (
);

FILL FILL_5__1916_ (
);

FILL FILL_0_CLKBUF1_insert26 (
);

FILL FILL_0_CLKBUF1_insert27 (
);

FILL FILL_0_CLKBUF1_insert28 (
);

FILL FILL_0_CLKBUF1_insert29 (
);

FILL FILL_1__1908_ (
);

FILL FILL_4__2385_ (
);

FILL FILL_6__3672_ (
);

FILL FILL_0__2285_ (
);

FILL FILL_6__3252_ (
);

FILL FILL_2__3664_ (
);

FILL FILL_2__3244_ (
);

AND2X2 _2704_ (
    .A(_370_),
    .B(_374_),
    .Y(_375_)
);

FILL FILL_5__2874_ (
);

FILL FILL_5__2454_ (
);

FILL FILL_5__2034_ (
);

FILL FILL_1__2866_ (
);

FILL FILL_1__2446_ (
);

FILL FILL_1__2026_ (
);

FILL FILL_3__3313_ (
);

FILL FILL_5__3659_ (
);

FILL FILL_5__3239_ (
);

FILL FILL_0__1976_ (
);

FILL FILL_6__2943_ (
);

OAI21X1 _3662_ (
    .A(_1714__bF$buf1),
    .B(_1623_),
    .C(_1688_),
    .Y(_1518_)
);

FILL FILL_6__2523_ (
);

FILL FILL_6__2103_ (
);

OAI21X1 _3242_ (
    .A(_931__bF$buf1),
    .B(_928_),
    .C(_1027__bF$buf1),
    .Y(_818_)
);

FILL FILL_2__2935_ (
);

FILL FILL_2__2515_ (
);

FILL FILL_6__3308_ (
);

FILL FILL_0__3702_ (
);

FILL FILL_4__2194_ (
);

FILL FILL_6__3481_ (
);

FILL FILL_0__2094_ (
);

FILL FILL_6__3061_ (
);

FILL FILL_2__3473_ (
);

FILL FILL_2__3053_ (
);

NAND2X1 _2933_ (
    .A(_1327_),
    .B(_1395_),
    .Y(_576_)
);

NOR2X1 _2513_ (
    .A(_1464_),
    .B(_207_),
    .Y(_208_)
);

FILL FILL_1__1890_ (
);

FILL FILL_0__3299_ (
);

FILL FILL_5__2683_ (
);

FILL FILL_5__2263_ (
);

FILL FILL_1__2675_ (
);

FILL FILL_7__3642_ (
);

FILL FILL_1__2255_ (
);

FILL FILL_7__3222_ (
);

FILL FILL_3__3542_ (
);

FILL FILL_3__3122_ (
);

FILL FILL_5__3468_ (
);

FILL FILL_5__3048_ (
);

FILL FILL_4__1885_ (
);

FILL FILL_0__1785_ (
);

FILL FILL_6__2752_ (
);

NAND2X1 _3471_ (
    .A(alu_op[0]),
    .B(_1716_),
    .Y(_1717_)
);

FILL FILL_6__2332_ (
);

NAND2X1 _3051_ (
    .A(plp),
    .B(ADD[6]),
    .Y(_666_)
);

FILL FILL_2__2744_ (
);

FILL FILL_2__2324_ (
);

FILL FILL169650x158550 (
);

FILL FILL_4__3611_ (
);

FILL FILL_6__3537_ (
);

FILL FILL_6__3117_ (
);

FILL FILL_2__3529_ (
);

FILL FILL_0__3511_ (
);

FILL FILL_2__3109_ (
);

FILL FILL_5__1954_ (
);

FILL FILL_1__1946_ (
);

FILL FILL_3__2813_ (
);

FILL FILL_5__2739_ (
);

FILL FILL_5__2319_ (
);

FILL FILL_6__3290_ (
);

FILL FILL_2__3282_ (
);

OAI21X1 _2742_ (
    .A(_268_),
    .B(_352_),
    .C(_408_),
    .Y(_409_)
);

NAND3X1 _2322_ (
    .A(_1426_),
    .B(_1428_),
    .C(_1425_),
    .Y(_1429_)
);

FILL FILL_5__2492_ (
);

FILL FILL_5__2072_ (
);

FILL FILL_6__2808_ (
);

OAI22X1 _3527_ (
    .A(_1722_),
    .B(_1539_),
    .C(_1556_),
    .D(_1552_),
    .Y(_1557_)
);

NAND2X1 _3107_ (
    .A(RDY_bF$buf9),
    .B(DI[7]),
    .Y(_716_)
);

FILL FILL_1__2484_ (
);

FILL FILL_7__3451_ (
);

FILL FILL_1__2064_ (
);

FILL FILL_5__3697_ (
);

FILL FILL_5__3277_ (
);

FILL FILL_1__3269_ (
);

FILL FILL_6__2981_ (
);

FILL FILL_6__2561_ (
);

OAI21X1 _3280_ (
    .A(_903__bF$buf0),
    .B(_969_),
    .C(_977_),
    .Y(_856_)
);

FILL FILL_6__2141_ (
);

FILL FILL_2__2973_ (
);

FILL FILL_2__2553_ (
);

FILL FILL_2__2133_ (
);

FILL FILL_4__2899_ (
);

FILL FILL_4__2479_ (
);

FILL FILL_4__2059_ (
);

FILL FILL_4__3000_ (
);

FILL FILL_0__2799_ (
);

FILL FILL_0__2379_ (
);

FILL FILL_5__1763_ (
);

FILL FILL_1__1755_ (
);

FILL FILL_7__2722_ (
);

FILL FILL_3__2622_ (
);

FILL FILL_3__2202_ (
);

FILL FILL_5__2968_ (
);

FILL FILL_5__2548_ (
);

FILL FILL_5__2128_ (
);

FILL FILL_2__3091_ (
);

FILL FILL_6__1832_ (
);

NOR2X1 _2971_ (
    .A(_1172_),
    .B(_1214_),
    .Y(_603_)
);

INVX1 _2551_ (
    .A(_242_),
    .Y(_1741_[3])
);

NOR2X1 _2131_ (
    .A(_1239_),
    .B(_1237_),
    .Y(_1240_)
);

FILL FILL_2__1824_ (
);

FILL FILL_6__2617_ (
);

DFFSR _3336_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_14_),
    .CLK(clk_bF$buf2),
    .Q(PC[12])
);

FILL FILL_1__2293_ (
);

FILL FILL_2__2609_ (
);

FILL FILL_3__3580_ (
);

FILL FILL_3__3160_ (
);

FILL FILL_5__3086_ (
);

FILL FILL_1__3498_ (
);

FILL FILL_1__3078_ (
);

FILL FILL_5__1819_ (
);

FILL FILL_6__2790_ (
);

FILL FILL_6__2370_ (
);

FILL FILL_2__2782_ (
);

FILL FILL_2__2362_ (
);

FILL FILL_4__2288_ (
);

NOR2X1 _1822_ (
    .A(state[0]),
    .B(_905_),
    .Y(_948_)
);

FILL FILL_6__3575_ (
);

FILL FILL_0__2188_ (
);

FILL FILL_6__3155_ (
);

FILL FILL_2__3567_ (
);

FILL FILL_2__3147_ (
);

FILL FILL_5__1992_ (
);

INVX1 _2607_ (
    .A(PC[12]),
    .Y(_290_)
);

FILL FILL_1__1984_ (
);

FILL FILL_7__2951_ (
);

FILL FILL_7__2111_ (
);

FILL FILL169350x144150 (
);

FILL FILL_3__2851_ (
);

FILL FILL_3__2431_ (
);

FILL FILL_3__2011_ (
);

FILL FILL_5__2777_ (
);

FILL FILL_5__2357_ (
);

FILL FILL_1__2769_ (
);

FILL FILL_1__2349_ (
);

FILL FILL_1__3710_ (
);

FILL FILL_3__3636_ (
);

FILL FILL_3__3216_ (
);

OAI22X1 _2780_ (
    .A(RDY_bF$buf4),
    .B(_280_),
    .C(_444_),
    .D(_439_),
    .Y(_12_)
);

AND2X2 _2360_ (
    .A(_1463_),
    .B(_1465_),
    .Y(_1466_)
);

FILL FILL_4__1979_ (
);

FILL FILL_4__2920_ (
);

FILL FILL_4__2500_ (
);

FILL FILL_0__1879_ (
);

FILL FILL_6__2846_ (
);

OAI21X1 _3565_ (
    .A(_1594_),
    .B(_1593_),
    .C(_1571_),
    .Y(_1595_)
);

FILL FILL_6__2426_ (
);

FILL FILL_6__2006_ (
);

NAND2X1 _3145_ (
    .A(_748_),
    .B(_749_),
    .Y(_750_)
);

FILL FILL_2__2838_ (
);

FILL FILL_0__2820_ (
);

FILL FILL_2__2418_ (
);

FILL FILL_0__2400_ (
);

FILL FILL_4__3705_ (
);

FILL FILL_0__3605_ (
);

FILL FILL_2__2591_ (
);

FILL FILL_2__2171_ (
);

FILL FILL_4__2097_ (
);

FILL FILL_3__2907_ (
);

FILL FILL_6_BUFX2_insert40 (
);

FILL FILL_6_BUFX2_insert41 (
);

FILL FILL_6_BUFX2_insert42 (
);

FILL FILL_6_BUFX2_insert43 (
);

FILL FILL_6_BUFX2_insert44 (
);

FILL FILL_6_BUFX2_insert45 (
);

FILL FILL_6_BUFX2_insert46 (
);

FILL FILL_6_BUFX2_insert47 (
);

FILL FILL_6_BUFX2_insert48 (
);

FILL FILL_6_BUFX2_insert49 (
);

NOR3X1 _2836_ (
    .A(_465_),
    .B(_497_),
    .C(_485_),
    .Y(_498_)
);

NOR2X1 _2416_ (
    .A(_121_),
    .B(_124_),
    .Y(_125_)
);

FILL FILL_1__1793_ (
);

FILL FILL_7__2340_ (
);

FILL FILL_3__2660_ (
);

FILL FILL_3__2240_ (
);

FILL FILL_5__2586_ (
);

FILL FILL_5__2166_ (
);

FILL FILL_1__2998_ (
);

FILL FILL_1__2578_ (
);

FILL FILL_7__3545_ (
);

FILL FILL_1__2158_ (
);

FILL FILL_7__3125_ (
);

FILL FILL_3__3025_ (
);

FILL FILL_6__1870_ (
);

FILL FILL_2__1862_ (
);

FILL FILL_4__1788_ (
);

FILL FILL_6__2655_ (
);

DFFSR _3374_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_51_),
    .CLK(clk_bF$buf10),
    .Q(load_reg)
);

FILL FILL_6__2235_ (
);

FILL FILL_2__2647_ (
);

FILL FILL_2__2227_ (
);

FILL FILL_4__3514_ (
);

FILL FILL_3__1931_ (
);

FILL FILL_5__1857_ (
);

FILL FILL_1__1849_ (
);

FILL FILL_7__2816_ (
);

FILL FILL_3__2716_ (
);

OAI21X1 _1860_ (
    .A(_914__bF$buf4),
    .B(_984_),
    .C(_983_),
    .Y(_985_)
);

FILL FILL_6__3193_ (
);

FILL FILL_2__3185_ (
);

FILL FILL_6__1926_ (
);

NAND3X1 _2645_ (
    .A(_1432_),
    .B(_316_),
    .C(_319_),
    .Y(_320_)
);

AOI22X1 _2225_ (
    .A(_886__bF$buf1),
    .B(_943_),
    .C(_1332_),
    .D(_1330_),
    .Y(_1333_)
);

FILL FILL_2__1918_ (
);

FILL FILL_0__1900_ (
);

FILL FILL_5__2395_ (
);

FILL FILL_1__2387_ (
);

FILL FILL_3__3674_ (
);

FILL FILL_3__3254_ (
);

FILL FILL_6__2884_ (
);

FILL FILL_6__2464_ (
);

INVX1 _3183_ (
    .A(_783_),
    .Y(_784_)
);

FILL FILL_6__2044_ (
);

FILL FILL_2__2876_ (
);

FILL FILL_2__2456_ (
);

FILL FILL_2__2036_ (
);

OAI21X1 _1916_ (
    .A(_914__bF$buf0),
    .B(_942_),
    .C(_1032_),
    .Y(_1033_)
);

FILL FILL_7__1840_ (
);

FILL FILL_6__3669_ (
);

FILL FILL_6__3249_ (
);

FILL FILL_0__3643_ (
);

FILL FILL_0__3223_ (
);

FILL FILL_7__2625_ (
);

FILL FILL_3__2945_ (
);

FILL FILL_3__2525_ (
);

FILL FILL_3__2105_ (
);

INVX1 _2874_ (
    .A(plp),
    .Y(_529_)
);

AOI22X1 _2454_ (
    .A(PC[1]),
    .B(_1080_),
    .C(_144_),
    .D(ADD[1]),
    .Y(_156_)
);

INVX1 _2034_ (
    .A(ABH[7]),
    .Y(_1144_)
);

OAI21X1 _3659_ (
    .A(_1612_),
    .B(_1686_),
    .C(RDY_bF$buf9),
    .Y(_1687_)
);

OAI21X1 _3239_ (
    .A(_720__bF$buf3),
    .B(_808_),
    .C(\AXYS[3] [7]),
    .Y(_816_)
);

FILL FILL_7__3583_ (
);

FILL FILL_1__2196_ (
);

FILL FILL_0__2914_ (
);

FILL FILL_3__3483_ (
);

FILL FILL_3__3063_ (
);

FILL FILL_6__2693_ (
);

FILL FILL_6__2273_ (
);

FILL FILL_2__2685_ (
);

FILL FILL_2__2265_ (
);

FILL FILL_4__3552_ (
);

FILL FILL_4__3132_ (
);

FILL FILL_6__3478_ (
);

FILL FILL_6__3058_ (
);

FILL FILL169650x18150 (
);

FILL FILL_0__3452_ (
);

FILL FILL_0__3032_ (
);

FILL FILL_5__1895_ (
);

FILL FILL_1__1887_ (
);

FILL FILL_7__2854_ (
);

FILL FILL_7__2014_ (
);

FILL FILL_3__2754_ (
);

FILL FILL_3__2334_ (
);

FILL FILL_5__3621_ (
);

FILL FILL_5__3201_ (
);

FILL FILL_7__3219_ (
);

FILL FILL_1__3613_ (
);

FILL FILL_3__3539_ (
);

FILL FILL_3__3119_ (
);

FILL FILL_6__1964_ (
);

INVX1 _2683_ (
    .A(ADD[3]),
    .Y(_355_)
);

NAND3X1 _2263_ (
    .A(_1150__bF$buf3),
    .B(_1365_),
    .C(_1370_),
    .Y(_1371_)
);

FILL FILL_2__1956_ (
);

FILL FILL_4__2823_ (
);

FILL FILL_4__2403_ (
);

FILL FILL_6__2749_ (
);

INVX4 _3468_ (
    .A(RDY_bF$buf7),
    .Y(_1714_)
);

FILL FILL_6__2329_ (
);

NOR2X1 _3048_ (
    .A(clv),
    .B(_662_),
    .Y(_663_)
);

FILL FILL_0__2723_ (
);

FILL FILL_0__2303_ (
);

FILL FILL_3__3292_ (
);

FILL FILL_4__3608_ (
);

FILL FILL_0__3508_ (
);

FILL FILL_6__2082_ (
);

FILL FILL_2__2494_ (
);

FILL FILL_2__2074_ (
);

NOR2X1 _1954_ (
    .A(_1068_),
    .B(_1070_),
    .Y(_1071_)
);

FILL FILL_6__3287_ (
);

FILL FILL_2__3699_ (
);

FILL FILL_0__3261_ (
);

FILL FILL_2__3279_ (
);

NAND2X1 _2739_ (
    .A(ABH[0]),
    .B(_323_),
    .Y(_406_)
);

OAI21X1 _2319_ (
    .A(_908_),
    .B(_1031_),
    .C(_903__bF$buf0),
    .Y(_1426_)
);

FILL FILL_7__2243_ (
);

FILL FILL_3__2983_ (
);

FILL FILL_3__2563_ (
);

FILL FILL_3__2143_ (
);

FILL FILL_5__2489_ (
);

FILL FILL_5__2069_ (
);

FILL FILL_7__3028_ (
);

FILL FILL_5__3010_ (
);

FILL FILL_1__3002_ (
);

FILL FILL_6__1773_ (
);

OAI21X1 _2492_ (
    .A(_1319__bF$buf0),
    .B(_1263_),
    .C(PC[15]),
    .Y(_188_)
);

AOI21X1 _2072_ (
    .A(_1168_),
    .B(_1013_),
    .C(_1180_),
    .Y(_1181_)
);

FILL FILL_2__1765_ (
);

FILL FILL_4__2632_ (
);

FILL FILL_4__2212_ (
);

FILL FILL_6__2978_ (
);

BUFX2 _3697_ (
    .A(_1741_[14]),
    .Y(AB[14])
);

FILL FILL_6__2558_ (
);

AND2X2 _3277_ (
    .A(_836_),
    .B(_824_),
    .Y(_853_)
);

FILL FILL_6__2138_ (
);

FILL FILL_0__2952_ (
);

FILL FILL_0__2532_ (
);

FILL FILL_0__2112_ (
);

FILL FILL_7__1934_ (
);

FILL FILL_3__1834_ (
);

FILL FILL_0__3317_ (
);

FILL FILL_7__2719_ (
);

FILL FILL_5__2701_ (
);

FILL FILL_3__2619_ (
);

INVX1 _1763_ (
    .A(DIHOLD[6]),
    .Y(_891_)
);

FILL FILL_4__3590_ (
);

FILL FILL_4__3170_ (
);

FILL FILL_6__3096_ (
);

FILL FILL_0__3490_ (
);

FILL FILL_2__3088_ (
);

FILL FILL_0__3070_ (
);

FILL FILL_4__1903_ (
);

FILL FILL_6__1829_ (
);

OAI22X1 _2968_ (
    .A(_1207_),
    .B(_1150__bF$buf0),
    .C(_550_),
    .D(_600_),
    .Y(_44_)
);

AOI21X1 _2548_ (
    .A(_237_),
    .B(ADD[3]),
    .C(_239_),
    .Y(_240_)
);

OAI21X1 _2128_ (
    .A(_886__bF$buf0),
    .B(_1234_),
    .C(_1236_),
    .Y(_1237_)
);

FILL FILL_7__2472_ (
);

FILL FILL_0__1803_ (
);

FILL FILL_3__2792_ (
);

FILL FILL_3__2372_ (
);

FILL FILL_5__2298_ (
);

FILL FILL_7__3677_ (
);

FILL FILL_7__3257_ (
);

FILL FILL_1__3651_ (
);

FILL FILL_1__3231_ (
);

FILL FILL_3__3577_ (
);

FILL FILL_3__3157_ (
);

FILL FILL_2__1994_ (
);

FILL FILL_4__2861_ (
);

FILL FILL_4__2441_ (
);

FILL FILL_4__2021_ (
);

FILL FILL_6__2787_ (
);

FILL FILL_6__2367_ (
);

INVX1 _3086_ (
    .A(Z),
    .Y(_697_)
);

FILL FILL_2__2779_ (
);

FILL FILL_0__2761_ (
);

FILL FILL_2__2359_ (
);

FILL FILL_0__2341_ (
);

FILL FILL_2__3300_ (
);

NAND3X1 _1819_ (
    .A(_940_),
    .B(_936_),
    .C(_944_),
    .Y(_945_)
);

FILL FILL_4__3646_ (
);

FILL FILL_4__3226_ (
);

FILL FILL_0__3546_ (
);

FILL FILL_0__3126_ (
);

FILL FILL_5__1989_ (
);

FILL FILL_7__2948_ (
);

FILL FILL_5__2930_ (
);

FILL FILL_5__2510_ (
);

FILL FILL_7__2108_ (
);

FILL FILL_1__2922_ (
);

FILL FILL_1__2502_ (
);

FILL FILL_3__2848_ (
);

FILL FILL_3__2428_ (
);

FILL FILL_3__2008_ (
);

AOI22X1 _1992_ (
    .A(_1049_),
    .B(\AXYS[3] [3]),
    .C(\AXYS[2] [3]),
    .D(_1057_),
    .Y(_1106_)
);

FILL FILL_5__3715_ (
);

FILL FILL_1__3707_ (
);

NAND2X1 _2777_ (
    .A(_433_),
    .B(_436_),
    .Y(_442_)
);

AOI22X1 _2357_ (
    .A(_886__bF$buf1),
    .B(_1268_),
    .C(_1283_),
    .D(_1330_),
    .Y(_1463_)
);

FILL FILL_3__2181_ (
);

FILL FILL_4__2917_ (
);

FILL FILL_1__2099_ (
);

FILL FILL_0__2817_ (
);

FILL FILL_1__3460_ (
);

FILL FILL_1__3040_ (
);

FILL FILL169350x150 (
);

FILL FILL_4__2670_ (
);

FILL FILL_4__2250_ (
);

FILL FILL_6__2596_ (
);

FILL FILL_6__2176_ (
);

FILL FILL_0__2990_ (
);

FILL FILL_2__2588_ (
);

FILL FILL_0__2570_ (
);

FILL FILL_2__2168_ (
);

FILL FILL_0__2150_ (
);

FILL FILL_7__1972_ (
);

FILL FILL_4__3455_ (
);

FILL FILL_4__3035_ (
);

FILL FILL_3__1872_ (
);

FILL FILL_5__1798_ (
);

FILL FILL_7__2337_ (
);

FILL FILL_1__2731_ (
);

FILL FILL_1__2311_ (
);

FILL FILL_3__2657_ (
);

FILL FILL_3__2237_ (
);

FILL FILL_5__3524_ (
);

FILL FILL_5__3104_ (
);

FILL FILL_1__3516_ (
);

FILL FILL_4__1941_ (
);

FILL FILL_6__1867_ (
);

AOI22X1 _2586_ (
    .A(ADD[0]),
    .B(_198_),
    .C(_272_),
    .D(DIMUX[0]),
    .Y(_273_)
);

NOR2X1 _2166_ (
    .A(_914__bF$buf1),
    .B(_974_),
    .Y(_1275_)
);

FILL FILL_7__2090_ (
);

FILL FILL_0__1841_ (
);

FILL FILL_2__1859_ (
);

FILL FILL_2__2800_ (
);

FILL FILL_4__2726_ (
);

FILL FILL_4__2306_ (
);

FILL FILL_0__2626_ (
);

FILL FILL_0__2206_ (
);

FILL FILL_3__3195_ (
);

FILL FILL_3__1928_ (
);

FILL FILL_2__2397_ (
);

NOR2X1 _1857_ (
    .A(_902__bF$buf2),
    .B(_981_),
    .Y(_982_)
);

FILL FILL_4__3264_ (
);

FILL FILL_0__3584_ (
);

FILL FILL_0__3164_ (
);

FILL FILL_7__2986_ (
);

FILL FILL_7__2566_ (
);

FILL FILL_7__2146_ (
);

FILL FILL_1__2960_ (
);

FILL FILL_1__2540_ (
);

FILL FILL_1__2120_ (
);

FILL FILL_3__2886_ (
);

FILL FILL_3__2466_ (
);

FILL FILL_3__2046_ (
);

FILL FILL_4__1750_ (
);

NAND3X1 _2395_ (
    .A(_1262_),
    .B(_1308_),
    .C(_1274_),
    .Y(_1500_)
);

FILL FILL_4__2955_ (
);

FILL FILL_4__2535_ (
);

FILL FILL_4__2115_ (
);

FILL FILL_0__2855_ (
);

FILL FILL_0__2435_ (
);

FILL FILL_0__2015_ (
);

FILL FILL_7__1837_ (
);

FILL FILL_1__1811_ (
);

FILL FILL_5__2604_ (
);

FILL FILL_4__3493_ (
);

FILL FILL_4__3073_ (
);

FILL FILL_4__1806_ (
);

FILL FILL_7__2795_ (
);

FILL FILL_7__2375_ (
);

FILL FILL_3__2695_ (
);

FILL FILL_3__2275_ (
);

FILL FILL_5__3562_ (
);

FILL FILL_5__3142_ (
);

FILL FILL_1__3554_ (
);

FILL FILL_1__3134_ (
);

FILL FILL_2__1897_ (
);

FILL FILL_4__2764_ (
);

FILL FILL_4__2344_ (
);

FILL FILL_0__2664_ (
);

FILL FILL_6__3631_ (
);

FILL FILL_0__2244_ (
);

FILL FILL_6__3211_ (
);

FILL FILL_2__3623_ (
);

FILL FILL_2__3203_ (
);

FILL FILL_4__3549_ (
);

FILL FILL_4__3129_ (
);

FILL FILL_3__1966_ (
);

FILL FILL_0__3449_ (
);

FILL FILL_0__3029_ (
);

FILL FILL_5__2833_ (
);

FILL FILL_5__2413_ (
);

FILL FILL_1__2825_ (
);

FILL FILL_1__2405_ (
);

FILL FILL168450x158550 (
);

INVX2 _1895_ (
    .A(PC[6]),
    .Y(_1014_)
);

FILL FILL_5__3618_ (
);

FILL FILL_7__2184_ (
);

FILL FILL_0__1935_ (
);

FILL FILL_6__2902_ (
);

OAI21X1 _3621_ (
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1647_),
    .Y(_1651_)
);

OAI21X1 _3201_ (
    .A(_767_),
    .B(_789_),
    .C(_795_),
    .Y(_82_)
);

FILL FILL_3__2084_ (
);

FILL FILL_3__3289_ (
);

FILL FILL_4__2993_ (
);

FILL FILL_4__2573_ (
);

FILL FILL_4__2153_ (
);

FILL FILL_6__2499_ (
);

FILL FILL_6__2079_ (
);

FILL FILL_0__2893_ (
);

FILL FILL_0__2473_ (
);

FILL FILL_0__2053_ (
);

FILL FILL_6__3020_ (
);

FILL FILL_2__3012_ (
);

FILL FILL_0__3678_ (
);

FILL FILL_3__1775_ (
);

FILL FILL_0__3258_ (
);

FILL FILL_5__2642_ (
);

FILL FILL_5__2222_ (
);

FILL FILL_1__2634_ (
);

FILL FILL_7__3601_ (
);

FILL FILL_1__2214_ (
);

FILL FILL_3__3501_ (
);

FILL FILL_5__3007_ (
);

FILL FILL_4__1844_ (
);

OAI21X1 _2489_ (
    .A(_1374_),
    .B(_165_),
    .C(_185_),
    .Y(_186_)
);

NAND2X1 _2069_ (
    .A(_1167_),
    .B(_1177_),
    .Y(_1178_)
);

FILL FILL_0__1744_ (
);

FILL FILL_6__2711_ (
);

DFFSR _3430_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_98_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[3] [5])
);

OAI21X1 _3010_ (
    .A(_1394_),
    .B(_578_),
    .C(_635_),
    .Y(_636_)
);

FILL FILL_2__2703_ (
);

FILL FILL_4__2629_ (
);

FILL FILL_4__2209_ (
);

FILL FILL_1_BUFX2_insert10 (
);

FILL FILL_1_BUFX2_insert11 (
);

FILL FILL_1_BUFX2_insert12 (
);

FILL FILL_1_BUFX2_insert13 (
);

FILL FILL_5__3180_ (
);

FILL FILL_7__3198_ (
);

FILL FILL_1_BUFX2_insert14 (
);

FILL FILL_1_BUFX2_insert15 (
);

FILL FILL_1_BUFX2_insert16 (
);

FILL FILL_1_BUFX2_insert17 (
);

FILL FILL_1_BUFX2_insert18 (
);

FILL FILL_1_BUFX2_insert19 (
);

FILL FILL_0__2949_ (
);

FILL FILL_0__2529_ (
);

FILL FILL_0__2109_ (
);

FILL FILL_1__3592_ (
);

FILL FILL_1__3172_ (
);

FILL FILL_3__3098_ (
);

FILL FILL_5__1913_ (
);

FILL FILL_1__1905_ (
);

FILL FILL_4__2382_ (
);

FILL FILL_0__2282_ (
);

FILL FILL_2__3661_ (
);

FILL FILL_2__3241_ (
);

FILL FILL_4__3587_ (
);

FILL FILL_4__3167_ (
);

AOI21X1 _2701_ (
    .A(ABL[4]),
    .B(_323_),
    .C(_1334_),
    .Y(_372_)
);

FILL FILL_0__3487_ (
);

FILL FILL_0__3067_ (
);

FILL FILL_5__2871_ (
);

FILL FILL_5__2451_ (
);

FILL FILL_7__2469_ (
);

FILL FILL_5__2031_ (
);

FILL FILL_1__2863_ (
);

FILL FILL_1__2443_ (
);

FILL FILL_1__2023_ (
);

FILL FILL_3__2789_ (
);

FILL FILL_3__2369_ (
);

FILL FILL_3__3310_ (
);

FILL FILL_5__3656_ (
);

FILL FILL_5__3236_ (
);

FILL FILL169350x64950 (
);

FILL FILL_1__3648_ (
);

FILL FILL_1__3228_ (
);

FILL FILL_6__1999_ (
);

NOR2X1 _2298_ (
    .A(_1159_),
    .B(_1404_),
    .Y(_1405_)
);

FILL FILL168150x144150 (
);

FILL FILL_0__1973_ (
);

FILL FILL_6__2940_ (
);

FILL FILL_6__2520_ (
);

FILL FILL_6__2100_ (
);

FILL FILL_2__2932_ (
);

FILL FILL_2__2512_ (
);

FILL FILL_4__2858_ (
);

FILL FILL_4__2438_ (
);

FILL FILL_4__2018_ (
);

FILL FILL_0__2758_ (
);

FILL FILL_0__2338_ (
);

FILL FILL_6__3305_ (
);

FILL FILL_4__2191_ (
);

FILL FILL_5__2927_ (
);

FILL FILL_5__2507_ (
);

FILL FILL_0__2091_ (
);

FILL FILL_1__2919_ (
);

FILL FILL_2__3470_ (
);

AOI21X1 _1989_ (
    .A(_1082_),
    .B(ADD[2]),
    .C(_1103_),
    .Y(_1104_)
);

FILL FILL_2__3050_ (
);

NAND2X1 _2930_ (
    .A(_1164_),
    .B(_1178_),
    .Y(_573_)
);

NAND3X1 _2510_ (
    .A(_1077_),
    .B(_204_),
    .C(_1081_),
    .Y(_205_)
);

FILL FILL_0__3296_ (
);

FILL FILL_7__2698_ (
);

FILL FILL_5__2680_ (
);

FILL FILL_5__2260_ (
);

BUFX2 _3715_ (
    .A(_1743_),
    .Y(WE)
);

FILL FILL_1__2672_ (
);

FILL FILL_1__2252_ (
);

FILL FILL_3__2598_ (
);

FILL FILL_3__2178_ (
);

FILL FILL_5__3465_ (
);

FILL FILL_5__3045_ (
);

FILL FILL_1__3457_ (
);

FILL FILL_1__3037_ (
);

FILL FILL_4__1882_ (
);

FILL FILL_0__1782_ (
);

FILL FILL_2__2741_ (
);

FILL FILL_2__2321_ (
);

FILL FILL_4__2667_ (
);

FILL FILL_4__2247_ (
);

FILL FILL_0__2987_ (
);

FILL FILL_0__2567_ (
);

FILL FILL_6__3534_ (
);

FILL FILL_0__2147_ (
);

FILL FILL_6__3114_ (
);

FILL FILL167850x61350 (
);

FILL FILL_2__3526_ (
);

FILL FILL_2__3106_ (
);

FILL FILL_7__1969_ (
);

FILL FILL_5__1951_ (
);

FILL FILL_1__1943_ (
);

FILL FILL_3__1869_ (
);

FILL FILL_3__2810_ (
);

FILL FILL_5__2736_ (
);

FILL FILL_5__2316_ (
);

FILL FILL_2_BUFX2_insert60 (
);

FILL FILL_2_BUFX2_insert61 (
);

FILL FILL_2_BUFX2_insert62 (
);

FILL FILL_2_BUFX2_insert63 (
);

FILL FILL_2_BUFX2_insert64 (
);

FILL FILL_2_BUFX2_insert65 (
);

FILL FILL_2_BUFX2_insert66 (
);

FILL FILL_1__2728_ (
);

FILL FILL_2_BUFX2_insert67 (
);

FILL FILL_2_BUFX2_insert68 (
);

FILL FILL_1__2308_ (
);

FILL FILL_2_BUFX2_insert69 (
);

NAND2X1 _1798_ (
    .A(state[1]),
    .B(_906_),
    .Y(_924_)
);

FILL FILL_4__1938_ (
);

FILL FILL_7__2087_ (
);

FILL FILL_0__1838_ (
);

FILL FILL_6__2805_ (
);

INVX1 _3524_ (
    .A(AI[2]),
    .Y(_1554_)
);

MUX2X1 _3104_ (
    .A(_713_),
    .B(DIMUX[0]),
    .S(_956_),
    .Y(_714_)
);

FILL FILL_1__2481_ (
);

FILL FILL_1__2061_ (
);

FILL FILL_5__3694_ (
);

FILL FILL_5__3274_ (
);

FILL FILL_1__3266_ (
);

FILL FILL_2__2970_ (
);

FILL FILL_2__2550_ (
);

FILL FILL_2__2130_ (
);

FILL FILL_4__2896_ (
);

FILL FILL_4__2476_ (
);

FILL FILL_4__2056_ (
);

FILL FILL_0__2796_ (
);

FILL FILL_0__2376_ (
);

FILL FILL_5__1760_ (
);

FILL FILL_1__1752_ (
);

FILL FILL_5__2965_ (
);

FILL FILL_5__2545_ (
);

FILL FILL_5__2125_ (
);

FILL FILL_1__2957_ (
);

FILL FILL_1__2537_ (
);

FILL FILL_7__3504_ (
);

FILL FILL_1__2117_ (
);

FILL FILL_2__1821_ (
);

FILL FILL_4__1747_ (
);

FILL FILL_6__2614_ (
);

DFFSR _3333_ (
    .R(_1__bF$buf4),
    .S(vdd),
    .D(_11_),
    .CLK(clk_bF$buf2),
    .Q(PC[9])
);

FILL FILL_1__2290_ (
);

FILL FILL_2__2606_ (
);

FILL FILL_5__3083_ (
);

FILL FILL_1__3495_ (
);

FILL FILL_1__3075_ (
);

FILL FILL_5__1816_ (
);

FILL FILL_1__1808_ (
);

FILL FILL_4__2285_ (
);

FILL FILL_6__3572_ (
);

FILL FILL_0__2185_ (
);

FILL FILL_6__3152_ (
);

FILL FILL_2__3564_ (
);

FILL FILL_2__3144_ (
);

NAND2X1 _2604_ (
    .A(_287_),
    .B(_286_),
    .Y(_288_)
);

FILL FILL_1__1981_ (
);

FILL FILL_5__2774_ (
);

FILL FILL_5__2354_ (
);

FILL FILL_1__2766_ (
);

FILL FILL_1__2346_ (
);

FILL FILL_3__3633_ (
);

FILL FILL_3__3213_ (
);

FILL FILL_5__3559_ (
);

FILL FILL_5__3139_ (
);

FILL FILL_4__1976_ (
);

FILL FILL_0__1876_ (
);

FILL FILL_6__2843_ (
);

NAND3X1 _3562_ (
    .A(_1579_),
    .B(_1583_),
    .C(_1591_),
    .Y(_1592_)
);

FILL FILL_6__2423_ (
);

FILL FILL_6__2003_ (
);

NOR2X1 _3142_ (
    .A(_739_),
    .B(_746_),
    .Y(_747_)
);

FILL FILL_2__2835_ (
);

FILL FILL_2__2415_ (
);

FILL FILL_4__3702_ (
);

FILL FILL_6__3628_ (
);

FILL FILL_6__3208_ (
);

FILL FILL_0__3602_ (
);

FILL FILL_4__2094_ (
);

FILL FILL_3__2904_ (
);

FILL FILL169950x158550 (
);

FILL FILL_6_BUFX2_insert10 (
);

FILL FILL_6_BUFX2_insert11 (
);

FILL FILL_6_BUFX2_insert12 (
);

FILL FILL_6_BUFX2_insert13 (
);

FILL FILL_6_BUFX2_insert14 (
);

FILL FILL_6_BUFX2_insert15 (
);

FILL FILL_6_BUFX2_insert16 (
);

FILL FILL_6_BUFX2_insert17 (
);

FILL FILL_6_BUFX2_insert18 (
);

FILL FILL_6_BUFX2_insert19 (
);

FILL FILL_4__3299_ (
);

NOR2X1 _2833_ (
    .A(_494_),
    .B(_493_),
    .Y(_495_)
);

OAI21X1 _2413_ (
    .A(RDY_bF$buf5),
    .B(_1227_),
    .C(_1359_),
    .Y(_122_)
);

FILL FILL_1__1790_ (
);

FILL FILL_0__3199_ (
);

FILL FILL_5__2583_ (
);

FILL FILL_5__2163_ (
);

NAND2X1 _3618_ (
    .A(_1647_),
    .B(_1645_),
    .Y(_1648_)
);

FILL FILL_1__2995_ (
);

FILL FILL_1__2575_ (
);

FILL FILL_7__3542_ (
);

FILL FILL_1__2155_ (
);

FILL FILL_7__3122_ (
);

FILL FILL_3__3022_ (
);

FILL FILL_4__1785_ (
);

FILL FILL_6__2652_ (
);

FILL FILL_6__2232_ (
);

DFFSR _3371_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_48_),
    .CLK(clk_bF$buf10),
    .Q(src_reg[1])
);

FILL FILL_2__2644_ (
);

FILL FILL_2__2224_ (
);

FILL FILL_4__3511_ (
);

FILL FILL_6__3017_ (
);

FILL FILL_2__3009_ (
);

FILL FILL_5__1854_ (
);

FILL FILL_1__1846_ (
);

FILL FILL_3__2713_ (
);

FILL FILL_5__2639_ (
);

FILL FILL_5__2219_ (
);

FILL FILL_6__3190_ (
);

FILL FILL_2__3182_ (
);

FILL FILL_6__1923_ (
);

AOI21X1 _2642_ (
    .A(_901_),
    .B(_1221_),
    .C(_967_),
    .Y(_317_)
);

NOR2X1 _2222_ (
    .A(_1149__bF$buf3),
    .B(_1178_),
    .Y(_1330_)
);

FILL FILL_2__1915_ (
);

FILL FILL_5__2392_ (
);

FILL FILL_6__2708_ (
);

DFFSR _3427_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_95_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[3] [2])
);

INVX1 _3007_ (
    .A(load_reg),
    .Y(_633_)
);

FILL FILL_1__2384_ (
);

FILL FILL_3__3671_ (
);

FILL FILL_3__3251_ (
);

FILL FILL_5__3597_ (
);

FILL FILL_5__3177_ (
);

FILL FILL_1__3589_ (
);

FILL FILL_1__3169_ (
);

FILL FILL_6__2881_ (
);

FILL FILL_6__2461_ (
);

OAI21X1 _3180_ (
    .A(CO),
    .B(_728_),
    .C(_692_),
    .Y(_781_)
);

FILL FILL_6__2041_ (
);

FILL FILL_2__2873_ (
);

FILL FILL_2__2453_ (
);

FILL FILL_2__2033_ (
);

FILL FILL_4__2799_ (
);

FILL FILL_4__2379_ (
);

NOR2X1 _1913_ (
    .A(_913_),
    .B(_901_),
    .Y(_1030_)
);

FILL FILL_0__2699_ (
);

FILL FILL_6__3666_ (
);

FILL FILL_0__2279_ (
);

FILL FILL_6__3246_ (
);

FILL FILL_2__3658_ (
);

FILL FILL_0__3640_ (
);

FILL FILL_0__3220_ (
);

FILL FILL_2__3238_ (
);

FILL FILL_7__2622_ (
);

FILL FILL_3__2942_ (
);

FILL FILL_3__2522_ (
);

FILL FILL_3__2102_ (
);

FILL FILL_5__2868_ (
);

FILL FILL_5__2448_ (
);

FILL FILL_5__2028_ (
);

FILL FILL_3__3307_ (
);

OAI21X1 _2871_ (
    .A(_886__bF$buf5),
    .B(_1412_),
    .C(_527_),
    .Y(_20_)
);

FILL FILL169050x118950 (
);

OAI21X1 _2451_ (
    .A(_1319__bF$buf2),
    .B(_1263_),
    .C(PC[9]),
    .Y(_153_)
);

NAND3X1 _2031_ (
    .A(\AXYS[0] [7]),
    .B(_1051_),
    .C(_1053_),
    .Y(_1141_)
);

FILL FILL169650x144150 (
);

FILL FILL_6__2937_ (
);

NAND2X1 _3656_ (
    .A(ADD[0]),
    .B(_1714__bF$buf3),
    .Y(_1684_)
);

FILL FILL_6__2517_ (
);

OAI21X1 _3236_ (
    .A(_767_),
    .B(_807_),
    .C(_814_),
    .Y(_98_)
);

FILL FILL_7__3580_ (
);

FILL FILL_1__2193_ (
);

FILL FILL_0__2911_ (
);

FILL FILL_2__2929_ (
);

FILL FILL_2__2509_ (
);

FILL FILL_3__3480_ (
);

FILL FILL_3__3060_ (
);

FILL FILL_6__2690_ (
);

FILL FILL_6__2270_ (
);

FILL FILL_2__2682_ (
);

FILL FILL_2__2262_ (
);

FILL FILL_4__2188_ (
);

FILL FILL_6__3475_ (
);

FILL FILL_0__2088_ (
);

FILL FILL_6__3055_ (
);

FILL FILL_2__3467_ (
);

FILL FILL_2__3047_ (
);

FILL FILL_5__1892_ (
);

AOI22X1 _2927_ (
    .A(_132_),
    .B(_1149__bF$buf2),
    .C(_567_),
    .D(_570_),
    .Y(_33_)
);

NAND2X1 _2507_ (
    .A(_201_),
    .B(_194_),
    .Y(_202_)
);

FILL FILL_1__1884_ (
);

FILL FILL_7__2851_ (
);

FILL FILL_7__2011_ (
);

FILL FILL_3__2751_ (
);

FILL FILL_3__2331_ (
);

FILL FILL_5__2677_ (
);

FILL FILL_5__2257_ (
);

FILL FILL_1__2669_ (
);

FILL FILL_1__2249_ (
);

FILL FILL_1__3610_ (
);

FILL FILL_3__3536_ (
);

FILL FILL_3__3116_ (
);

FILL FILL_6__1961_ (
);

NAND3X1 _2680_ (
    .A(_1092_),
    .B(_328_),
    .C(_351_),
    .Y(_352_)
);

NAND3X1 _2260_ (
    .A(_1150__bF$buf0),
    .B(_1365_),
    .C(_1367_),
    .Y(_1368_)
);

FILL FILL_2__1953_ (
);

FILL FILL_4__1879_ (
);

FILL FILL_4__2820_ (
);

FILL FILL_4__2400_ (
);

FILL FILL_0__1779_ (
);

FILL FILL_6__2746_ (
);

OAI21X1 _3465_ (
    .A(_1704_),
    .B(_1705_),
    .C(_1712_),
    .Y(_1713_)
);

FILL FILL_6__2326_ (
);

INVX1 _3045_ (
    .A(_659_),
    .Y(_660_)
);

FILL FILL169650x39750 (
);

FILL FILL_2__2738_ (
);

FILL FILL_0__2720_ (
);

FILL FILL_2__2318_ (
);

FILL FILL_0__2300_ (
);

FILL FILL_4__3605_ (
);

FILL FILL_0__3505_ (
);

FILL FILL_5__1948_ (
);

FILL FILL_7__2907_ (
);

FILL FILL_2__2491_ (
);

FILL FILL_2__2071_ (
);

FILL FILL_3__2807_ (
);

INVX1 _1951_ (
    .A(_1067_),
    .Y(_1068_)
);

FILL FILL_6__3284_ (
);

FILL FILL_2__3696_ (
);

FILL FILL_2__3276_ (
);

AOI21X1 _2736_ (
    .A(_211_),
    .B(_321_),
    .C(_966_),
    .Y(_403_)
);

AND2X2 _2316_ (
    .A(_1231_),
    .B(_1229_),
    .Y(_1423_)
);

FILL FILL_7__2240_ (
);

FILL FILL_3__2980_ (
);

FILL FILL_3__2560_ (
);

FILL FILL_3__2140_ (
);

FILL FILL_5__2486_ (
);

FILL FILL_5__2066_ (
);

FILL FILL_1__2898_ (
);

FILL FILL_1__2478_ (
);

FILL FILL_1__2058_ (
);

FILL FILL_7__3025_ (
);

FILL FILL_6__1770_ (
);

FILL FILL_2__1762_ (
);

FILL FILL_6__2975_ (
);

BUFX2 _3694_ (
    .A(_1741_[11]),
    .Y(AB[11])
);

FILL FILL_6__2555_ (
);

OR2X2 _3274_ (
    .A(_846_),
    .B(_849_),
    .Y(_850_)
);

FILL FILL_6__2135_ (
);

FILL FILL_2__2967_ (
);

FILL FILL_2__2547_ (
);

FILL FILL_2__2127_ (
);

FILL FILL_3__1831_ (
);

FILL FILL_0__3314_ (
);

FILL FILL_5__1757_ (
);

FILL FILL_1__1749_ (
);

FILL FILL_7__2716_ (
);

FILL FILL_3__2616_ (
);

INVX1 _1760_ (
    .A(DIHOLD[5]),
    .Y(_889_)
);

FILL FILL_6__3093_ (
);

FILL FILL_2__3085_ (
);

FILL FILL_4__1900_ (
);

FILL FILL_6__1826_ (
);

OAI21X1 _2965_ (
    .A(_886__bF$buf4),
    .B(_1027__bF$buf1),
    .C(load_only),
    .Y(_599_)
);

OR2X2 _2545_ (
    .A(_209_),
    .B(_216_),
    .Y(_237_)
);

INVX1 _2125_ (
    .A(_1233_),
    .Y(_1234_)
);

FILL FILL_2__1818_ (
);

FILL FILL_0__1800_ (
);

FILL FILL_5__2295_ (
);

FILL FILL_7__3674_ (
);

FILL FILL_1__2287_ (
);

FILL FILL_7__3254_ (
);

FILL FILL_7_BUFX2_insert80 (
);

FILL FILL_7_BUFX2_insert82 (
);

FILL FILL_3__3574_ (
);

FILL FILL_7_BUFX2_insert83 (
);

FILL FILL_3__3154_ (
);

FILL FILL_2__1991_ (
);

FILL FILL_6__2784_ (
);

FILL FILL_6__2364_ (
);

AOI21X1 _3083_ (
    .A(_1227_),
    .B(_694_),
    .C(_691_),
    .Y(_695_)
);

FILL FILL_2__2776_ (
);

FILL FILL_2__2356_ (
);

INVX2 _1816_ (
    .A(_941_),
    .Y(_942_)
);

FILL FILL_4__3643_ (
);

FILL FILL_4__3223_ (
);

FILL FILL_6__3569_ (
);

FILL FILL_6__3149_ (
);

FILL FILL_0__3543_ (
);

FILL FILL_0__3123_ (
);

FILL FILL_5__1986_ (
);

FILL FILL_1__1978_ (
);

FILL FILL_7__2945_ (
);

FILL FILL_7__2525_ (
);

FILL FILL_7__2105_ (
);

FILL FILL_3__2845_ (
);

FILL FILL_3__2425_ (
);

FILL FILL_3__2005_ (
);

FILL FILL_5__3712_ (
);

FILL FILL_1__3704_ (
);

NOR2X1 _2774_ (
    .A(_438_),
    .B(_430_),
    .Y(_439_)
);

NOR2X1 _2354_ (
    .A(_1459_),
    .B(_1458_),
    .Y(_1460_)
);

FILL FILL_4__2914_ (
);

NAND2X1 _3559_ (
    .A(_1588_),
    .B(_1587_),
    .Y(_1589_)
);

NAND2X1 _3139_ (
    .A(\AXYS[0] [2]),
    .B(_722_),
    .Y(_745_)
);

FILL FILL_1__2096_ (
);

FILL FILL_0__2814_ (
);

FILL FILL_6__2593_ (
);

FILL FILL_6__2173_ (
);

FILL FILL_2__2585_ (
);

FILL FILL_2__2165_ (
);

FILL FILL_4__3452_ (
);

FILL FILL_4__3032_ (
);

FILL FILL_5__1795_ (
);

FILL FILL_1__1787_ (
);

FILL FILL_7__2754_ (
);

FILL FILL_3__2654_ (
);

FILL FILL_3__2234_ (
);

FILL FILL_5__3521_ (
);

FILL FILL_7__3119_ (
);

FILL FILL_5__3101_ (
);

FILL FILL_1__3513_ (
);

FILL FILL_3__3019_ (
);

FILL FILL_6__1864_ (
);

INVX2 _2583_ (
    .A(_196_),
    .Y(_270_)
);

INVX2 _2163_ (
    .A(_1031_),
    .Y(_1272_)
);

FILL FILL_2__1856_ (
);

FILL FILL_4__2723_ (
);

FILL FILL_4__2303_ (
);

FILL FILL_6__2649_ (
);

FILL FILL_6__2229_ (
);

DFFSR _3368_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_45_),
    .CLK(clk_bF$buf10),
    .Q(store)
);

FILL FILL_0__2623_ (
);

FILL FILL_0__2203_ (
);

FILL FILL_3__3192_ (
);

FILL FILL_4__3508_ (
);

FILL FILL_3__1925_ (
);

FILL FILL_2__2394_ (
);

OAI21X1 _1854_ (
    .A(_902__bF$buf0),
    .B(_974_),
    .C(_978_),
    .Y(_979_)
);

FILL FILL_4__3261_ (
);

FILL FILL_6__3187_ (
);

FILL FILL_0__3581_ (
);

FILL FILL_2__3599_ (
);

FILL FILL_0__3161_ (
);

FILL FILL_2__3179_ (
);

OAI21X1 _2639_ (
    .A(_913_),
    .B(_901_),
    .C(_1427_),
    .Y(_314_)
);

AND2X2 _2219_ (
    .A(_1171_),
    .B(_1167_),
    .Y(_1327_)
);

FILL FILL_7__2983_ (
);

FILL FILL_7__2143_ (
);

FILL FILL_3__2883_ (
);

FILL FILL_3__2463_ (
);

FILL FILL_3__2043_ (
);

FILL FILL_5__2389_ (
);

FILL FILL_3__3668_ (
);

FILL FILL_3__3248_ (
);

INVX1 _2392_ (
    .A(_1293_),
    .Y(_1497_)
);

FILL FILL_4__2952_ (
);

FILL FILL_4__2532_ (
);

FILL FILL_4__2112_ (
);

FILL FILL_6__2878_ (
);

OAI21X1 _3597_ (
    .A(_1725_),
    .B(alu_op[2]),
    .C(_1535_),
    .Y(_1627_)
);

FILL FILL_6__2458_ (
);

FILL FILL_6__2038_ (
);

NAND2X1 _3177_ (
    .A(\AXYS[0] [6]),
    .B(_722_),
    .Y(_779_)
);

FILL FILL_0__2852_ (
);

FILL FILL_0__2432_ (
);

FILL FILL_0__2012_ (
);

FILL FILL_7__1834_ (
);

FILL FILL_4__3317_ (
);

FILL FILL_0__3637_ (
);

FILL FILL_0__3217_ (
);

FILL FILL_5__2601_ (
);

FILL FILL_7__2619_ (
);

FILL FILL_3__2939_ (
);

FILL FILL_3__2519_ (
);

FILL FILL_4__3490_ (
);

FILL FILL_4__3070_ (
);

FILL FILL_4__1803_ (
);

NAND2X1 _2868_ (
    .A(RDY_bF$buf2),
    .B(_1181_),
    .Y(_526_)
);

NAND3X1 _2448_ (
    .A(_145_),
    .B(_146_),
    .C(_150_),
    .Y(_151_)
);

OAI21X1 _2028_ (
    .A(_1074_),
    .B(_1133_),
    .C(_1138_),
    .Y(AI[6])
);

FILL FILL_7__2372_ (
);

FILL FILL_3__2692_ (
);

FILL FILL_3__2272_ (
);

FILL FILL_5__2198_ (
);

FILL FILL_7__3577_ (
);

FILL FILL_7__3157_ (
);

FILL FILL_0__2908_ (
);

FILL FILL_1__3551_ (
);

FILL FILL_1__3131_ (
);

FILL FILL_3__3477_ (
);

FILL FILL_3__3057_ (
);

FILL FILL_2__1894_ (
);

FILL FILL_4__2761_ (
);

FILL FILL_4__2341_ (
);

FILL FILL_6__2687_ (
);

FILL FILL_6__2267_ (
);

FILL FILL_2__2679_ (
);

FILL FILL_0__2661_ (
);

FILL FILL_2__2259_ (
);

FILL FILL_0__2241_ (
);

FILL FILL_2__3620_ (
);

FILL FILL_2__3200_ (
);

FILL FILL_4__3546_ (
);

FILL FILL_4__3126_ (
);

FILL FILL_3__1963_ (
);

FILL FILL_0__3026_ (
);

FILL FILL_5__1889_ (
);

FILL FILL_7__2848_ (
);

FILL FILL_5__2830_ (
);

FILL FILL_5__2410_ (
);

FILL FILL_7__2008_ (
);

FILL FILL_1__2822_ (
);

FILL FILL_1__2402_ (
);

FILL FILL_3__2748_ (
);

FILL FILL_3__2328_ (
);

INVX2 _1892_ (
    .A(PC[5]),
    .Y(_1012_)
);

FILL FILL_5__3615_ (
);

FILL FILL_1__3607_ (
);

FILL FILL_6__1958_ (
);

OAI21X1 _2677_ (
    .A(_340_),
    .B(_349_),
    .C(RDY_bF$buf3),
    .Y(_350_)
);

NOR2X1 _2257_ (
    .A(_1160_),
    .B(_1173_),
    .Y(_1365_)
);

FILL FILL_0__1932_ (
);

FILL FILL_3__2081_ (
);

FILL FILL_4__2817_ (
);

FILL FILL_0__2717_ (
);

FILL FILL_3__3286_ (
);

FILL FILL_4__2990_ (
);

FILL FILL_4__2570_ (
);

FILL FILL_4__2150_ (
);

FILL FILL_6__2496_ (
);

FILL FILL_6__2076_ (
);

FILL FILL_0__2890_ (
);

FILL FILL_2__2488_ (
);

FILL FILL_0__2470_ (
);

FILL FILL_2__2068_ (
);

FILL FILL_0__2050_ (
);

NAND2X1 _1948_ (
    .A(_1064_),
    .B(_951_),
    .Y(_1065_)
);

FILL FILL_7__1872_ (
);

FILL FILL_0__3675_ (
);

FILL FILL_3__1772_ (
);

FILL FILL_0__3255_ (
);

FILL FILL_7__2237_ (
);

FILL FILL_1__2631_ (
);

FILL FILL_1__2211_ (
);

FILL FILL_3__2977_ (
);

FILL FILL_3__2557_ (
);

FILL FILL_3__2137_ (
);

FILL FILL_5__3004_ (
);

FILL FILL_4__1841_ (
);

FILL FILL_6__1767_ (
);

OAI21X1 _2486_ (
    .A(_1319__bF$buf0),
    .B(_1263_),
    .C(PC[14]),
    .Y(_183_)
);

NAND2X1 _2066_ (
    .A(_1161_),
    .B(_1174_),
    .Y(_1175_)
);

FILL FILL_2__1759_ (
);

FILL FILL_2__2700_ (
);

FILL FILL_4__2626_ (
);

FILL FILL_4__2206_ (
);

FILL FILL_0__2946_ (
);

FILL FILL_0__2526_ (
);

FILL FILL_0__2106_ (
);

FILL FILL_3__3095_ (
);

FILL FILL_5__1910_ (
);

FILL FILL_1__1902_ (
);

FILL FILL_3__1828_ (
);

FILL FILL_2__2297_ (
);

OR2X2 _1757_ (
    .A(RDY_bF$buf9),
    .B(DIHOLD[4]),
    .Y(_887_)
);

FILL FILL_4__3584_ (
);

FILL FILL_4__3164_ (
);

FILL FILL_0__3484_ (
);

FILL FILL_0__3064_ (
);

FILL FILL_7__2466_ (
);

FILL FILL_7__2046_ (
);

FILL FILL_1__2860_ (
);

FILL FILL_1__2440_ (
);

FILL FILL_1__2020_ (
);

FILL FILL_3__2786_ (
);

FILL FILL_3__2366_ (
);

FILL FILL_5__3653_ (
);

FILL FILL_5__3233_ (
);

FILL FILL_1__3645_ (
);

FILL FILL_1__3225_ (
);

FILL FILL_6__1996_ (
);

NOR2X1 _2295_ (
    .A(_1185_),
    .B(_1179_),
    .Y(_1402_)
);

FILL FILL_2__1988_ (
);

FILL FILL_0__1970_ (
);

FILL FILL_4__2855_ (
);

FILL FILL_4__2435_ (
);

FILL FILL_4__2015_ (
);

FILL FILL_0__2755_ (
);

FILL FILL_0__2335_ (
);

FILL FILL_6__3302_ (
);

FILL FILL_2__3714_ (
);

FILL FILL_5__2924_ (
);

FILL FILL_5__2504_ (
);

FILL FILL_1__2916_ (
);

INVX1 _1986_ (
    .A(_1100_),
    .Y(_1101_)
);

FILL FILL_5_BUFX2_insert0 (
);

FILL FILL_5_BUFX2_insert1 (
);

FILL FILL_5_BUFX2_insert2 (
);

FILL FILL_5_BUFX2_insert3 (
);

FILL FILL_5_BUFX2_insert4 (
);

FILL FILL_5_BUFX2_insert5 (
);

FILL FILL_5_BUFX2_insert6 (
);

FILL FILL_5_BUFX2_insert7 (
);

FILL FILL_5_BUFX2_insert8 (
);

FILL FILL_5_BUFX2_insert9 (
);

FILL FILL_5__3709_ (
);

FILL FILL_0__3293_ (
);

FILL FILL_7__2695_ (
);

FILL FILL_7__2275_ (
);

BUFX2 _3712_ (
    .A(_1742_[5]),
    .Y(DO[5])
);

FILL FILL_3__2595_ (
);

FILL FILL_3__2175_ (
);

FILL FILL_5__3462_ (
);

FILL FILL_5__3042_ (
);

FILL FILL168750x158550 (
);

FILL FILL_1__3454_ (
);

FILL FILL_1__3034_ (
);

FILL FILL_2__1797_ (
);

FILL FILL_4__2664_ (
);

FILL FILL_4__2244_ (
);

FILL FILL_0__2984_ (
);

FILL FILL_0__2564_ (
);

FILL FILL_6__3531_ (
);

FILL FILL_0__2144_ (
);

FILL FILL_6__3111_ (
);

FILL FILL_2__3523_ (
);

FILL FILL_2__3103_ (
);

FILL FILL_7__1966_ (
);

FILL FILL_4__3449_ (
);

FILL FILL_4__3029_ (
);

FILL FILL_1__1940_ (
);

FILL FILL_3__1866_ (
);

FILL FILL_5__2733_ (
);

FILL FILL_5__2313_ (
);

FILL FILL_1__2725_ (
);

FILL FILL_2_BUFX2_insert37 (
);

FILL FILL_2_BUFX2_insert38 (
);

FILL FILL_1__2305_ (
);

FILL FILL_2_BUFX2_insert39 (
);

INVX1 _1795_ (
    .A(compare),
    .Y(_921_)
);

FILL FILL_5__3518_ (
);

FILL FILL_4__1935_ (
);

FILL FILL_7__2084_ (
);

FILL FILL_0__1835_ (
);

FILL FILL_6__2802_ (
);

NAND3X1 _3521_ (
    .A(BI[2]),
    .B(AI[2]),
    .C(_1718_),
    .Y(_1551_)
);

AOI21X1 _3101_ (
    .A(plp),
    .B(ADD[0]),
    .C(_706_),
    .Y(_711_)
);

FILL FILL_5__3691_ (
);

FILL FILL_5__3271_ (
);

FILL FILL_1__3263_ (
);

FILL FILL_3__3189_ (
);

FILL FILL_4__2893_ (
);

FILL FILL_4__2473_ (
);

FILL FILL_4__2053_ (
);

FILL FILL_6__2399_ (
);

FILL FILL_0__2793_ (
);

FILL FILL_0__2373_ (
);

FILL FILL_4__3678_ (
);

FILL FILL_4__3258_ (
);

FILL FILL_0__3578_ (
);

FILL FILL_0__3158_ (
);

FILL FILL_5__2962_ (
);

FILL FILL_5__2542_ (
);

FILL FILL_5__2122_ (
);

FILL FILL_1__2954_ (
);

FILL FILL_1__2534_ (
);

FILL FILL_7__3501_ (
);

FILL FILL_1__2114_ (
);

FILL FILL_4__1744_ (
);

NAND3X1 _2389_ (
    .A(_1475_),
    .B(_1476_),
    .C(_1333_),
    .Y(_1494_)
);

FILL FILL_6__2611_ (
);

DFFSR _3330_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(_8_),
    .CLK(clk_bF$buf5),
    .Q(PC[6])
);

FILL FILL_2__2603_ (
);

FILL FILL_4__2949_ (
);

FILL FILL_4__2529_ (
);

FILL FILL_4__2109_ (
);

FILL FILL_5__3080_ (
);

FILL FILL_7__3098_ (
);

FILL FILL_0__2849_ (
);

FILL FILL_0__2429_ (
);

FILL FILL_0__2009_ (
);

FILL FILL_1__3492_ (
);

FILL FILL_1__3072_ (
);

FILL FILL_5__1813_ (
);

FILL FILL_1__1805_ (
);

FILL FILL168450x144150 (
);

FILL FILL_4__2282_ (
);

FILL FILL_0__2182_ (
);

FILL FILL_2__3561_ (
);

FILL FILL_2__3141_ (
);

FILL FILL_4__3487_ (
);

FILL FILL_4__3067_ (
);

INVX2 _2601_ (
    .A(PC[11]),
    .Y(_285_)
);

FILL FILL_5__2771_ (
);

FILL FILL_7__2369_ (
);

FILL FILL_5__2351_ (
);

FILL FILL_1__2763_ (
);

FILL FILL_1__2343_ (
);

FILL FILL_3__2689_ (
);

FILL FILL_3__2269_ (
);

FILL FILL_3__3630_ (
);

FILL FILL_3__3210_ (
);

FILL FILL_5__3556_ (
);

FILL FILL_5__3136_ (
);

FILL FILL_1__3548_ (
);

FILL FILL_1__3128_ (
);

FILL FILL_4__1973_ (
);

FILL FILL_6__1899_ (
);

OAI21X1 _2198_ (
    .A(_931__bF$buf4),
    .B(_949_),
    .C(RDY_bF$buf6),
    .Y(_1307_)
);

FILL FILL_0__1873_ (
);

FILL FILL_6__2840_ (
);

FILL FILL_6__2420_ (
);

FILL FILL_6__2000_ (
);

FILL FILL_2__2832_ (
);

FILL FILL_2__2412_ (
);

FILL FILL_4__2758_ (
);

FILL FILL_4__2338_ (
);

FILL FILL_0__2658_ (
);

FILL FILL_6__3625_ (
);

FILL FILL_0__2238_ (
);

FILL FILL_6__3205_ (
);

FILL FILL_2__3617_ (
);

FILL FILL_4__2091_ (
);

FILL FILL_3__2901_ (
);

FILL FILL_5__2827_ (
);

FILL FILL_5__2407_ (
);

FILL FILL_1__2819_ (
);

OAI22X1 _1889_ (
    .A(_1009_),
    .B(_968_),
    .C(_1010_),
    .D(_1004_),
    .Y(BI[3])
);

FILL FILL_4__3296_ (
);

NOR2X1 _2830_ (
    .A(_489_),
    .B(_491_),
    .Y(_492_)
);

NOR2X1 _2410_ (
    .A(_1237_),
    .B(_1339_),
    .Y(_119_)
);

FILL FILL_0__3196_ (
);

FILL FILL_7_BUFX2_insert0 (
);

FILL FILL_7_BUFX2_insert1 (
);

FILL FILL_7_BUFX2_insert3 (
);

FILL FILL_7_BUFX2_insert4 (
);

FILL FILL_7_BUFX2_insert6 (
);

FILL FILL_7_BUFX2_insert8 (
);

FILL FILL_7_BUFX2_insert9 (
);

FILL FILL_7__2598_ (
);

FILL FILL_5__2580_ (
);

FILL FILL_5__2160_ (
);

FILL FILL_0__1929_ (
);

OAI21X1 _3615_ (
    .A(_1644_),
    .B(_1643_),
    .C(_1640_),
    .Y(_1645_)
);

FILL FILL_1__2992_ (
);

FILL FILL_1__2572_ (
);

FILL FILL_1__2152_ (
);

FILL FILL_3__2498_ (
);

FILL FILL_3__2078_ (
);

FILL FILL_4__1782_ (
);

FILL FILL_2__2641_ (
);

FILL FILL_2__2221_ (
);

FILL FILL_4__2987_ (
);

FILL FILL_4__2567_ (
);

FILL FILL_4__2147_ (
);

FILL FILL_0__2887_ (
);

FILL FILL_0__2467_ (
);

FILL FILL_0__2047_ (
);

FILL FILL_6__3014_ (
);

FILL FILL_2__3006_ (
);

FILL FILL_7__1869_ (
);

FILL FILL_5__1851_ (
);

FILL FILL_1__1843_ (
);

FILL FILL_3__1769_ (
);

FILL FILL_3__2710_ (
);

FILL FILL_5__2636_ (
);

FILL FILL_5__2216_ (
);

FILL FILL_1__2628_ (
);

FILL FILL_1__2208_ (
);

FILL FILL_6__1920_ (
);

FILL FILL_2__1912_ (
);

FILL FILL_4__1838_ (
);

FILL FILL_6__2705_ (
);

DFFSR _3424_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_0_),
    .CLK(clk_bF$buf4),
    .Q(adj_bcd)
);

INVX1 _3004_ (
    .A(_621_),
    .Y(_631_)
);

FILL FILL_1__2381_ (
);

FILL FILL_5__3594_ (
);

FILL FILL_5__3174_ (
);

FILL FILL_1__3586_ (
);

FILL FILL_1__3166_ (
);

FILL FILL_5__1907_ (
);

FILL FILL_2__2870_ (
);

FILL FILL_2__2450_ (
);

FILL FILL_2__2030_ (
);

FILL FILL168150x32550 (
);

FILL FILL_4__2796_ (
);

FILL FILL_4__2376_ (
);

NAND3X1 _1910_ (
    .A(_927_),
    .B(_910_),
    .C(_929_),
    .Y(_1027_)
);

FILL FILL_0__2696_ (
);

FILL FILL_6__3663_ (
);

FILL FILL_0__2276_ (
);

FILL FILL_6__3243_ (
);

FILL FILL_2__3655_ (
);

FILL FILL_2__3235_ (
);

FILL FILL_3__1998_ (
);

FILL FILL_5__2865_ (
);

FILL FILL_5__2445_ (
);

FILL FILL_5__2025_ (
);

FILL FILL_1__2857_ (
);

FILL FILL_1__2437_ (
);

FILL FILL_1__2017_ (
);

FILL FILL_3__3304_ (
);

FILL FILL_0__1967_ (
);

FILL FILL_6__2934_ (
);

OAI21X1 _3653_ (
    .A(_1714__bF$buf2),
    .B(_1682_),
    .C(_1732_),
    .Y(_1515_)
);

FILL FILL_6__2514_ (
);

OAI21X1 _3233_ (
    .A(_720__bF$buf1),
    .B(_808_),
    .C(\AXYS[3] [4]),
    .Y(_813_)
);

FILL FILL_1__2190_ (
);

FILL FILL_2__2926_ (
);

FILL FILL_2__2506_ (
);

FILL FILL_4__2185_ (
);

FILL FILL_6__3472_ (
);

FILL FILL_0__2085_ (
);

FILL FILL_6__3052_ (
);

FILL FILL_2__3464_ (
);

FILL FILL_2__3044_ (
);

NAND2X1 _2924_ (
    .A(_1187_),
    .B(_1348_),
    .Y(_568_)
);

NOR2X1 _2504_ (
    .A(_196_),
    .B(_198_),
    .Y(_199_)
);

FILL FILL_1__1881_ (
);

FILL FILL_5__2674_ (
);

FILL FILL_5__2254_ (
);

BUFX2 _3709_ (
    .A(_1742_[2]),
    .Y(DO[2])
);

FILL FILL_1__2666_ (
);

FILL FILL_7__3633_ (
);

FILL FILL_1__2246_ (
);

FILL FILL_3__3533_ (
);

FILL FILL_3__3113_ (
);

FILL FILL_5__3459_ (
);

FILL FILL_5__3039_ (
);

FILL FILL_2__1950_ (
);

FILL FILL_4__1876_ (
);

FILL FILL_0__1776_ (
);

FILL FILL_6__2743_ (
);

INVX1 _3462_ (
    .A(_1709_),
    .Y(_1710_)
);

FILL FILL_6__2323_ (
);

OAI21X1 _3042_ (
    .A(_902__bF$buf1),
    .B(_954_),
    .C(_1027__bF$buf3),
    .Y(_657_)
);

FILL FILL_2__2735_ (
);

FILL FILL_2__2315_ (
);

FILL FILL_4__3602_ (
);

FILL FILL_6__3528_ (
);

FILL FILL_6__3108_ (
);

FILL FILL_0__3502_ (
);

FILL FILL_5__1945_ (
);

FILL FILL_1__1937_ (
);

FILL FILL_7__2904_ (
);

FILL FILL_3__2804_ (
);

FILL FILL_6__3281_ (
);

FILL FILL_2__3693_ (
);

FILL FILL_2__3273_ (
);

FILL FILL_4__3199_ (
);

NAND3X1 _2733_ (
    .A(_392_),
    .B(_399_),
    .C(_386_),
    .Y(_401_)
);

AOI21X1 _2313_ (
    .A(_1251_),
    .B(_1356_),
    .C(_1255_),
    .Y(_1420_)
);

FILL FILL_0__3099_ (
);

FILL FILL_5__2483_ (
);

FILL FILL_5__2063_ (
);

OAI21X1 _3518_ (
    .A(BI[3]),
    .B(_1739_),
    .C(_1547_),
    .Y(_1548_)
);

FILL FILL_1__2895_ (
);

FILL FILL_1__2475_ (
);

FILL FILL_1__2055_ (
);

FILL FILL_7__3022_ (
);

FILL FILL_5__3268_ (
);

FILL FILL_6__2972_ (
);

FILL FILL_6__2552_ (
);

BUFX2 _3691_ (
    .A(_1741_[0]),
    .Y(AB[0])
);

NOR2X1 _3271_ (
    .A(_1021_),
    .B(_1235_),
    .Y(_847_)
);

FILL FILL_6__2132_ (
);

FILL FILL_2__2964_ (
);

FILL FILL_2__2544_ (
);

FILL FILL_2__2124_ (
);

FILL FILL168450x75750 (
);

FILL FILL_0__3311_ (
);

FILL FILL_5__1754_ (
);

FILL FILL_1__1746_ (
);

FILL FILL_3__2613_ (
);

FILL FILL_5__2959_ (
);

FILL FILL_5__2539_ (
);

FILL FILL_5__2119_ (
);

FILL FILL_6__3090_ (
);

FILL FILL_2__3082_ (
);

FILL FILL_6__1823_ (
);

NAND3X1 _2962_ (
    .A(_1181_),
    .B(_543_),
    .C(_596_),
    .Y(_597_)
);

OAI21X1 _2542_ (
    .A(_1007_),
    .B(_218_),
    .C(_234_),
    .Y(_235_)
);

NOR2X1 _2122_ (
    .A(_886__bF$buf6),
    .B(_1205_),
    .Y(_1231_)
);

FILL FILL_2__1815_ (
);

FILL FILL_5__2292_ (
);

FILL FILL_6__2608_ (
);

DFFSR _3327_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(_5_),
    .CLK(clk_bF$buf3),
    .Q(PC[3])
);

FILL FILL_7__3671_ (
);

FILL FILL_1__2284_ (
);

FILL FILL_7__3251_ (
);

FILL FILL_7_BUFX2_insert50 (
);

FILL FILL_7_BUFX2_insert51 (
);

FILL FILL_3__3571_ (
);

FILL FILL_7_BUFX2_insert53 (
);

FILL FILL_3__3151_ (
);

FILL FILL_7_BUFX2_insert54 (
);

FILL FILL_7_BUFX2_insert56 (
);

FILL FILL_5__3497_ (
);

FILL FILL_7_BUFX2_insert58 (
);

FILL FILL_5__3077_ (
);

FILL FILL_7_BUFX2_insert59 (
);

FILL FILL_1__3489_ (
);

FILL FILL_1__3069_ (
);

FILL FILL169350x118950 (
);

FILL FILL_6__2781_ (
);

FILL FILL_6__2361_ (
);

INVX1 _3080_ (
    .A(AN),
    .Y(_692_)
);

FILL FILL169950x144150 (
);

FILL FILL_2__2773_ (
);

FILL FILL_2__2353_ (
);

FILL FILL_4__2699_ (
);

FILL FILL_4__2279_ (
);

INVX1 _1813_ (
    .A(_938_),
    .Y(_939_)
);

FILL FILL_4__3640_ (
);

FILL FILL_4__3220_ (
);

FILL FILL_0__2599_ (
);

FILL FILL_6__3566_ (
);

FILL FILL_0__2179_ (
);

FILL FILL_6__3146_ (
);

FILL FILL_0__3540_ (
);

FILL FILL_2__3558_ (
);

FILL FILL_0__3120_ (
);

FILL FILL_2__3138_ (
);

FILL FILL_5__1983_ (
);

FILL FILL_1__1975_ (
);

FILL FILL_7__2522_ (
);

FILL FILL_3__2842_ (
);

FILL FILL_3__2422_ (
);

FILL FILL_3__2002_ (
);

FILL FILL_5__2768_ (
);

FILL FILL_5__2348_ (
);

FILL FILL_7__3307_ (
);

FILL FILL_1__3701_ (
);

FILL FILL_3__3627_ (
);

FILL FILL_3__3207_ (
);

AND2X2 _2771_ (
    .A(_434_),
    .B(_435_),
    .Y(_436_)
);

INVX1 _2351_ (
    .A(_1401_),
    .Y(_1457_)
);

FILL FILL_4__2911_ (
);

FILL FILL_6__2837_ (
);

NOR2X1 _3556_ (
    .A(alu_shift_right),
    .B(_1585_),
    .Y(_1586_)
);

FILL FILL_6__2417_ (
);

OAI21X1 _3136_ (
    .A(_732_),
    .B(_741_),
    .C(_1018_),
    .Y(_742_)
);

FILL FILL_7__3480_ (
);

FILL FILL_1__2093_ (
);

FILL FILL_0__2811_ (
);

FILL FILL_2__2829_ (
);

FILL FILL_2__2409_ (
);

FILL FILL_1__3298_ (
);

FILL FILL_6__2590_ (
);

FILL FILL_6__2170_ (
);

FILL FILL_2__2582_ (
);

FILL FILL_2__2162_ (
);

FILL FILL_4__2088_ (
);

FILL FILL_5__1792_ (
);

OAI21X1 _2827_ (
    .A(_295_),
    .B(_313_),
    .C(_1126_),
    .Y(_489_)
);

AND2X2 _2407_ (
    .A(_1510_),
    .B(_1463_),
    .Y(_1511_)
);

FILL FILL_1__1784_ (
);

FILL FILL_7__2751_ (
);

FILL FILL_3__2651_ (
);

FILL FILL_3__2231_ (
);

FILL FILL_5__2997_ (
);

FILL FILL_5__2577_ (
);

FILL FILL_5__2157_ (
);

FILL FILL_1__2989_ (
);

FILL FILL_1__2569_ (
);

FILL FILL_1__2149_ (
);

FILL FILL_1__3510_ (
);

FILL FILL_3__3016_ (
);

FILL FILL_6__1861_ (
);

INVX1 _2580_ (
    .A(_267_),
    .Y(_1741_[7])
);

NAND2X1 _2160_ (
    .A(RDY_bF$buf6),
    .B(_1268_),
    .Y(_1269_)
);

FILL FILL_2__1853_ (
);

FILL FILL_4__1779_ (
);

FILL FILL_4__2720_ (
);

FILL FILL_4__2300_ (
);

FILL FILL_6__2646_ (
);

FILL FILL_6__2226_ (
);

DFFSR _3365_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_42_),
    .CLK(clk_bF$buf10),
    .Q(inc)
);

FILL FILL_2__2638_ (
);

FILL FILL_0__2620_ (
);

FILL FILL_0__2200_ (
);

FILL FILL_2__2218_ (
);

FILL FILL_4__3505_ (
);

FILL FILL_3__1922_ (
);

FILL FILL_5__1848_ (
);

FILL FILL_2__2391_ (
);

FILL FILL_3__2707_ (
);

NAND2X1 _1851_ (
    .A(state[0]),
    .B(_905_),
    .Y(_976_)
);

FILL FILL_6__3184_ (
);

FILL FILL_2__3596_ (
);

FILL FILL_2__3176_ (
);

FILL FILL_6__1917_ (
);

OAI21X1 _2636_ (
    .A(_914__bF$buf2),
    .B(_942_),
    .C(_1470_),
    .Y(_311_)
);

NOR2X1 _2216_ (
    .A(_1280_),
    .B(_1324_),
    .Y(_1325_)
);

FILL FILL_7__2980_ (
);

FILL FILL_7__2140_ (
);

FILL FILL_2__1909_ (
);

FILL FILL_3__2880_ (
);

FILL FILL_3__2460_ (
);

FILL FILL_3__2040_ (
);

FILL FILL_5__2386_ (
);

FILL FILL_1__2798_ (
);

FILL FILL_1__2378_ (
);

FILL FILL_3__3665_ (
);

FILL FILL_3__3245_ (
);

FILL FILL_6__2875_ (
);

AOI21X1 _3594_ (
    .A(_1620_),
    .B(_1623_),
    .C(_1608_),
    .Y(_1624_)
);

FILL FILL_6__2455_ (
);

FILL FILL_6__2035_ (
);

OAI21X1 _3174_ (
    .A(_765_),
    .B(_772_),
    .C(_775_),
    .Y(_776_)
);

FILL FILL_2__2867_ (
);

FILL FILL_2__2447_ (
);

FILL FILL_2__2027_ (
);

NAND2X1 _1907_ (
    .A(_901_),
    .B(_993_),
    .Y(_1024_)
);

FILL FILL_4__3314_ (
);

FILL FILL_0__3634_ (
);

FILL FILL_0__3214_ (
);

FILL FILL_7__2616_ (
);

FILL FILL_3__2936_ (
);

FILL FILL_3__2516_ (
);

FILL FILL_4__1800_ (
);

INVX1 _2865_ (
    .A(NMI_1),
    .Y(_524_)
);

NAND2X1 _2445_ (
    .A(_929_),
    .B(_935_),
    .Y(_148_)
);

INVX1 _2025_ (
    .A(_1135_),
    .Y(_1136_)
);

FILL FILL_5__2195_ (
);

FILL FILL_7__3574_ (
);

FILL FILL_1__2187_ (
);

FILL FILL_7__3154_ (
);

FILL FILL_0__2905_ (
);

FILL FILL_3__3474_ (
);

FILL FILL_3__3054_ (
);

FILL FILL_2__1891_ (
);

FILL FILL_6__2684_ (
);

FILL FILL_6__2264_ (
);

FILL FILL_2__2676_ (
);

FILL FILL_2__2256_ (
);

FILL FILL_4__3543_ (
);

FILL FILL_4__3123_ (
);

FILL FILL_6__3469_ (
);

FILL FILL_6__3049_ (
);

FILL FILL_3__1960_ (
);

FILL FILL_0__3023_ (
);

FILL FILL_5__1886_ (
);

FILL FILL_1__1878_ (
);

FILL FILL_7__2845_ (
);

FILL FILL_7__2425_ (
);

FILL FILL_7__2005_ (
);

FILL FILL_3__2745_ (
);

FILL FILL_3__2325_ (
);

FILL FILL_5__3612_ (
);

FILL FILL_1__3604_ (
);

FILL FILL_6__1955_ (
);

OAI21X1 _2674_ (
    .A(_1007_),
    .B(_330_),
    .C(_346_),
    .Y(_347_)
);

NAND2X1 _2254_ (
    .A(_1284_),
    .B(_1332_),
    .Y(_1362_)
);

FILL FILL_2__1947_ (
);

FILL FILL_4__2814_ (
);

INVX1 _3459_ (
    .A(AN),
    .Y(_1707_)
);

OAI21X1 _3039_ (
    .A(_893_),
    .B(_647_),
    .C(_655_),
    .Y(_60_)
);

FILL FILL_0__2714_ (
);

FILL FILL_3__3283_ (
);

FILL FILL_6__2493_ (
);

FILL FILL_6__2073_ (
);

FILL FILL_2__2485_ (
);

FILL FILL_2__2065_ (
);

INVX1 _1945_ (
    .A(_1061_),
    .Y(_1062_)
);

FILL FILL_6__3698_ (
);

FILL FILL_6__3278_ (
);

FILL FILL_0__3672_ (
);

FILL FILL_0__3252_ (
);

FILL FILL_7__2654_ (
);

FILL FILL_7__2234_ (
);

FILL FILL_3__2974_ (
);

FILL FILL_3__2554_ (
);

FILL FILL_3__2134_ (
);

FILL FILL_7__3019_ (
);

FILL FILL_5__3001_ (
);

FILL FILL_6__1764_ (
);

OAI21X1 _2483_ (
    .A(_179_),
    .B(_174_),
    .C(_180_),
    .Y(_181_)
);

NAND2X1 _2063_ (
    .A(_1167_),
    .B(_1171_),
    .Y(_1172_)
);

FILL FILL_2__1756_ (
);

FILL FILL_4__2623_ (
);

FILL FILL_4__2203_ (
);

FILL FILL_6__2969_ (
);

DFFSR _3688_ (
    .R(_1513_),
    .S(vdd),
    .D(_1523_),
    .CLK(clk_bF$buf3),
    .Q(ADD[6])
);

FILL FILL_6__2549_ (
);

OAI21X1 _3268_ (
    .A(_977_),
    .B(_1427_),
    .C(_929_),
    .Y(_844_)
);

FILL FILL_6__2129_ (
);

FILL FILL_0__2943_ (
);

FILL FILL_0__2523_ (
);

FILL FILL_0__2103_ (
);

FILL FILL_3__3092_ (
);

FILL FILL_3__1825_ (
);

FILL FILL_0__3308_ (
);

FILL FILL_2__2294_ (
);

NAND2X1 _1754_ (
    .A(RDY_bF$buf9),
    .B(DI[3]),
    .Y(_885_)
);

FILL FILL_4__3581_ (
);

FILL FILL_4__3161_ (
);

FILL FILL_6__3087_ (
);

FILL FILL_2__3499_ (
);

FILL FILL_0__3481_ (
);

FILL FILL_2__3079_ (
);

FILL FILL_0__3061_ (
);

OAI22X1 _2959_ (
    .A(_309_),
    .B(_593_),
    .C(_594_),
    .D(_595_),
    .Y(_40_)
);

OAI21X1 _2539_ (
    .A(_216_),
    .B(_209_),
    .C(ADD[2]),
    .Y(_232_)
);

NAND3X1 _2119_ (
    .A(_1227_),
    .B(_1224_),
    .C(_1226_),
    .Y(_1228_)
);

FILL FILL_7__2883_ (
);

FILL FILL_7__2043_ (
);

FILL FILL_3__2783_ (
);

FILL FILL_3__2363_ (
);

FILL FILL_5__2289_ (
);

FILL FILL_5__3650_ (
);

FILL FILL_5__3230_ (
);

FILL FILL_7__3248_ (
);

FILL FILL_1__3642_ (
);

FILL FILL_1__3222_ (
);

FILL FILL_3__3568_ (
);

FILL FILL_3__3148_ (
);

FILL FILL_6__1993_ (
);

OAI21X1 _2292_ (
    .A(_1213_),
    .B(_1215_),
    .C(_1328_),
    .Y(_1399_)
);

FILL FILL_2__1985_ (
);

FILL FILL_4__2852_ (
);

FILL FILL_4__2432_ (
);

FILL FILL_4__2012_ (
);

FILL FILL_6__2778_ (
);

OAI21X1 _3497_ (
    .A(BI[5]),
    .B(_1739_),
    .C(_1526_),
    .Y(_1527_)
);

FILL FILL_6__2358_ (
);

AOI21X1 _3077_ (
    .A(_687_),
    .B(load_reg),
    .C(_688_),
    .Y(_689_)
);

FILL FILL_0__2752_ (
);

FILL FILL_0__2332_ (
);

FILL FILL_2__3711_ (
);

FILL FILL_4__3637_ (
);

FILL FILL_4__3217_ (
);

FILL FILL_0__3537_ (
);

FILL FILL_0__3117_ (
);

FILL FILL_5__2921_ (
);

FILL FILL_7__2519_ (
);

FILL FILL_5__2501_ (
);

FILL FILL_1__2913_ (
);

FILL FILL_3__2839_ (
);

FILL FILL_3__2419_ (
);

AOI22X1 _1983_ (
    .A(_1049_),
    .B(\AXYS[3] [2]),
    .C(\AXYS[2] [2]),
    .D(_1057_),
    .Y(_1098_)
);

FILL FILL_5__3706_ (
);

FILL FILL_0__3290_ (
);

AOI21X1 _2768_ (
    .A(ABH[2]),
    .B(_323_),
    .C(_432_),
    .Y(_433_)
);

NAND3X1 _2348_ (
    .A(_1308_),
    .B(_1256_),
    .C(_1302_),
    .Y(_1455_)
);

FILL FILL_7__2272_ (
);

FILL FILL_3__2592_ (
);

FILL FILL_3__2172_ (
);

FILL FILL_5__2098_ (
);

FILL FILL_4__2908_ (
);

FILL FILL_7__3477_ (
);

FILL FILL_7__3057_ (
);

FILL FILL_0__2808_ (
);

FILL FILL_1__3451_ (
);

FILL FILL_1__3031_ (
);

FILL FILL_2__1794_ (
);

FILL FILL_4__2661_ (
);

FILL FILL_4__2241_ (
);

FILL FILL_6__2587_ (
);

FILL FILL_6__2167_ (
);

FILL FILL_2__2999_ (
);

FILL FILL_0__2981_ (
);

FILL FILL_0__2561_ (
);

FILL FILL_2__2579_ (
);

FILL FILL_2__2159_ (
);

FILL FILL_0__2141_ (
);

FILL FILL_2__3520_ (
);

FILL FILL_2__3100_ (
);

FILL FILL_7__1963_ (
);

FILL FILL_4__3026_ (
);

FILL FILL_3__1863_ (
);

FILL FILL_5__1789_ (
);

FILL FILL_7__2748_ (
);

FILL FILL_5__2730_ (
);

FILL FILL_5__2310_ (
);

FILL FILL_1__2722_ (
);

FILL FILL_1__2302_ (
);

FILL FILL_3__2648_ (
);

FILL FILL_3__2228_ (
);

NOR2X1 _1792_ (
    .A(load_only),
    .B(_917_),
    .Y(_918_)
);

FILL FILL_5__3515_ (
);

FILL FILL_1__3507_ (
);

FILL FILL_4__1932_ (
);

FILL FILL_6__1858_ (
);

OAI21X1 _2997_ (
    .A(_1327_),
    .B(_1178_),
    .C(_1161_),
    .Y(_625_)
);

AND2X2 _2577_ (
    .A(_263_),
    .B(_264_),
    .Y(_265_)
);

NAND3X1 _2157_ (
    .A(_1262_),
    .B(_1265_),
    .C(_1259_),
    .Y(_1266_)
);

FILL FILL_0__1832_ (
);

FILL FILL_4__2717_ (
);

FILL FILL_7__3286_ (
);

FILL FILL_0__2617_ (
);

FILL FILL_1__3260_ (
);

FILL FILL_3__3186_ (
);

FILL FILL_3__1919_ (
);

FILL FILL_4__2890_ (
);

FILL FILL_4__2470_ (
);

FILL FILL_4__2050_ (
);

FILL FILL_6__2396_ (
);

FILL FILL_0__2790_ (
);

FILL FILL_0__2370_ (
);

FILL FILL_2__2388_ (
);

NOR2X1 _1848_ (
    .A(state[2]),
    .B(state[3]),
    .Y(_973_)
);

FILL FILL_4__3675_ (
);

FILL FILL_7__1772_ (
);

FILL FILL_4__3255_ (
);

FILL FILL_0__3575_ (
);

FILL FILL_0__3155_ (
);

FILL FILL_7__2977_ (
);

FILL FILL_7__2137_ (
);

FILL FILL_1__2951_ (
);

FILL FILL_1__2531_ (
);

FILL FILL_1__2111_ (
);

FILL FILL_3__2877_ (
);

FILL FILL_3__2457_ (
);

FILL FILL_3__2037_ (
);

FILL FILL_1__3316_ (
);

NAND3X1 _2386_ (
    .A(_1485_),
    .B(_1486_),
    .C(_1491_),
    .Y(_1492_)
);

FILL FILL_2__2600_ (
);

FILL FILL_4__2946_ (
);

FILL FILL_4__2526_ (
);

FILL FILL_4__2106_ (
);

FILL FILL_7__3095_ (
);

FILL FILL_0__2846_ (
);

FILL FILL_0__2426_ (
);

FILL FILL_0__2006_ (
);

FILL FILL_5__1810_ (
);

FILL FILL_1__1802_ (
);

FILL FILL_2__2197_ (
);

FILL FILL_4__3484_ (
);

FILL FILL_4__3064_ (
);

FILL FILL_7__2366_ (
);

FILL FILL_1__2760_ (
);

FILL FILL_1__2340_ (
);

FILL FILL_3__2686_ (
);

FILL FILL_3__2266_ (
);

FILL FILL_5__3553_ (
);

FILL FILL_5__3133_ (
);

FILL FILL_1__3545_ (
);

FILL FILL_1__3125_ (
);

FILL FILL_4__1970_ (
);

FILL FILL_6__1896_ (
);

INVX1 _2195_ (
    .A(_1303_),
    .Y(_1304_)
);

FILL FILL_2__1888_ (
);

FILL FILL_0__1870_ (
);

FILL FILL_4__2755_ (
);

FILL FILL_4__2335_ (
);

FILL FILL_0__2655_ (
);

FILL FILL_6__3622_ (
);

FILL FILL_0__2235_ (
);

FILL FILL_6__3202_ (
);

FILL FILL_2__3614_ (
);

FILL FILL_3__1957_ (
);

FILL FILL_5__2824_ (
);

FILL FILL_5__2404_ (
);

FILL FILL_1__2816_ (
);

OAI22X1 _1886_ (
    .A(_1007_),
    .B(_968_),
    .C(_1008_),
    .D(_1004_),
    .Y(BI[2])
);

FILL FILL_4__3293_ (
);

FILL FILL_5__3609_ (
);

FILL FILL_0__3193_ (
);

FILL FILL_7__2595_ (
);

FILL FILL_7__2175_ (
);

FILL FILL_0__1926_ (
);

NAND2X1 _3612_ (
    .A(AI[6]),
    .B(_1641_),
    .Y(_1642_)
);

FILL FILL_3__2495_ (
);

FILL FILL_3__2075_ (
);

FILL FILL_4__2984_ (
);

FILL FILL_4__2564_ (
);

FILL FILL_4__2144_ (
);

FILL FILL_0__2884_ (
);

FILL FILL_0__2464_ (
);

FILL FILL_0__2044_ (
);

FILL FILL_6__3011_ (
);

FILL FILL_2__3003_ (
);

FILL FILL_7__1866_ (
);

FILL FILL_1__1840_ (
);

FILL FILL_0__3669_ (
);

FILL FILL_3__1766_ (
);

FILL FILL_0__3249_ (
);

FILL FILL_5__2633_ (
);

FILL FILL_5__2213_ (
);

FILL FILL_1__2625_ (
);

FILL FILL_1__2205_ (
);

FILL FILL_4__1835_ (
);

FILL FILL_6__2702_ (
);

DFFSR _3421_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_90_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[2] [5])
);

OAI21X1 _3001_ (
    .A(_1042_),
    .B(_1150__bF$buf4),
    .C(_628_),
    .Y(_49_)
);

FILL FILL_5__3591_ (
);

FILL FILL_5__3171_ (
);

FILL FILL_1__3583_ (
);

FILL FILL_1__3163_ (
);

FILL FILL_3__3089_ (
);

FILL FILL_5__1904_ (
);

FILL FILL_4__2793_ (
);

FILL FILL_4__2373_ (
);

FILL FILL_6__2299_ (
);

FILL FILL_0__2693_ (
);

FILL FILL_6__3660_ (
);

FILL FILL_0__2273_ (
);

FILL FILL_6__3240_ (
);

FILL FILL_2__3652_ (
);

FILL FILL_2__3232_ (
);

FILL FILL_4__3578_ (
);

FILL FILL_4__3158_ (
);

FILL FILL_3__1995_ (
);

FILL FILL_0__3478_ (
);

FILL FILL_0__3058_ (
);

FILL FILL_5__2862_ (
);

FILL FILL_5__2442_ (
);

FILL FILL_5__2022_ (
);

FILL FILL168750x144150 (
);

FILL FILL_1__2854_ (
);

FILL FILL_1__2434_ (
);

FILL FILL_1__2014_ (
);

FILL FILL_3__3301_ (
);

FILL FILL_5__3647_ (
);

FILL FILL_5__3227_ (
);

FILL FILL_1__3639_ (
);

FILL FILL_1__3219_ (
);

INVX1 _2289_ (
    .A(_1395_),
    .Y(_1396_)
);

FILL FILL_0__1964_ (
);

FILL FILL_6__2931_ (
);

NAND2X1 _3650_ (
    .A(_1679_),
    .B(_1673_),
    .Y(_1680_)
);

FILL FILL_6__2511_ (
);

OAI21X1 _3230_ (
    .A(_744_),
    .B(_807_),
    .C(_811_),
    .Y(_95_)
);

FILL FILL_3_BUFX2_insert70 (
);

FILL FILL_3_BUFX2_insert71 (
);

FILL FILL_3_BUFX2_insert72 (
);

FILL FILL_2__2923_ (
);

FILL FILL_3_BUFX2_insert73 (
);

FILL FILL_2__2503_ (
);

FILL FILL_3_BUFX2_insert74 (
);

FILL FILL_3_BUFX2_insert75 (
);

FILL FILL_3_BUFX2_insert76 (
);

FILL FILL_3_BUFX2_insert77 (
);

FILL FILL_4__2849_ (
);

FILL FILL_3_BUFX2_insert78 (
);

FILL FILL_4__2429_ (
);

FILL FILL_3_BUFX2_insert79 (
);

FILL FILL_4__2009_ (
);

FILL FILL_0__2749_ (
);

FILL FILL_0__2329_ (
);

FILL FILL_2__3708_ (
);

FILL FILL_4__2182_ (
);

FILL FILL_5__2918_ (
);

FILL FILL_0__2082_ (
);

FILL FILL_2__3461_ (
);

FILL FILL_2__3041_ (
);

NOR2X1 _2921_ (
    .A(_556_),
    .B(_561_),
    .Y(_566_)
);

OAI21X1 _2501_ (
    .A(_902__bF$buf1),
    .B(_949_),
    .C(_909_),
    .Y(_196_)
);

FILL FILL_0__3287_ (
);

FILL FILL_5__2671_ (
);

FILL FILL_7__2269_ (
);

FILL FILL_5__2251_ (
);

BUFX2 _3706_ (
    .A(_1741_[9]),
    .Y(AB[9])
);

FILL FILL_1__2663_ (
);

FILL FILL_7__3630_ (
);

FILL FILL_1__2243_ (
);

FILL FILL_3__2589_ (
);

FILL FILL_3__2169_ (
);

FILL FILL_3__3530_ (
);

FILL FILL_3__3110_ (
);

FILL FILL_5__3456_ (
);

FILL FILL_5__3036_ (
);

FILL FILL_1__3028_ (
);

FILL FILL_4__1873_ (
);

FILL FILL_6__1799_ (
);

INVX1 _2098_ (
    .A(write_back),
    .Y(_1207_)
);

FILL FILL_0__1773_ (
);

FILL FILL_6__2740_ (
);

FILL FILL_6__2320_ (
);

FILL FILL_2__2732_ (
);

FILL FILL_2__2312_ (
);

FILL FILL_4__2658_ (
);

FILL FILL_4__2238_ (
);

FILL FILL_0__2978_ (
);

FILL FILL_0__2558_ (
);

FILL FILL_6__3525_ (
);

FILL FILL_0__2138_ (
);

FILL FILL_6__3105_ (
);

FILL FILL_2__3517_ (
);

FILL FILL_5__1942_ (
);

FILL FILL_1__1934_ (
);

FILL FILL_7__2901_ (
);

FILL FILL_3__2801_ (
);

FILL FILL_5__2727_ (
);

FILL FILL_5__2307_ (
);

FILL FILL_1__2719_ (
);

FILL FILL_2__3270_ (
);

OAI21X1 _1789_ (
    .A(_912_),
    .B(_914__bF$buf2),
    .C(_909_),
    .Y(_915_)
);

FILL FILL_4__3196_ (
);

AOI21X1 _2730_ (
    .A(_322_),
    .B(AN),
    .C(_397_),
    .Y(_398_)
);

OAI21X1 _2310_ (
    .A(_1172_),
    .B(_1212_),
    .C(_1150__bF$buf0),
    .Y(_1417_)
);

FILL FILL_0__3096_ (
);

FILL FILL_4__1929_ (
);

FILL FILL_5__2480_ (
);

FILL FILL_7__2498_ (
);

FILL FILL_5__2060_ (
);

FILL FILL_0__1829_ (
);

OAI21X1 _3515_ (
    .A(_1722_),
    .B(_1537_),
    .C(_1544_),
    .Y(_1545_)
);

FILL FILL_1__2892_ (
);

FILL FILL_1__2472_ (
);

FILL FILL_1__2052_ (
);

FILL FILL_3__2398_ (
);

FILL FILL_5__3265_ (
);

FILL FILL_1__3677_ (
);

FILL FILL_1__3257_ (
);

FILL FILL_2__2961_ (
);

FILL FILL_2__2541_ (
);

FILL FILL_2__2121_ (
);

FILL FILL_4__2887_ (
);

FILL FILL_4__2467_ (
);

FILL FILL_4__2047_ (
);

FILL FILL_0__2787_ (
);

FILL FILL_0__2367_ (
);

FILL FILL_5__1751_ (
);

FILL FILL_7__1769_ (
);

FILL FILL_3__2610_ (
);

FILL FILL_5__2956_ (
);

FILL FILL_5__2536_ (
);

FILL FILL_5__2116_ (
);

FILL FILL_1__2948_ (
);

FILL FILL_1__2528_ (
);

FILL FILL_1__2108_ (
);

FILL FILL_6__1820_ (
);

FILL FILL_2__1812_ (
);

FILL FILL_6__2605_ (
);

DFFSR _3324_ (
    .R(_1__bF$buf7),
    .S(vdd),
    .D(_2_),
    .CLK(clk_bF$buf3),
    .Q(PC[0])
);

FILL FILL_1__2281_ (
);

FILL FILL_7_BUFX2_insert21 (
);

FILL FILL_7_BUFX2_insert22 (
);

FILL FILL_7_BUFX2_insert24 (
);

FILL FILL_7_BUFX2_insert25 (
);

FILL FILL_5__3494_ (
);

FILL FILL_5__3074_ (
);

FILL FILL_1__3486_ (
);

FILL FILL_1__3066_ (
);

FILL FILL_5__1807_ (
);

FILL FILL_2__2770_ (
);

FILL FILL_2__2350_ (
);

FILL FILL_4__2696_ (
);

FILL FILL_4__2276_ (
);

NAND2X1 _1810_ (
    .A(_903__bF$buf3),
    .B(_935_),
    .Y(_936_)
);

FILL FILL_0__2596_ (
);

FILL FILL_6__3563_ (
);

FILL FILL_0__2176_ (
);

FILL FILL_6__3143_ (
);

FILL FILL_2__3555_ (
);

FILL FILL_2__3135_ (
);

FILL FILL_5__1980_ (
);

FILL FILL_7__1998_ (
);

FILL FILL_1__1972_ (
);

FILL FILL_3__1898_ (
);

FILL FILL_5__2765_ (
);

FILL FILL_5__2345_ (
);

FILL FILL_1__2757_ (
);

FILL FILL_1__2337_ (
);

FILL FILL_7__3304_ (
);

FILL FILL_3__3624_ (
);

FILL FILL_3__3204_ (
);

FILL FILL169950x165750 (
);

FILL FILL_4__1967_ (
);

FILL FILL_0__1867_ (
);

FILL FILL_6__2834_ (
);

OAI21X1 _3553_ (
    .A(_1740_),
    .B(_1575_),
    .C(_1582_),
    .Y(_1583_)
);

FILL FILL_6__2414_ (
);

NOR2X1 _3133_ (
    .A(_431_),
    .B(_727_),
    .Y(_739_)
);

FILL FILL_1__2090_ (
);

FILL FILL_2__2826_ (
);

FILL FILL_2__2406_ (
);

FILL FILL_6__3619_ (
);

FILL FILL_1__3295_ (
);

FILL FILL_4__2085_ (
);

AND2X2 _2824_ (
    .A(_467_),
    .B(_486_),
    .Y(_487_)
);

INVX1 _2404_ (
    .A(_1478_),
    .Y(_1508_)
);

FILL FILL_1__1781_ (
);

FILL FILL_5__2994_ (
);

FILL FILL_5__2574_ (
);

FILL FILL_5__2154_ (
);

INVX1 _3609_ (
    .A(_1638_),
    .Y(_1639_)
);

FILL FILL_1__2986_ (
);

FILL FILL_1__2566_ (
);

FILL FILL_7__3533_ (
);

FILL FILL_1__2146_ (
);

FILL FILL_3__3013_ (
);

FILL FILL_2__1850_ (
);

FILL FILL_4__1776_ (
);

FILL FILL_6__2643_ (
);

DFFSR _3362_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_39_),
    .CLK(clk_bF$buf10),
    .Q(shift)
);

FILL FILL_6__2223_ (
);

FILL FILL_2__2635_ (
);

FILL FILL_2__2215_ (
);

FILL FILL_4__3502_ (
);

FILL FILL_6__3008_ (
);

FILL FILL_5__1845_ (
);

FILL FILL_1__1837_ (
);

FILL FILL_7__2804_ (
);

FILL FILL_3__2704_ (
);

FILL FILL_6__3181_ (
);

FILL FILL_2__3593_ (
);

FILL FILL_2__3173_ (
);

FILL FILL_4__3099_ (
);

FILL FILL_6__1914_ (
);

INVX1 _2633_ (
    .A(shift_right),
    .Y(_310_)
);

NAND3X1 _2213_ (
    .A(_1314_),
    .B(_1321_),
    .C(_1318_),
    .Y(_1322_)
);

FILL FILL_2__1906_ (
);

FILL FILL_5__2383_ (
);

DFFSR _3418_ (
    .R(_1__bF$buf8),
    .S(vdd),
    .D(_87_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[2] [2])
);

FILL FILL_1__2795_ (
);

FILL FILL_1__2375_ (
);

FILL FILL_3__3662_ (
);

FILL FILL_3__3242_ (
);

FILL FILL_5__3588_ (
);

FILL FILL_5__3168_ (
);

FILL FILL169650x150 (
);

FILL FILL_6__2872_ (
);

OAI21X1 _3591_ (
    .A(_1568_),
    .B(_1570_),
    .C(_1571_),
    .Y(_1621_)
);

FILL FILL_6__2452_ (
);

NAND2X1 _3171_ (
    .A(_765_),
    .B(_772_),
    .Y(_773_)
);

FILL FILL_6__2032_ (
);

FILL FILL_2__2864_ (
);

FILL FILL_2__2444_ (
);

FILL FILL_2__2024_ (
);

NOR2X1 _1904_ (
    .A(_914__bF$buf3),
    .B(_958_),
    .Y(_1021_)
);

FILL FILL_4__3311_ (
);

FILL FILL_6__3657_ (
);

FILL FILL_6__3237_ (
);

FILL FILL_2__3649_ (
);

FILL FILL_0__3631_ (
);

FILL FILL_2__3229_ (
);

FILL FILL_0__3211_ (
);

FILL FILL169650x118950 (
);

FILL FILL_3__2933_ (
);

FILL FILL_3__2513_ (
);

FILL FILL_5__2859_ (
);

FILL FILL_5__2439_ (
);

FILL FILL_5__2019_ (
);

NAND3X1 _2862_ (
    .A(_500_),
    .B(_509_),
    .C(_466_),
    .Y(_522_)
);

NAND2X1 _2442_ (
    .A(ADD[0]),
    .B(_144_),
    .Y(_145_)
);

INVX1 _2022_ (
    .A(_1132_),
    .Y(_1133_)
);

FILL FILL_5__2192_ (
);

FILL FILL_6__2928_ (
);

FILL FILL_6__2508_ (
);

NAND2X1 _3647_ (
    .A(_1634_),
    .B(_1671_),
    .Y(_1677_)
);

OAI21X1 _3227_ (
    .A(_720__bF$buf3),
    .B(_808_),
    .C(\AXYS[3] [1]),
    .Y(_810_)
);

FILL FILL_7__3571_ (
);

FILL FILL_1__2184_ (
);

FILL FILL_7__3151_ (
);

FILL FILL_0__2902_ (
);

FILL FILL_3__3471_ (
);

FILL FILL_3__3051_ (
);

FILL FILL_6__2681_ (
);

FILL FILL_6__2261_ (
);

FILL FILL_2__2673_ (
);

FILL FILL_2__2253_ (
);

FILL FILL_4__2599_ (
);

FILL FILL_4__2179_ (
);

FILL FILL_4__3540_ (
);

FILL FILL_4__3120_ (
);

FILL FILL_0__2499_ (
);

FILL FILL_6__3466_ (
);

FILL FILL_0__2079_ (
);

FILL FILL_6__3046_ (
);

FILL FILL_2__3458_ (
);

FILL FILL_0__3020_ (
);

FILL FILL_2__3038_ (
);

FILL FILL_5__1883_ (
);

AOI21X1 _2918_ (
    .A(_1181_),
    .B(_561_),
    .C(_562_),
    .Y(_563_)
);

FILL FILL_1__1875_ (
);

FILL FILL_7__2422_ (
);

FILL FILL_3__2742_ (
);

FILL FILL_3__2322_ (
);

FILL FILL_5__2668_ (
);

FILL FILL_5__2248_ (
);

FILL FILL_7__3627_ (
);

FILL FILL_7__3207_ (
);

FILL FILL_1__3601_ (
);

FILL FILL_3__3527_ (
);

FILL FILL_3__3107_ (
);

FILL FILL_6__1952_ (
);

AOI22X1 _2671_ (
    .A(ABL[2]),
    .B(_323_),
    .C(_322_),
    .D(ADD[2]),
    .Y(_344_)
);

NAND2X1 _2251_ (
    .A(RDY_bF$buf5),
    .B(_982_),
    .Y(_1359_)
);

FILL FILL_2__1944_ (
);

FILL FILL168450x61350 (
);

FILL FILL_4__2811_ (
);

FILL FILL_6__2737_ (
);

AND2X2 _3456_ (
    .A(_1703_),
    .B(CO),
    .Y(_1704_)
);

FILL FILL_6__2317_ (
);

OAI21X1 _3036_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[6]),
    .Y(_654_)
);

FILL FILL_0__2711_ (
);

FILL FILL_2__2729_ (
);

FILL FILL_2__2309_ (
);

FILL FILL_3__3280_ (
);

FILL FILL_1__3198_ (
);

FILL FILL_5__1939_ (
);

FILL FILL_6__2490_ (
);

FILL FILL_6__2070_ (
);

FILL FILL_2__2482_ (
);

FILL FILL_2__2062_ (
);

NAND3X1 _1942_ (
    .A(_1054_),
    .B(_1058_),
    .C(_1050_),
    .Y(_1059_)
);

FILL FILL_6__3695_ (
);

FILL FILL_6__3275_ (
);

FILL FILL_2__3267_ (
);

OAI22X1 _2727_ (
    .A(RDY_bF$buf0),
    .B(_1014_),
    .C(_393_),
    .D(_395_),
    .Y(_8_)
);

OAI21X1 _2307_ (
    .A(_1175_),
    .B(_1413_),
    .C(_1411_),
    .Y(_1414_)
);

FILL FILL_7__2651_ (
);

FILL FILL_3__2971_ (
);

FILL FILL_3__2551_ (
);

FILL FILL_3__2131_ (
);

FILL FILL_5__2897_ (
);

FILL FILL_5__2477_ (
);

FILL FILL_5__2057_ (
);

FILL FILL_1__2889_ (
);

FILL FILL_1__2469_ (
);

FILL FILL_1__2049_ (
);

FILL FILL_7__3016_ (
);

FILL FILL_6__1761_ (
);

OAI21X1 _2480_ (
    .A(_1012_),
    .B(_136_),
    .C(_165_),
    .Y(_178_)
);

INVX1 _2060_ (
    .A(IRHOLD[2]),
    .Y(_1169_)
);

FILL FILL_2__1753_ (
);

FILL FILL_4__2620_ (
);

FILL FILL_4__2200_ (
);

FILL FILL_0__1999_ (
);

FILL FILL_6__2966_ (
);

DFFSR _3685_ (
    .R(_1513_),
    .S(vdd),
    .D(_1520_),
    .CLK(clk_bF$buf5),
    .Q(ADD[3])
);

FILL FILL_6__2546_ (
);

NAND3X1 _3265_ (
    .A(_314_),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

FILL FILL_6__2126_ (
);

FILL FILL_2__2958_ (
);

FILL FILL_0__2940_ (
);

FILL FILL_0__2520_ (
);

FILL FILL_2__2538_ (
);

FILL FILL_2__2118_ (
);

FILL FILL_0__2100_ (
);

FILL FILL_7__1922_ (
);

FILL FILL_3__1822_ (
);

FILL FILL_0__3305_ (
);

FILL FILL_5__1748_ (
);

FILL FILL_2__2291_ (
);

FILL FILL_3__2607_ (
);

NAND2X1 _1751_ (
    .A(RDY_bF$buf9),
    .B(DI[2]),
    .Y(_883_)
);

FILL FILL_6__3084_ (
);

FILL FILL_2__3496_ (
);

FILL FILL_2__3076_ (
);

INVX1 _2956_ (
    .A(_592_),
    .Y(_593_)
);

FILL FILL_6__1817_ (
);

OAI21X1 _2536_ (
    .A(_1005_),
    .B(_218_),
    .C(_229_),
    .Y(_230_)
);

INVX1 _2116_ (
    .A(_974_),
    .Y(_1225_)
);

FILL FILL_7__2880_ (
);

FILL FILL_7__2040_ (
);

FILL FILL_2__1809_ (
);

FILL FILL_3__2780_ (
);

FILL FILL_3__2360_ (
);

FILL FILL_5__2286_ (
);

FILL FILL_1__2698_ (
);

FILL FILL_1__2278_ (
);

FILL FILL_3__3565_ (
);

FILL FILL_3__3145_ (
);

FILL FILL_6__1990_ (
);

FILL FILL_2__1982_ (
);

FILL FILL_6__2775_ (
);

NAND2X1 _3494_ (
    .A(alu_op[2]),
    .B(_1725_),
    .Y(_1739_)
);

FILL FILL_6__2355_ (
);

OAI21X1 _3074_ (
    .A(_1055_),
    .B(_1036_),
    .C(_1045_),
    .Y(_686_)
);

FILL FILL_2__2767_ (
);

FILL FILL_2__2347_ (
);

OAI21X1 _1807_ (
    .A(_925_),
    .B(_932_),
    .C(CO),
    .Y(_933_)
);

FILL FILL_4__3634_ (
);

FILL FILL_4__3214_ (
);

FILL FILL_0__3534_ (
);

FILL FILL_0__3114_ (
);

FILL FILL_5__1977_ (
);

FILL FILL_1__1969_ (
);

FILL FILL_7__2516_ (
);

FILL FILL_1__2910_ (
);

FILL FILL_3__2836_ (
);

FILL FILL_3__2416_ (
);

AOI21X1 _1980_ (
    .A(_1082_),
    .B(ADD[1]),
    .C(_1095_),
    .Y(_1096_)
);

FILL FILL_5__3703_ (
);

NOR2X1 _2765_ (
    .A(_428_),
    .B(_401_),
    .Y(_430_)
);

OR2X2 _2345_ (
    .A(_1358_),
    .B(_1363_),
    .Y(_1452_)
);

FILL FILL_5__2095_ (
);

FILL FILL_4__2905_ (
);

FILL FILL_7__3474_ (
);

FILL FILL_1__2087_ (
);

FILL FILL_7__3054_ (
);

FILL FILL_0__2805_ (
);

FILL FILL_2__1791_ (
);

FILL FILL_6__2584_ (
);

FILL FILL_6__2164_ (
);

FILL FILL_2__2996_ (
);

FILL FILL_2__2576_ (
);

FILL FILL_2__2156_ (
);

FILL FILL_4__3023_ (
);

FILL FILL_3__1860_ (
);

FILL FILL_5__1786_ (
);

FILL FILL_1__1778_ (
);

FILL FILL_7__2745_ (
);

FILL FILL_7__2325_ (
);

FILL FILL_3__2645_ (
);

FILL FILL_3__2225_ (
);

FILL FILL_5__3512_ (
);

FILL FILL_1__3504_ (
);

FILL FILL_6__1855_ (
);

OAI21X1 _2994_ (
    .A(_1160_),
    .B(_621_),
    .C(_622_),
    .Y(_623_)
);

INVX1 _2574_ (
    .A(_262_),
    .Y(_1741_[6])
);

NOR2X1 _2154_ (
    .A(_914__bF$buf2),
    .B(_1069_),
    .Y(_1263_)
);

FILL FILL_2__1847_ (
);

FILL FILL_4__2714_ (
);

DFFSR _3359_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_36_),
    .CLK(clk_bF$buf9),
    .Q(rotate)
);

FILL FILL_7__3283_ (
);

FILL FILL_0__2614_ (
);

FILL FILL_3__3183_ (
);

FILL FILL_3__1916_ (
);

FILL FILL_6__2393_ (
);

FILL FILL_2__2385_ (
);

NAND2X1 _1845_ (
    .A(state[2]),
    .B(state[3]),
    .Y(_970_)
);

FILL FILL_4__3672_ (
);

FILL FILL_4__3252_ (
);

FILL FILL_6__3598_ (
);

FILL FILL_6__3178_ (
);

FILL FILL_0__3572_ (
);

FILL FILL_0__3152_ (
);

FILL FILL_7__2974_ (
);

FILL FILL_7__2554_ (
);

FILL FILL_7__2134_ (
);

FILL FILL_3__2874_ (
);

FILL FILL_3__2454_ (
);

FILL FILL_3__2034_ (
);

FILL FILL_1__3313_ (
);

FILL FILL_3__3659_ (
);

FILL FILL_3__3239_ (
);

NAND3X1 _2383_ (
    .A(_1308_),
    .B(_1336_),
    .C(_1488_),
    .Y(_1489_)
);

FILL FILL_4__2943_ (
);

FILL FILL_4__2523_ (
);

FILL FILL_4__2103_ (
);

FILL FILL_6__2869_ (
);

NAND2X1 _3588_ (
    .A(_1617_),
    .B(_1614_),
    .Y(_1618_)
);

FILL FILL_6__2449_ (
);

NOR2X1 _3168_ (
    .A(_769_),
    .B(_759_),
    .Y(_770_)
);

FILL FILL_6__2029_ (
);

FILL FILL_0__2843_ (
);

FILL FILL_0__2423_ (
);

FILL FILL_0__2003_ (
);

FILL FILL_4__3308_ (
);

FILL FILL_0__3628_ (
);

FILL FILL_0__3208_ (
);

FILL FILL_2__2194_ (
);

FILL FILL_4__3481_ (
);

FILL FILL_4__3061_ (
);

NOR2X1 _2859_ (
    .A(_518_),
    .B(_514_),
    .Y(_519_)
);

NAND3X1 _2439_ (
    .A(_1227_),
    .B(_142_),
    .C(_138_),
    .Y(_1743_)
);

AOI22X1 _2019_ (
    .A(_1049_),
    .B(\AXYS[3] [6]),
    .C(\AXYS[2] [6]),
    .D(_1057_),
    .Y(_1130_)
);

FILL FILL_7__2783_ (
);

FILL FILL_3__2683_ (
);

FILL FILL_3__2263_ (
);

FILL FILL_5__2189_ (
);

FILL FILL_5__3550_ (
);

FILL FILL_7__3148_ (
);

FILL FILL_5__3130_ (
);

FILL FILL_1__3542_ (
);

FILL FILL_1__3122_ (
);

FILL FILL_3__3468_ (
);

FILL FILL_3__3048_ (
);

FILL FILL_6__1893_ (
);

NAND2X1 _2192_ (
    .A(_1300_),
    .B(_1294_),
    .Y(_1301_)
);

FILL FILL_2__1885_ (
);

FILL FILL_4__2752_ (
);

FILL FILL_4__2332_ (
);

FILL FILL_6__2678_ (
);

DFFSR _3397_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_66_),
    .CLK(clk_bF$buf1),
    .Q(Z)
);

FILL FILL_6__2258_ (
);

FILL FILL_0__2652_ (
);

FILL FILL_0__2232_ (
);

FILL FILL_2__3611_ (
);

FILL FILL_4__3537_ (
);

FILL FILL_4__3117_ (
);

FILL FILL_3__1954_ (
);

FILL FILL_0__3017_ (
);

FILL FILL_5__2821_ (
);

FILL FILL_7__2419_ (
);

FILL FILL_5__2401_ (
);

FILL FILL_1__2813_ (
);

FILL FILL_3__2739_ (
);

FILL FILL_3__2319_ (
);

OAI22X1 _1883_ (
    .A(_1005_),
    .B(_968_),
    .C(_1006_),
    .D(_1004_),
    .Y(BI[1])
);

FILL FILL_4__3290_ (
);

FILL FILL_5__3606_ (
);

FILL FILL_0__3190_ (
);

FILL FILL_6__1949_ (
);

OAI22X1 _2668_ (
    .A(RDY_bF$buf3),
    .B(_1005_),
    .C(_341_),
    .D(_339_),
    .Y(_3_)
);

NOR2X1 _2248_ (
    .A(_1217_),
    .B(_1355_),
    .Y(_1356_)
);

FILL FILL_7__2172_ (
);

FILL FILL_0__1923_ (
);

FILL FILL_3__2492_ (
);

FILL FILL_3__2072_ (
);

FILL FILL_4__2808_ (
);

FILL FILL_0__2708_ (
);

FILL FILL_3__3697_ (
);

FILL FILL_3__3277_ (
);

FILL FILL_4__2981_ (
);

FILL FILL_4__2561_ (
);

FILL FILL_4__2141_ (
);

FILL FILL_6__2487_ (
);

FILL FILL_6__2067_ (
);

FILL FILL_0__2881_ (
);

FILL FILL_2__2899_ (
);

FILL FILL_2__2479_ (
);

FILL FILL_0__2461_ (
);

FILL FILL_2__2059_ (
);

FILL FILL_0__2041_ (
);

NAND3X1 _1939_ (
    .A(_1055_),
    .B(_1035_),
    .C(_1026_),
    .Y(_1056_)
);

FILL FILL_2__3000_ (
);

FILL FILL_7__1863_ (
);

FILL FILL_0__3666_ (
);

FILL FILL_3__1763_ (
);

FILL FILL_0__3246_ (
);

FILL FILL_7__2648_ (
);

FILL FILL_5__2630_ (
);

FILL FILL_5__2210_ (
);

FILL FILL_1__2622_ (
);

FILL FILL_1__2202_ (
);

FILL FILL_3__2968_ (
);

FILL FILL_3__2548_ (
);

FILL FILL_3__2128_ (
);

FILL FILL_4__1832_ (
);

FILL FILL_6__1758_ (
);

OAI21X1 _2897_ (
    .A(_886__bF$buf1),
    .B(_1027__bF$buf1),
    .C(cli),
    .Y(_546_)
);

OAI21X1 _2477_ (
    .A(_173_),
    .B(_174_),
    .C(_175_),
    .Y(_176_)
);

NAND2X1 _2057_ (
    .A(_1152_),
    .B(_1153_),
    .Y(_1166_)
);

FILL FILL_4__2617_ (
);

FILL FILL_7__3186_ (
);

FILL FILL_0__2937_ (
);

FILL FILL_0__2517_ (
);

FILL FILL_1__3580_ (
);

FILL FILL_1__3160_ (
);

FILL FILL_3__3086_ (
);

FILL FILL_5__1901_ (
);

FILL FILL_7__1919_ (
);

FILL FILL_3__1819_ (
);

FILL FILL_4__2790_ (
);

FILL FILL_4__2370_ (
);

FILL FILL_6__2296_ (
);

FILL FILL_0__2690_ (
);

FILL FILL_0__2270_ (
);

FILL FILL_2__2288_ (
);

NAND2X1 _1748_ (
    .A(RDY_bF$buf9),
    .B(DI[1]),
    .Y(_881_)
);

FILL FILL_4__3575_ (
);

FILL FILL_4__3155_ (
);

FILL FILL_3__1992_ (
);

FILL FILL_0__3475_ (
);

FILL FILL_0__3055_ (
);

FILL FILL_7__2877_ (
);

FILL FILL_7__2037_ (
);

FILL FILL_1__2851_ (
);

FILL FILL_1__2431_ (
);

FILL FILL_1__2011_ (
);

FILL FILL_3__2777_ (
);

FILL FILL_3__2357_ (
);

FILL FILL_5__3644_ (
);

FILL FILL_5__3224_ (
);

FILL FILL_1__3636_ (
);

FILL FILL_1__3216_ (
);

FILL FILL_6__1987_ (
);

OAI21X1 _2286_ (
    .A(_1184_),
    .B(_1177_),
    .C(_1167_),
    .Y(_1393_)
);

FILL FILL_2__1979_ (
);

FILL FILL_0__1961_ (
);

FILL FILL_3_BUFX2_insert40 (
);

FILL FILL_3_BUFX2_insert41 (
);

FILL FILL_3_BUFX2_insert42 (
);

FILL FILL_3_BUFX2_insert43 (
);

FILL FILL_2__2920_ (
);

FILL FILL_2__2500_ (
);

FILL FILL_3_BUFX2_insert44 (
);

FILL FILL_3_BUFX2_insert45 (
);

FILL FILL_3_BUFX2_insert46 (
);

FILL FILL_3_BUFX2_insert47 (
);

FILL FILL_4__2846_ (
);

FILL FILL_3_BUFX2_insert48 (
);

FILL FILL_4__2426_ (
);

FILL FILL_3_BUFX2_insert49 (
);

FILL FILL_4__2006_ (
);

FILL FILL_0__2746_ (
);

FILL FILL_6__3713_ (
);

FILL FILL_0__2326_ (
);

FILL FILL_2__3705_ (
);

FILL FILL_5__2915_ (
);

FILL FILL_2__2097_ (
);

FILL FILL_1__2907_ (
);

NOR2X1 _1977_ (
    .A(_1091_),
    .B(_1092_),
    .Y(_1093_)
);

FILL FILL_0__3284_ (
);

FILL FILL_7__2266_ (
);

BUFX2 _3703_ (
    .A(_1741_[6]),
    .Y(AB[6])
);

FILL FILL_1__2660_ (
);

FILL FILL_1__2240_ (
);

FILL FILL_3__2586_ (
);

FILL FILL_3__2166_ (
);

FILL FILL_5__3453_ (
);

FILL FILL_5__3033_ (
);

FILL FILL_1__3025_ (
);

FILL FILL_4__1870_ (
);

FILL FILL_6__1796_ (
);

NOR2X1 _2095_ (
    .A(_1201_),
    .B(_1203_),
    .Y(_1204_)
);

FILL FILL_2__1788_ (
);

FILL FILL_0__1770_ (
);

FILL FILL_4__2655_ (
);

FILL FILL_4__2235_ (
);

FILL FILL_0__2975_ (
);

FILL FILL_0__2555_ (
);

FILL FILL_6__3522_ (
);

FILL FILL_0__2135_ (
);

FILL FILL_6__3102_ (
);

FILL FILL_2__3514_ (
);

FILL FILL_1__1931_ (
);

FILL FILL_3__1857_ (
);

FILL FILL_5__2724_ (
);

FILL FILL_5__2304_ (
);

FILL FILL_1__2716_ (
);

NAND2X1 _1786_ (
    .A(_910_),
    .B(_911_),
    .Y(_912_)
);

FILL FILL_4__3193_ (
);

FILL FILL_5__3509_ (
);

FILL FILL_0__3093_ (
);

FILL FILL_4__1926_ (
);

FILL FILL_7__2495_ (
);

FILL FILL_7__2075_ (
);

FILL FILL_0__1826_ (
);

OAI21X1 _3512_ (
    .A(alu_op[1]),
    .B(_1538_),
    .C(_1541_),
    .Y(_1542_)
);

FILL FILL_3__2395_ (
);

FILL FILL_5__3262_ (
);

FILL FILL_1__3674_ (
);

FILL FILL_1__3254_ (
);

FILL FILL_4__2884_ (
);

FILL FILL_4__2464_ (
);

FILL FILL_4__2044_ (
);

FILL FILL_0__2784_ (
);

FILL FILL_0__2364_ (
);

FILL FILL_4__3669_ (
);

FILL FILL_7__1766_ (
);

FILL FILL_4__3249_ (
);

FILL FILL_0__3569_ (
);

FILL FILL_0__3149_ (
);

FILL FILL_5__2953_ (
);

FILL FILL_5__2533_ (
);

FILL FILL_5__2113_ (
);

FILL FILL_1__2945_ (
);

FILL FILL_1__2525_ (
);

FILL FILL_1__2105_ (
);

FILL FILL168450x118950 (
);

FILL FILL_6__2602_ (
);

DFFSR _3321_ (
    .R(vdd),
    .S(_1__bF$buf9),
    .D(_1512_[3]),
    .CLK(clk_bF$buf6),
    .Q(state[3])
);

FILL FILL_5__3491_ (
);

FILL FILL_5__3071_ (
);

FILL FILL_1__3483_ (
);

FILL FILL_1__3063_ (
);

FILL FILL_5__1804_ (
);

FILL FILL_4__2693_ (
);

FILL FILL_4__2273_ (
);

FILL FILL_6__2199_ (
);

FILL FILL_0__2593_ (
);

FILL FILL_6__3560_ (
);

FILL FILL_0__2173_ (
);

FILL FILL_6__3140_ (
);

FILL FILL_2__3552_ (
);

FILL FILL_2__3132_ (
);

FILL FILL_7__1995_ (
);

FILL FILL_4__3478_ (
);

FILL FILL_4__3058_ (
);

FILL FILL_3__1895_ (
);

FILL FILL_5__2762_ (
);

FILL FILL_5__2342_ (
);

FILL FILL_1__2754_ (
);

FILL FILL_1__2334_ (
);

FILL FILL_7__3301_ (
);

FILL FILL_3__3621_ (
);

FILL FILL_3__3201_ (
);

FILL FILL_5__3547_ (
);

FILL FILL_5__3127_ (
);

FILL FILL_1__3539_ (
);

FILL FILL_1__3119_ (
);

FILL FILL_4__1964_ (
);

OAI21X1 _2189_ (
    .A(_1297_),
    .B(_1092_),
    .C(RDY_bF$buf7),
    .Y(_1298_)
);

FILL FILL_0__1864_ (
);

FILL FILL_6__2831_ (
);

OAI21X1 _3550_ (
    .A(_1574_),
    .B(_1578_),
    .C(_1579_),
    .Y(_1580_)
);

FILL FILL_6__2411_ (
);

INVX1 _3130_ (
    .A(_736_),
    .Y(_737_)
);

FILL FILL_2__2823_ (
);

FILL FILL_2__2403_ (
);

FILL FILL_4__2749_ (
);

FILL FILL_4__2329_ (
);

FILL FILL_0__2649_ (
);

FILL FILL_6__3616_ (
);

FILL FILL_0__2229_ (
);

FILL FILL_1__3292_ (
);

FILL FILL_2__3608_ (
);

FILL FILL_4__2082_ (
);

FILL FILL_5__2818_ (
);

FILL FILL_4__3287_ (
);

NOR3X1 _2821_ (
    .A(_478_),
    .B(_443_),
    .C(_483_),
    .Y(_484_)
);

NAND3X1 _2401_ (
    .A(_1495_),
    .B(_1505_),
    .C(_1503_),
    .Y(_1512_[4])
);

FILL FILL_0__3187_ (
);

FILL FILL_5__2991_ (
);

FILL FILL_5__2571_ (
);

FILL FILL_5__2151_ (
);

FILL FILL_7__2169_ (
);

AOI22X1 _3606_ (
    .A(_1738_),
    .B(_1527_),
    .C(_1630_),
    .D(_1635_),
    .Y(_1636_)
);

FILL FILL_1__2983_ (
);

FILL FILL_1__2563_ (
);

FILL FILL_7__3530_ (
);

FILL FILL_1__2143_ (
);

FILL FILL_3__2489_ (
);

FILL FILL_3__2069_ (
);

FILL FILL_3__3010_ (
);

FILL FILL_4__1773_ (
);

FILL FILL_6__2640_ (
);

FILL FILL_6__2220_ (
);

FILL FILL_2__2632_ (
);

FILL FILL_2__2212_ (
);

FILL FILL_4__2978_ (
);

FILL FILL_4__2558_ (
);

FILL FILL_4__2138_ (
);

FILL FILL_0__2878_ (
);

FILL FILL_0__2458_ (
);

FILL FILL_0__2038_ (
);

FILL FILL_6__3005_ (
);

FILL FILL_5__1842_ (
);

FILL FILL_1__1834_ (
);

FILL FILL_7__2801_ (
);

FILL FILL_3__2701_ (
);

FILL FILL_5__2627_ (
);

FILL FILL_5__2207_ (
);

FILL FILL_1__2619_ (
);

FILL FILL_2__3590_ (
);

FILL FILL_2__3170_ (
);

FILL FILL_4__3096_ (
);

FILL FILL_6__1911_ (
);

NOR2X1 _2630_ (
    .A(_308_),
    .B(_164_),
    .Y(_0_)
);

INVX4 _2210_ (
    .A(_1018_),
    .Y(_1319_)
);

FILL FILL_2__1903_ (
);

FILL FILL_4__1829_ (
);

FILL FILL_7__2398_ (
);

FILL FILL_5__2380_ (
);

DFFSR _3415_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_84_),
    .CLK(clk_bF$buf7),
    .Q(\AXYS[1] [7])
);

FILL FILL_1__2792_ (
);

FILL FILL_1__2372_ (
);

FILL FILL_3__2298_ (
);

FILL FILL_5__3585_ (
);

FILL FILL_5__3165_ (
);

FILL FILL_1__3577_ (
);

FILL FILL_1__3157_ (
);

FILL FILL_2__2861_ (
);

FILL FILL_2__2441_ (
);

FILL FILL_2__2021_ (
);

FILL FILL_4__2787_ (
);

FILL FILL_4__2367_ (
);

NAND2X1 _1901_ (
    .A(_969_),
    .B(_935_),
    .Y(_1018_)
);

FILL FILL_0__2687_ (
);

FILL FILL_6__3654_ (
);

FILL FILL_0__2267_ (
);

FILL FILL_6__3234_ (
);

FILL FILL_2__3646_ (
);

FILL FILL_2__3226_ (
);

FILL FILL_3__1989_ (
);

FILL FILL_3__2930_ (
);

FILL FILL_3__2510_ (
);

FILL FILL_5__2856_ (
);

FILL FILL_5__2436_ (
);

FILL FILL_5__2016_ (
);

FILL FILL_1__2848_ (
);

FILL FILL_1__2428_ (
);

FILL FILL_1__2008_ (
);

FILL FILL_3__3715_ (
);

FILL FILL_0__1958_ (
);

FILL FILL_6__2925_ (
);

NAND3X1 _3644_ (
    .A(_1638_),
    .B(_1648_),
    .C(_1673_),
    .Y(_1674_)
);

FILL FILL_6__2505_ (
);

INVX2 _3224_ (
    .A(_1049_),
    .Y(_808_)
);

FILL FILL_1__2181_ (
);

FILL FILL_2__2917_ (
);

FILL FILL_2__2670_ (
);

FILL FILL_2__2250_ (
);

FILL FILL_4__2596_ (
);

FILL FILL_4__2176_ (
);

FILL FILL_0__2496_ (
);

FILL FILL_6__3463_ (
);

FILL FILL_0__2076_ (
);

FILL FILL_6__3043_ (
);

FILL FILL_2__3455_ (
);

FILL FILL_2__3035_ (
);

FILL FILL_7__1898_ (
);

FILL FILL_5__1880_ (
);

NOR2X1 _2915_ (
    .A(_1217_),
    .B(_559_),
    .Y(_560_)
);

FILL FILL_1__1872_ (
);

FILL FILL_3__1798_ (
);

FILL FILL_5__2665_ (
);

FILL FILL_5__2245_ (
);

FILL FILL_1__2657_ (
);

FILL FILL_7__3624_ (
);

FILL FILL_1__2237_ (
);

FILL FILL_7__3204_ (
);

FILL FILL_3__3524_ (
);

FILL FILL_3__3104_ (
);

FILL FILL_2__1941_ (
);

FILL FILL_4__1867_ (
);

FILL FILL_0__1767_ (
);

FILL FILL_6__2734_ (
);

NAND3X1 _3453_ (
    .A(_1699_),
    .B(_1700_),
    .C(_1701_),
    .Y(_1702_)
);

FILL FILL_6__2314_ (
);

OAI21X1 _3033_ (
    .A(_888_),
    .B(_647_),
    .C(_652_),
    .Y(_57_)
);

FILL FILL_2__2726_ (
);

FILL FILL_2__2306_ (
);

FILL FILL_6__3519_ (
);

FILL FILL_1__3195_ (
);

FILL FILL_5__1936_ (
);

FILL FILL_1__1928_ (
);

FILL FILL_6__3692_ (
);

FILL FILL_6__3272_ (
);

FILL FILL_2__3264_ (
);

NOR2X1 _2724_ (
    .A(_392_),
    .B(_386_),
    .Y(_393_)
);

NAND2X1 _2304_ (
    .A(_1370_),
    .B(_1351_),
    .Y(_1411_)
);

FILL FILL_5__2894_ (
);

FILL FILL_5__2474_ (
);

FILL FILL_5__2054_ (
);

INVX1 _3509_ (
    .A(AI[3]),
    .Y(_1539_)
);

FILL FILL_1__2886_ (
);

FILL FILL_1__2466_ (
);

FILL FILL_1__2046_ (
);

FILL FILL_5__3259_ (
);

FILL FILL_2__1750_ (
);

FILL FILL_0__1996_ (
);

FILL FILL_6__2963_ (
);

DFFSR _3682_ (
    .R(_1513_),
    .S(vdd),
    .D(_1517_),
    .CLK(clk_bF$buf5),
    .Q(ADD[0])
);

FILL FILL_6__2543_ (
);

NAND3X1 _3262_ (
    .A(_1022_),
    .B(_317_),
    .C(_837_),
    .Y(_838_)
);

FILL FILL_6__2123_ (
);

FILL FILL_2__2955_ (
);

FILL FILL_2__2535_ (
);

FILL FILL_2__2115_ (
);

FILL FILL_0__3302_ (
);

FILL FILL_5__1745_ (
);

FILL FILL_7__2704_ (
);

FILL FILL_3__2604_ (
);

FILL FILL_6__3081_ (
);

FILL FILL169950x151350 (
);

FILL FILL_2__3493_ (
);

FILL FILL_2__3073_ (
);

FILL FILL_6__1814_ (
);

NAND2X1 _2953_ (
    .A(_1150__bF$buf1),
    .B(_564_),
    .Y(_591_)
);

INVX1 _2533_ (
    .A(_201_),
    .Y(_227_)
);

NAND2X1 _2113_ (
    .A(_969_),
    .B(_1221_),
    .Y(_1222_)
);

FILL FILL_2__1806_ (
);

FILL FILL169950x118950 (
);

FILL FILL_5__2283_ (
);

DFFSR _3318_ (
    .R(_1__bF$buf9),
    .S(vdd),
    .D(_1512_[0]),
    .CLK(clk_bF$buf6),
    .Q(state[0])
);

FILL FILL_1__2695_ (
);

FILL FILL_7__3662_ (
);

FILL FILL_1__2275_ (
);

FILL FILL_3__3562_ (
);

FILL FILL_3__3142_ (
);

FILL FILL_5__3488_ (
);

FILL FILL_5__3068_ (
);

FILL FILL_6__2772_ (
);

AOI22X1 _3491_ (
    .A(_1716_),
    .B(BI[5]),
    .C(_1735_),
    .D(_1717_),
    .Y(_1736_)
);

FILL FILL_6__2352_ (
);

NOR2X1 _3071_ (
    .A(_1021_),
    .B(_683_),
    .Y(_684_)
);

FILL FILL_2__2764_ (
);

FILL FILL_2__2344_ (
);

NAND2X1 _1804_ (
    .A(_929_),
    .B(_900_),
    .Y(_930_)
);

FILL FILL_4__3631_ (
);

FILL FILL_4__3211_ (
);

FILL FILL_6__3557_ (
);

FILL FILL_6__3137_ (
);

FILL FILL_0__3531_ (
);

FILL FILL_2__3549_ (
);

FILL FILL_2__3129_ (
);

FILL FILL_0__3111_ (
);

FILL FILL_5__1974_ (
);

FILL FILL_1__1966_ (
);

FILL FILL_7__2933_ (
);

FILL FILL_3__2833_ (
);

FILL FILL_3__2413_ (
);

FILL FILL_5__2759_ (
);

FILL FILL_5__2339_ (
);

FILL FILL_5__3700_ (
);

FILL FILL_3__3618_ (
);

OAI21X1 _2762_ (
    .A(_426_),
    .B(_427_),
    .C(_423_),
    .Y(_428_)
);

OR2X2 _2342_ (
    .A(_1202_),
    .B(RDY_bF$buf8),
    .Y(_1449_)
);

FILL FILL_5__2092_ (
);

FILL FILL_4__2902_ (
);

FILL FILL_6__2828_ (
);

OAI21X1 _3547_ (
    .A(alu_op[0]),
    .B(_1575_),
    .C(_1576_),
    .Y(_1577_)
);

FILL FILL_6__2408_ (
);

NOR2X1 _3127_ (
    .A(_1319__bF$buf3),
    .B(_733_),
    .Y(_734_)
);

FILL FILL_7__3471_ (
);

FILL FILL_1__2084_ (
);

FILL FILL_7__3051_ (
);

FILL FILL_0__2802_ (
);

FILL FILL_5__3297_ (
);

FILL FILL_1__3289_ (
);

FILL FILL_6__2581_ (
);

FILL FILL_6__2161_ (
);

FILL FILL_2__2993_ (
);

FILL FILL_2__2573_ (
);

FILL FILL_2__2153_ (
);

FILL FILL_4__2499_ (
);

FILL FILL_4__2079_ (
);

FILL FILL_4__3020_ (
);

FILL FILL_0__2399_ (
);

FILL FILL_5__1783_ (
);

NAND3X1 _2818_ (
    .A(_446_),
    .B(_480_),
    .C(_479_),
    .Y(_481_)
);

FILL FILL_1__1775_ (
);

FILL FILL_7__2322_ (
);

FILL FILL_3__2642_ (
);

FILL FILL_3__2222_ (
);

FILL FILL_5__2988_ (
);

FILL FILL_5__2568_ (
);

FILL FILL_5__2148_ (
);

FILL FILL_7__3527_ (
);

FILL FILL_7__3107_ (
);

FILL FILL_1__3501_ (
);

FILL FILL_3__3007_ (
);

OAI21X1 _2991_ (
    .A(_579_),
    .B(_578_),
    .C(_1150__bF$buf4),
    .Y(_620_)
);

FILL FILL_6__1852_ (
);

AND2X2 _2571_ (
    .A(_258_),
    .B(_259_),
    .Y(_260_)
);

NOR2X1 _2151_ (
    .A(_931__bF$buf4),
    .B(_1069_),
    .Y(_1260_)
);

FILL FILL_2__1844_ (
);

FILL FILL_4__2711_ (
);

FILL FILL_6__2637_ (
);

DFFSR _3356_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_33_),
    .CLK(clk_bF$buf9),
    .Q(op[1])
);

FILL FILL_6__2217_ (
);

FILL FILL_7__3280_ (
);

FILL FILL_0__2611_ (
);

FILL FILL_2__2629_ (
);

FILL FILL_2__2209_ (
);

FILL FILL_3__3180_ (
);

FILL FILL_1__3098_ (
);

FILL FILL_3__1913_ (
);

FILL FILL_5__1839_ (
);

FILL FILL_6__2390_ (
);

CLKBUF1 CLKBUF1_insert30 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert31 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert32 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert33 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert34 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert35 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert36 (
    .A(clk),
    .Y(clk_bF$buf0)
);

FILL FILL_2__2382_ (
);

NOR2X1 _1842_ (
    .A(_914__bF$buf4),
    .B(_946_),
    .Y(_967_)
);

FILL FILL_6__3595_ (
);

FILL FILL_6__3175_ (
);

FILL FILL_2__3587_ (
);

FILL FILL_2__3167_ (
);

FILL FILL_6__1908_ (
);

AOI21X1 _2627_ (
    .A(_272_),
    .B(DIMUX[7]),
    .C(_306_),
    .Y(_307_)
);

OAI21X1 _2207_ (
    .A(_902__bF$buf2),
    .B(_958_),
    .C(_886__bF$buf0),
    .Y(_1316_)
);

FILL FILL_7__2551_ (
);

FILL FILL_3__2871_ (
);

FILL FILL_3__2451_ (
);

FILL FILL_3__2031_ (
);

FILL FILL_5__2797_ (
);

FILL FILL_5__2377_ (
);

FILL FILL_1__2789_ (
);

FILL FILL_1__2369_ (
);

FILL FILL_1__3310_ (
);

FILL FILL_3__3656_ (
);

FILL FILL_3__3236_ (
);

NOR2X1 _2380_ (
    .A(_1479_),
    .B(_1452_),
    .Y(_1486_)
);

FILL FILL_4__1999_ (
);

FILL FILL_4__2940_ (
);

FILL FILL_4__2520_ (
);

FILL FILL_4__2100_ (
);

FILL FILL_0__1899_ (
);

FILL FILL_6__2866_ (
);

INVX1 _3585_ (
    .A(_1570_),
    .Y(_1615_)
);

FILL FILL_6__2446_ (
);

FILL FILL_6__2026_ (
);

NAND2X1 _3165_ (
    .A(\AXYS[0] [5]),
    .B(_722_),
    .Y(_768_)
);

FILL FILL_0__2840_ (
);

FILL FILL_2__2858_ (
);

FILL FILL169650x32550 (
);

FILL FILL_2__2438_ (
);

FILL FILL_0__2420_ (
);

FILL FILL_2__2018_ (
);

FILL FILL_0__2000_ (
);

FILL FILL_7__1822_ (
);

FILL FILL_4__3305_ (
);

FILL FILL_0__3625_ (
);

FILL FILL_0__3205_ (
);

FILL FILL_2__2191_ (
);

FILL FILL_3__2927_ (
);

FILL FILL_3__2507_ (
);

AOI22X1 _2856_ (
    .A(AN),
    .B(_1299_),
    .C(_323_),
    .D(ABH[7]),
    .Y(_516_)
);

NOR2X1 _2436_ (
    .A(_140_),
    .B(_129_),
    .Y(alu_op[3])
);

AOI21X1 _2016_ (
    .A(_1082_),
    .B(ADD[5]),
    .C(_1127_),
    .Y(_1128_)
);

FILL FILL_7__2780_ (
);

FILL FILL_3__2680_ (
);

FILL FILL_3__2260_ (
);

FILL FILL_5__2186_ (
);

FILL FILL168450x14550 (
);

FILL FILL_1__2598_ (
);

FILL FILL_1__2178_ (
);

FILL FILL_7__3145_ (
);

FILL FILL_3__3465_ (
);

FILL FILL_3__3045_ (
);

FILL FILL_6__1890_ (
);

FILL FILL_2__1882_ (
);

FILL FILL_6__2675_ (
);

DFFSR _3394_ (
    .R(_1__bF$buf5),
    .S(vdd),
    .D(_63_),
    .CLK(clk_bF$buf1),
    .Q(D)
);

FILL FILL_6__2255_ (
);

FILL FILL_2__2667_ (
);

FILL FILL_2__2247_ (
);

FILL FILL_4__3534_ (
);

FILL FILL_4__3114_ (
);

FILL FILL_3__1951_ (
);

FILL FILL_0__3014_ (
);

FILL FILL_5__1877_ (
);

FILL FILL_1__1869_ (
);

FILL FILL_7__2416_ (
);

FILL FILL_1__2810_ (
);

FILL FILL_3__2736_ (
);

FILL FILL_3__2316_ (
);

OAI22X1 _1880_ (
    .A(_965_),
    .B(_968_),
    .C(_966_),
    .D(_1004_),
    .Y(BI[0])
);

FILL FILL_5__3603_ (
);

FILL FILL_6__1946_ (
);

NOR2X1 _2665_ (
    .A(_338_),
    .B(_333_),
    .Y(_339_)
);

NAND3X1 _2245_ (
    .A(_1347_),
    .B(_1352_),
    .C(_1346_),
    .Y(_1353_)
);

FILL FILL_0__1920_ (
);

FILL FILL_2__1938_ (
);

FILL FILL_4__2805_ (
);

FILL FILL_0__2705_ (
);

FILL FILL_3__3694_ (
);

FILL FILL_3__3274_ (
);

FILL FILL_6__2484_ (
);

FILL FILL_6__2064_ (
);

FILL FILL_2__2896_ (
);

FILL FILL_2__2476_ (
);

FILL FILL_2__2056_ (
);

OAI21X1 _1936_ (
    .A(src_reg[0]),
    .B(_1036_),
    .C(_1052_),
    .Y(_1053_)
);

FILL FILL_6__3269_ (
);

FILL FILL_3__1760_ (
);

FILL FILL_0__3663_ (
);

FILL FILL_0__3243_ (
);

FILL FILL_7__2645_ (
);

FILL FILL_7__2225_ (
);

FILL FILL_3__2965_ (
);

FILL FILL_3__2545_ (
);

FILL FILL_3__2125_ (
);

FILL FILL_6__1755_ (
);

OAI21X1 _2894_ (
    .A(_537_),
    .B(_544_),
    .C(_542_),
    .Y(_26_)
);

INVX1 _2474_ (
    .A(ADD[4]),
    .Y(_173_)
);

AOI21X1 _2054_ (
    .A(IRHOLD_valid),
    .B(_1162_),
    .C(_1154_),
    .Y(_1163_)
);

FILL FILL_2__1747_ (
);

FILL FILL_4__2614_ (
);

DFFSR _3679_ (
    .R(_1513_),
    .S(vdd),
    .D(_1514_),
    .CLK(clk_bF$buf6),
    .Q(\u_ALU8.BI7 )
);

OAI21X1 _3259_ (
    .A(_834_),
    .B(_831_),
    .C(_826_),
    .Y(_835_)
);

FILL FILL_7__3183_ (
);

FILL FILL_0__2934_ (
);

FILL FILL_0__2514_ (
);

FILL FILL_3__3083_ (
);

FILL FILL169950x75750 (
);

FILL FILL_7__1916_ (
);

FILL FILL_3__1816_ (
);

FILL FILL_6__2293_ (
);

FILL FILL_2__2285_ (
);

NAND2X1 _1745_ (
    .A(DI[0]),
    .B(RDY_bF$buf0),
    .Y(_879_)
);

FILL FILL_4__3572_ (
);

FILL FILL_4__3152_ (
);

FILL FILL_6__3498_ (
);

FILL FILL_6__3078_ (
);

FILL FILL_0__3472_ (
);

FILL FILL_0__3052_ (
);

FILL FILL_7__2874_ (
);

FILL FILL_7__2454_ (
);

FILL FILL_7__2034_ (
);

FILL FILL_3__2774_ (
);

FILL FILL_3__2354_ (
);

FILL FILL_7__3659_ (
);

FILL FILL_5__3641_ (
);

FILL FILL_5__3221_ (
);

FILL FILL168750x57750 (
);

FILL FILL_1__3633_ (
);

FILL FILL_1__3213_ (
);

FILL FILL_3__3559_ (
);

FILL FILL_3__3139_ (
);

FILL FILL_6__1984_ (
);

NAND3X1 _2283_ (
    .A(_1364_),
    .B(_1390_),
    .C(_1354_),
    .Y(_1391_)
);

FILL FILL_2__1976_ (
);

FILL FILL_3_BUFX2_insert10 (
);

FILL FILL_3_BUFX2_insert11 (
);

FILL FILL_3_BUFX2_insert12 (
);

FILL FILL_3_BUFX2_insert13 (
);

FILL FILL_3_BUFX2_insert14 (
);

FILL FILL_3_BUFX2_insert15 (
);

FILL FILL_3_BUFX2_insert16 (
);

FILL FILL_3_BUFX2_insert17 (
);

FILL FILL_4__2843_ (
);

FILL FILL_3_BUFX2_insert18 (
);

FILL FILL_3_BUFX2_insert19 (
);

FILL FILL_4__2423_ (
);

FILL FILL_4__2003_ (
);

FILL FILL_6__2769_ (
);

NAND2X1 _3488_ (
    .A(alu_shift_right),
    .B(AI[6]),
    .Y(_1733_)
);

FILL FILL_6__2349_ (
);

NOR2X1 _3068_ (
    .A(_431_),
    .B(_988_),
    .Y(_681_)
);

FILL FILL_0__2743_ (
);

FILL FILL_6__3710_ (
);

FILL FILL_0__2323_ (
);

FILL FILL_2__3702_ (
);

FILL FILL_4__3628_ (
);

FILL FILL_4__3208_ (
);

FILL FILL_0__3528_ (
);

FILL FILL_0__3108_ (
);

FILL FILL_5__2912_ (
);

FILL FILL_2__2094_ (
);

FILL FILL_1__2904_ (
);

INVX1 _1974_ (
    .A(_1089_),
    .Y(_1090_)
);

FILL FILL_2__3299_ (
);

FILL FILL_0__3281_ (
);

NOR2X1 _2759_ (
    .A(_404_),
    .B(_407_),
    .Y(_425_)
);

OAI21X1 _2339_ (
    .A(write_back),
    .B(_1241_),
    .C(_1243_),
    .Y(_1446_)
);

FILL FILL_7__2683_ (
);

FILL FILL_7__2263_ (
);

BUFX2 _3700_ (
    .A(_1741_[3]),
    .Y(AB[3])
);

FILL FILL_3__2583_ (
);

FILL FILL_3__2163_ (
);

FILL FILL_5__2089_ (
);

FILL FILL_5__3450_ (
);

FILL FILL_7__3048_ (
);

FILL FILL_5__3030_ (
);

FILL FILL_1__3022_ (
);

FILL FILL_6__1793_ (
);

NOR2X1 _2092_ (
    .A(_902__bF$buf3),
    .B(_938_),
    .Y(_1201_)
);

FILL FILL_2__1785_ (
);

FILL FILL_4__2652_ (
);

FILL FILL_4__2232_ (
);

FILL FILL_6__2998_ (
);

FILL FILL_6__2578_ (
);

NAND2X1 _3297_ (
    .A(ABL[6]),
    .B(_860_),
    .Y(_867_)
);

FILL FILL_6__2158_ (
);

FILL FILL_0__2972_ (
);

FILL FILL_0__2552_ (
);

FILL FILL_0__2132_ (
);

FILL FILL_2__3511_ (
);

FILL FILL_4__3017_ (
);

FILL FILL_3__1854_ (
);

FILL FILL_5__2721_ (
);

FILL FILL_7__2319_ (
);

FILL FILL_5__2301_ (
);

FILL FILL_1__2713_ (
);

FILL FILL_3__2639_ (
);

FILL FILL_3__2219_ (
);

OAI21X1 _1783_ (
    .A(_900_),
    .B(_908_),
    .C(_903__bF$buf0),
    .Y(_909_)
);

FILL FILL_4__3190_ (
);

FILL FILL_5__3506_ (
);

FILL FILL_0__3090_ (
);

FILL FILL_4__1923_ (
);

FILL FILL_6__1849_ (
);

OAI21X1 _2988_ (
    .A(_578_),
    .B(_553_),
    .C(_617_),
    .Y(_618_)
);

INVX1 _2568_ (
    .A(_257_),
    .Y(_1741_[5])
);

NOR2X1 _2148_ (
    .A(_902__bF$buf3),
    .B(_1069_),
    .Y(_1257_)
);

FILL FILL_7__2072_ (
);

FILL FILL_0__1823_ (
);

FILL FILL_3__2392_ (
);

FILL FILL_4__2708_ (
);

FILL FILL_7__3697_ (
);

FILL FILL_7__3277_ (
);

FILL FILL_0__2608_ (
);

FILL FILL_1__3671_ (
);

FILL FILL_1__3251_ (
);

FILL FILL_3__3597_ (
);

FILL FILL_3__3177_ (
);

FILL FILL_4__2881_ (
);

FILL FILL_4__2461_ (
);

FILL FILL_4__2041_ (
);

FILL FILL_6__2387_ (
);

FILL FILL_2__2799_ (
);

FILL FILL_0__2781_ (
);

FILL FILL_0__2361_ (
);

FILL FILL_2__2379_ (
);

OAI21X1 _1839_ (
    .A(_894_),
    .B(_919_),
    .C(_964_),
    .Y(CI)
);

FILL FILL_4__3666_ (
);

FILL FILL_7__1763_ (
);

FILL FILL_4__3246_ (
);

FILL FILL_0__3566_ (
);

FILL FILL_0__3146_ (
);

FILL FILL_4_BUFX2_insert60 (
);

FILL FILL_4_BUFX2_insert61 (
);

FILL FILL_4_BUFX2_insert62 (
);

FILL FILL_4_BUFX2_insert63 (
);

FILL FILL_4_BUFX2_insert64 (
);

FILL FILL_4_BUFX2_insert65 (
);

FILL FILL_4_BUFX2_insert66 (
);

FILL FILL_4_BUFX2_insert67 (
);

FILL FILL_4_BUFX2_insert68 (
);

FILL FILL_5__2950_ (
);

FILL FILL_4_BUFX2_insert69 (
);

FILL FILL_7__2548_ (
);

FILL FILL_5__2530_ (
);

FILL FILL_5__2110_ (
);

FILL FILL_1__2942_ (
);

FILL FILL_1__2522_ (
);

FILL FILL_1__2102_ (
);

FILL FILL_3__2868_ (
);

FILL FILL_3__2448_ (
);

FILL FILL_3__2028_ (
);

FILL FILL_5__3315_ (
);

FILL FILL_1__3307_ (
);

AOI21X1 _2797_ (
    .A(ADD[4]),
    .B(_1299_),
    .C(_1334_),
    .Y(_460_)
);

NOR2X1 _2377_ (
    .A(_1391_),
    .B(_1482_),
    .Y(_1483_)
);

FILL FILL_4__2937_ (
);

FILL FILL_4__2517_ (
);

FILL FILL_7__3086_ (
);

FILL FILL_0__2837_ (
);

FILL FILL_0__2417_ (
);

FILL FILL_1__3480_ (
);

FILL FILL_1__3060_ (
);

FILL FILL_7__1819_ (
);

FILL FILL_5__1801_ (
);

FILL FILL_4__2690_ (
);

FILL FILL_4__2270_ (
);

FILL FILL_6__2196_ (
);

FILL FILL_0__2590_ (
);

FILL FILL_2__2188_ (
);

FILL FILL_0__2170_ (
);

FILL FILL_7__1992_ (
);

FILL FILL_4__3475_ (
);

FILL FILL_4__3055_ (
);

FILL FILL_3__1892_ (
);

FILL FILL_7__2777_ (
);

FILL FILL_1__2751_ (
);

FILL FILL_1__2331_ (
);

FILL FILL_3__2677_ (
);

FILL FILL_3__2257_ (
);

FILL FILL_5__3544_ (
);

FILL FILL_5__3124_ (
);

FILL FILL_1__3536_ (
);

FILL FILL_1__3116_ (
);

FILL FILL_4__1961_ (
);

FILL FILL_6__1887_ (
);

NAND2X1 _2186_ (
    .A(CO),
    .B(backwards),
    .Y(_1295_)
);

FILL FILL_2__1879_ (
);

FILL FILL_0__1861_ (
);

FILL FILL_2__2820_ (
);

FILL FILL_2__2400_ (
);

FILL FILL_4__2746_ (
);

FILL FILL_4__2326_ (
);

FILL FILL_0__2646_ (
);

FILL FILL_6__3613_ (
);

FILL FILL_0__2226_ (
);

FILL FILL_2__3605_ (
);

FILL FILL_3__1948_ (
);

FILL FILL_5__2815_ (
);

FILL FILL_1__2807_ (
);

NAND3X1 _1877_ (
    .A(_996_),
    .B(_997_),
    .C(_1001_),
    .Y(_1002_)
);

FILL FILL_4__3284_ (
);

FILL FILL_0__3184_ (
);

FILL FILL_7__2166_ (
);

FILL FILL_0__1917_ (
);

INVX1 _3603_ (
    .A(_1632_),
    .Y(_1633_)
);

FILL FILL_1__2980_ (
);

FILL FILL_1__2560_ (
);

FILL FILL_1__2140_ (
);

FILL FILL_3__2486_ (
);

FILL FILL_3__2066_ (
);

FILL FILL_4__1770_ (
);

FILL FILL_4__2975_ (
);

FILL FILL_4__2555_ (
);

FILL FILL_4__2135_ (
);

FILL FILL_0__2875_ (
);

FILL FILL_0__2455_ (
);

FILL FILL_0__2035_ (
);

FILL FILL_6__3002_ (
);

FILL FILL_1__1831_ (
);

FILL FILL_3__1757_ (
);

FILL FILL_5__2624_ (
);

FILL FILL_5__2204_ (
);

FILL FILL_1__2616_ (
);

FILL FILL_4__3093_ (
);

FILL FILL_2__1900_ (
);

FILL FILL_4__1826_ (
);

FILL FILL_7__2395_ (
);

DFFSR _3412_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_81_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[1] [4])
);

FILL FILL_3__2295_ (
);

FILL FILL_5__3582_ (
);

FILL FILL_5__3162_ (
);

FILL FILL_1__3574_ (
);

FILL FILL_1__3154_ (
);

FILL FILL168750x118950 (
);

FILL FILL_4__2784_ (
);

FILL FILL_4__2364_ (
);

FILL FILL_0__2684_ (
);

FILL FILL_6__3651_ (
);

FILL FILL_0__2264_ (
);

FILL FILL_6__3231_ (
);

FILL FILL_2__3643_ (
);

FILL FILL_2__3223_ (
);

FILL FILL_4__3569_ (
);

FILL FILL_4__3149_ (
);

FILL FILL_3__1986_ (
);

FILL FILL_0__3469_ (
);

FILL FILL_0__3049_ (
);

FILL FILL_5__2853_ (
);

FILL FILL_5__2433_ (
);

FILL FILL_5__2013_ (
);

FILL FILL_1__2845_ (
);

FILL FILL_1__2425_ (
);

FILL FILL_1__2005_ (
);

FILL FILL_3__3712_ (
);

FILL FILL_5__3638_ (
);

FILL FILL_5__3218_ (
);

FILL FILL_0__1955_ (
);

FILL FILL_6__2922_ (
);

AOI22X1 _3641_ (
    .A(_1533_),
    .B(_1535_),
    .C(_1669_),
    .D(_1670_),
    .Y(_1671_)
);

FILL FILL_6__2502_ (
);

NOR2X1 _3221_ (
    .A(\AXYS[2] [7]),
    .B(_798_),
    .Y(_806_)
);

FILL FILL_2__2914_ (
);

FILL FILL_6__3707_ (
);

FILL FILL_4__2593_ (
);

FILL FILL_4__2173_ (
);

FILL FILL_6__2099_ (
);

FILL FILL_5__2909_ (
);

FILL FILL_0__2493_ (
);

FILL FILL_6__3460_ (
);

FILL FILL_0__2073_ (
);

FILL FILL_6__3040_ (
);

FILL FILL169050x57750 (
);

FILL FILL_2__3452_ (
);

FILL FILL_2__3032_ (
);

FILL FILL_7__1895_ (
);

OAI21X1 _2912_ (
    .A(_886__bF$buf5),
    .B(_1027__bF$buf2),
    .C(bit_ins),
    .Y(_558_)
);

FILL FILL_0__3698_ (
);

FILL FILL_3__1795_ (
);

FILL FILL_0__3278_ (
);

FILL FILL_5__2662_ (
);

FILL FILL_5__2242_ (
);

FILL FILL_1__2654_ (
);

FILL FILL_7__3621_ (
);

FILL FILL_1__2234_ (
);

FILL FILL_7__3201_ (
);

FILL FILL_3__3521_ (
);

FILL FILL_3__3101_ (
);

FILL FILL_5__3027_ (
);

FILL FILL_1__3019_ (
);

FILL FILL_4__1864_ (
);

NAND2X1 _2089_ (
    .A(_1197_),
    .B(_1192_),
    .Y(_1198_)
);

FILL FILL_0__1764_ (
);

FILL FILL_6__2731_ (
);

NOR2X1 _3450_ (
    .A(ADD[5]),
    .B(ADD[4]),
    .Y(_1699_)
);

FILL FILL_6__2311_ (
);

OAI21X1 _3030_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[3]),
    .Y(_651_)
);

FILL FILL_2__2723_ (
);

FILL FILL_2__2303_ (
);

FILL FILL_4__2649_ (
);

FILL FILL_4__2229_ (
);

FILL FILL_0__2969_ (
);

FILL FILL_0__2549_ (
);

FILL FILL_6__3516_ (
);

FILL FILL_0__2129_ (
);

FILL FILL_1__3192_ (
);

FILL FILL_2__3508_ (
);

FILL FILL_5__1933_ (
);

FILL FILL_1__1925_ (
);

FILL FILL_5__2718_ (
);

FILL FILL_2__3261_ (
);

FILL FILL_4__3187_ (
);

OAI21X1 _2721_ (
    .A(_389_),
    .B(_378_),
    .C(_148_),
    .Y(_390_)
);

AND2X2 _2301_ (
    .A(_1403_),
    .B(_1407_),
    .Y(_1408_)
);

FILL FILL_0__3087_ (
);

FILL FILL_5__2891_ (
);

FILL FILL_5__2471_ (
);

FILL FILL_7__2069_ (
);

FILL FILL_5__2051_ (
);

NAND2X1 _3506_ (
    .A(_1535_),
    .B(_1533_),
    .Y(_1536_)
);

FILL FILL_1__2883_ (
);

FILL FILL_1__2463_ (
);

FILL FILL_1__2043_ (
);

FILL FILL_3__2389_ (
);

FILL FILL_5__3676_ (
);

FILL FILL_5__3256_ (
);

FILL FILL_1__3668_ (
);

FILL FILL_1__3248_ (
);

FILL FILL_0__1993_ (
);

FILL FILL_6__2960_ (
);

FILL FILL_6__2540_ (
);

FILL FILL_6__2120_ (
);

FILL FILL_2__2952_ (
);

FILL FILL_2__2532_ (
);

FILL FILL_2__2112_ (
);

FILL FILL_4__2878_ (
);

FILL FILL_4__2458_ (
);

FILL FILL_4__2038_ (
);

FILL FILL_0__2778_ (
);

FILL FILL_0__2358_ (
);

FILL FILL_2__3317_ (
);

FILL FILL_7__2701_ (
);

FILL FILL_3__2601_ (
);

FILL FILL_5__2947_ (
);

FILL FILL_5__2527_ (
);

FILL FILL_5__2107_ (
);

FILL FILL_1__2939_ (
);

FILL FILL_1__2519_ (
);

FILL FILL_2__3490_ (
);

FILL FILL_2__3070_ (
);

NOR2X1 _2950_ (
    .A(_1185_),
    .B(_1149__bF$buf4),
    .Y(_589_)
);

FILL FILL_6__1811_ (
);

AOI21X1 _2530_ (
    .A(_1059_),
    .B(_195_),
    .C(_224_),
    .Y(_225_)
);

OAI22X1 _2110_ (
    .A(_1216_),
    .B(_1218_),
    .C(_1213_),
    .D(_1215_),
    .Y(_1219_)
);

FILL FILL_2__1803_ (
);

FILL FILL_5__2280_ (
);

FILL FILL_7__2298_ (
);

OAI21X1 _3315_ (
    .A(_1134_),
    .B(_869_),
    .C(_876_),
    .Y(_115_)
);

FILL FILL_1__2692_ (
);

FILL FILL_1__2272_ (
);

FILL FILL_3__2198_ (
);

FILL FILL_5__3485_ (
);

FILL FILL_5__3065_ (
);

FILL FILL_1__3477_ (
);

FILL FILL_1__3057_ (
);

FILL FILL_2__2761_ (
);

FILL FILL_2__2341_ (
);

FILL FILL_4__2687_ (
);

FILL FILL_4__2267_ (
);

NOR2X1 _1801_ (
    .A(state[1]),
    .B(state[0]),
    .Y(_927_)
);

FILL FILL_0__2587_ (
);

FILL FILL_6__3554_ (
);

FILL FILL_0__2167_ (
);

FILL FILL_6__3134_ (
);

FILL FILL_2__3546_ (
);

FILL FILL_2__3126_ (
);

FILL FILL_5__1971_ (
);

FILL FILL_1__1963_ (
);

FILL FILL_7__2930_ (
);

FILL FILL_3__1889_ (
);

FILL FILL_3__2830_ (
);

FILL FILL_3__2410_ (
);

FILL FILL_5__2756_ (
);

FILL FILL_5__2336_ (
);

FILL FILL_1__2748_ (
);

FILL FILL_7__3715_ (
);

FILL FILL_1__2328_ (
);

FILL FILL_3__3615_ (
);

FILL FILL_4__1958_ (
);

FILL FILL_0__1858_ (
);

FILL FILL_6__2825_ (
);

AOI22X1 _3544_ (
    .A(BI[0]),
    .B(_1573_),
    .C(_1717_),
    .D(_1572_),
    .Y(_1574_)
);

FILL FILL_6__2405_ (
);

NOR2X1 _3124_ (
    .A(HC),
    .B(_728_),
    .Y(_731_)
);

FILL FILL_1__2081_ (
);

FILL FILL_2__2817_ (
);

FILL FILL_5__3294_ (
);

FILL FILL_1__3286_ (
);

FILL FILL169650x7350 (
);

FILL FILL_2__2990_ (
);

FILL FILL_2__2570_ (
);

FILL FILL_2__2150_ (
);

FILL FILL_4__2496_ (
);

FILL FILL_4__2076_ (
);

FILL FILL_0__2396_ (
);

FILL FILL_7__1798_ (
);

FILL FILL_5__1780_ (
);

OAI21X1 _2815_ (
    .A(_365_),
    .B(_477_),
    .C(_471_),
    .Y(_478_)
);

FILL FILL_1__1772_ (
);

FILL FILL_5__2985_ (
);

FILL FILL_5__2565_ (
);

FILL FILL_5__2145_ (
);

FILL FILL_1__2977_ (
);

FILL FILL_1__2557_ (
);

FILL FILL_7__3524_ (
);

FILL FILL_1__2137_ (
);

FILL FILL_7__3104_ (
);

FILL FILL_3__3004_ (
);

FILL FILL_2__1841_ (
);

FILL FILL_4__1767_ (
);

FILL FILL_6__2634_ (
);

DFFSR _3353_ (
    .R(_1__bF$buf2),
    .S(vdd),
    .D(_30_),
    .CLK(clk_bF$buf10),
    .Q(clv)
);

FILL FILL_6__2214_ (
);

FILL FILL_2__2626_ (
);

FILL FILL_2__2206_ (
);

FILL FILL_1__3095_ (
);

FILL FILL_3__1910_ (
);

FILL FILL_5__1836_ (
);

FILL FILL_1__1828_ (
);

FILL FILL_6__3592_ (
);

FILL FILL_6__3172_ (
);

FILL FILL_2__3584_ (
);

FILL FILL_2__3164_ (
);

FILL FILL_6__1905_ (
);

INVX1 _2624_ (
    .A(PC[15]),
    .Y(_304_)
);

OAI21X1 _2204_ (
    .A(_914__bF$buf1),
    .B(_1075_),
    .C(RDY_bF$buf1),
    .Y(_1313_)
);

FILL FILL_5__2794_ (
);

FILL FILL_5__2374_ (
);

DFFSR _3409_ (
    .R(_1__bF$buf10),
    .S(vdd),
    .D(_78_),
    .CLK(clk_bF$buf8),
    .Q(\AXYS[1] [1])
);

FILL FILL_1__2786_ (
);

FILL FILL_1__2366_ (
);

FILL FILL_3__3653_ (
);

FILL FILL_3__3233_ (
);

FILL FILL_5__3579_ (
);

FILL FILL_5__3159_ (
);

FILL FILL_4__1996_ (
);

FILL FILL_0__1896_ (
);

FILL FILL_6__2863_ (
);

INVX1 _3582_ (
    .A(_1586_),
    .Y(_1612_)
);

FILL FILL_6__2443_ (
);

FILL FILL_6__2023_ (
);

INVX1 _3162_ (
    .A(_764_),
    .Y(_765_)
);

FILL FILL_2__2855_ (
);

FILL FILL_2__2435_ (
);

FILL FILL_2__2015_ (
);

FILL FILL_4__3302_ (
);

FILL FILL_6__3648_ (
);

FILL FILL_6__3228_ (
);

FILL FILL_0__3622_ (
);

FILL FILL_0__3202_ (
);

FILL FILL_7__2604_ (
);

FILL FILL_3__2924_ (
);

FILL FILL_3__2504_ (
);

FILL FILL_3__3709_ (
);

NOR3X1 _2853_ (
    .A(_456_),
    .B(_508_),
    .C(_401_),
    .Y(_513_)
);

AOI22X1 _2433_ (
    .A(backwards),
    .B(_925_),
    .C(_915_),
    .D(op[2]),
    .Y(_139_)
);

INVX1 _2013_ (
    .A(_1124_),
    .Y(_1125_)
);

FILL FILL_0_BUFX2_insert0 (
);

FILL FILL_0_BUFX2_insert1 (
);

FILL FILL_0_BUFX2_insert2 (
);

FILL FILL_0_BUFX2_insert3 (
);

FILL FILL_0_BUFX2_insert4 (
);

FILL FILL_0_BUFX2_insert5 (
);

FILL FILL_0_BUFX2_insert6 (
);

FILL FILL_0_BUFX2_insert7 (
);

FILL FILL_0_BUFX2_insert8 (
);

FILL FILL_0_BUFX2_insert9 (
);

FILL FILL_5__2183_ (
);

FILL FILL_6__2919_ (
);

OAI21X1 _3638_ (
    .A(_1545_),
    .B(_1549_),
    .C(_1625_),
    .Y(_1668_)
);

AOI21X1 _3218_ (
    .A(_767_),
    .B(_798_),
    .C(_804_),
    .Y(_90_)
);

FILL FILL_1__2595_ (
);

FILL FILL_1__2175_ (
);

FILL FILL_3__3462_ (
);

FILL FILL_3__3042_ (
);

FILL FILL_6__2672_ (
);

DFFPOSX1 _3391_ (
    .D(_60_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD[7])
);

FILL FILL_6__2252_ (
);

FILL FILL_2__2664_ (
);

FILL FILL_2__2244_ (
);

FILL FILL_4__3531_ (
);

FILL FILL_4__3111_ (
);

FILL FILL_6__3457_ (
);

FILL FILL_6__3037_ (
);

FILL FILL_2__3449_ (
);

FILL FILL_2__3029_ (
);

FILL FILL_0__3011_ (
);

FILL FILL_5__1874_ (
);

NAND3X1 _2909_ (
    .A(_1185_),
    .B(_1412_),
    .C(_1181_),
    .Y(_555_)
);

FILL FILL_1__1866_ (
);

FILL FILL_7__2833_ (
);

FILL FILL_3__2733_ (
);

FILL FILL_3__2313_ (
);

FILL FILL_5__2659_ (
);

FILL FILL_5__2239_ (
);

FILL FILL_5__3600_ (
);

FILL FILL_3__3518_ (
);

FILL FILL_6__1943_ (
);

OAI21X1 _2662_ (
    .A(res),
    .B(_148_),
    .C(_335_),
    .Y(_336_)
);

NOR2X1 _2242_ (
    .A(_1188_),
    .B(_1349_),
    .Y(_1350_)
);

FILL FILL_2__1935_ (
);

FILL FILL_4__2802_ (
);

FILL FILL_6__2728_ (
);

DFFSR _3447_ (
    .R(_1__bF$buf0),
    .S(vdd),
    .D(_115_),
    .CLK(clk_bF$buf0),
    .Q(ABH[6])
);

FILL FILL_6__2308_ (
);

OAI21X1 _3027_ (
    .A(_1006_),
    .B(_647_),
    .C(_649_),
    .Y(_54_)
);

FILL FILL_0__2702_ (
);

FILL FILL_3__3691_ (
);

FILL FILL_3__3271_ (
);

FILL FILL_5__3197_ (
);

FILL FILL_1__3189_ (
);

FILL FILL_6__2481_ (
);

FILL FILL_6__2061_ (
);

FILL FILL_2__2893_ (
);

FILL FILL_2__2473_ (
);

FILL FILL_2__2053_ (
);

FILL FILL_4__2399_ (
);

AOI22X1 _1933_ (
    .A(\AXYS[3] [0]),
    .B(_1049_),
    .C(_1047_),
    .D(\AXYS[1] [0]),
    .Y(_1050_)
);

FILL FILL_0__2299_ (
);

FILL FILL_6__3266_ (
);

FILL FILL169950x104550 (
);

FILL FILL_0__3660_ (
);

FILL FILL_2__3678_ (
);

FILL FILL_0__3240_ (
);

FILL FILL_2__3258_ (
);

NAND3X1 _2718_ (
    .A(RDY_bF$buf0),
    .B(_387_),
    .C(_383_),
    .Y(_388_)
);

FILL FILL_7__2222_ (
);

FILL FILL_3__2962_ (
);

FILL FILL_3__2542_ (
);

FILL FILL_3__2122_ (
);

FILL FILL_5__2888_ (
);

FILL FILL_5__2468_ (
);

FILL FILL_5__2048_ (
);

FILL FILL_7__3007_ (
);

FILL FILL_6__1752_ (
);

OAI21X1 _2891_ (
    .A(_886__bF$buf5),
    .B(_1027__bF$buf2),
    .C(cld),
    .Y(_542_)
);

OAI21X1 _2471_ (
    .A(_143_),
    .B(_1109_),
    .C(_170_),
    .Y(_1742_[3])
);

NAND2X1 _2051_ (
    .A(_1156_),
    .B(_1159_),
    .Y(_1160_)
);

FILL FILL_2__1744_ (
);

FILL FILL_4__2611_ (
);

FILL FILL_6__2957_ (
);

OAI21X1 _3676_ (
    .A(_1707_),
    .B(RDY_bF$buf7),
    .C(_1696_),
    .Y(_1524_)
);

FILL FILL_6__2537_ (
);

FILL FILL_6__2117_ (
);

OAI21X1 _3256_ (
    .A(_931__bF$buf2),
    .B(_942_),
    .C(_974_),
    .Y(_832_)
);

FILL FILL_7__3180_ (
);

FILL FILL_2__2949_ (
);

FILL FILL_0__2931_ (
);

FILL FILL_2__2529_ (
);

FILL FILL_0__2511_ (
);

FILL FILL_2__2109_ (
);

FILL FILL_3__3080_ (
);

FILL FILL_7__1913_ (
);

FILL FILL_3__1813_ (
);

FILL FILL_6__2290_ (
);

FILL FILL_2__2282_ (
);

FILL FILL_6__3495_ (
);

FILL FILL_6__3075_ (
);

FILL FILL_0_BUFX2_insert80 (
);

FILL FILL_0_BUFX2_insert81 (
);

FILL FILL_0_BUFX2_insert82 (
);

FILL FILL_2__3487_ (
);

FILL FILL_0_BUFX2_insert83 (
);

FILL FILL_2__3067_ (
);

OAI21X1 _2947_ (
    .A(_1212_),
    .B(_1327_),
    .C(_540_),
    .Y(_588_)
);

FILL FILL_6__1808_ (
);

AOI21X1 _2527_ (
    .A(_216_),
    .B(ADD[0]),
    .C(_221_),
    .Y(_222_)
);

NAND2X1 _2107_ (
    .A(_1159_),
    .B(_1164_),
    .Y(_1216_)
);

FILL FILL_7__2451_ (
);

FILL FILL_3__2771_ (
);

FILL FILL_3__2351_ (
);

FILL FILL_5__2697_ (
);

FILL FILL_5__2277_ (
);

FILL FILL_1__2689_ (
);

FILL FILL_7__3656_ (
);

FILL FILL_1__2269_ (
);

FILL FILL_7__3236_ (
);

FILL FILL_1__3630_ (
);

FILL FILL_1__3210_ (
);

FILL FILL_3__3556_ (
);

FILL FILL_3__3136_ (
);

FILL FILL_6__1981_ (
);

AOI21X1 _2280_ (
    .A(_1383_),
    .B(_1384_),
    .C(_1387_),
    .Y(_1388_)
);

FILL FILL_2__1973_ (
);

FILL FILL_4__1899_ (
);

FILL FILL_4__2840_ (
);

FILL FILL_4__2420_ (
);

FILL FILL_4__2000_ (
);

FILL FILL_0__1799_ (
);

FILL FILL_6__2766_ (
);

NAND2X1 _3485_ (
    .A(\u_ALU8.BI7 ),
    .B(_1714__bF$buf2),
    .Y(_1731_)
);

FILL FILL_6__2346_ (
);

NAND2X1 _3065_ (
    .A(_548_),
    .B(_677_),
    .Y(_678_)
);

FILL FILL_2__2758_ (
);

FILL FILL_0__2740_ (
);

FILL FILL_2__2338_ (
);

FILL FILL_0__2320_ (
);

FILL FILL_4__3625_ (
);

FILL FILL_4__3205_ (
);

FILL FILL_0__3525_ (
);

FILL FILL_0__3105_ (
);

FILL FILL_5__1968_ (
);

FILL FILL_7__2927_ (
);

FILL FILL_2__2091_ (
);

FILL FILL_1__2901_ (
);

FILL FILL_3__2827_ (
);

FILL FILL_3__2407_ (
);

AOI22X1 _1971_ (
    .A(_1049_),
    .B(\AXYS[3] [1]),
    .C(\AXYS[2] [1]),
    .D(_1057_),
    .Y(_1087_)
);

FILL FILL_2__3296_ (
);

AOI21X1 _2756_ (
    .A(DIMUX[1]),
    .B(_419_),
    .C(_421_),
    .Y(_422_)
);

INVX1 _2336_ (
    .A(_1442_),
    .Y(_1443_)
);

FILL FILL_7__2680_ (
);

FILL FILL_3__2580_ (
);

FILL FILL_3__2160_ (
);

FILL FILL_5__2086_ (
);

FILL FILL_2_BUFX2_insert0 (
);

FILL FILL_1__2498_ (
);

FILL FILL_2_BUFX2_insert1 (
);

FILL FILL_2_BUFX2_insert2 (
);

FILL FILL_1__2078_ (
);

FILL FILL_7__3045_ (
);

FILL FILL_2_BUFX2_insert3 (
);

FILL FILL_2_BUFX2_insert4 (
);

FILL FILL_2_BUFX2_insert5 (
);

FILL FILL_2_BUFX2_insert6 (
);

FILL FILL_2_BUFX2_insert7 (
);

FILL FILL_2_BUFX2_insert8 (
);

FILL FILL_2_BUFX2_insert9 (
);

FILL FILL_6__1790_ (
);

FILL FILL_2__1782_ (
);

FILL FILL_6__2995_ (
);

FILL FILL_6__2575_ (
);

OAI21X1 _3294_ (
    .A(_860_),
    .B(_249_),
    .C(_865_),
    .Y(_105_)
);

FILL FILL_6__2155_ (
);

FILL FILL_2__2987_ (
);

FILL FILL_2__2567_ (
);

FILL FILL_2__2147_ (
);

FILL FILL_7__1951_ (
);

FILL FILL_4__3014_ (
);

FILL FILL_3__1851_ (
);

FILL FILL_5__1777_ (
);

FILL FILL_1__1769_ (
);

FILL FILL_7__2316_ (
);

FILL FILL_1__2710_ (
);

FILL FILL_3__2636_ (
);

FILL FILL_3__2216_ (
);

INVX1 _1780_ (
    .A(state[0]),
    .Y(_906_)
);

FILL FILL_5__3503_ (
);

FILL FILL_4__1920_ (
);

FILL FILL_6__1846_ (
);

INVX1 _2985_ (
    .A(_614_),
    .Y(_615_)
);

INVX1 _2565_ (
    .A(_254_),
    .Y(_255_)
);

AOI22X1 _2145_ (
    .A(_886__bF$buf1),
    .B(_1063_),
    .C(_1253_),
    .D(_1150__bF$buf3),
    .Y(_1254_)
);

FILL FILL_2__1838_ (
);

FILL FILL_0__1820_ (
);

FILL FILL_4__2705_ (
);

FILL FILL_7__3694_ (
);

FILL FILL_0__2605_ (
);

FILL FILL_3__3594_ (
);

FILL FILL_3__3174_ (
);

FILL FILL_3__1907_ (
);

FILL FILL_6__2384_ (
);

FILL FILL_2__2796_ (
);

FILL FILL_2__2376_ (
);

NOR2X1 _1836_ (
    .A(_961_),
    .B(_945_),
    .Y(_962_)
);

FILL FILL_4__3663_ (
);

FILL FILL_4__3243_ (
);

FILL FILL_6__3589_ (
);

FILL FILL_6__3169_ (
);

FILL FILL_0__3563_ (
);

FILL FILL_0__3143_ (
);

FILL FILL_4_BUFX2_insert37 (
);

FILL FILL_1__1998_ (
);

FILL FILL_4_BUFX2_insert38 (
);

FILL FILL_4_BUFX2_insert39 (
);

FILL FILL_7__2545_ (
);

FILL FILL_7__2125_ (
);

FILL FILL_3__2865_ (
);

FILL FILL_3__2445_ (
);

FILL FILL_3__2025_ (
);

FILL FILL_5__3312_ (
);

FILL FILL_1__3304_ (
);

OAI22X1 _2794_ (
    .A(RDY_bF$buf4),
    .B(_285_),
    .C(_457_),
    .D(_452_),
    .Y(_13_)
);

INVX1 _2374_ (
    .A(_1479_),
    .Y(_1480_)
);

FILL FILL_4__2934_ (
);

FILL FILL_4__2514_ (
);

NAND2X1 _3579_ (
    .A(_1599_),
    .B(_1595_),
    .Y(_1609_)
);

INVX1 _3159_ (
    .A(_759_),
    .Y(_762_)
);

FILL FILL_7__3083_ (
);

FILL FILL_0__2834_ (
);

FILL FILL_0__2414_ (
);

FILL FILL_7__1816_ (
);

FILL FILL_0__3619_ (
);

FILL FILL_6__2193_ (
);

FILL FILL_2__2185_ (
);

FILL FILL_4__3472_ (
);

FILL FILL_4__3052_ (
);

FILL FILL_7__2774_ (
);

FILL FILL_7__2354_ (
);

FILL FILL_3__2674_ (
);

FILL FILL_3__2254_ (
);

FILL FILL_5__3541_ (
);

FILL FILL_7__3559_ (
);

FILL FILL_5__3121_ (
);

FILL FILL168450x3750 (
);

FILL FILL_1__3533_ (
);

FILL FILL_1__3113_ (
);

FILL FILL_3__3459_ (
);

FILL FILL_3__3039_ (
);

FILL FILL_6__1884_ (
);

NAND2X1 _2183_ (
    .A(_886__bF$buf4),
    .B(_1291_),
    .Y(_1292_)
);

FILL FILL_2__1876_ (
);

FILL FILL_4__2743_ (
);

FILL FILL_4__2323_ (
);

FILL FILL_6__2669_ (
);

DFFPOSX1 _3388_ (
    .D(_57_),
    .CLK(clk_bF$buf8),
    .Q(IRHOLD[4])
);

FILL FILL_6__2249_ (
);

FILL FILL_0__2643_ (
);

FILL FILL_6__3610_ (
);

FILL FILL_0__2223_ (
);

FILL FILL_2__3602_ (
);

FILL FILL_4__3528_ (
);

FILL FILL_4__3108_ (
);

FILL FILL_3__1945_ (
);

FILL FILL_0__3008_ (
);

FILL FILL_5__2812_ (
);

FILL FILL_1__2804_ (
);

OAI21X1 _1874_ (
    .A(_931__bF$buf0),
    .B(_958_),
    .C(_960_),
    .Y(_999_)
);

FILL FILL_4__3281_ (
);

FILL FILL_0__3181_ (
);

FILL FILL_2__3199_ (
);

OR2X2 _2659_ (
    .A(_333_),
    .B(_886__bF$buf3),
    .Y(_334_)
);

OR2X2 _2239_ (
    .A(_1290_),
    .B(RDY_bF$buf5),
    .Y(_1347_)
);

FILL FILL_7__2583_ (
);

FILL FILL_7__2163_ (
);

FILL FILL_0__1914_ (
);

OAI21X1 _3600_ (
    .A(_1629_),
    .B(_1626_),
    .C(_1536_),
    .Y(_1630_)
);

FILL FILL_3__2483_ (
);

FILL FILL_3__2063_ (
);

FILL FILL169950x61350 (
);

FILL FILL_3__3268_ (
);

FILL FILL_4_BUFX2_insert0 (
);

FILL FILL169950x28950 (
);

FILL FILL_4_BUFX2_insert1 (
);

FILL FILL_4_BUFX2_insert2 (
);

FILL FILL_4_BUFX2_insert3 (
);

FILL FILL_4_BUFX2_insert4 (
);

FILL FILL_4_BUFX2_insert5 (
);

FILL FILL_4_BUFX2_insert6 (
);

FILL FILL_4_BUFX2_insert7 (
);

FILL FILL_4_BUFX2_insert8 (
);

FILL FILL_4_BUFX2_insert9 (
);

FILL FILL_4__2972_ (
);

FILL FILL_4__2552_ (
);

FILL FILL_4__2132_ (
);

FILL FILL_6__2898_ (
);

FILL FILL_6__2478_ (
);

FILL FILL_6__2058_ (
);

OAI21X1 _3197_ (
    .A(_754_),
    .B(_789_),
    .C(_793_),
    .Y(_80_)
);

FILL FILL_0__2872_ (
);

FILL FILL_0__2452_ (
);

FILL FILL_0__2032_ (
);

FILL FILL_3__1754_ (
);

FILL FILL_0__3657_ (
);

FILL FILL_0__3237_ (
);

FILL FILL_5__2621_ (
);

FILL FILL_7__2219_ (
);

FILL FILL_5__2201_ (
);

FILL FILL_1__2613_ (
);

FILL FILL_3__2959_ (
);

FILL FILL_3__2539_ (
);

FILL FILL_3__2119_ (
);

FILL FILL_4__3090_ (
);

FILL FILL_4__1823_ (
);

FILL FILL_6__1749_ (
);

NOR2X1 _2888_ (
    .A(_1027__bF$buf2),
    .B(_526_),
    .Y(_540_)
);

AOI21X1 _2468_ (
    .A(ADD[3]),
    .B(_144_),
    .C(_167_),
    .Y(_168_)
);

INVX1 _2048_ (
    .A(IRHOLD[0]),
    .Y(_1157_)
);

FILL FILL_7__2392_ (
);

FILL FILL_3__2292_ (
);

FILL FILL_4__2608_ (
);

FILL FILL_7__3177_ (
);

FILL FILL_0__2928_ (
);

FILL FILL_0__2508_ (
);

FILL FILL_1__3571_ (
);

FILL FILL_1__3151_ (
);

FILL FILL_3__3497_ (
);

FILL FILL_3__3077_ (
);

FILL FILL_4__2781_ (
);

FILL FILL_4__2361_ (
);

FILL FILL_6__2287_ (
);

FILL FILL_2__2699_ (
);

FILL FILL_0__2681_ (
);

FILL FILL_2__2279_ (
);

FILL FILL_0__2261_ (
);

FILL FILL_2__3640_ (
);

FILL FILL_2__3220_ (
);

FILL FILL_4__3566_ (
);

FILL FILL_4__3146_ (
);

FILL FILL_3__1983_ (
);

FILL FILL_0__3466_ (
);

FILL FILL_0__3046_ (
);

FILL FILL_5__2850_ (
);

FILL FILL_7__2448_ (
);

FILL FILL_5__2430_ (
);

FILL FILL_5__2010_ (
);

FILL FILL_1__2842_ (
);

FILL FILL_1__2422_ (
);

FILL FILL_1__2002_ (
);

FILL FILL_3__2768_ (
);

FILL FILL_3__2348_ (
);

FILL FILL_5__3635_ (
);

FILL FILL_5__3215_ (
);

FILL FILL_1__3627_ (
);

FILL FILL_1__3207_ (
);

FILL FILL_6__1978_ (
);

INVX1 _2697_ (
    .A(_357_),
    .Y(_368_)
);

NOR2X1 _2277_ (
    .A(_886__bF$buf2),
    .B(_978_),
    .Y(_1385_)
);

FILL FILL_0__1952_ (
);

FILL FILL_2__2911_ (
);

FILL FILL_4__2837_ (
);

FILL FILL_4__2417_ (
);

FILL FILL_0__2737_ (
);

FILL FILL_0__2317_ (
);

FILL FILL_6__3704_ (
);

FILL FILL_4__2590_ (
);

FILL FILL_4__2170_ (
);

FILL FILL_6__2096_ (
);

FILL FILL_5__2906_ (
);

FILL FILL_0__2490_ (
);

FILL FILL_2__2088_ (
);

FILL FILL_0__2070_ (
);

AOI21X1 _1968_ (
    .A(_1082_),
    .B(ADD[0]),
    .C(_1084_),
    .Y(_1085_)
);

FILL FILL_7__1892_ (
);

FILL FILL_0__3695_ (
);

FILL FILL_3__1792_ (
);

FILL FILL_0__3275_ (
);

FILL FILL_7__2677_ (
);

FILL FILL_1__2651_ (
);

FILL FILL_1__2231_ (
);

FILL FILL_3__2997_ (
);

FILL FILL_3__2577_ (
);

FILL FILL_3__2157_ (
);

FILL FILL_5__3024_ (
);

FILL FILL_1__3016_ (
);

FILL FILL_4__1861_ (
);

FILL FILL_6__1787_ (
);

NAND2X1 _2086_ (
    .A(RDY_bF$buf8),
    .B(_1194_),
    .Y(_1195_)
);

FILL FILL_0__1761_ (
);

FILL FILL_2__1779_ (
);

FILL FILL169950x150 (
);

FILL FILL_2__2720_ (
);

FILL FILL_2__2300_ (
);

FILL FILL_4__2646_ (
);

FILL FILL_4__2226_ (
);

FILL FILL_0__2966_ (
);

FILL FILL_0__2546_ (
);

FILL FILL_6__3513_ (
);

FILL FILL_0__2126_ (
);

FILL FILL_2__3505_ (
);

FILL FILL_7__1948_ (
);

FILL FILL_5__1930_ (
);

FILL FILL_1__1922_ (
);

FILL FILL_3__1848_ (
);

FILL FILL_5__2715_ (
);

FILL FILL_1__2707_ (
);

INVX4 _1777_ (
    .A(_902__bF$buf0),
    .Y(_903_)
);

FILL FILL_4__3184_ (
);

FILL FILL_0__3084_ (
);

FILL FILL_4__1917_ (
);

FILL FILL_7__2066_ (
);

FILL FILL_0__1817_ (
);

OAI21X1 _3503_ (
    .A(_1532_),
    .B(_1531_),
    .C(_1528_),
    .Y(_1533_)
);

FILL FILL_1__2880_ (
);

FILL FILL_1__2460_ (
);

FILL FILL_1__2040_ (
);

FILL FILL_3__2386_ (
);

FILL FILL_5__3673_ (
);

FILL FILL_5__3253_ (
);

FILL FILL_1__3665_ (
);

FILL FILL_1__3245_ (
);

FILL FILL_0__1990_ (
);

FILL FILL_6_BUFX2_insert0 (
);

FILL FILL_6_BUFX2_insert1 (
);

FILL FILL_6_BUFX2_insert2 (
);

FILL FILL_6_BUFX2_insert3 (
);

FILL FILL_4__2875_ (
);

FILL FILL_4__2455_ (
);

FILL FILL_6_BUFX2_insert4 (
);

FILL FILL_6_BUFX2_insert5 (
);

FILL FILL_4__2035_ (
);

FILL FILL_6_BUFX2_insert6 (
);

FILL FILL_6_BUFX2_insert7 (
);

FILL FILL_6_BUFX2_insert8 (
);

FILL FILL_6_BUFX2_insert9 (
);

FILL FILL_0__2775_ (
);

FILL FILL_0__2355_ (
);

FILL FILL_2__3314_ (
);

FILL FILL167550x75750 (
);

FILL FILL_5__2944_ (
);

FILL FILL_5__2524_ (
);

FILL FILL_5__2104_ (
);

FILL FILL_1__2936_ (
);

FILL FILL_1__2516_ (
);

FILL FILL_5__3309_ (
);

FILL FILL_2__1800_ (
);

FILL FILL_7__2295_ (
);

NAND2X1 _3312_ (
    .A(_1741_[13]),
    .B(_869_),
    .Y(_875_)
);

FILL FILL_3__2195_ (
);

FILL FILL_5__3482_ (
);

FILL FILL_5__3062_ (
);

FILL FILL_1__3474_ (
);

FILL FILL_1__3054_ (
);

FILL FILL_5_CLKBUF1_insert26 (
);

FILL FILL_5_CLKBUF1_insert27 (
);

FILL FILL_5_CLKBUF1_insert28 (
);

FILL FILL_5_CLKBUF1_insert29 (
);

FILL FILL_4__2684_ (
);

FILL FILL_4__2264_ (
);

FILL FILL_0__2584_ (
);

FILL FILL_6__3551_ (
);

FILL FILL_0__2164_ (
);

FILL FILL_6__3131_ (
);

FILL FILL_2__3543_ (
);

FILL FILL_2__3123_ (
);

FILL FILL_4__3469_ (
);

FILL FILL_4__3049_ (
);

FILL FILL_1__1960_ (
);

FILL FILL_3__1886_ (
);

FILL FILL_5__2753_ (
);

FILL FILL_5__2333_ (
);

FILL FILL_1__2745_ (
);

FILL FILL_7__3712_ (
);

FILL FILL_1__2325_ (
);

FILL FILL_3__3612_ (
);

FILL FILL_5__3538_ (
);

FILL FILL_5__3118_ (
);

FILL FILL_4__1955_ (
);

FILL FILL_0__1855_ (
);

FILL FILL_6__2822_ (
);

OAI21X1 _3541_ (
    .A(_1728_),
    .B(_1570_),
    .C(_1568_),
    .Y(_1571_)
);

FILL FILL_6__2402_ (
);

NAND2X1 _3121_ (
    .A(adj_bcd),
    .B(_309_),
    .Y(_728_)
);

FILL FILL_2__2814_ (
);

FILL FILL_5__3291_ (
);

FILL FILL_6__3607_ (
);

FILL FILL_1__3283_ (
);

FILL FILL_4__2493_ (
);

FILL FILL_4__2073_ (
);

FILL FILL_5__2809_ (
);

FILL FILL_0__2393_ (
);

FILL FILL_4__3698_ (
);

FILL FILL_7__1795_ (
);

FILL FILL_4__3278_ (
);

AOI21X1 _2812_ (
    .A(ABH[1]),
    .B(_323_),
    .C(_474_),
    .Y(_475_)
);

FILL FILL_0__3598_ (
);

FILL FILL_0__3178_ (
);

FILL FILL_5__2982_ (
);

FILL FILL_5__2562_ (
);

FILL FILL_5__2142_ (
);

FILL FILL_1__2974_ (
);

FILL FILL_1__2554_ (
);

FILL FILL_7__3521_ (
);

FILL FILL_1__2134_ (
);

FILL FILL_7__3101_ (
);

FILL FILL_3__3001_ (
);

FILL FILL_4__1764_ (
);

FILL FILL_6__2631_ (
);

FILL FILL_6__2211_ (
);

DFFSR _3350_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_27_),
    .CLK(clk_bF$buf9),
    .Q(sed)
);

FILL FILL_2__2623_ (
);

FILL FILL_2__2203_ (
);

FILL FILL_4__2969_ (
);

FILL FILL_4__2549_ (
);

FILL FILL_4__2129_ (
);

FILL FILL_0__2869_ (
);

FILL FILL_0__2449_ (
);

FILL FILL_0__2029_ (
);

FILL FILL_1__3092_ (
);

FILL FILL_5__1833_ (
);

FILL FILL_1__1825_ (
);

FILL FILL_5__2618_ (
);

FILL FILL_2__3581_ (
);

FILL FILL_2__3161_ (
);

FILL FILL_4__3087_ (
);

FILL FILL_6__1902_ (
);

OAI21X1 _2621_ (
    .A(_1134_),
    .B(_270_),
    .C(_301_),
    .Y(_302_)
);

OAI21X1 _2201_ (
    .A(_931__bF$buf4),
    .B(_942_),
    .C(RDY_bF$buf1),
    .Y(_1310_)
);

FILL FILL_5__2791_ (
);

FILL FILL_5__2371_ (
);

DFFSR _3406_ (
    .R(_1__bF$buf3),
    .S(vdd),
    .D(_75_),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[0] [6])
);

FILL FILL_1__2783_ (
);

FILL FILL_1__2363_ (
);

FILL FILL_3__2289_ (
);

FILL FILL_3__3650_ (
);

FILL FILL_3__3230_ (
);

FILL FILL_5__3576_ (
);

FILL FILL_5__3156_ (
);

FILL FILL_1__3568_ (
);

FILL FILL_1__3148_ (
);

FILL FILL_4__1993_ (
);

FILL FILL_0__1893_ (
);

FILL FILL_6__2860_ (
);

FILL FILL_6__2440_ (
);

FILL FILL_6__2020_ (
);

FILL FILL_2__2852_ (
);

FILL FILL_2__2432_ (
);

FILL FILL_2__2012_ (
);

FILL FILL_4__2778_ (
);

FILL FILL_4__2358_ (
);

FILL FILL_0__2678_ (
);

FILL FILL_6__3645_ (
);

FILL FILL_0__2258_ (
);

FILL FILL_6__3225_ (
);

FILL FILL_2__3637_ (
);

FILL FILL_2__3217_ (
);

FILL FILL_7__2601_ (
);

FILL FILL_3__2921_ (
);

FILL FILL_3__2501_ (
);

FILL FILL_5__2847_ (
);

FILL FILL_5__2427_ (
);

FILL FILL_5__2007_ (
);

FILL FILL_1__2839_ (
);

FILL FILL_1__2419_ (
);

FILL FILL_3__3706_ (
);

NAND3X1 _2850_ (
    .A(RDY_bF$buf4),
    .B(_510_),
    .C(_507_),
    .Y(_511_)
);

INVX2 _2430_ (
    .A(_1080_),
    .Y(_136_)
);

AOI22X1 _2010_ (
    .A(_1049_),
    .B(\AXYS[3] [5]),
    .C(\AXYS[2] [5]),
    .D(_1057_),
    .Y(_1122_)
);

FILL FILL_5__2180_ (
);

FILL FILL_7__2198_ (
);

FILL FILL_0__1949_ (
);

FILL FILL_6__2916_ (
);

NOR2X1 _3635_ (
    .A(_1599_),
    .B(_1595_),
    .Y(_1665_)
);

NOR2X1 _3215_ (
    .A(\AXYS[2] [4]),
    .B(_798_),
    .Y(_803_)
);

FILL FILL_1__2592_ (
);

FILL FILL_1__2172_ (
);

FILL FILL_3__2098_ (
);

FILL FILL_2__2908_ (
);

FILL FILL_2__2661_ (
);

FILL FILL_2__2241_ (
);

FILL FILL_4__2587_ (
);

FILL FILL_4__2167_ (
);

FILL FILL_0__2487_ (
);

FILL FILL_6__3454_ (
);

FILL FILL_0__2067_ (
);

FILL FILL_6__3034_ (
);

FILL FILL_2__3026_ (
);

FILL FILL_5__1871_ (
);

INVX1 _2906_ (
    .A(_552_),
    .Y(_553_)
);

FILL FILL_1__1863_ (
);

FILL FILL_7__2830_ (
);

FILL FILL_3__1789_ (
);

FILL FILL_3__2730_ (
);

FILL FILL_3__2310_ (
);

FILL FILL_5__2656_ (
);

FILL FILL_5__2236_ (
);

FILL FILL_1__2648_ (
);

FILL FILL_1__2228_ (
);

FILL FILL_3__3515_ (
);

FILL FILL_6__1940_ (
);

FILL FILL_2__1932_ (
);

FILL FILL_4__1858_ (
);

FILL FILL_0__1758_ (
);

FILL FILL_6__2725_ (
);

DFFSR _3444_ (
    .R(_1__bF$buf1),
    .S(vdd),
    .D(_112_),
    .CLK(clk_bF$buf2),
    .Q(ABH[3])
);

FILL FILL_6__2305_ (
);

OAI21X1 _3024_ (
    .A(reset),
    .B(_645_),
    .C(IRHOLD[0]),
    .Y(_648_)
);

FILL FILL_2__2717_ (
);

FILL FILL_5__3194_ (
);

FILL FILL_1__3186_ (
);

FILL FILL_5__1927_ (
);

FILL FILL_1__1919_ (
);

FILL FILL_2__2890_ (
);

FILL FILL_2__2470_ (
);

FILL FILL_2__2050_ (
);

FILL FILL_4__2396_ (
);

AOI21X1 _1930_ (
    .A(_1045_),
    .B(_1046_),
    .C(_1040_),
    .Y(_1047_)
);

FILL FILL_0__2296_ (
);

FILL FILL_6__3263_ (
);

FILL FILL_2__3675_ (
);

FILL FILL_2__3255_ (
);

OAI22X1 _2715_ (
    .A(_373_),
    .B(_384_),
    .C(_377_),
    .D(_381_),
    .Y(_385_)
);

FILL FILL_5__2885_ (
);

FILL FILL_5__2465_ (
);

FILL FILL_5__2045_ (
);

FILL FILL_1__2877_ (
);

FILL FILL_1__2457_ (
);

FILL FILL_1__2037_ (
);

FILL FILL_7__3004_ (
);

FILL FILL_4_CLKBUF1_insert30 (
);

FILL FILL_4_CLKBUF1_insert31 (
);

FILL FILL_4_CLKBUF1_insert32 (
);

FILL FILL_4_CLKBUF1_insert33 (
);

FILL FILL_4_CLKBUF1_insert34 (
);

FILL FILL_4_CLKBUF1_insert35 (
);

FILL FILL_4_CLKBUF1_insert36 (
);

FILL FILL_0__1987_ (
);

FILL FILL_6__2954_ (
);

NAND2X1 _3673_ (
    .A(ADD[6]),
    .B(_1714__bF$buf0),
    .Y(_1695_)
);

FILL FILL_6__2534_ (
);

OAI21X1 _3253_ (
    .A(state[5]),
    .B(_1272_),
    .C(_1061_),
    .Y(_829_)
);

FILL FILL_6__2114_ (
);

FILL FILL_2__2946_ (
);

FILL FILL_2__2526_ (
);

FILL FILL_2__2106_ (
);

FILL FILL_0__3713_ (
);

FILL FILL_3__1810_ (
);

FILL FILL_6__3492_ (
);

FILL FILL_6__3072_ (
);

FILL FILL_0_BUFX2_insert50 (
);

FILL FILL_0_BUFX2_insert51 (
);

FILL FILL_2__3484_ (
);

FILL FILL_0_BUFX2_insert52 (
);

FILL FILL_0_BUFX2_insert53 (
);

FILL FILL_2__3064_ (
);

FILL FILL_0_BUFX2_insert54 (
);

FILL FILL_0_BUFX2_insert55 (
);

FILL FILL_0_BUFX2_insert56 (
);

FILL FILL_0_BUFX2_insert57 (
);

FILL FILL_0_BUFX2_insert58 (
);

FILL FILL_0_BUFX2_insert59 (
);

FILL FILL_6__1805_ (
);

AOI22X1 _2944_ (
    .A(_571_),
    .B(_1149__bF$buf1),
    .C(_584_),
    .D(_586_),
    .Y(_34_)
);

NAND2X1 _2524_ (
    .A(ADD[0]),
    .B(_209_),
    .Y(_219_)
);

NAND2X1 _2104_ (
    .A(_1172_),
    .B(_1212_),
    .Y(_1213_)
);

FILL FILL_5__2694_ (
);

FILL FILL_5__2274_ (
);

OAI21X1 _3309_ (
    .A(_448_),
    .B(_869_),
    .C(_873_),
    .Y(_112_)
);

FILL FILL_1__2686_ (
);

FILL FILL_7__3653_ (
);

FILL FILL_1__2266_ (
);

FILL FILL_7__3233_ (
);

FILL FILL_3__3553_ (
);

FILL FILL_3__3133_ (
);

FILL FILL_5__3479_ (
);

FILL FILL_5__3059_ (
);

FILL FILL_2__1970_ (
);

FILL FILL_4__1896_ (
);

FILL FILL_0__1796_ (
);

FILL FILL_6__2763_ (
);

NOR2X1 _3482_ (
    .A(alu_op[2]),
    .B(_1725_),
    .Y(_1728_)
);

FILL FILL_6__2343_ (
);

MUX2X1 _3062_ (
    .A(_675_),
    .B(DIMUX[3]),
    .S(_956_),
    .Y(_676_)
);

FILL FILL_2__2755_ (
);

FILL FILL_2__2335_ (
);

FILL FILL_4__3622_ (
);

FILL FILL_4__3202_ (
);

FILL FILL_6__3548_ (
);

FILL FILL_6__3128_ (
);

FILL FILL_0__3522_ (
);

FILL FILL_0__3102_ (
);

FILL FILL_5__1965_ (
);

FILL FILL_1__1957_ (
);

FILL FILL_7__2924_ (
);

FILL FILL_7__2504_ (
);

FILL FILL_3__2824_ (
);

FILL FILL_3__2404_ (
);

FILL FILL_2__3293_ (
);

FILL FILL_3__3609_ (
);

INVX1 _2753_ (
    .A(_351_),
    .Y(_419_)
);

OR2X2 _2333_ (
    .A(_1431_),
    .B(_1439_),
    .Y(_1440_)
);

FILL FILL_5__2083_ (
);

FILL FILL_6__2819_ (
);

OAI22X1 _3538_ (
    .A(_1722_),
    .B(_1554_),
    .C(_1564_),
    .D(_1567_),
    .Y(_1568_)
);

OAI21X1 _3118_ (
    .A(_722_),
    .B(_724_),
    .C(_725_),
    .Y(_69_)
);

FILL FILL_1__2495_ (
);

FILL FILL_1__2075_ (
);

FILL FILL_5__3288_ (
);

FILL FILL_6__2992_ (
);

FILL FILL_6__2572_ (
);

NAND2X1 _3291_ (
    .A(ABL[3]),
    .B(_860_),
    .Y(_864_)
);

FILL FILL_6__2152_ (
);

FILL FILL_2__2984_ (
);

FILL FILL_2__2564_ (
);

FILL FILL_2__2144_ (
);

FILL FILL_4__3011_ (
);

FILL FILL_5__1774_ (
);

OAI21X1 _2809_ (
    .A(_1291_),
    .B(_325_),
    .C(DIMUX[1]),
    .Y(_472_)
);

FILL FILL_1__1766_ (
);

FILL FILL_7__2733_ (
);

FILL FILL_7__2313_ (
);

FILL FILL_3__2633_ (
);

FILL FILL_3__2213_ (
);

FILL FILL_5__2979_ (
);

FILL FILL_5__2559_ (
);

FILL FILL_5__2139_ (
);

FILL FILL_5__3500_ (
);

FILL FILL_6__1843_ (
);

NAND2X1 _2982_ (
    .A(_1348_),
    .B(_606_),
    .Y(_612_)
);

OAI22X1 _2562_ (
    .A(_1013_),
    .B(_201_),
    .C(_251_),
    .D(_199_),
    .Y(_252_)
);

NOR2X1 _2142_ (
    .A(_1160_),
    .B(_1213_),
    .Y(_1251_)
);

FILL FILL_2__1835_ (
);

FILL FILL_4__2702_ (
);

FILL FILL_6__2628_ (
);

DFFSR _3347_ (
    .R(_1__bF$buf6),
    .S(vdd),
    .D(_24_),
    .CLK(clk_bF$buf9),
    .Q(clc)
);

FILL FILL_6__2208_ (
);

FILL FILL_7__3691_ (
);

FILL FILL_0__2602_ (
);

FILL FILL_3__3591_ (
);

FILL FILL_3__3171_ (
);

FILL FILL_5__3097_ (
);

FILL FILL_1__3089_ (
);

FILL FILL_3__1904_ (
);

FILL FILL_6__2381_ (
);

FILL FILL_2__2793_ (
);

FILL FILL_2__2373_ (
);

FILL FILL_4__2299_ (
);

OAI21X1 _1833_ (
    .A(_902__bF$buf1),
    .B(_958_),
    .C(_956_),
    .Y(_959_)
);

FILL FILL_4__3660_ (
);

FILL FILL_4__3240_ (
);

FILL FILL_6__3586_ (
);

FILL FILL_0__2199_ (
);

FILL FILL_6__3166_ (
);

FILL FILL_2__3578_ (
);

FILL FILL_0__3560_ (
);

FILL FILL_2__3158_ (
);

FILL FILL_0__3140_ (
);

OAI21X1 _2618_ (
    .A(_295_),
    .B(_218_),
    .C(_299_),
    .Y(_1741_[13])
);

FILL FILL_1__1995_ (
);

FILL FILL_7__2962_ (
);

FILL FILL_7__2122_ (
);

FILL FILL_3__2862_ (
);

FILL FILL_3__2442_ (
);

FILL FILL_3__2022_ (
);

FILL FILL_5__2788_ (
);

FILL FILL_5__2368_ (
);

BUFX2 BUFX2_insert60 (
    .A(_1714_),
    .Y(_1714__bF$buf3)
);

BUFX2 BUFX2_insert61 (
    .A(_1714_),
    .Y(_1714__bF$buf2)
);

BUFX2 BUFX2_insert62 (
    .A(_1714_),
    .Y(_1714__bF$buf1)
);

BUFX2 BUFX2_insert63 (
    .A(_1714_),
    .Y(_1714__bF$buf0)
);

BUFX2 BUFX2_insert64 (
    .A(_886_),
    .Y(_886__bF$buf6)
);

FILL FILL_1__3301_ (
);

BUFX2 BUFX2_insert65 (
    .A(_886_),
    .Y(_886__bF$buf5)
);

BUFX2 BUFX2_insert66 (
    .A(_886_),
    .Y(_886__bF$buf4)
);

BUFX2 BUFX2_insert67 (
    .A(_886_),
    .Y(_886__bF$buf3)
);

BUFX2 BUFX2_insert68 (
    .A(_886_),
    .Y(_886__bF$buf2)
);

BUFX2 BUFX2_insert69 (
    .A(_886_),
    .Y(_886__bF$buf1)
);

FILL FILL_3__3647_ (
);

FILL FILL_3__3227_ (
);

AOI22X1 _2791_ (
    .A(_408_),
    .B(_453_),
    .C(_450_),
    .D(_454_),
    .Y(_455_)
);

OAI21X1 _2371_ (
    .A(_902__bF$buf2),
    .B(_954_),
    .C(RDY_bF$buf1),
    .Y(_1477_)
);

FILL FILL_4__2931_ (
);

FILL FILL_4__2511_ (
);

FILL FILL_6__2857_ (
);

FILL FILL_6__2437_ (
);

NAND2X1 _3576_ (
    .A(_1605_),
    .B(_1604_),
    .Y(_1606_)
);

FILL FILL_6__2017_ (
);

NAND2X1 _3156_ (
    .A(CO),
    .B(_726_),
    .Y(_759_)
);

FILL FILL_7__3080_ (
);

FILL FILL_2__2849_ (
);

FILL FILL_0__2831_ (
);

FILL FILL_2__2429_ (
);

FILL FILL_0__2411_ (
);

FILL FILL_2__2009_ (
);

FILL FILL_7__1813_ (
);

FILL FILL_0__3616_ (
);

FILL FILL_6__2190_ (
);

FILL FILL_2__2182_ (
);

FILL FILL_3__2918_ (
);

OAI21X1 _2847_ (
    .A(_493_),
    .B(_494_),
    .C(_488_),
    .Y(_508_)
);

INVX1 _2427_ (
    .A(_1337_),
    .Y(_133_)
);

AOI21X1 _2007_ (
    .A(_1082_),
    .B(ADD[4]),
    .C(_1119_),
    .Y(_1120_)
);

FILL FILL_7__2351_ (
);

FILL FILL_3__2671_ (
);

FILL FILL_3__2251_ (
);

FILL FILL_5__2597_ (
);

FILL FILL_5__2177_ (
);

FILL FILL_1__2589_ (
);

FILL FILL_7__3556_ (
);

FILL FILL_1__2169_ (
);

FILL FILL_7__3136_ (
);

FILL FILL_1__3530_ (
);

FILL FILL_1__3110_ (
);

FILL FILL_3__3456_ (
);

FILL FILL_3__3036_ (
);

FILL FILL_6__1881_ (
);

MUX2X1 _2180_ (
    .A(_956_),
    .B(_953_),
    .S(_886__bF$buf4),
    .Y(_1289_)
);

FILL FILL_2__1873_ (
);

FILL FILL_4__1799_ (
);

FILL FILL_4__2740_ (
);

FILL FILL_4__2320_ (
);

FILL FILL_6__2666_ (
);

DFFPOSX1 _3385_ (
    .D(_54_),
    .CLK(clk_bF$buf4),
    .Q(IRHOLD[1])
);

FILL FILL_6__2246_ (
);

FILL FILL_2__2658_ (
);

FILL FILL_0__2640_ (
);

FILL FILL_2__2238_ (
);

FILL FILL_0__2220_ (
);

FILL FILL_4__3525_ (
);

FILL FILL_4__3105_ (
);

FILL FILL169350x18150 (
);

FILL FILL_3__1942_ (
);

FILL FILL_0__3005_ (
);

FILL FILL_5__1868_ (
);

FILL FILL_7__2827_ (
);

FILL FILL_1__2801_ (
);

FILL FILL_3__2727_ (
);

FILL FILL_3__2307_ (
);

NAND2X1 _1871_ (
    .A(_901_),
    .B(_952_),
    .Y(_996_)
);

FILL FILL_2__3196_ (
);

FILL FILL_6__1937_ (
);

OAI21X1 _2656_ (
    .A(_965_),
    .B(_330_),
    .C(_324_),
    .Y(_331_)
);

NAND2X1 _2236_ (
    .A(_929_),
    .B(_1078_),
    .Y(_1344_)
);

FILL FILL_7__2580_ (
);

FILL FILL_0__1911_ (
);

FILL FILL_2__1929_ (
);

FILL FILL_3__2480_ (
);

FILL FILL_3__2060_ (
);

FILL FILL_1__2398_ (
);

FILL FILL_3__3265_ (
);

FILL FILL_6__2895_ (
);

FILL FILL_6__2475_ (
);

OAI21X1 _3194_ (
    .A(_720__bF$buf0),
    .B(_687_),
    .C(\AXYS[1] [2]),
    .Y(_792_)
);

FILL FILL_6__2055_ (
);

FILL FILL_2__2887_ (
);

FILL FILL_2__2467_ (
);

FILL FILL_2__2047_ (
);

NOR3X1 _1927_ (
    .A(_1043_),
    .B(_1023_),
    .C(_1025_),
    .Y(_1044_)
);

FILL FILL_7__1851_ (
);

FILL FILL_3__1751_ (
);

FILL FILL_0__3654_ (
);

FILL FILL_0__3234_ (
);

FILL FILL169950x82950 (
);

FILL FILL_7__2216_ (
);

FILL FILL_1__2610_ (
);

FILL FILL_3__2956_ (
);

FILL FILL_3__2536_ (
);

FILL FILL_3__2116_ (
);

FILL FILL_4__1820_ (
);

FILL FILL_6__1746_ (
);

OR2X2 _2885_ (
    .A(_530_),
    .B(_1366_),
    .Y(_538_)
);

INVX1 _2465_ (
    .A(_149_),
    .Y(_165_)
);

OAI21X1 _2045_ (
    .A(I),
    .B(_1152_),
    .C(_1153_),
    .Y(_1154_)
);

FILL FILL_4__2605_ (
);

FILL FILL_7__3174_ (
);

FILL FILL_0__2925_ (
);

FILL FILL_0__2505_ (
);

FILL FILL_3__3494_ (
);

FILL FILL_3__3074_ (
);

FILL FILL168750x64950 (
);

FILL FILL_3__1807_ (
);

FILL FILL_6__2284_ (
);

FILL FILL_2__2696_ (
);

FILL FILL_2__2276_ (
);

FILL FILL_4__3563_ (
);

FILL FILL_4__3143_ (
);

FILL FILL_6__3489_ (
);

FILL FILL_6__3069_ (
);

FILL FILL_3__1980_ (
);

FILL FILL_0__3463_ (
);

FILL FILL_0__3043_ (
);

FILL FILL_1__1898_ (
);

FILL FILL_7__2445_ (
);

FILL FILL_3__2765_ (
);

FILL FILL_3__2345_ (
);

FILL FILL_5__3632_ (
);

FILL FILL_5__3212_ (
);

FILL FILL_1__3624_ (
);

FILL FILL_1__3204_ (
);

FILL FILL_6__1975_ (
);

NOR2X1 _2694_ (
    .A(_364_),
    .B(_322_),
    .Y(_365_)
);

NAND2X1 _2274_ (
    .A(_1373_),
    .B(_1380_),
    .Y(_1382_)
);

FILL FILL_2__1967_ (
);

FILL FILL_4__2834_ (
);

FILL FILL_4__2414_ (
);

INVX4 _3479_ (
    .A(alu_op[3]),
    .Y(_1725_)
);

NAND2X1 _3059_ (
    .A(D),
    .B(_672_),
    .Y(_673_)
);

FILL FILL_0__2734_ (
);

FILL FILL_6__3701_ (
);

FILL FILL_0__2314_ (
);

FILL FILL_4__3619_ (
);

FILL FILL_0__3519_ (
);

FILL FILL_6__2093_ (
);

FILL FILL_5__2903_ (
);

FILL FILL_2__2085_ (
);

NAND3X1 _1965_ (
    .A(_940_),
    .B(_1077_),
    .C(_1081_),
    .Y(_1082_)
);

FILL FILL_6__3298_ (
);

FILL FILL_0__3692_ (
);

FILL FILL_0__3272_ (
);

FILL FILL_7__2674_ (
);

FILL FILL_7__2254_ (
);

FILL FILL_3__2994_ (
);

FILL FILL_3__2574_ (
);

FILL FILL_3__2154_ (
);

FILL FILL_7__3459_ (
);

FILL FILL_5__3021_ (
);

FILL FILL_1__3013_ (
);

FILL FILL_6__1784_ (
);

AOI22X1 _2083_ (
    .A(_886__bF$buf1),
    .B(_947_),
    .C(_1191_),
    .D(_1150__bF$buf3),
    .Y(_1192_)
);

FILL FILL_5_BUFX2_insert70 (
);

FILL FILL_5_BUFX2_insert71 (
);

FILL FILL_5_BUFX2_insert72 (
);

FILL FILL_5_BUFX2_insert73 (
);

FILL FILL_5_BUFX2_insert74 (
);

FILL FILL_2__1776_ (
);

FILL FILL_5_BUFX2_insert75 (
);

FILL FILL_5_BUFX2_insert76 (
);

FILL FILL_5_BUFX2_insert77 (
);

FILL FILL_5_BUFX2_insert78 (
);

FILL FILL_5_BUFX2_insert79 (
);

FILL FILL_4__2643_ (
);

FILL FILL_4__2223_ (
);

FILL FILL_6__2989_ (
);

FILL FILL_6__2569_ (
);

OAI21X1 _3288_ (
    .A(_231_),
    .B(_860_),
    .C(_862_),
    .Y(_102_)
);

FILL FILL_6__2149_ (
);

FILL FILL_0__2963_ (
);

FILL FILL_0__2543_ (
);

FILL FILL_6__3510_ (
);

FILL FILL_0__2123_ (
);

FILL FILL_2__3502_ (
);

FILL FILL_7__1945_ (
);

FILL FILL_4__3008_ (
);

FILL FILL_3__1845_ (
);

FILL FILL_5__2712_ (
);

FILL FILL_1__2704_ (
);

NOR2X1 _1774_ (
    .A(_899_),
    .B(_898_),
    .Y(_900_)
);

FILL FILL_4__3181_ (
);

FILL FILL_0__3081_ (
);

FILL FILL_2__3099_ (
);

FILL FILL_4__1914_ (
);

NOR2X1 _2979_ (
    .A(_1181_),
    .B(_605_),
    .Y(_609_)
);

INVX1 _2559_ (
    .A(_249_),
    .Y(_1741_[4])
);

NAND3X1 _2139_ (
    .A(_1220_),
    .B(_1247_),
    .C(_1210_),
    .Y(_1248_)
);

FILL FILL_7__2483_ (
);

FILL FILL_7__2063_ (
);

FILL FILL_0__1814_ (
);

NAND2X1 _3500_ (
    .A(AI[4]),
    .B(_1529_),
    .Y(_1530_)
);

FILL FILL_3__2383_ (
);

FILL FILL_5__3670_ (
);

FILL FILL_5__3250_ (
);

FILL FILL_1__3662_ (
);

FILL FILL_1__3242_ (
);

FILL FILL_3__3588_ (
);

FILL FILL_3__3168_ (
);

FILL FILL_4__2872_ (
);

FILL FILL_4__2452_ (
);

FILL FILL_4__2032_ (
);

FILL FILL_6__2798_ (
);

FILL FILL_6__2378_ (
);

NAND3X1 _3097_ (
    .A(_539_),
    .B(_706_),
    .C(_705_),
    .Y(_707_)
);

FILL FILL_0__2772_ (
);

FILL FILL_0__2352_ (
);

FILL FILL_2__3311_ (
);

FILL FILL_4__3657_ (
);

FILL FILL_4__3237_ (
);

FILL FILL_0__3557_ (
);

FILL FILL_0__3137_ (
);

FILL FILL_7__2959_ (
);

FILL FILL_5__2941_ (
);

FILL FILL_5__2521_ (
);

FILL FILL_7__2119_ (
);

FILL FILL_5__2101_ (
);

FILL FILL_1__2933_ (
);

FILL FILL_1__2513_ (
);

FILL FILL_3__2859_ (
);

FILL FILL_3__2439_ (
);

FILL FILL_3__2019_ (
);

FILL FILL_5__3306_ (
);

AOI21X1 _2788_ (
    .A(_430_),
    .B(_438_),
    .C(_451_),
    .Y(_452_)
);

NOR2X1 _2368_ (
    .A(_1473_),
    .B(_1342_),
    .Y(_1474_)
);

FILL FILL_7__2292_ (
);

FILL FILL_3__2192_ (
);

FILL FILL_4__2928_ (
);

FILL FILL_4__2508_ (
);

FILL FILL_7__3077_ (
);

FILL FILL_0__2828_ (
);

FILL FILL_0__2408_ (
);

FILL FILL_1__3471_ (
);

FILL FILL_1__3051_ (
);

FILL FILL_4__2681_ (
);

FILL FILL_4__2261_ (
);

FILL FILL_6__2187_ (
);

FILL FILL_0__2581_ (
);

FILL FILL_2__2599_ (
);

FILL FILL_0__2161_ (
);

FILL FILL_2__2179_ (
);

FILL FILL_2__3540_ (
);

FILL FILL_2__3120_ (
);

FILL FILL_4__3466_ (
);

FILL FILL_4__3046_ (
);

FILL FILL_3__1883_ (
);

FILL FILL_5__2750_ (
);

FILL FILL_5__2330_ (
);

FILL FILL_7__2348_ (
);

FILL FILL_1__2742_ (
);

FILL FILL_1__2322_ (
);

FILL FILL_3__2668_ (
);

FILL FILL_3__2248_ (
);

FILL FILL169950x14550 (
);

FILL FILL_5__3535_ (
);

FILL FILL_5__3115_ (
);

FILL FILL_1__3527_ (
);

FILL FILL_1__3107_ (
);

FILL FILL_4__1952_ (
);

FILL FILL_6__1878_ (
);

OAI21X1 _2597_ (
    .A(_925_),
    .B(_196_),
    .C(ABH[2]),
    .Y(_282_)
);

OAI21X1 _2177_ (
    .A(_914__bF$buf0),
    .B(_949_),
    .C(RDY_bF$buf5),
    .Y(_1286_)
);

FILL FILL_0__1852_ (
);

FILL FILL_2__2811_ (
);

FILL FILL_4__2737_ (
);

FILL FILL_4__2317_ (
);

FILL FILL_0__2637_ (
);

FILL FILL_6__3604_ (
);

FILL FILL_0__2217_ (
);

FILL FILL_1__3280_ (
);

FILL FILL_3__1939_ (
);

FILL FILL_4__2490_ (
);

FILL FILL_4__2070_ (
);

FILL FILL_5__2806_ (
);

FILL FILL_0__2390_ (
);

NOR2X1 _1868_ (
    .A(_934_),
    .B(_907_),
    .Y(_993_)
);

FILL FILL_4__3695_ (
);

FILL FILL_7__1792_ (
);

FILL FILL_4__3275_ (
);

FILL FILL_0__3595_ (
);

FILL FILL_0__3175_ (
);

FILL FILL_7__2577_ (
);

FILL FILL_0__1908_ (
);

FILL FILL_1__2971_ (
);

FILL FILL_1__2551_ (
);

FILL FILL_1__2131_ (
);

FILL FILL_3__2897_ (
);

FILL FILL_3__2477_ (
);

FILL FILL_3__2057_ (
);

FILL FILL_4__1761_ (
);

endmodule
